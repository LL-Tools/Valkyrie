

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9573, n9574, n9575, n9576, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839;

  AOI211_X1 U11006 ( .C1(n10524), .C2(n19639), .A(n19642), .B(n19481), .ZN(
        n19452) );
  NOR2_X1 U11007 ( .A1(n14345), .A2(n14347), .ZN(n14346) );
  CLKBUF_X2 U11008 ( .A(n18400), .Z(n9569) );
  INV_X2 U11009 ( .A(n14777), .ZN(n14764) );
  CLKBUF_X1 U11010 ( .A(n11330), .Z(n11393) );
  NAND2_X1 U11011 ( .A1(n11736), .A2(n11735), .ZN(n11774) );
  AND2_X1 U11012 ( .A1(n14104), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10361) );
  AND2_X1 U11013 ( .A1(n14093), .A2(n10334), .ZN(n14121) );
  AND2_X1 U11014 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10335), .ZN(
        n14122) );
  AND2_X1 U11015 ( .A1(n9589), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10437) );
  BUF_X2 U11016 ( .A(n11215), .Z(n16932) );
  CLKBUF_X2 U11017 ( .A(n14278), .Z(n14295) );
  INV_X2 U11018 ( .A(n16746), .ZN(n16953) );
  INV_X4 U11019 ( .A(n11392), .ZN(n9574) );
  NOR2_X1 U11020 ( .A1(n17546), .A2(n17534), .ZN(n16551) );
  CLKBUF_X3 U11021 ( .A(n11216), .Z(n16899) );
  NAND2_X1 U11022 ( .A1(n9642), .A2(n10686), .ZN(n11130) );
  INV_X2 U11023 ( .A(n10237), .ZN(n10767) );
  CLKBUF_X1 U11024 ( .A(n10214), .Z(n19050) );
  INV_X1 U11025 ( .A(n16696), .ZN(n16933) );
  NOR2_X1 U11026 ( .A1(n11183), .A2(n11182), .ZN(n11268) );
  CLKBUF_X2 U11027 ( .A(n11575), .Z(n13886) );
  CLKBUF_X1 U11028 ( .A(n11716), .Z(n13838) );
  INV_X1 U11029 ( .A(n11655), .ZN(n11675) );
  AND2_X1 U11030 ( .A1(n11587), .A2(n10101), .ZN(n11661) );
  AND2_X1 U11031 ( .A1(n9697), .A2(n11527), .ZN(n11826) );
  AND2_X1 U11032 ( .A1(n12802), .A2(n15559), .ZN(n11695) );
  AND2_X1 U11033 ( .A1(n9697), .A2(n14844), .ZN(n11709) );
  AND2_X2 U11034 ( .A1(n11528), .A2(n12813), .ZN(n11806) );
  CLKBUF_X1 U11035 ( .A(n18288), .Z(n9562) );
  NOR2_X1 U11036 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18224), .ZN(
        n18288) );
  INV_X1 U11037 ( .A(n17941), .ZN(n9563) );
  INV_X1 U11038 ( .A(n9563), .ZN(n9564) );
  AOI221_X1 U11039 ( .B1(n11445), .B2(n11444), .C1(n11443), .C2(n11444), .A(
        n18450), .ZN(n17941) );
  INV_X4 U11040 ( .A(n17852), .ZN(n9578) );
  CLKBUF_X2 U11044 ( .A(n11826), .Z(n13880) );
  AND2_X1 U11045 ( .A1(n9697), .A2(n11526), .ZN(n11576) );
  INV_X1 U11046 ( .A(n11974), .ZN(n12003) );
  NOR2_X1 U11047 ( .A1(n13436), .A2(n13437), .ZN(n15000) );
  INV_X1 U11048 ( .A(n9623), .ZN(n13195) );
  NAND2_X1 U11050 ( .A1(n18551), .A2(n18560), .ZN(n11186) );
  NOR2_X1 U11051 ( .A1(n11185), .A2(n11187), .ZN(n11271) );
  AND4_X1 U11052 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11544) );
  INV_X1 U11053 ( .A(n11130), .ZN(n14022) );
  NAND2_X1 U11054 ( .A1(n10549), .A2(n10548), .ZN(n11168) );
  AND2_X1 U11055 ( .A1(n9568), .A2(n10141), .ZN(n14115) );
  INV_X1 U11056 ( .A(n16746), .ZN(n9591) );
  AND3_X1 U11057 ( .A1(n9942), .A2(n9944), .A3(n9941), .ZN(n17565) );
  INV_X1 U11058 ( .A(n19778), .ZN(n19751) );
  INV_X1 U11059 ( .A(n12929), .ZN(n12528) );
  NOR2_X1 U11060 ( .A1(n14957), .A2(n13537), .ZN(n11015) );
  INV_X1 U11061 ( .A(n10468), .ZN(n13985) );
  NAND2_X1 U11062 ( .A1(n15173), .A2(n15029), .ZN(n13981) );
  NAND2_X1 U11063 ( .A1(n13160), .A2(n11167), .ZN(n13265) );
  BUF_X1 U11064 ( .A(n10222), .Z(n19043) );
  NOR2_X1 U11065 ( .A1(n16599), .A2(n17555), .ZN(n17535) );
  NAND2_X1 U11066 ( .A1(n18568), .A2(n18575), .ZN(n16657) );
  AND2_X1 U11067 ( .A1(n15302), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15268) );
  AND2_X1 U11068 ( .A1(n15340), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15327) );
  INV_X2 U11069 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12581) );
  INV_X1 U11070 ( .A(n10012), .ZN(n10001) );
  NOR2_X1 U11071 ( .A1(n17991), .A2(n17036), .ZN(n17033) );
  INV_X1 U11072 ( .A(n17991), .ZN(n17144) );
  INV_X1 U11073 ( .A(n17460), .ZN(n17473) );
  NOR2_X1 U11075 ( .A1(n18598), .A2(n16314), .ZN(n17612) );
  OR2_X1 U11077 ( .A1(n12420), .A2(n12991), .ZN(n14929) );
  XOR2_X1 U11078 ( .A(n14007), .B(n13987), .Z(n9565) );
  INV_X4 U11079 ( .A(n11661), .ZN(n11767) );
  NAND2_X2 U11080 ( .A1(n10337), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12645) );
  NAND2_X1 U11081 ( .A1(n10467), .A2(n10222), .ZN(n10212) );
  NOR2_X1 U11082 ( .A1(n10222), .A2(n10467), .ZN(n10168) );
  BUF_X4 U11086 ( .A(n10756), .Z(n9567) );
  NAND2_X1 U11087 ( .A1(n10219), .A2(n10217), .ZN(n10756) );
  INV_X2 U11088 ( .A(n10201), .ZN(n10705) );
  AND2_X1 U11089 ( .A1(n9579), .A2(n10141), .ZN(n10344) );
  INV_X1 U11090 ( .A(n12645), .ZN(n9568) );
  INV_X1 U11091 ( .A(n9567), .ZN(n10686) );
  AND2_X2 U11092 ( .A1(n15041), .A2(n9901), .ZN(n13523) );
  OAI22_X2 U11093 ( .A1(n12770), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11817), 
        .B2(n11800), .ZN(n11706) );
  NAND2_X4 U11094 ( .A1(n10100), .A2(n11544), .ZN(n19994) );
  AOI21_X1 U11095 ( .B1(n18389), .B2(n18415), .A(n18388), .ZN(n18400) );
  NOR3_X2 U11096 ( .A1(n17076), .A2(n17043), .A3(n16999), .ZN(n17037) );
  NOR2_X2 U11097 ( .A1(n18403), .A2(n18411), .ZN(n17836) );
  AOI21_X2 U11098 ( .B1(n11318), .B2(n10075), .A(n11317), .ZN(n12132) );
  AND2_X2 U11099 ( .A1(n10170), .A2(n10168), .ZN(n10718) );
  NOR2_X2 U11100 ( .A1(n14401), .A2(n13747), .ZN(n14391) );
  AOI21_X2 U11101 ( .B1(n11286), .B2(n9948), .A(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9947) );
  NOR2_X2 U11102 ( .A1(n16539), .A2(n17483), .ZN(n16492) );
  NAND2_X2 U11103 ( .A1(n9696), .A2(n9695), .ZN(n10222) );
  NAND2_X2 U11104 ( .A1(n10139), .A2(n10140), .ZN(n10214) );
  OAI21_X2 U11105 ( .B1(n15342), .B2(n15344), .A(n15048), .ZN(n15325) );
  NAND2_X2 U11106 ( .A1(n15052), .A2(n15051), .ZN(n15342) );
  NAND2_X2 U11107 ( .A1(n10803), .A2(n19639), .ZN(n10827) );
  XNOR2_X2 U11108 ( .A(n10485), .B(n10484), .ZN(n11140) );
  BUF_X4 U11109 ( .A(n9574), .Z(n9571) );
  NAND2_X1 U11110 ( .A1(n14625), .A2(n14634), .ZN(n14626) );
  AOI211_X1 U11111 ( .C1(n16358), .C2(n18452), .A(n16357), .B(n16356), .ZN(
        n16361) );
  AND3_X1 U11112 ( .A1(n13227), .A2(n9681), .A3(n13228), .ZN(n13409) );
  AOI21_X1 U11113 ( .B1(n10053), .B2(n9693), .A(n9648), .ZN(n10055) );
  AND2_X1 U11114 ( .A1(n9979), .A2(n17275), .ZN(n16380) );
  NOR2_X1 U11115 ( .A1(n12137), .A2(n17627), .ZN(n17524) );
  AND2_X1 U11116 ( .A1(n11299), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11301) );
  NAND2_X1 U11118 ( .A1(n11764), .A2(n11757), .ZN(n12510) );
  NAND2_X2 U11119 ( .A1(n10303), .A2(n9636), .ZN(n10423) );
  CLKBUF_X1 U11120 ( .A(n12251), .Z(n19970) );
  NAND2_X1 U11121 ( .A1(n9630), .A2(n9699), .ZN(n12814) );
  BUF_X1 U11122 ( .A(n10295), .Z(n9598) );
  BUF_X1 U11123 ( .A(n10294), .Z(n10297) );
  NOR2_X1 U11124 ( .A1(n16483), .A2(n10012), .ZN(n16475) );
  XNOR2_X1 U11125 ( .A(n11039), .B(n11040), .ZN(n10279) );
  NAND2_X1 U11126 ( .A1(n10267), .A2(n10266), .ZN(n11040) );
  AND2_X1 U11127 ( .A1(n9893), .A2(n9898), .ZN(n9897) );
  NOR2_X1 U11128 ( .A1(n11019), .A2(n10237), .ZN(n12585) );
  INV_X4 U11130 ( .A(n19683), .ZN(n9573) );
  NAND3_X2 U11131 ( .A1(n11653), .A2(n11652), .A3(n9750), .ZN(n19985) );
  AND2_X1 U11132 ( .A1(n10150), .A2(n10151), .ZN(n10202) );
  CLKBUF_X1 U11133 ( .A(n11661), .Z(n11937) );
  AND2_X2 U11134 ( .A1(n9579), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10432) );
  CLKBUF_X2 U11135 ( .A(n11806), .Z(n9594) );
  CLKBUF_X2 U11137 ( .A(n11709), .Z(n13937) );
  CLKBUF_X2 U11138 ( .A(n11710), .Z(n13821) );
  CLKBUF_X2 U11139 ( .A(n11576), .Z(n13878) );
  CLKBUF_X2 U11140 ( .A(n11574), .Z(n13806) );
  BUF_X2 U11141 ( .A(n11241), .Z(n16799) );
  INV_X8 U11142 ( .A(n16864), .ZN(n9575) );
  CLKBUF_X2 U11143 ( .A(n11241), .Z(n16952) );
  NOR2_X1 U11144 ( .A1(n16657), .A2(n11187), .ZN(n16845) );
  CLKBUF_X2 U11145 ( .A(n11695), .Z(n13881) );
  CLKBUF_X2 U11146 ( .A(n11597), .Z(n13887) );
  NOR2_X2 U11147 ( .A1(n11184), .A2(n11182), .ZN(n11215) );
  AND2_X1 U11148 ( .A1(n11528), .A2(n14844), .ZN(n13682) );
  NAND2_X1 U11149 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11187) );
  OAI21_X1 U11150 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(n14861) );
  OR2_X1 U11151 ( .A1(n14230), .A2(n14229), .ZN(n14231) );
  OR2_X1 U11152 ( .A1(n14206), .A2(n14205), .ZN(n10080) );
  NOR2_X1 U11153 ( .A1(n9807), .A2(n9806), .ZN(n16041) );
  AND2_X1 U11154 ( .A1(n14391), .A2(n9868), .ZN(n14355) );
  AOI21_X1 U11155 ( .B1(n15945), .B2(n16150), .A(n15138), .ZN(n15139) );
  OR2_X1 U11156 ( .A1(n11016), .A2(n14934), .ZN(n15969) );
  AND2_X1 U11157 ( .A1(n9843), .A2(n11910), .ZN(n14671) );
  INV_X1 U11158 ( .A(n9900), .ZN(n15952) );
  NOR2_X1 U11159 ( .A1(n14700), .A2(n9701), .ZN(n13484) );
  AND2_X1 U11160 ( .A1(n13261), .A2(n13262), .ZN(n10053) );
  AND2_X1 U11161 ( .A1(n13485), .A2(n11908), .ZN(n14685) );
  NAND2_X1 U11162 ( .A1(n13485), .A2(n9629), .ZN(n14700) );
  OR2_X1 U11163 ( .A1(n14699), .A2(n14695), .ZN(n9701) );
  NOR2_X2 U11164 ( .A1(n9622), .A2(n14924), .ZN(n14925) );
  OR2_X1 U11165 ( .A1(n11168), .A2(n9804), .ZN(n11171) );
  AND2_X1 U11166 ( .A1(n11881), .A2(n11880), .ZN(n13063) );
  AND2_X1 U11167 ( .A1(n11160), .A2(n11159), .ZN(n16110) );
  OR2_X1 U11168 ( .A1(n11160), .A2(n11159), .ZN(n11164) );
  NAND2_X1 U11169 ( .A1(n12837), .A2(n12844), .ZN(n12836) );
  NAND2_X1 U11170 ( .A1(n10504), .A2(n10503), .ZN(n12724) );
  OR2_X1 U11171 ( .A1(n11876), .A2(n11875), .ZN(n11897) );
  OAI21_X1 U11172 ( .B1(n19969), .B2(n13607), .A(n12880), .ZN(n12881) );
  NAND2_X1 U11173 ( .A1(n13385), .A2(n13384), .ZN(n13436) );
  NOR2_X2 U11174 ( .A1(n17118), .A2(n17627), .ZN(n17516) );
  INV_X1 U11175 ( .A(n17623), .ZN(n17582) );
  AND2_X1 U11176 ( .A1(n13207), .A2(n13248), .ZN(n13385) );
  OR2_X1 U11177 ( .A1(n11816), .A2(n11841), .ZN(n19969) );
  AND2_X1 U11178 ( .A1(n10445), .A2(n10444), .ZN(n10446) );
  NOR2_X1 U11179 ( .A1(n11153), .A2(n11152), .ZN(n10447) );
  NAND2_X1 U11180 ( .A1(n10547), .A2(n10546), .ZN(n11161) );
  CLKBUF_X1 U11181 ( .A(n17615), .Z(n9599) );
  OAI21_X1 U11182 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18605), .A(n16314), 
        .ZN(n17623) );
  AOI21_X1 U11183 ( .B1(n17447), .B2(n11296), .A(n17454), .ZN(n11303) );
  AND3_X1 U11184 ( .A1(n9737), .A2(n10421), .A3(n9651), .ZN(n9736) );
  NAND2_X1 U11185 ( .A1(n11298), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17452) );
  NOR2_X1 U11186 ( .A1(n17256), .A2(n17081), .ZN(n17077) );
  AOI21_X1 U11187 ( .B1(n10369), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A(n9735), .ZN(n9737) );
  OR2_X1 U11188 ( .A1(n13270), .A2(n9880), .ZN(n16134) );
  NOR2_X1 U11189 ( .A1(n17513), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17493) );
  XNOR2_X1 U11190 ( .A(n12510), .B(n12511), .ZN(n20053) );
  INV_X1 U11191 ( .A(n9952), .ZN(n17541) );
  AND2_X1 U11192 ( .A1(n12543), .A2(n12977), .ZN(n12556) );
  AOI211_X1 U11193 ( .C1(n10407), .C2(n19639), .A(n19642), .B(n19278), .ZN(
        n19252) );
  AND2_X1 U11194 ( .A1(n10296), .A2(n9598), .ZN(n10524) );
  INV_X1 U11196 ( .A(n10514), .ZN(n19022) );
  AND2_X1 U11197 ( .A1(n12464), .A2(n12544), .ZN(n12469) );
  AND2_X1 U11198 ( .A1(n12468), .A2(n12467), .ZN(n12470) );
  NOR2_X2 U11199 ( .A1(n10320), .A2(n10319), .ZN(n19308) );
  NAND2_X1 U11200 ( .A1(n10308), .A2(n9734), .ZN(n10418) );
  NAND2_X1 U11201 ( .A1(n10303), .A2(n10305), .ZN(n10516) );
  NAND2_X1 U11202 ( .A1(n10308), .A2(n10305), .ZN(n10426) );
  AND2_X1 U11203 ( .A1(n10308), .A2(n9608), .ZN(n19149) );
  NOR2_X2 U11204 ( .A1(n18919), .A2(n19496), .ZN(n13050) );
  OR2_X2 U11205 ( .A1(n12532), .A2(n12340), .ZN(n10320) );
  NOR2_X2 U11206 ( .A1(n18928), .A2(n19496), .ZN(n13025) );
  NOR2_X2 U11207 ( .A1(n19029), .A2(n19496), .ZN(n19030) );
  NOR2_X2 U11208 ( .A1(n19034), .A2(n19496), .ZN(n19035) );
  XNOR2_X1 U11209 ( .A(n12814), .B(n20134), .ZN(n20255) );
  NAND2_X1 U11210 ( .A1(n9847), .A2(n11761), .ZN(n12511) );
  INV_X2 U11211 ( .A(n15728), .ZN(n9576) );
  NAND2_X2 U11212 ( .A1(n19797), .A2(n20015), .ZN(n14530) );
  AND2_X1 U11213 ( .A1(n9976), .A2(n9975), .ZN(n16464) );
  XNOR2_X1 U11214 ( .A(n9798), .B(n10292), .ZN(n12456) );
  OR2_X1 U11215 ( .A1(n16313), .A2(n11488), .ZN(n9933) );
  NAND2_X1 U11216 ( .A1(n10286), .A2(n10287), .ZN(n10293) );
  XNOR2_X1 U11217 ( .A(n10261), .B(n9897), .ZN(n10294) );
  AOI21_X1 U11218 ( .B1(n11794), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11685), .ZN(n11689) );
  OR2_X1 U11219 ( .A1(n11684), .A2(n11683), .ZN(n11688) );
  OR2_X1 U11220 ( .A1(n10291), .A2(n11033), .ZN(n10278) );
  NAND2_X1 U11221 ( .A1(n9690), .A2(n10225), .ZN(n10261) );
  OR2_X1 U11222 ( .A1(n12434), .A2(n12433), .ZN(n12436) );
  NAND2_X1 U11223 ( .A1(n10276), .A2(n10275), .ZN(n11033) );
  NOR2_X1 U11224 ( .A1(n11490), .A2(n11486), .ZN(n11489) );
  INV_X2 U11225 ( .A(n12176), .ZN(n10012) );
  INV_X2 U11226 ( .A(n14026), .ZN(n13995) );
  OR2_X2 U11227 ( .A1(n18975), .A2(n18973), .ZN(n12392) );
  NAND2_X1 U11228 ( .A1(n10273), .A2(n10272), .ZN(n10291) );
  NAND2_X1 U11229 ( .A1(n12984), .A2(n9872), .ZN(n10821) );
  NAND2_X1 U11230 ( .A1(n11480), .A2(n11479), .ZN(n11490) );
  AND2_X1 U11231 ( .A1(n11483), .A2(n11497), .ZN(n11480) );
  NOR3_X1 U11232 ( .A1(n17144), .A2(n15416), .A3(n15612), .ZN(n11493) );
  NOR2_X2 U11233 ( .A1(n16333), .A2(n17270), .ZN(n16198) );
  NOR3_X1 U11234 ( .A1(n18390), .A2(n11485), .A3(n17969), .ZN(n11478) );
  CLKBUF_X1 U11235 ( .A(n11017), .Z(n12681) );
  AND2_X1 U11236 ( .A1(n12268), .A2(n10227), .ZN(n10232) );
  NAND2_X1 U11237 ( .A1(n12220), .A2(n12693), .ZN(n11017) );
  NOR2_X1 U11238 ( .A1(n16337), .A2(n17304), .ZN(n17285) );
  NOR2_X1 U11239 ( .A1(n17613), .A2(n11281), .ZN(n17604) );
  MUX2_X1 U11240 ( .A(n10230), .B(n10811), .S(n10759), .Z(n10231) );
  INV_X1 U11241 ( .A(n20669), .ZN(n19826) );
  AND2_X1 U11242 ( .A1(n10686), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10242) );
  INV_X1 U11243 ( .A(n12771), .ZN(n9721) );
  AND2_X1 U11244 ( .A1(n10220), .A2(n19050), .ZN(n10803) );
  NOR2_X1 U11245 ( .A1(n17345), .A2(n17346), .ZN(n17328) );
  XNOR2_X1 U11246 ( .A(n11451), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11452) );
  NAND2_X1 U11247 ( .A1(n12691), .A2(n10226), .ZN(n10761) );
  NOR2_X1 U11248 ( .A1(n10200), .A2(n10212), .ZN(n10218) );
  NOR2_X1 U11249 ( .A1(n17137), .A2(n11451), .ZN(n11450) );
  CLKBUF_X1 U11250 ( .A(n11673), .Z(n11999) );
  INV_X1 U11251 ( .A(n12367), .ZN(n19690) );
  INV_X1 U11252 ( .A(n10705), .ZN(n13054) );
  INV_X1 U11253 ( .A(n10219), .ZN(n10226) );
  NAND2_X1 U11254 ( .A1(n12345), .A2(n10467), .ZN(n10229) );
  AND3_X1 U11255 ( .A1(n12481), .A2(n11937), .A3(n12482), .ZN(n12381) );
  NAND2_X1 U11256 ( .A1(n10712), .A2(n10221), .ZN(n10237) );
  AND2_X1 U11257 ( .A1(n19043), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12341) );
  NOR2_X1 U11258 ( .A1(n16266), .A2(n16225), .ZN(n16268) );
  NAND3_X1 U11259 ( .A1(n11402), .A2(n11401), .A3(n11400), .ZN(n17960) );
  CLKBUF_X1 U11260 ( .A(n11702), .Z(n19999) );
  INV_X1 U11261 ( .A(n11702), .ZN(n12482) );
  AND2_X1 U11262 ( .A1(n11655), .A2(n20015), .ZN(n12494) );
  BUF_X2 U11263 ( .A(n10467), .Z(n10468) );
  INV_X1 U11264 ( .A(n19985), .ZN(n19827) );
  NAND2_X1 U11265 ( .A1(n10186), .A2(n10185), .ZN(n10219) );
  INV_X1 U11266 ( .A(n10704), .ZN(n10712) );
  CLKBUF_X1 U11267 ( .A(n10202), .Z(n10759) );
  NOR2_X1 U11268 ( .A1(n10704), .A2(n10201), .ZN(n9733) );
  INV_X2 U11269 ( .A(n10217), .ZN(n12691) );
  INV_X1 U11270 ( .A(n10202), .ZN(n10221) );
  INV_X2 U11271 ( .A(U214), .ZN(n16266) );
  NAND4_X1 U11272 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11702) );
  NAND2_X1 U11273 ( .A1(n10126), .A2(n10125), .ZN(n10467) );
  NAND2_X2 U11274 ( .A1(n10199), .A2(n9892), .ZN(n10217) );
  AND4_X1 U11275 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n11610) );
  AND4_X1 U11276 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(
        n11609) );
  AND4_X1 U11277 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(
        n11573) );
  AND4_X1 U11278 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n11630) );
  AND4_X1 U11279 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11631) );
  AND4_X1 U11280 ( .A1(n11616), .A2(n11615), .A3(n11614), .A4(n11613), .ZN(
        n11632) );
  AND2_X1 U11281 ( .A1(n11650), .A2(n11651), .ZN(n9750) );
  AND4_X1 U11282 ( .A1(n11641), .A2(n11640), .A3(n11639), .A4(n11638), .ZN(
        n11652) );
  AND4_X1 U11283 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11608) );
  NAND2_X1 U11284 ( .A1(n10198), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9892) );
  NAND2_X1 U11285 ( .A1(n10193), .A2(n10141), .ZN(n10199) );
  NAND4_X2 U11286 ( .A1(n11563), .A2(n11562), .A3(n10082), .A4(n11561), .ZN(
        n20015) );
  AND4_X1 U11287 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(
        n10100) );
  AND2_X1 U11288 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n9779) );
  OR2_X1 U11289 ( .A1(n11715), .A2(n11592), .ZN(n11596) );
  AND4_X1 U11290 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11607) );
  AOI21_X1 U11291 ( .B1(n11710), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n11564), .ZN(n11568) );
  AND4_X1 U11292 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n11587) );
  AND4_X1 U11293 ( .A1(n11628), .A2(n11627), .A3(n11626), .A4(n11625), .ZN(
        n11629) );
  INV_X2 U11294 ( .A(n11194), .ZN(n16926) );
  AND4_X1 U11295 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11653) );
  AND4_X1 U11296 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n11650) );
  AND4_X1 U11297 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11651) );
  AND2_X2 U11298 ( .A1(n14295), .A2(n10141), .ZN(n14120) );
  AND2_X2 U11299 ( .A1(n14297), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10864) );
  AND2_X2 U11300 ( .A1(n14297), .A2(n10141), .ZN(n14114) );
  AND2_X1 U11301 ( .A1(n10172), .A2(n10171), .ZN(n10176) );
  AND2_X1 U11302 ( .A1(n10179), .A2(n10178), .ZN(n10183) );
  INV_X2 U11303 ( .A(n11715), .ZN(n13861) );
  AND3_X1 U11304 ( .A1(n9802), .A2(n9801), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10149) );
  AND3_X1 U11305 ( .A1(n9964), .A2(n9963), .A3(n10141), .ZN(n10145) );
  AND4_X1 U11306 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n11563) );
  AND4_X1 U11307 ( .A1(n11552), .A2(n11551), .A3(n11550), .A4(n11549), .ZN(
        n11562) );
  AND4_X1 U11308 ( .A1(n11560), .A2(n11559), .A3(n11558), .A4(n11557), .ZN(
        n11561) );
  AND4_X1 U11309 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(
        n10082) );
  INV_X2 U11310 ( .A(n16298), .ZN(U215) );
  INV_X1 U11311 ( .A(n13682), .ZN(n11715) );
  CLKBUF_X1 U11312 ( .A(n14091), .Z(n14092) );
  AND2_X1 U11313 ( .A1(n9592), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11564) );
  BUF_X2 U11314 ( .A(n10329), .Z(n14297) );
  INV_X1 U11315 ( .A(n16845), .ZN(n16746) );
  CLKBUF_X3 U11316 ( .A(n11323), .Z(n16934) );
  INV_X1 U11317 ( .A(n11270), .ZN(n11392) );
  NAND2_X1 U11318 ( .A1(n9773), .A2(n9772), .ZN(n16696) );
  INV_X2 U11319 ( .A(n11251), .ZN(n15502) );
  NOR2_X1 U11320 ( .A1(n11184), .A2(n11185), .ZN(n11216) );
  NOR2_X1 U11321 ( .A1(n16657), .A2(n11186), .ZN(n11270) );
  OR2_X2 U11322 ( .A1(n11183), .A2(n16657), .ZN(n11251) );
  NOR2_X1 U11323 ( .A1(n18392), .A2(n11186), .ZN(n11330) );
  INV_X2 U11324 ( .A(n16303), .ZN(n16305) );
  AND2_X2 U11325 ( .A1(n11526), .A2(n11529), .ZN(n11574) );
  INV_X2 U11326 ( .A(n19695), .ZN(n19613) );
  NAND2_X1 U11327 ( .A1(n18396), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n18420) );
  NAND2_X1 U11328 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18457), .ZN(n16659) );
  BUF_X4 U11329 ( .A(n10128), .Z(n9579) );
  NAND2_X1 U11330 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18551), .ZN(
        n11184) );
  INV_X1 U11331 ( .A(n12205), .ZN(n9926) );
  NAND2_X1 U11332 ( .A1(n18560), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11183) );
  NAND2_X1 U11333 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18575), .ZN(
        n11182) );
  AND2_X1 U11334 ( .A1(n12648), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12650) );
  AND2_X1 U11335 ( .A1(n11520), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11526) );
  AND2_X1 U11336 ( .A1(n11519), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11527) );
  AND2_X1 U11337 ( .A1(n9710), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9697) );
  INV_X1 U11338 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18568) );
  NAND2_X1 U11339 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18392) );
  AND2_X1 U11340 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11525) );
  AND3_X1 U11341 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12802) );
  NOR2_X2 U11342 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11529) );
  NAND2_X1 U11343 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12205) );
  NOR2_X1 U11344 ( .A1(n13006), .A2(n10034), .ZN(n9580) );
  AND2_X1 U11345 ( .A1(n9581), .A2(n12626), .ZN(n12750) );
  NOR2_X1 U11346 ( .A1(n12867), .A2(n12624), .ZN(n9581) );
  NOR2_X1 U11347 ( .A1(n13006), .A2(n10034), .ZN(n13468) );
  NAND2_X1 U11348 ( .A1(n12750), .A2(n12749), .ZN(n13006) );
  AND2_X1 U11349 ( .A1(n10293), .A2(n10290), .ZN(n12340) );
  NOR2_X1 U11350 ( .A1(n11309), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16206) );
  NAND2_X1 U11351 ( .A1(n10048), .A2(n10045), .ZN(n9582) );
  NAND2_X1 U11352 ( .A1(n12902), .A2(n9586), .ZN(n9583) );
  AND2_X2 U11353 ( .A1(n9583), .A2(n9584), .ZN(n15785) );
  OR2_X1 U11354 ( .A1(n9585), .A2(n19903), .ZN(n9584) );
  INV_X1 U11355 ( .A(n11840), .ZN(n9585) );
  AND2_X1 U11356 ( .A1(n11821), .A2(n11840), .ZN(n9586) );
  NAND2_X1 U11357 ( .A1(n9587), .A2(n10042), .ZN(n11764) );
  NOR2_X1 U11358 ( .A1(n11755), .A2(n11740), .ZN(n9587) );
  NAND2_X1 U11359 ( .A1(n10048), .A2(n10045), .ZN(n14708) );
  NAND2_X2 U11360 ( .A1(n15738), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11920) );
  AND2_X2 U11361 ( .A1(n10336), .A2(n12581), .ZN(n9588) );
  AND2_X2 U11362 ( .A1(n10336), .A2(n12581), .ZN(n9589) );
  NOR2_X1 U11363 ( .A1(n9722), .A2(n9721), .ZN(n9720) );
  NAND3_X2 U11364 ( .A1(n9602), .A2(n9707), .A3(n9708), .ZN(n11662) );
  OR2_X1 U11365 ( .A1(n11186), .A2(n11182), .ZN(n10095) );
  OAI21_X2 U11366 ( .B1(n15015), .B2(n15018), .A(n10090), .ZN(n14018) );
  NAND2_X1 U11367 ( .A1(n19827), .A2(n19972), .ZN(n20669) );
  AND2_X4 U11368 ( .A1(n12802), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11582) );
  OAI21_X2 U11370 ( .B1(n13981), .B2(n10062), .A(n10060), .ZN(n14007) );
  AND2_X1 U11371 ( .A1(n11528), .A2(n14844), .ZN(n9592) );
  AND2_X1 U11372 ( .A1(n11528), .A2(n14844), .ZN(n9593) );
  XNOR2_X2 U11373 ( .A(n10509), .B(n11159), .ZN(n16108) );
  OR2_X1 U11374 ( .A1(n12246), .A2(n12025), .ZN(n12771) );
  NAND2_X2 U11375 ( .A1(n10483), .A2(n18811), .ZN(n10509) );
  NAND3_X2 U11376 ( .A1(n11379), .A2(n11378), .A3(n11377), .ZN(n17991) );
  INV_X1 U11377 ( .A(n17192), .ZN(n18598) );
  NOR2_X2 U11378 ( .A1(n11329), .A2(n11328), .ZN(n17192) );
  OAI21_X2 U11379 ( .B1(n15325), .B2(n10634), .A(n10633), .ZN(n15201) );
  NAND2_X2 U11380 ( .A1(n11975), .A2(n19827), .ZN(n12484) );
  NOR2_X4 U11381 ( .A1(n11664), .A2(n10098), .ZN(n11975) );
  AND2_X2 U11382 ( .A1(n12479), .A2(n12484), .ZN(n9602) );
  OR2_X1 U11383 ( .A1(n12532), .A2(n10316), .ZN(n10317) );
  AND2_X1 U11384 ( .A1(n12532), .A2(n12456), .ZN(n10308) );
  OR2_X1 U11385 ( .A1(n12532), .A2(n10314), .ZN(n10315) );
  AND2_X1 U11386 ( .A1(n10318), .A2(n12532), .ZN(n10303) );
  OAI21_X1 U11387 ( .B1(n12532), .B2(n12538), .A(n12537), .ZN(n12547) );
  NAND3_X4 U11388 ( .A1(n9797), .A2(n10284), .A3(n9796), .ZN(n12532) );
  XNOR2_X1 U11389 ( .A(n11820), .B(n19943), .ZN(n12904) );
  OAI211_X1 U11390 ( .C1(n11019), .C2(n10236), .A(n10235), .B(n10234), .ZN(
        n9596) );
  NAND2_X1 U11391 ( .A1(n12720), .A2(n11791), .ZN(n11820) );
  XNOR2_X1 U11392 ( .A(n10293), .B(n10297), .ZN(n10295) );
  OAI211_X2 U11393 ( .C1(n15787), .C2(n9728), .A(n15778), .B(n9726), .ZN(
        n13330) );
  OAI22_X2 U11394 ( .A1(n12835), .A2(n12834), .B1(n10508), .B2(n12844), .ZN(
        n16109) );
  AOI211_X2 U11395 ( .C1(n14742), .C2(n14741), .A(n14740), .B(n14739), .ZN(
        n14743) );
  XNOR2_X2 U11396 ( .A(n11708), .B(n11707), .ZN(n12253) );
  NAND3_X2 U11397 ( .A1(n10044), .A2(n11671), .A3(n9716), .ZN(n11708) );
  NAND2_X1 U11398 ( .A1(n9706), .A2(n9705), .ZN(n11876) );
  NOR3_X1 U11399 ( .A1(n12854), .A2(n9616), .A3(n11852), .ZN(n9705) );
  AOI21_X1 U11400 ( .B1(n20058), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11927), .ZN(n11926) );
  NAND2_X1 U11401 ( .A1(n11801), .A2(n11800), .ZN(n11936) );
  INV_X1 U11402 ( .A(n12494), .ZN(n11990) );
  INV_X1 U11403 ( .A(n11815), .ZN(n9706) );
  INV_X1 U11404 ( .A(n10467), .ZN(n10127) );
  NAND2_X1 U11405 ( .A1(n19994), .A2(n19985), .ZN(n12025) );
  AND2_X1 U11407 ( .A1(n19985), .A2(n19972), .ZN(n12929) );
  NAND2_X1 U11408 ( .A1(n11993), .A2(n11992), .ZN(n12018) );
  NAND2_X1 U11409 ( .A1(n11662), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11684) );
  NAND2_X1 U11410 ( .A1(n20255), .A2(n20571), .ZN(n11814) );
  CLKBUF_X1 U11411 ( .A(n11988), .Z(n12784) );
  XNOR2_X1 U11412 ( .A(n10478), .B(n10475), .ZN(n10720) );
  OR2_X1 U11413 ( .A1(n10564), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10565) );
  NOR2_X1 U11414 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14093) );
  NAND2_X1 U11415 ( .A1(n10029), .A2(n10030), .ZN(n14181) );
  NAND2_X1 U11416 ( .A1(n14892), .A2(n9619), .ZN(n10030) );
  NOR2_X1 U11417 ( .A1(n12564), .A2(n9971), .ZN(n9970) );
  INV_X1 U11418 ( .A(n12550), .ZN(n9971) );
  AND4_X1 U11419 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(
        n10461) );
  OAI21_X1 U11420 ( .B1(n11140), .B2(n12727), .A(n11151), .ZN(n11156) );
  INV_X1 U11421 ( .A(n10241), .ZN(n9898) );
  NAND2_X1 U11422 ( .A1(n10810), .A2(n10226), .ZN(n10978) );
  AOI22_X1 U11423 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15525), .B1(
        n11406), .B2(n18551), .ZN(n11416) );
  NOR2_X1 U11424 ( .A1(n11406), .A2(n18551), .ZN(n11415) );
  NAND2_X1 U11425 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18404), .ZN(
        n11410) );
  INV_X2 U11426 ( .A(n11194), .ZN(n16944) );
  NOR2_X1 U11427 ( .A1(n17121), .A2(n11290), .ZN(n11262) );
  AND2_X1 U11428 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11291), .ZN(
        n11292) );
  NOR2_X1 U11429 ( .A1(n20015), .A2(n20573), .ZN(n12512) );
  AND2_X1 U11430 ( .A1(n20573), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13953) );
  NOR2_X1 U11431 ( .A1(n9862), .A2(n14328), .ZN(n9861) );
  INV_X1 U11432 ( .A(n13903), .ZN(n9862) );
  NAND2_X1 U11433 ( .A1(n14346), .A2(n13903), .ZN(n14327) );
  NAND2_X1 U11434 ( .A1(n12040), .A2(n12114), .ZN(n12121) );
  OR2_X1 U11435 ( .A1(n15737), .A2(n9715), .ZN(n9609) );
  INV_X1 U11436 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9714) );
  OAI21_X1 U11437 ( .B1(n14613), .B2(n14615), .A(n15769), .ZN(n14634) );
  INV_X1 U11438 ( .A(n12018), .ZN(n12126) );
  NAND2_X1 U11439 ( .A1(n9791), .A2(n11962), .ZN(n12822) );
  OAI21_X1 U11440 ( .B1(n11960), .B2(n11959), .A(n9792), .ZN(n9791) );
  NAND2_X1 U11441 ( .A1(n10696), .A2(n10695), .ZN(n10737) );
  NAND2_X1 U11442 ( .A1(n12555), .A2(n10039), .ZN(n10038) );
  NOR2_X1 U11443 ( .A1(n12548), .A2(n10040), .ZN(n10039) );
  INV_X1 U11444 ( .A(n12546), .ZN(n10040) );
  INV_X1 U11445 ( .A(n16174), .ZN(n12989) );
  NAND2_X1 U11446 ( .A1(n12683), .A2(n9573), .ZN(n12574) );
  AND2_X1 U11447 ( .A1(n9632), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15021) );
  AND2_X1 U11448 ( .A1(n11014), .A2(n14933), .ZN(n9876) );
  NAND2_X1 U11449 ( .A1(n10647), .A2(n9652), .ZN(n9748) );
  AND2_X1 U11450 ( .A1(n15039), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15175) );
  NAND2_X1 U11451 ( .A1(n11038), .A2(n10281), .ZN(n9965) );
  NAND2_X1 U11452 ( .A1(n17471), .A2(n9936), .ZN(n16177) );
  INV_X1 U11453 ( .A(n12133), .ZN(n9936) );
  AND2_X1 U11454 ( .A1(n14677), .A2(n12714), .ZN(n19916) );
  AND2_X1 U11455 ( .A1(n19824), .A2(n15572), .ZN(n19917) );
  OR2_X1 U11456 ( .A1(n14313), .A2(n13998), .ZN(n15146) );
  AND2_X1 U11457 ( .A1(n13997), .A2(n13996), .ZN(n13998) );
  NAND2_X1 U11458 ( .A1(n9606), .A2(n19827), .ZN(n9723) );
  NAND2_X1 U11459 ( .A1(n11659), .A2(n11972), .ZN(n9708) );
  NAND2_X1 U11460 ( .A1(n11936), .A2(n11941), .ZN(n9790) );
  AOI22_X1 U11461 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11937), .B1(n11936), 
        .B2(n19985), .ZN(n11948) );
  NAND2_X1 U11462 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10171) );
  NAND2_X1 U11463 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n10072) );
  NAND2_X1 U11464 ( .A1(n19149), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n9689) );
  AOI22_X1 U11465 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10329), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10165) );
  BUF_X1 U11466 ( .A(n11612), .Z(n13843) );
  NAND2_X1 U11467 ( .A1(n20571), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9795) );
  NAND2_X1 U11468 ( .A1(n10474), .A2(n10473), .ZN(n10478) );
  AND2_X1 U11469 ( .A1(n9871), .A2(n14378), .ZN(n9870) );
  NOR2_X1 U11470 ( .A1(n13799), .A2(n14392), .ZN(n9871) );
  INV_X1 U11471 ( .A(n14462), .ZN(n13799) );
  NAND2_X1 U11472 ( .A1(n9852), .A2(n9850), .ZN(n14401) );
  AND2_X1 U11473 ( .A1(n13710), .A2(n9851), .ZN(n9850) );
  INV_X1 U11474 ( .A(n9853), .ZN(n9851) );
  INV_X1 U11475 ( .A(n13949), .ZN(n13896) );
  NAND2_X1 U11476 ( .A1(n14840), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13949) );
  AND2_X1 U11477 ( .A1(n9620), .A2(n13592), .ZN(n9855) );
  INV_X1 U11478 ( .A(n13498), .ZN(n9857) );
  INV_X1 U11479 ( .A(n13296), .ZN(n13295) );
  NAND2_X1 U11480 ( .A1(n9706), .A2(n9704), .ZN(n11853) );
  NOR2_X1 U11481 ( .A1(n12854), .A2(n9616), .ZN(n9704) );
  CLKBUF_X1 U11482 ( .A(n13797), .Z(n13946) );
  NOR2_X1 U11483 ( .A1(n11920), .A2(n9715), .ZN(n9712) );
  INV_X1 U11484 ( .A(n14474), .ZN(n9759) );
  NAND2_X1 U11485 ( .A1(n13484), .A2(n9719), .ZN(n9718) );
  INV_X1 U11486 ( .A(n14683), .ZN(n9719) );
  NAND2_X1 U11487 ( .A1(n12067), .A2(n9768), .ZN(n9767) );
  INV_X1 U11488 ( .A(n14525), .ZN(n9768) );
  NAND2_X1 U11489 ( .A1(n19985), .A2(n11767), .ZN(n11963) );
  NOR2_X1 U11490 ( .A1(n13299), .A2(n9755), .ZN(n9754) );
  INV_X1 U11491 ( .A(n13231), .ZN(n9755) );
  NAND2_X1 U11492 ( .A1(n12929), .A2(n14331), .ZN(n12120) );
  NAND2_X1 U11493 ( .A1(n12929), .A2(n12114), .ZN(n12113) );
  OR2_X1 U11494 ( .A1(n11733), .A2(n11732), .ZN(n11780) );
  NAND2_X1 U11495 ( .A1(n10042), .A2(n11895), .ZN(n11756) );
  NAND2_X1 U11496 ( .A1(n12926), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11801) );
  OR2_X1 U11497 ( .A1(n19999), .A2(n20571), .ZN(n11800) );
  AND2_X1 U11498 ( .A1(n9845), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11794) );
  NAND2_X1 U11499 ( .A1(n9846), .A2(n11669), .ZN(n9700) );
  INV_X1 U11500 ( .A(n12824), .ZN(n19968) );
  OAI21_X1 U11501 ( .B1(n20670), .B2(n12829), .A(n14857), .ZN(n19971) );
  AOI221_X1 U11502 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11926), 
        .C1(n15917), .C2(n11926), .A(n11925), .ZN(n11970) );
  AND2_X1 U11503 ( .A1(n10655), .A2(n14889), .ZN(n10658) );
  NOR2_X1 U11504 ( .A1(n10649), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10655) );
  NOR2_X1 U11505 ( .A1(n10610), .A2(n10585), .ZN(n9837) );
  AND2_X1 U11506 ( .A1(n10560), .A2(n9833), .ZN(n9832) );
  INV_X1 U11507 ( .A(n13004), .ZN(n9960) );
  INV_X1 U11508 ( .A(n14867), .ZN(n10026) );
  NOR2_X1 U11509 ( .A1(n14863), .A2(n10025), .ZN(n10024) );
  INV_X1 U11510 ( .A(n10027), .ZN(n10025) );
  NAND2_X1 U11511 ( .A1(n9886), .A2(n13322), .ZN(n9885) );
  INV_X1 U11512 ( .A(n13269), .ZN(n9886) );
  NOR2_X1 U11513 ( .A1(n16035), .A2(n9903), .ZN(n9902) );
  INV_X1 U11514 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9903) );
  AND2_X1 U11515 ( .A1(n13472), .A2(n9974), .ZN(n9973) );
  INV_X1 U11516 ( .A(n12230), .ZN(n9974) );
  AND2_X1 U11517 ( .A1(n9615), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9911) );
  INV_X1 U11518 ( .A(n12604), .ZN(n9969) );
  NAND2_X1 U11519 ( .A1(n13983), .A2(n10065), .ZN(n10064) );
  NOR2_X1 U11520 ( .A1(n15965), .A2(n9804), .ZN(n13982) );
  NAND2_X1 U11521 ( .A1(n9808), .A2(n9621), .ZN(n9807) );
  NAND2_X1 U11522 ( .A1(n9809), .A2(n10055), .ZN(n9808) );
  INV_X1 U11523 ( .A(n13265), .ZN(n9809) );
  NAND2_X1 U11524 ( .A1(n10055), .A2(n10054), .ZN(n9810) );
  INV_X1 U11525 ( .A(n12961), .ZN(n9962) );
  NAND2_X1 U11526 ( .A1(n9905), .A2(n15269), .ZN(n15339) );
  INV_X1 U11527 ( .A(n15358), .ZN(n9905) );
  NAND2_X1 U11528 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  INV_X1 U11529 ( .A(n15382), .ZN(n9883) );
  INV_X1 U11530 ( .A(n9885), .ZN(n9884) );
  NAND2_X1 U11531 ( .A1(n9693), .A2(n13262), .ZN(n10054) );
  NAND2_X1 U11532 ( .A1(n15378), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15358) );
  NOR2_X1 U11533 ( .A1(n15392), .A2(n10058), .ZN(n10057) );
  INV_X1 U11534 ( .A(n10563), .ZN(n10058) );
  XNOR2_X1 U11535 ( .A(n11168), .B(n9804), .ZN(n11170) );
  OR2_X1 U11536 ( .A1(n10545), .A2(n10544), .ZN(n10853) );
  NAND2_X1 U11537 ( .A1(n10256), .A2(n10242), .ZN(n9691) );
  OR2_X1 U11538 ( .A1(n10343), .A2(n10342), .ZN(n10492) );
  AND2_X1 U11539 ( .A1(n13054), .A2(n19050), .ZN(n10227) );
  NAND2_X1 U11540 ( .A1(n10218), .A2(n12691), .ZN(n12693) );
  NOR2_X1 U11541 ( .A1(n10320), .A2(n10318), .ZN(n10296) );
  AOI21_X1 U11542 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18405), .A(
        n11404), .ZN(n11413) );
  AOI21_X1 U11543 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18426), .A(
        n11408), .ZN(n11417) );
  NOR2_X1 U11544 ( .A1(n10001), .A2(n17297), .ZN(n9998) );
  NOR2_X1 U11545 ( .A1(n16371), .A2(n17618), .ZN(n9986) );
  INV_X1 U11546 ( .A(n17384), .ZN(n9991) );
  NOR2_X1 U11547 ( .A1(n17414), .A2(n9993), .ZN(n9992) );
  INV_X1 U11548 ( .A(n17981), .ZN(n11479) );
  NOR2_X1 U11549 ( .A1(n11359), .A2(n11358), .ZN(n11435) );
  NOR2_X1 U11550 ( .A1(n11347), .A2(n9779), .ZN(n9778) );
  OR2_X1 U11551 ( .A1(n14512), .A2(n14501), .ZN(n14503) );
  NOR2_X1 U11552 ( .A1(n13363), .A2(n19727), .ZN(n13405) );
  NOR2_X2 U11553 ( .A1(n15769), .A2(n11901), .ZN(n13331) );
  NAND2_X1 U11554 ( .A1(n13100), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13099) );
  AND2_X1 U11555 ( .A1(n13559), .A2(n9822), .ZN(n9821) );
  INV_X1 U11556 ( .A(n14733), .ZN(n9822) );
  AND2_X1 U11557 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  INV_X1 U11558 ( .A(n13447), .ZN(n10046) );
  AND2_X1 U11559 ( .A1(n9631), .A2(n13073), .ZN(n13232) );
  NAND2_X1 U11560 ( .A1(n9729), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15778) );
  OR2_X1 U11561 ( .A1(n12126), .A2(n12776), .ZN(n19946) );
  NOR2_X1 U11562 ( .A1(n12611), .A2(n10093), .ZN(n14823) );
  INV_X1 U11563 ( .A(n20356), .ZN(n20283) );
  AND2_X1 U11564 ( .A1(n20473), .A2(n20001), .ZN(n20315) );
  INV_X1 U11565 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20507) );
  INV_X1 U11566 ( .A(n20287), .ZN(n20426) );
  AND2_X1 U11567 ( .A1(n12824), .A2(n12853), .ZN(n20475) );
  AND2_X1 U11568 ( .A1(n10723), .A2(n10737), .ZN(n12679) );
  NOR3_X1 U11569 ( .A1(n10778), .A2(n10777), .A3(n10776), .ZN(n12684) );
  NOR2_X1 U11570 ( .A1(n10672), .A2(n10673), .ZN(n14009) );
  NAND2_X1 U11571 ( .A1(n14015), .A2(n10660), .ZN(n9830) );
  INV_X1 U11572 ( .A(n15071), .ZN(n9917) );
  NOR2_X1 U11573 ( .A1(n10612), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10614) );
  INV_X1 U11574 ( .A(n18814), .ZN(n12216) );
  NOR2_X1 U11575 ( .A1(n9567), .A2(n12317), .ZN(n10071) );
  NOR2_X1 U11576 ( .A1(n10237), .A2(n9567), .ZN(n10073) );
  XNOR2_X1 U11577 ( .A(n14181), .B(n14177), .ZN(n14884) );
  INV_X1 U11578 ( .A(n13208), .ZN(n9888) );
  AND2_X1 U11579 ( .A1(n13167), .A2(n10860), .ZN(n13270) );
  XNOR2_X1 U11580 ( .A(n12193), .B(n12192), .ZN(n14031) );
  CLKBUF_X1 U11581 ( .A(n12210), .Z(n12213) );
  NAND2_X1 U11582 ( .A1(n12198), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12209) );
  AND4_X1 U11583 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        n10460) );
  AND4_X1 U11584 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10463) );
  NAND2_X1 U11585 ( .A1(n14007), .A2(n14006), .ZN(n15015) );
  AND2_X1 U11586 ( .A1(n15158), .A2(n10800), .ZN(n15149) );
  NOR2_X1 U11587 ( .A1(n15168), .A2(n9747), .ZN(n9746) );
  INV_X1 U11588 ( .A(n10652), .ZN(n9747) );
  NAND2_X1 U11589 ( .A1(n9881), .A2(n15371), .ZN(n9880) );
  INV_X1 U11590 ( .A(n9882), .ZN(n9881) );
  NOR2_X1 U11591 ( .A1(n11170), .A2(n11169), .ZN(n13261) );
  NAND2_X1 U11592 ( .A1(n10505), .A2(n12724), .ZN(n12835) );
  AND2_X1 U11593 ( .A1(n10834), .A2(n9879), .ZN(n9878) );
  INV_X1 U11594 ( .A(n12730), .ZN(n9879) );
  INV_X1 U11595 ( .A(n12848), .ZN(n11047) );
  NAND2_X1 U11596 ( .A1(n9895), .A2(n9897), .ZN(n9894) );
  INV_X1 U11597 ( .A(n10261), .ZN(n9895) );
  NAND2_X1 U11598 ( .A1(n9803), .A2(n10368), .ZN(n10485) );
  NAND2_X1 U11599 ( .A1(n9686), .A2(n10395), .ZN(n10484) );
  AND2_X1 U11600 ( .A1(n10755), .A2(n12989), .ZN(n11174) );
  BUF_X4 U11601 ( .A(n12216), .Z(n18830) );
  NOR2_X1 U11602 ( .A1(n19636), .A2(n19663), .ZN(n19087) );
  NAND2_X1 U11603 ( .A1(n13034), .A2(n19663), .ZN(n19229) );
  NAND2_X1 U11604 ( .A1(n16167), .A2(n12317), .ZN(n13017) );
  OR2_X1 U11605 ( .A1(n19647), .A2(n18847), .ZN(n19394) );
  NAND2_X1 U11606 ( .A1(n19636), .A2(n19663), .ZN(n19395) );
  NAND2_X1 U11607 ( .A1(n19636), .A2(n13040), .ZN(n19446) );
  NAND2_X1 U11608 ( .A1(n10706), .A2(n10703), .ZN(n12683) );
  INV_X1 U11609 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13184) );
  OR2_X1 U11610 ( .A1(n16380), .A2(n10012), .ZN(n9978) );
  NAND2_X1 U11611 ( .A1(n9613), .A2(n10000), .ZN(n9999) );
  INV_X1 U11612 ( .A(n17297), .ZN(n10000) );
  NOR2_X1 U11613 ( .A1(n16412), .A2(n16413), .ZN(n16411) );
  OAI21_X1 U11614 ( .B1(n10012), .B2(n10016), .A(n10015), .ZN(n10014) );
  INV_X1 U11615 ( .A(n17370), .ZN(n10016) );
  INV_X1 U11616 ( .A(n17353), .ZN(n10015) );
  OR2_X1 U11617 ( .A1(n16474), .A2(n10012), .ZN(n9976) );
  INV_X1 U11618 ( .A(n17985), .ZN(n11390) );
  AND2_X2 U11619 ( .A1(n11229), .A2(n11228), .ZN(n11451) );
  NOR2_X1 U11620 ( .A1(n11227), .A2(n11226), .ZN(n11228) );
  AOI211_X1 U11621 ( .C1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .C2(n11215), .A(
        n11223), .B(n11222), .ZN(n11229) );
  NOR2_X1 U11622 ( .A1(n17283), .A2(n11308), .ZN(n11309) );
  NAND2_X1 U11623 ( .A1(n11307), .A2(n10087), .ZN(n11308) );
  OR2_X1 U11624 ( .A1(n17301), .A2(n17528), .ZN(n11307) );
  NAND2_X1 U11625 ( .A1(n11309), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11310) );
  NOR3_X1 U11626 ( .A1(n17308), .A2(n17331), .A3(n17672), .ZN(n17301) );
  AND2_X1 U11627 ( .A1(n17454), .A2(n17423), .ZN(n11300) );
  AND2_X1 U11628 ( .A1(n11295), .A2(n17838), .ZN(n9955) );
  NOR2_X1 U11629 ( .A1(n11297), .A2(n9951), .ZN(n9950) );
  NAND2_X1 U11630 ( .A1(n17528), .A2(n17862), .ZN(n9951) );
  INV_X1 U11631 ( .A(n17452), .ZN(n17430) );
  AND2_X2 U11632 ( .A1(n12527), .A2(n19701), .ZN(n19797) );
  OAI21_X1 U11633 ( .B1(n12526), .B2(n12528), .A(n12792), .ZN(n12527) );
  NAND2_X1 U11634 ( .A1(n15730), .A2(n12496), .ZN(n15721) );
  AND2_X1 U11635 ( .A1(n13909), .A2(n19966), .ZN(n15723) );
  INV_X1 U11636 ( .A(n15730), .ZN(n14604) );
  INV_X1 U11637 ( .A(n14601), .ZN(n15727) );
  AND2_X1 U11638 ( .A1(n12489), .A2(n19701), .ZN(n15730) );
  XNOR2_X1 U11639 ( .A(n9865), .B(n9864), .ZN(n14533) );
  INV_X1 U11640 ( .A(n9865), .ZN(n14326) );
  OR2_X1 U11641 ( .A1(n19917), .A2(n12249), .ZN(n14677) );
  XNOR2_X1 U11642 ( .A(n12123), .B(n12122), .ZN(n14453) );
  AND2_X1 U11643 ( .A1(n14626), .A2(n9816), .ZN(n9824) );
  NOR2_X1 U11644 ( .A1(n9825), .A2(n14734), .ZN(n9816) );
  NOR3_X1 U11645 ( .A1(n14728), .A2(n14719), .A3(n9785), .ZN(n14717) );
  AND2_X1 U11646 ( .A1(n15889), .A2(n14723), .ZN(n9785) );
  XNOR2_X1 U11647 ( .A(n14333), .B(n9782), .ZN(n14721) );
  INV_X1 U11648 ( .A(n14332), .ZN(n9782) );
  XNOR2_X1 U11649 ( .A(n9730), .B(n13560), .ZN(n14730) );
  OAI21_X1 U11650 ( .B1(n14626), .B2(n14733), .A(n9731), .ZN(n9730) );
  OAI21_X1 U11651 ( .B1(n15819), .B2(n14787), .A(n15866), .ZN(n14790) );
  OR2_X1 U11652 ( .A1(n12126), .A2(n12125), .ZN(n19955) );
  OR2_X1 U11653 ( .A1(n12126), .A2(n11998), .ZN(n19925) );
  INV_X1 U11654 ( .A(n20568), .ZN(n20498) );
  AND2_X1 U11655 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12596) );
  NOR2_X1 U11656 ( .A1(n14306), .A2(n14307), .ZN(n14042) );
  XNOR2_X1 U11657 ( .A(n14935), .B(n14307), .ZN(n15945) );
  NAND2_X1 U11658 ( .A1(n15931), .A2(n18988), .ZN(n14034) );
  NOR2_X1 U11659 ( .A1(n14003), .A2(n18992), .ZN(n10067) );
  INV_X1 U11660 ( .A(n15233), .ZN(n9688) );
  NAND2_X1 U11661 ( .A1(n12324), .A2(n12318), .ZN(n16121) );
  NAND2_X1 U11662 ( .A1(n10068), .A2(n9644), .ZN(n15155) );
  INV_X1 U11663 ( .A(n15021), .ZN(n10068) );
  AOI21_X1 U11664 ( .B1(n15951), .B2(n19004), .A(n9656), .ZN(n9875) );
  NAND2_X1 U11665 ( .A1(n14306), .A2(n9877), .ZN(n15152) );
  OR2_X1 U11666 ( .A1(n14934), .A2(n14933), .ZN(n9877) );
  AND2_X1 U11667 ( .A1(n11174), .A2(n19671), .ZN(n18999) );
  INV_X1 U11668 ( .A(n16158), .ZN(n19004) );
  AND2_X1 U11669 ( .A1(n11174), .A2(n19669), .ZN(n16154) );
  NOR2_X1 U11670 ( .A1(n16464), .A2(n10012), .ZN(n16454) );
  NAND2_X1 U11671 ( .A1(n9931), .A2(n9637), .ZN(n9928) );
  NAND2_X1 U11672 ( .A1(n12135), .A2(n9983), .ZN(n9931) );
  NOR2_X1 U11673 ( .A1(n16196), .A2(n16197), .ZN(n9935) );
  NOR2_X1 U11674 ( .A1(n17583), .A2(n17585), .ZN(n17560) );
  INV_X1 U11675 ( .A(n17615), .ZN(n17627) );
  INV_X1 U11676 ( .A(n17612), .ZN(n17628) );
  NOR3_X2 U11677 ( .A1(n17118), .A2(n18590), .A3(n9563), .ZN(n17850) );
  NOR2_X1 U11679 ( .A1(n10418), .A2(n10419), .ZN(n9735) );
  INV_X1 U11680 ( .A(n19149), .ZN(n10526) );
  NAND2_X1 U11681 ( .A1(n11924), .A2(n11923), .ZN(n11933) );
  XNOR2_X1 U11682 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U11683 ( .A1(n11933), .A2(n11932), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20256), .ZN(n11928) );
  NOR2_X1 U11684 ( .A1(n11928), .A2(n11929), .ZN(n11927) );
  OR2_X1 U11685 ( .A1(n11851), .A2(n11850), .ZN(n11877) );
  NOR2_X1 U11686 ( .A1(n15559), .A2(n20571), .ZN(n9717) );
  NOR2_X1 U11687 ( .A1(n11664), .A2(n11663), .ZN(n12013) );
  AND2_X1 U11688 ( .A1(n11978), .A2(n11977), .ZN(n12011) );
  NOR2_X1 U11689 ( .A1(n11948), .A2(n11945), .ZN(n11946) );
  NAND2_X1 U11690 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10179) );
  AOI22_X1 U11691 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10173) );
  AND2_X1 U11692 ( .A1(n19666), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10679) );
  INV_X1 U11693 ( .A(n10168), .ZN(n10213) );
  INV_X1 U11694 ( .A(n10553), .ZN(n9833) );
  AND4_X1 U11695 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n10535) );
  INV_X1 U11696 ( .A(n10853), .ZN(n10552) );
  INV_X1 U11697 ( .A(n11161), .ZN(n10548) );
  AOI21_X1 U11698 ( .B1(n10247), .B2(P2_EBX_REG_3__SCAN_IN), .A(n10096), .ZN(
        n10264) );
  NOR2_X1 U11699 ( .A1(n9567), .A2(n10072), .ZN(n10070) );
  OR2_X1 U11700 ( .A1(n10367), .A2(n10366), .ZN(n10824) );
  OAI22_X1 U11701 ( .A1(n10299), .A2(n10417), .B1(n10423), .B2(n10298), .ZN(
        n10302) );
  OAI21_X1 U11702 ( .B1(n10300), .B2(n10418), .A(n9689), .ZN(n10301) );
  INV_X1 U11703 ( .A(n11130), .ZN(n10248) );
  AND2_X1 U11704 ( .A1(n10229), .A2(n10226), .ZN(n10766) );
  NAND2_X1 U11705 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n9964) );
  NAND2_X1 U11706 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n9963) );
  NAND2_X1 U11707 ( .A1(n9568), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9802) );
  NAND2_X1 U11708 ( .A1(n14104), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n9801) );
  NAND2_X1 U11709 ( .A1(n10051), .A2(n10049), .ZN(n10201) );
  NAND2_X1 U11710 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18568), .ZN(
        n11185) );
  INV_X1 U11711 ( .A(n13378), .ZN(n9866) );
  NAND2_X1 U11712 ( .A1(n11655), .A2(n11661), .ZN(n12481) );
  NAND2_X1 U11713 ( .A1(n9855), .A2(n9854), .ZN(n9853) );
  INV_X1 U11714 ( .A(n14599), .ZN(n9854) );
  NOR2_X1 U11715 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13797) );
  OR2_X1 U11716 ( .A1(n11722), .A2(n11721), .ZN(n11899) );
  AND2_X1 U11717 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12873), .ZN(
        n12915) );
  OR2_X1 U11718 ( .A1(n11812), .A2(n11811), .ZN(n11856) );
  NAND2_X1 U11719 ( .A1(n14488), .A2(n9756), .ZN(n9761) );
  NOR2_X1 U11720 ( .A1(n12101), .A2(n9758), .ZN(n9756) );
  NOR2_X1 U11721 ( .A1(n14467), .A2(n14381), .ZN(n12108) );
  NOR2_X1 U11722 ( .A1(n15769), .A2(n9683), .ZN(n14695) );
  OR2_X1 U11723 ( .A1(n11750), .A2(n11749), .ZN(n11779) );
  INV_X1 U11724 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20058) );
  AND2_X1 U11725 ( .A1(n9653), .A2(n11526), .ZN(n10041) );
  INV_X1 U11726 ( .A(n20427), .ZN(n20505) );
  AND2_X1 U11727 ( .A1(n11961), .A2(n9793), .ZN(n9792) );
  INV_X1 U11728 ( .A(n9794), .ZN(n9793) );
  OAI21_X1 U11729 ( .B1(n9789), .B2(n11968), .A(n9795), .ZN(n9794) );
  AOI21_X1 U11730 ( .B1(n10478), .B2(n10477), .A(n10476), .ZN(n10694) );
  OR2_X1 U11731 ( .A1(n10406), .A2(n10405), .ZN(n10480) );
  NAND2_X1 U11732 ( .A1(n10658), .A2(n11124), .ZN(n10662) );
  INV_X1 U11733 ( .A(n9837), .ZN(n10600) );
  NOR2_X1 U11734 ( .A1(n10605), .A2(n10603), .ZN(n10608) );
  NOR2_X1 U11735 ( .A1(n16056), .A2(n9913), .ZN(n9912) );
  INV_X1 U11736 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9913) );
  AND2_X1 U11737 ( .A1(n11066), .A2(n9839), .ZN(n9838) );
  NOR2_X1 U11738 ( .A1(n9836), .A2(n9835), .ZN(n9834) );
  INV_X1 U11739 ( .A(n10482), .ZN(n9835) );
  MUX2_X1 U11740 ( .A(n10733), .B(P2_EBX_REG_3__SCAN_IN), .S(n13985), .Z(
        n10486) );
  CLKBUF_X1 U11741 ( .A(n9579), .Z(n14279) );
  CLKBUF_X1 U11742 ( .A(n9568), .Z(n14296) );
  NAND2_X1 U11743 ( .A1(n14885), .A2(n14182), .ZN(n14204) );
  INV_X1 U11744 ( .A(n14227), .ZN(n14201) );
  NAND2_X1 U11745 ( .A1(n14903), .A2(n14904), .ZN(n10032) );
  INV_X1 U11746 ( .A(n15315), .ZN(n9887) );
  NAND2_X1 U11747 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9925) );
  AND2_X1 U11748 ( .A1(n13983), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9743) );
  AND2_X1 U11749 ( .A1(n10660), .A2(n10858), .ZN(n9827) );
  AND2_X1 U11750 ( .A1(n14983), .A2(n16012), .ZN(n9891) );
  NAND2_X1 U11751 ( .A1(n11158), .A2(n9804), .ZN(n10483) );
  INV_X1 U11752 ( .A(n16110), .ZN(n9899) );
  NAND2_X1 U11753 ( .A1(n10274), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9690) );
  AOI22_X1 U11754 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n19088), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10380) );
  AND4_X1 U11755 ( .A1(n10373), .A2(n10372), .A3(n10371), .A4(n10370), .ZN(
        n10383) );
  OAI211_X2 U11756 ( .C1(n11019), .C2(n10236), .A(n10235), .B(n10234), .ZN(
        n11022) );
  NAND2_X1 U11757 ( .A1(n10767), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10236) );
  NAND2_X1 U11758 ( .A1(n11017), .A2(n10233), .ZN(n10235) );
  OR2_X1 U11759 ( .A1(n10356), .A2(n10355), .ZN(n11141) );
  NAND2_X1 U11760 ( .A1(n9608), .A2(n10303), .ZN(n10514) );
  INV_X1 U11761 ( .A(n10516), .ZN(n19058) );
  NAND2_X1 U11762 ( .A1(n10303), .A2(n9734), .ZN(n10417) );
  NAND2_X1 U11763 ( .A1(n10296), .A2(n12447), .ZN(n10411) );
  NAND3_X1 U11764 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19642), .A3(n19392), 
        .ZN(n13022) );
  INV_X1 U11765 ( .A(n11265), .ZN(n16844) );
  NOR2_X1 U11766 ( .A1(n11184), .A2(n18392), .ZN(n11323) );
  NOR2_X1 U11767 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15523), .ZN(
        n11265) );
  NOR2_X1 U11768 ( .A1(n11184), .A2(n16657), .ZN(n11241) );
  INV_X1 U11769 ( .A(n18392), .ZN(n9772) );
  INV_X1 U11770 ( .A(n11183), .ZN(n9773) );
  INV_X1 U11771 ( .A(n17960), .ZN(n12179) );
  OR2_X1 U11772 ( .A1(n11492), .A2(n18443), .ZN(n15516) );
  INV_X1 U11773 ( .A(n9933), .ZN(n11492) );
  OR2_X1 U11774 ( .A1(n17542), .A2(n17874), .ZN(n9952) );
  NAND2_X1 U11775 ( .A1(n9945), .A2(n9938), .ZN(n9942) );
  NAND2_X1 U11776 ( .A1(n9947), .A2(n17580), .ZN(n9944) );
  XNOR2_X1 U11777 ( .A(n11451), .B(n17137), .ZN(n11282) );
  INV_X1 U11778 ( .A(n17973), .ZN(n11484) );
  INV_X1 U11779 ( .A(n9848), .ZN(n12001) );
  INV_X1 U11780 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U11781 ( .A1(n12028), .A2(n9769), .ZN(n12031) );
  OR3_X1 U11782 ( .A1(n20664), .A2(n12914), .A3(n12913), .ZN(n13915) );
  AND2_X1 U11783 ( .A1(n19824), .A2(n12474), .ZN(n19802) );
  AND2_X1 U11784 ( .A1(n12920), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13929) );
  NOR2_X1 U11785 ( .A1(n13852), .A2(n20813), .ZN(n13855) );
  AND2_X1 U11786 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n12919), .ZN(
        n13818) );
  INV_X1 U11787 ( .A(n13815), .ZN(n12919) );
  NAND2_X1 U11788 ( .A1(n13818), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13852) );
  AND2_X1 U11789 ( .A1(n9870), .A2(n9869), .ZN(n9868) );
  INV_X1 U11790 ( .A(n14364), .ZN(n9869) );
  NAND2_X1 U11791 ( .A1(n14391), .A2(n9870), .ZN(n14377) );
  NOR2_X1 U11792 ( .A1(n13773), .A2(n14396), .ZN(n13777) );
  NAND2_X1 U11793 ( .A1(n13777), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13815) );
  NOR2_X1 U11794 ( .A1(n13742), .A2(n12918), .ZN(n13711) );
  INV_X1 U11795 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12918) );
  INV_X1 U11796 ( .A(n14391), .ZN(n15633) );
  NAND2_X1 U11797 ( .A1(n14666), .A2(n9634), .ZN(n11917) );
  OAI21_X1 U11798 ( .B1(n14666), .B2(n11918), .A(n15769), .ZN(n15737) );
  NOR2_X1 U11799 ( .A1(n13644), .A2(n15655), .ZN(n13610) );
  NAND2_X1 U11800 ( .A1(n13610), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13742) );
  NOR2_X1 U11801 ( .A1(n13676), .A2(n14425), .ZN(n13643) );
  NAND2_X1 U11802 ( .A1(n13643), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13644) );
  AND2_X1 U11803 ( .A1(n13673), .A2(n13672), .ZN(n14414) );
  OR2_X1 U11804 ( .A1(n14503), .A2(n14414), .ZN(n14491) );
  NOR2_X1 U11805 ( .A1(n13694), .A2(n12917), .ZN(n13675) );
  INV_X1 U11806 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12917) );
  NAND2_X1 U11807 ( .A1(n13675), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13676) );
  NAND2_X1 U11808 ( .A1(n13593), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13694) );
  NOR2_X1 U11809 ( .A1(n13562), .A2(n14437), .ZN(n13593) );
  OR2_X1 U11810 ( .A1(n13587), .A2(n15699), .ZN(n13562) );
  AND3_X1 U11811 ( .A1(n13591), .A2(n13590), .A3(n13589), .ZN(n14523) );
  NAND2_X1 U11812 ( .A1(n13494), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13587) );
  NAND2_X1 U11813 ( .A1(n12916), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13363) );
  AND3_X1 U11814 ( .A1(n13294), .A2(n13293), .A3(n13292), .ZN(n13296) );
  NAND2_X1 U11815 ( .A1(n13227), .A2(n13228), .ZN(n13297) );
  NOR2_X1 U11816 ( .A1(n13099), .A2(n13114), .ZN(n13221) );
  AND2_X1 U11817 ( .A1(n13097), .A2(n12881), .ZN(n9867) );
  AOI21_X1 U11818 ( .B1(n13104), .B2(n13706), .A(n13103), .ZN(n13118) );
  AND2_X1 U11819 ( .A1(n12915), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13100) );
  NAND2_X1 U11820 ( .A1(n12882), .A2(n12881), .ZN(n13095) );
  AOI21_X1 U11821 ( .B1(n13607), .B2(n9860), .A(n9859), .ZN(n9858) );
  INV_X1 U11822 ( .A(n12871), .ZN(n9859) );
  AND2_X1 U11823 ( .A1(n12822), .A2(n19701), .ZN(n19824) );
  NAND2_X1 U11824 ( .A1(n13558), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9825) );
  AND2_X1 U11825 ( .A1(n14357), .A2(n14342), .ZN(n14344) );
  NOR2_X1 U11826 ( .A1(n14365), .A2(n14358), .ZN(n14357) );
  NAND2_X1 U11827 ( .A1(n12108), .A2(n9770), .ZN(n14365) );
  INV_X1 U11828 ( .A(n14367), .ZN(n9770) );
  OR2_X1 U11829 ( .A1(n9761), .A2(n9760), .ZN(n14467) );
  INV_X1 U11830 ( .A(n14464), .ZN(n9760) );
  INV_X1 U11831 ( .A(n12108), .ZN(n14383) );
  NAND2_X1 U11832 ( .A1(n14488), .A2(n9757), .ZN(n15636) );
  INV_X1 U11833 ( .A(n14790), .ZN(n15810) );
  AND2_X1 U11834 ( .A1(n12088), .A2(n12087), .ZN(n14486) );
  AND2_X1 U11835 ( .A1(n14495), .A2(n14486), .ZN(n14488) );
  NOR2_X1 U11836 ( .A1(n14494), .A2(n14493), .ZN(n14495) );
  NAND2_X1 U11837 ( .A1(n9718), .A2(n9844), .ZN(n9843) );
  INV_X1 U11838 ( .A(n14809), .ZN(n9844) );
  OR2_X1 U11839 ( .A1(n14506), .A2(n14422), .ZN(n14494) );
  NOR2_X1 U11840 ( .A1(n14526), .A2(n9765), .ZN(n14518) );
  NAND2_X1 U11841 ( .A1(n9766), .A2(n12073), .ZN(n9765) );
  INV_X1 U11842 ( .A(n9767), .ZN(n9766) );
  NAND2_X1 U11843 ( .A1(n14518), .A2(n14504), .ZN(n14506) );
  NAND2_X1 U11844 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13485) );
  NOR2_X1 U11845 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14699) );
  NOR2_X1 U11846 ( .A1(n14526), .A2(n9767), .ZN(n10083) );
  NAND2_X1 U11847 ( .A1(n13232), .A2(n9752), .ZN(n15881) );
  NOR2_X1 U11848 ( .A1(n9753), .A2(n15879), .ZN(n9752) );
  INV_X1 U11849 ( .A(n9754), .ZN(n9753) );
  AND2_X1 U11850 ( .A1(n12061), .A2(n12060), .ZN(n13476) );
  NOR2_X1 U11851 ( .A1(n15881), .A2(n13476), .ZN(n13510) );
  NAND2_X1 U11852 ( .A1(n11904), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10047) );
  AND2_X1 U11853 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13447) );
  AND3_X1 U11854 ( .A1(n12054), .A2(n12090), .A3(n12053), .ZN(n13299) );
  NOR2_X1 U11855 ( .A1(n12998), .A2(n13121), .ZN(n9771) );
  AND2_X1 U11856 ( .A1(n12639), .A2(n12640), .ZN(n12884) );
  NAND2_X1 U11857 ( .A1(n12884), .A2(n12039), .ZN(n12999) );
  AND2_X1 U11858 ( .A1(n19946), .A2(n14823), .ZN(n12895) );
  NOR2_X1 U11859 ( .A1(n12126), .A2(n15558), .ZN(n12611) );
  AND2_X1 U11860 ( .A1(n12018), .A2(n12017), .ZN(n10093) );
  INV_X1 U11861 ( .A(n19946), .ZN(n14784) );
  NAND2_X1 U11862 ( .A1(n20094), .A2(n11758), .ZN(n20024) );
  INV_X1 U11863 ( .A(n12510), .ZN(n11763) );
  NAND2_X1 U11864 ( .A1(n11799), .A2(n11798), .ZN(n20134) );
  NAND2_X1 U11865 ( .A1(n20094), .A2(n11688), .ZN(n9699) );
  BUF_X1 U11866 ( .A(n11667), .Z(n14061) );
  AND2_X1 U11867 ( .A1(n12824), .A2(n12854), .ZN(n20232) );
  NAND2_X1 U11868 ( .A1(n12855), .A2(n19968), .ZN(n20356) );
  AND3_X1 U11869 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20571), .A3(n19971), 
        .ZN(n20016) );
  AND2_X1 U11870 ( .A1(n20053), .A2(n20052), .ZN(n20474) );
  NOR2_X2 U11871 ( .A1(n19965), .A2(n19967), .ZN(n20013) );
  NOR2_X2 U11872 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20518) );
  NAND2_X1 U11873 ( .A1(n20570), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15584) );
  NOR2_X1 U11874 ( .A1(n20573), .A2(n20570), .ZN(n12829) );
  AND2_X1 U11875 ( .A1(n20577), .A2(n11660), .ZN(n11972) );
  OR2_X1 U11876 ( .A1(n15953), .A2(n15954), .ZN(n9900) );
  NOR2_X1 U11877 ( .A1(n15960), .A2(n18830), .ZN(n15953) );
  INV_X1 U11878 ( .A(n15975), .ZN(n9910) );
  AND2_X1 U11879 ( .A1(n11009), .A2(n11008), .ZN(n13537) );
  NAND2_X1 U11880 ( .A1(n10635), .A2(n9674), .ZN(n10649) );
  INV_X1 U11881 ( .A(n10642), .ZN(n9841) );
  NAND2_X1 U11882 ( .A1(n10614), .A2(n11112), .ZN(n10638) );
  NAND2_X1 U11883 ( .A1(n9837), .A2(n9673), .ZN(n10612) );
  NAND2_X1 U11884 ( .A1(n10578), .A2(n10581), .ZN(n9840) );
  AND2_X1 U11885 ( .A1(n10567), .A2(n9838), .ZN(n10572) );
  NAND2_X1 U11886 ( .A1(n10567), .A2(n11066), .ZN(n10570) );
  NAND2_X1 U11887 ( .A1(n9834), .A2(n10507), .ZN(n10554) );
  NOR2_X1 U11888 ( .A1(n13997), .A2(n13996), .ZN(n14313) );
  AND2_X1 U11889 ( .A1(n10028), .A2(n14867), .ZN(n10027) );
  INV_X1 U11890 ( .A(n14872), .ZN(n10028) );
  OR2_X1 U11891 ( .A1(n13536), .A2(n11132), .ZN(n13997) );
  NAND2_X1 U11892 ( .A1(n13533), .A2(n13534), .ZN(n13536) );
  NAND2_X1 U11893 ( .A1(n9957), .A2(n9956), .ZN(n14897) );
  INV_X1 U11894 ( .A(n14895), .ZN(n9956) );
  INV_X1 U11895 ( .A(n14901), .ZN(n9957) );
  INV_X1 U11896 ( .A(n13338), .ZN(n11100) );
  NOR2_X1 U11897 ( .A1(n9655), .A2(n9959), .ZN(n9958) );
  NAND2_X1 U11898 ( .A1(n9960), .A2(n13029), .ZN(n9959) );
  INV_X1 U11899 ( .A(n14231), .ZN(n10022) );
  NAND2_X1 U11900 ( .A1(n14234), .A2(n10024), .ZN(n10023) );
  INV_X1 U11901 ( .A(n10031), .ZN(n10033) );
  INV_X1 U11902 ( .A(n10032), .ZN(n14905) );
  NAND2_X1 U11903 ( .A1(n9614), .A2(n13189), .ZN(n10034) );
  AND2_X1 U11904 ( .A1(n10981), .A2(n10980), .ZN(n15293) );
  NAND2_X1 U11905 ( .A1(n15349), .A2(n15350), .ZN(n15351) );
  OAI21_X1 U11906 ( .B1(n12165), .B2(n12164), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12166) );
  AND2_X1 U11907 ( .A1(n10894), .A2(n10893), .ZN(n15382) );
  INV_X1 U11908 ( .A(n10214), .ZN(n12991) );
  AND2_X1 U11909 ( .A1(n12273), .A2(n12232), .ZN(n18973) );
  AND2_X1 U11910 ( .A1(n9618), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9901) );
  NAND2_X1 U11911 ( .A1(n15041), .A2(n9618), .ZN(n15031) );
  AND2_X1 U11912 ( .A1(n14925), .A2(n9668), .ZN(n14913) );
  INV_X1 U11913 ( .A(n14914), .ZN(n9972) );
  NAND2_X1 U11914 ( .A1(n14925), .A2(n13472), .ZN(n13471) );
  NAND2_X1 U11915 ( .A1(n14925), .A2(n9973), .ZN(n14915) );
  INV_X1 U11916 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15098) );
  CLKBUF_X1 U11917 ( .A(n12197), .Z(n12208) );
  NOR2_X1 U11918 ( .A1(n9627), .A2(n9968), .ZN(n9967) );
  INV_X1 U11919 ( .A(n12598), .ZN(n9968) );
  NOR2_X1 U11920 ( .A1(n13964), .A2(n9627), .ZN(n12605) );
  NOR2_X1 U11921 ( .A1(n12760), .A2(n12205), .ZN(n12207) );
  OR3_X1 U11922 ( .A1(n15943), .A2(n9804), .A3(n14044), .ZN(n15016) );
  AOI21_X1 U11923 ( .B1(n14012), .B2(n10858), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15018) );
  AND2_X1 U11924 ( .A1(n11015), .A2(n11014), .ZN(n14934) );
  AOI22_X1 U11925 ( .A1(n13982), .A2(n10063), .B1(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U11926 ( .A1(n10064), .A2(n10061), .ZN(n10060) );
  AND2_X1 U11927 ( .A1(n13982), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10061) );
  OAI21_X1 U11928 ( .B1(n13986), .B2(n9804), .A(n15147), .ZN(n14006) );
  NOR2_X1 U11929 ( .A1(n9812), .A2(n13984), .ZN(n9811) );
  INV_X1 U11930 ( .A(n9813), .ZN(n9812) );
  INV_X1 U11931 ( .A(n10671), .ZN(n9740) );
  NOR2_X1 U11932 ( .A1(n13543), .A2(n9814), .ZN(n9813) );
  NAND2_X1 U11933 ( .A1(n15175), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15028) );
  NAND2_X1 U11934 ( .A1(n12233), .A2(n9889), .ZN(n14977) );
  AND2_X1 U11935 ( .A1(n9891), .A2(n9890), .ZN(n9889) );
  INV_X1 U11936 ( .A(n14975), .ZN(n9890) );
  NOR2_X2 U11937 ( .A1(n14977), .A2(n14964), .ZN(n14965) );
  NAND2_X1 U11938 ( .A1(n9810), .A2(n10790), .ZN(n9806) );
  NAND2_X1 U11939 ( .A1(n12233), .A2(n9891), .ZN(n16013) );
  AND2_X1 U11940 ( .A1(n12233), .A2(n14983), .ZN(n16011) );
  OR2_X1 U11941 ( .A1(n9807), .A2(n9805), .ZN(n15198) );
  INV_X1 U11942 ( .A(n9810), .ZN(n9805) );
  NAND2_X1 U11943 ( .A1(n9810), .A2(n9643), .ZN(n15085) );
  NAND2_X1 U11944 ( .A1(n9694), .A2(n10055), .ZN(n15378) );
  INV_X1 U11945 ( .A(n10054), .ZN(n10056) );
  NAND2_X1 U11946 ( .A1(n16147), .A2(n10854), .ZN(n13169) );
  NOR2_X1 U11947 ( .A1(n13964), .A2(n12564), .ZN(n12565) );
  NAND2_X1 U11948 ( .A1(n12836), .A2(n11157), .ZN(n16112) );
  NAND2_X1 U11949 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  INV_X1 U11950 ( .A(n10502), .ZN(n10504) );
  NAND2_X1 U11951 ( .A1(n10246), .A2(n10245), .ZN(n10286) );
  OAI22_X1 U11952 ( .A1(n10274), .A2(n10244), .B1(n10247), .B2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10246) );
  OAI211_X1 U11953 ( .C1(n10978), .C2(n11142), .A(n10826), .B(n10814), .ZN(
        n9872) );
  AND2_X1 U11954 ( .A1(n12317), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12455) );
  NAND2_X1 U11955 ( .A1(n12342), .A2(n19639), .ZN(n12536) );
  AND2_X1 U11956 ( .A1(n19647), .A2(n19654), .ZN(n19064) );
  INV_X1 U11957 ( .A(n10412), .ZN(n13023) );
  NAND2_X1 U11958 ( .A1(n10318), .A2(n12447), .ZN(n10313) );
  INV_X1 U11959 ( .A(n19064), .ZN(n19066) );
  AND2_X1 U11960 ( .A1(n19647), .A2(n18847), .ZN(n19632) );
  OR2_X1 U11961 ( .A1(n19647), .A2(n19654), .ZN(n19445) );
  INV_X1 U11962 ( .A(n19445), .ZN(n19500) );
  NOR2_X1 U11963 ( .A1(n13034), .A2(n19633), .ZN(n19499) );
  INV_X1 U11964 ( .A(n19033), .ZN(n19049) );
  NOR2_X2 U11965 ( .A1(n13211), .A2(n13022), .ZN(n19047) );
  NOR2_X2 U11966 ( .A1(n13021), .A2(n13022), .ZN(n19048) );
  AND2_X1 U11967 ( .A1(n12579), .A2(n12578), .ZN(n12702) );
  NOR2_X1 U11968 ( .A1(n11429), .A2(n18414), .ZN(n11487) );
  OAI211_X1 U11969 ( .C1(n11411), .C2(n11410), .A(n11417), .B(n11409), .ZN(
        n11425) );
  OAI21_X1 U11970 ( .B1(n11418), .B2(n11422), .A(n11417), .ZN(n11426) );
  NOR2_X1 U11971 ( .A1(n15611), .A2(n15516), .ZN(n18431) );
  INV_X1 U11972 ( .A(n17259), .ZN(n9977) );
  INV_X1 U11973 ( .A(n9997), .ZN(n9994) );
  NOR2_X1 U11974 ( .A1(n16412), .A2(n9999), .ZN(n9995) );
  AOI21_X1 U11975 ( .B1(n9613), .B2(n9998), .A(n10012), .ZN(n9997) );
  NOR2_X1 U11976 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16494), .ZN(n16486) );
  NOR2_X1 U11977 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16515), .ZN(n16505) );
  NOR2_X1 U11978 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16546), .ZN(n16525) );
  NAND2_X1 U11979 ( .A1(n9985), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9980) );
  OR2_X1 U11980 ( .A1(n16198), .A2(n9983), .ZN(n9982) );
  NAND2_X1 U11981 ( .A1(n16198), .A2(n9663), .ZN(n9981) );
  NOR2_X1 U11982 ( .A1(n18616), .A2(n12179), .ZN(n12181) );
  NAND2_X1 U11983 ( .A1(n18598), .A2(n17960), .ZN(n15419) );
  INV_X4 U11984 ( .A(n16844), .ZN(n16945) );
  BUF_X4 U11985 ( .A(n11267), .Z(n16954) );
  INV_X1 U11986 ( .A(n18399), .ZN(n15616) );
  NOR2_X1 U11987 ( .A1(n15520), .A2(n15519), .ZN(n15417) );
  AND2_X1 U11988 ( .A1(n18597), .A2(n15516), .ZN(n17152) );
  INV_X1 U11989 ( .A(n17151), .ZN(n17190) );
  NAND2_X1 U11990 ( .A1(n17473), .A2(n10001), .ZN(n9930) );
  INV_X1 U11991 ( .A(n12136), .ZN(n9929) );
  NAND2_X1 U11992 ( .A1(n16198), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16195) );
  AOI21_X1 U11993 ( .B1(n16204), .B2(n17266), .A(n17529), .ZN(n17267) );
  OAI211_X1 U11994 ( .C1(n17301), .C2(n17653), .A(n17300), .B(n10077), .ZN(
        n17284) );
  NOR2_X1 U11995 ( .A1(n17284), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17283) );
  NOR2_X1 U11996 ( .A1(n9628), .A2(n9990), .ZN(n9989) );
  NOR2_X1 U11997 ( .A1(n17415), .A2(n9628), .ZN(n17366) );
  INV_X1 U11998 ( .A(n17471), .ZN(n17383) );
  OAI21_X1 U11999 ( .B1(n17399), .B2(n17618), .A(n17995), .ZN(n17471) );
  NAND2_X1 U12000 ( .A1(n17296), .A2(n9597), .ZN(n17399) );
  NOR2_X1 U12001 ( .A1(n17528), .A2(n11310), .ZN(n16207) );
  OR2_X1 U12002 ( .A1(n17454), .A2(n17308), .ZN(n17300) );
  NOR2_X1 U12003 ( .A1(n17315), .A2(n17767), .ZN(n17665) );
  NAND2_X1 U12004 ( .A1(n17330), .A2(n11305), .ZN(n17309) );
  AND2_X1 U12005 ( .A1(n9955), .A2(n9954), .ZN(n9953) );
  NAND2_X1 U12006 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17527), .ZN(
        n17466) );
  NOR2_X1 U12007 ( .A1(n17466), .A2(n17755), .ZN(n17446) );
  INV_X1 U12008 ( .A(n17488), .ZN(n17451) );
  NAND2_X1 U12009 ( .A1(n17493), .A2(n17838), .ZN(n17488) );
  NOR2_X1 U12010 ( .A1(n11473), .A2(n17525), .ZN(n17821) );
  NOR2_X1 U12011 ( .A1(n17526), .A2(n17862), .ZN(n17525) );
  XNOR2_X1 U12012 ( .A(n11294), .B(n11293), .ZN(n17542) );
  NAND2_X1 U12013 ( .A1(n17836), .A2(n9569), .ZN(n17859) );
  AND2_X1 U12014 ( .A1(n11451), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11281) );
  NAND2_X1 U12015 ( .A1(n18431), .A2(n9780), .ZN(n18403) );
  INV_X1 U12016 ( .A(n11493), .ZN(n9780) );
  NOR2_X1 U12017 ( .A1(n11489), .A2(n11493), .ZN(n9932) );
  NOR2_X1 U12018 ( .A1(n18615), .A2(n15519), .ZN(n18411) );
  NAND3_X1 U12019 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15523) );
  NAND2_X1 U12020 ( .A1(n18394), .A2(n18415), .ZN(n15522) );
  NOR2_X1 U12021 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17958), .ZN(n18247) );
  NAND3_X1 U12022 ( .A1(n11340), .A2(n11339), .A3(n11338), .ZN(n17969) );
  AOI211_X1 U12023 ( .C1(n11393), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n11337), .B(n11336), .ZN(n11338) );
  NAND3_X1 U12024 ( .A1(n11369), .A2(n11368), .A3(n11367), .ZN(n17981) );
  AOI211_X1 U12025 ( .C1(n16881), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n11366), .B(n11365), .ZN(n11367) );
  OR2_X1 U12026 ( .A1(n9777), .A2(n11346), .ZN(n17985) );
  NOR2_X1 U12027 ( .A1(n11443), .A2(n11430), .ZN(n18427) );
  NOR2_X1 U12028 ( .A1(n11491), .A2(n11490), .ZN(n18443) );
  NAND2_X1 U12029 ( .A1(n12154), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19966)
         );
  NOR2_X1 U12030 ( .A1(n15584), .A2(n20571), .ZN(n19701) );
  NAND2_X1 U12031 ( .A1(n12376), .A2(n10043), .ZN(n12377) );
  INV_X1 U12032 ( .A(n11659), .ZN(n10043) );
  INV_X1 U12033 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20813) );
  INV_X1 U12034 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14396) );
  INV_X1 U12035 ( .A(n19747), .ZN(n15639) );
  INV_X1 U12036 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13114) );
  AND2_X1 U12037 ( .A1(n13915), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19779) );
  XNOR2_X1 U12038 ( .A(n12031), .B(n12614), .ZN(n12958) );
  INV_X2 U12039 ( .A(n15629), .ZN(n19774) );
  AND2_X1 U12040 ( .A1(n15657), .A2(n12924), .ZN(n19766) );
  INV_X1 U12041 ( .A(n14530), .ZN(n19793) );
  INV_X1 U12042 ( .A(n14528), .ZN(n19792) );
  INV_X1 U12043 ( .A(n19797), .ZN(n14520) );
  INV_X1 U12044 ( .A(n15723), .ZN(n14589) );
  INV_X1 U12045 ( .A(n15726), .ZN(n14593) );
  AND2_X1 U12046 ( .A1(n15730), .A2(n12491), .ZN(n15728) );
  AND2_X1 U12047 ( .A1(n12497), .A2(n15721), .ZN(n14601) );
  NOR2_X1 U12048 ( .A1(n15922), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19817) );
  BUF_X1 U12049 ( .A(n19817), .Z(n20667) );
  BUF_X1 U12050 ( .A(n19898), .Z(n19895) );
  OR2_X1 U12051 ( .A1(n14632), .A2(n19967), .ZN(n9711) );
  AND2_X1 U12052 ( .A1(n14401), .A2(n14479), .ZN(n15749) );
  OR2_X1 U12053 ( .A1(n14485), .A2(n14484), .ZN(n15658) );
  AND2_X1 U12054 ( .A1(n14503), .A2(n14502), .ZN(n15754) );
  INV_X1 U12055 ( .A(n13450), .ZN(n19794) );
  NAND2_X1 U12056 ( .A1(n9823), .A2(n9821), .ZN(n9819) );
  NAND2_X1 U12057 ( .A1(n9703), .A2(n9702), .ZN(n14627) );
  NAND2_X1 U12058 ( .A1(n14625), .A2(n14777), .ZN(n9702) );
  NAND2_X1 U12059 ( .A1(n14626), .A2(n14764), .ZN(n9703) );
  AND2_X1 U12060 ( .A1(n15801), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14756) );
  AOI21_X1 U12061 ( .B1(n15889), .B2(n15813), .A(n15810), .ZN(n15809) );
  NAND2_X1 U12062 ( .A1(n9787), .A2(n9786), .ZN(n15819) );
  NAND2_X1 U12063 ( .A1(n19950), .A2(n9675), .ZN(n9786) );
  INV_X1 U12064 ( .A(n12022), .ZN(n9787) );
  NAND2_X1 U12065 ( .A1(n13062), .A2(n11882), .ZN(n9815) );
  INV_X1 U12066 ( .A(n19955), .ZN(n19936) );
  INV_X1 U12067 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20428) );
  INV_X1 U12068 ( .A(n19970), .ZN(n20052) );
  INV_X1 U12069 ( .A(n20518), .ZN(n20509) );
  INV_X1 U12070 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20256) );
  INV_X1 U12071 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19964) );
  OAI21_X1 U12072 ( .B1(n12823), .B2(n15926), .A(n20140), .ZN(n19963) );
  NAND2_X1 U12073 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n12822), .ZN(n14857) );
  NAND2_X1 U12074 ( .A1(n20100), .A2(n20474), .ZN(n20128) );
  INV_X1 U12075 ( .A(n20137), .ZN(n20158) );
  INV_X1 U12076 ( .A(n20218), .ZN(n20182) );
  OAI211_X1 U12077 ( .C1(n10078), .C2(n20386), .A(n20315), .B(n20262), .ZN(
        n20279) );
  INV_X1 U12078 ( .A(n20254), .ZN(n20278) );
  OAI22_X1 U12079 ( .A1(n20320), .A2(n20319), .B1(n20318), .B2(n20472), .ZN(
        n20344) );
  INV_X1 U12080 ( .A(n20378), .ZN(n20367) );
  OAI211_X1 U12081 ( .C1(n20496), .C2(n20481), .A(n20480), .B(n20479), .ZN(
        n20499) );
  INV_X1 U12082 ( .A(n20380), .ZN(n20510) );
  INV_X1 U12083 ( .A(n20394), .ZN(n20523) );
  INV_X1 U12084 ( .A(n20402), .ZN(n20535) );
  AND2_X1 U12085 ( .A1(n20002), .A2(n20001), .ZN(n20541) );
  INV_X1 U12086 ( .A(n20406), .ZN(n20542) );
  INV_X1 U12087 ( .A(n20414), .ZN(n20553) );
  AND2_X1 U12088 ( .A1(n20475), .A2(n20231), .ZN(n20564) );
  INV_X1 U12089 ( .A(n20419), .ZN(n20560) );
  NAND2_X1 U12090 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20666) );
  INV_X2 U12091 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20573) );
  INV_X1 U12092 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20570) );
  INV_X1 U12093 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19698) );
  NOR2_X1 U12094 ( .A1(n12220), .A2(n12272), .ZN(n12273) );
  AND2_X1 U12095 ( .A1(n10745), .A2(n10744), .ZN(n19670) );
  NOR2_X1 U12096 ( .A1(n18830), .A2(n15974), .ZN(n15961) );
  INV_X1 U12097 ( .A(n9909), .ZN(n15974) );
  OAI21_X1 U12098 ( .B1(n15994), .B2(n18830), .A(n9907), .ZN(n9909) );
  INV_X1 U12099 ( .A(n9908), .ZN(n9907) );
  OAI21_X1 U12100 ( .B1(n18830), .B2(n15933), .A(n9910), .ZN(n9908) );
  NOR2_X1 U12101 ( .A1(n15994), .A2(n18830), .ZN(n15982) );
  NOR2_X1 U12102 ( .A1(n15982), .A2(n15983), .ZN(n15981) );
  INV_X1 U12103 ( .A(n9828), .ZN(n15984) );
  NOR2_X1 U12104 ( .A1(n18830), .A2(n16015), .ZN(n16001) );
  OAI21_X1 U12105 ( .B1(n18644), .B2(n18830), .A(n9915), .ZN(n9918) );
  INV_X1 U12106 ( .A(n9916), .ZN(n9915) );
  OAI21_X1 U12107 ( .B1(n18830), .B2(n9917), .A(n16051), .ZN(n9916) );
  NOR2_X1 U12108 ( .A1(n18644), .A2(n18830), .ZN(n12219) );
  NOR2_X1 U12109 ( .A1(n12219), .A2(n15071), .ZN(n15545) );
  AND2_X1 U12110 ( .A1(n18814), .A2(n12211), .ZN(n18656) );
  OR2_X1 U12111 ( .A1(n18623), .A2(n12225), .ZN(n18792) );
  INV_X1 U12112 ( .A(n18742), .ZN(n18859) );
  INV_X1 U12113 ( .A(n19654), .ZN(n18847) );
  AND2_X1 U12114 ( .A1(n18623), .A2(n12707), .ZN(n18855) );
  INV_X1 U12115 ( .A(n18792), .ZN(n18853) );
  INV_X1 U12116 ( .A(n13006), .ZN(n10035) );
  OR2_X1 U12117 ( .A1(n10931), .A2(n10930), .ZN(n12751) );
  NOR2_X1 U12118 ( .A1(n10904), .A2(n10903), .ZN(n12867) );
  OR2_X1 U12119 ( .A1(n10874), .A2(n10873), .ZN(n12602) );
  AND2_X1 U12120 ( .A1(n12975), .A2(n9685), .ZN(n10037) );
  NAND2_X1 U12121 ( .A1(n10038), .A2(n12975), .ZN(n13961) );
  AND2_X1 U12122 ( .A1(n12348), .A2(n12989), .ZN(n14918) );
  NOR2_X1 U12123 ( .A1(n13212), .A2(n12166), .ZN(n18865) );
  NOR2_X1 U12124 ( .A1(n13212), .A2(n13211), .ZN(n18864) );
  INV_X1 U12125 ( .A(n18865), .ZN(n15006) );
  INV_X1 U12126 ( .A(n18864), .ZN(n15008) );
  NAND2_X1 U12127 ( .A1(n18892), .A2(n12993), .ZN(n15005) );
  NOR2_X1 U12128 ( .A1(n13270), .A2(n13269), .ZN(n13321) );
  AND2_X1 U12129 ( .A1(n12990), .A2(n12989), .ZN(n18892) );
  NAND2_X1 U12130 ( .A1(n18892), .A2(n10811), .ZN(n18868) );
  INV_X1 U12131 ( .A(n18868), .ZN(n18922) );
  AND2_X1 U12132 ( .A1(n18892), .A2(n12991), .ZN(n18921) );
  OAI21_X1 U12133 ( .B1(n12574), .B2(n12365), .A(n12432), .ZN(n12366) );
  NAND2_X1 U12134 ( .A1(n12273), .A2(n19683), .ZN(n12432) );
  INV_X1 U12135 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20721) );
  NAND2_X1 U12136 ( .A1(n16055), .A2(n9684), .ZN(n9922) );
  INV_X1 U12137 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16067) );
  NAND2_X1 U12138 ( .A1(n10059), .A2(n9603), .ZN(n16074) );
  INV_X1 U12139 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16094) );
  INV_X1 U12140 ( .A(n16121), .ZN(n18979) );
  AOI21_X1 U12141 ( .B1(n15930), .B2(n16150), .A(n14052), .ZN(n14053) );
  OR2_X1 U12142 ( .A1(n14051), .A2(n14050), .ZN(n14052) );
  OR2_X1 U12143 ( .A1(n15137), .A2(n15136), .ZN(n15138) );
  NAND2_X1 U12144 ( .A1(n9831), .A2(n13983), .ZN(n13532) );
  NAND2_X1 U12145 ( .A1(n15175), .A2(n9813), .ZN(n13553) );
  NAND2_X1 U12146 ( .A1(n9748), .A2(n10652), .ZN(n15171) );
  OR2_X1 U12147 ( .A1(n10798), .A2(n12842), .ZN(n15385) );
  AND2_X1 U12148 ( .A1(n10788), .A2(n15400), .ZN(n15365) );
  NAND2_X1 U12149 ( .A1(n15286), .A2(n9923), .ZN(n16052) );
  NAND2_X1 U12150 ( .A1(n10059), .A2(n10563), .ZN(n15390) );
  OAI21_X1 U12151 ( .B1(n13265), .B2(n13261), .A(n13262), .ZN(n13308) );
  CLKBUF_X1 U12152 ( .A(n13163), .Z(n13164) );
  AND2_X1 U12153 ( .A1(n9878), .A2(n12982), .ZN(n12838) );
  NAND2_X1 U12154 ( .A1(n9965), .A2(n11043), .ZN(n12847) );
  INV_X1 U12155 ( .A(n12727), .ZN(n9692) );
  AND2_X1 U12156 ( .A1(n19006), .A2(n15258), .ZN(n15400) );
  NOR2_X1 U12157 ( .A1(n12414), .A2(n12347), .ZN(n19663) );
  AND4_X1 U12158 ( .A1(n12345), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12346), 
        .A4(n19639), .ZN(n12347) );
  INV_X1 U12159 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10817) );
  INV_X1 U12160 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19651) );
  NAND2_X1 U12161 ( .A1(n12982), .A2(n10834), .ZN(n12731) );
  OAI21_X1 U12162 ( .B1(n12469), .B2(n12470), .A(n12545), .ZN(n19647) );
  AND2_X1 U12163 ( .A1(n12555), .A2(n12558), .ZN(n19636) );
  AND2_X1 U12164 ( .A1(n19087), .A2(n19632), .ZN(n19142) );
  INV_X1 U12165 ( .A(n19154), .ZN(n19172) );
  NOR2_X1 U12166 ( .A1(n19147), .A2(n19394), .ZN(n19197) );
  INV_X1 U12167 ( .A(n19505), .ZN(n19453) );
  INV_X1 U12168 ( .A(n19510), .ZN(n19461) );
  INV_X1 U12169 ( .A(n19520), .ZN(n19467) );
  INV_X1 U12170 ( .A(n19526), .ZN(n19470) );
  INV_X1 U12171 ( .A(n19532), .ZN(n19474) );
  INV_X1 U12172 ( .A(n19538), .ZN(n19477) );
  OAI21_X1 U12173 ( .B1(n19457), .B2(n19456), .A(n19455), .ZN(n19484) );
  NOR2_X2 U12174 ( .A1(n19395), .A2(n19394), .ZN(n19483) );
  INV_X1 U12175 ( .A(n19549), .ZN(n19482) );
  INV_X1 U12176 ( .A(n19398), .ZN(n19502) );
  AND2_X1 U12177 ( .A1(n9573), .A2(n19049), .ZN(n19506) );
  INV_X1 U12178 ( .A(n19404), .ZN(n19507) );
  INV_X1 U12179 ( .A(n19410), .ZN(n19512) );
  AND2_X1 U12180 ( .A1(n10704), .A2(n19049), .ZN(n19511) );
  INV_X1 U12181 ( .A(n19416), .ZN(n19517) );
  INV_X1 U12182 ( .A(n19422), .ZN(n19523) );
  INV_X1 U12183 ( .A(n19417), .ZN(n19521) );
  INV_X1 U12184 ( .A(n19418), .ZN(n19522) );
  INV_X1 U12185 ( .A(n19428), .ZN(n19529) );
  AND2_X1 U12186 ( .A1(n10468), .A2(n19049), .ZN(n19527) );
  INV_X1 U12187 ( .A(n19434), .ZN(n19535) );
  NOR2_X2 U12188 ( .A1(n19446), .A2(n19445), .ZN(n19544) );
  INV_X1 U12189 ( .A(n19444), .ZN(n19543) );
  AND2_X1 U12190 ( .A1(n19050), .A2(n19049), .ZN(n19539) );
  AND2_X1 U12191 ( .A1(n12683), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16167) );
  INV_X1 U12192 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19639) );
  AND2_X1 U12193 ( .A1(n12709), .A2(n12708), .ZN(n19550) );
  INV_X1 U12194 ( .A(n18620), .ZN(n18616) );
  NOR2_X1 U12195 ( .A1(n11489), .A2(n11487), .ZN(n16313) );
  NAND2_X1 U12196 ( .A1(n18606), .A2(n18430), .ZN(n17151) );
  NAND2_X1 U12197 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18608) );
  INV_X1 U12198 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18603) );
  NAND2_X1 U12199 ( .A1(n9774), .A2(n18606), .ZN(n16314) );
  OAI21_X1 U12200 ( .B1(n9776), .B2(n15520), .A(n9775), .ZN(n9774) );
  NAND2_X1 U12201 ( .A1(n18427), .A2(n18589), .ZN(n9775) );
  NAND2_X1 U12202 ( .A1(n18475), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18612) );
  NAND2_X1 U12203 ( .A1(n16369), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n10004) );
  NOR2_X1 U12204 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  NOR2_X1 U12205 ( .A1(n16658), .A2(n16371), .ZN(n10006) );
  INV_X1 U12206 ( .A(n16370), .ZN(n10007) );
  NOR2_X1 U12207 ( .A1(n16366), .A2(n16367), .ZN(n16365) );
  AOI21_X1 U12208 ( .B1(n16366), .B2(n16367), .A(n16659), .ZN(n10009) );
  INV_X1 U12209 ( .A(n16664), .ZN(n16590) );
  NOR2_X1 U12210 ( .A1(n16411), .A2(n10012), .ZN(n16402) );
  NOR2_X1 U12211 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16424), .ZN(n16414) );
  NAND2_X1 U12212 ( .A1(n10014), .A2(n10001), .ZN(n10011) );
  NOR2_X1 U12214 ( .A1(n16348), .A2(n10012), .ZN(n16443) );
  NOR2_X1 U12215 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16455), .ZN(n16445) );
  NOR2_X1 U12216 ( .A1(n12178), .A2(n17370), .ZN(n16348) );
  INV_X1 U12217 ( .A(n17389), .ZN(n9975) );
  INV_X1 U12218 ( .A(n9976), .ZN(n16465) );
  NOR2_X1 U12219 ( .A1(n16475), .A2(n17404), .ZN(n16474) );
  NOR2_X1 U12220 ( .A1(n17417), .A2(n10085), .ZN(n16483) );
  NOR2_X1 U12221 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16594), .ZN(n16577) );
  INV_X1 U12222 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20785) );
  NOR3_X1 U12223 ( .A1(n16855), .A2(n16974), .A3(n16973), .ZN(n16978) );
  NOR3_X2 U12224 ( .A1(n15419), .A2(n18450), .A3(n15614), .ZN(n16995) );
  NOR2_X1 U12225 ( .A1(n17220), .A2(n17013), .ZN(n17007) );
  INV_X1 U12226 ( .A(n17017), .ZN(n17014) );
  NAND2_X1 U12227 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17014), .ZN(n17013) );
  NOR2_X1 U12228 ( .A1(n17214), .A2(n17026), .ZN(n17022) );
  INV_X1 U12229 ( .A(n17032), .ZN(n17027) );
  NAND2_X1 U12230 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17027), .ZN(n17026) );
  NOR2_X1 U12231 ( .A1(n17200), .A2(n17064), .ZN(n17059) );
  NAND2_X1 U12232 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17077), .ZN(n17076) );
  NOR2_X2 U12233 ( .A1(n11390), .A2(n17136), .ZN(n17074) );
  NOR3_X1 U12234 ( .A1(n17143), .A2(n17111), .A3(n16997), .ZN(n16998) );
  AOI22_X1 U12235 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U12236 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11378) );
  AOI211_X1 U12237 ( .C1(n16934), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n11376), .B(n11375), .ZN(n11377) );
  NOR2_X1 U12238 ( .A1(n17245), .A2(n17106), .ZN(n17102) );
  INV_X1 U12239 ( .A(n12137), .ZN(n17118) );
  NOR2_X1 U12240 ( .A1(n11193), .A2(n11192), .ZN(n17121) );
  NAND2_X1 U12241 ( .A1(n15616), .A2(n17000), .ZN(n17138) );
  NAND2_X2 U12242 ( .A1(n17000), .A2(n17991), .ZN(n17136) );
  INV_X1 U12243 ( .A(n17147), .ZN(n17141) );
  INV_X1 U12244 ( .A(n17000), .ZN(n17143) );
  NAND2_X1 U12245 ( .A1(n17144), .A2(n17000), .ZN(n17142) );
  NOR2_X1 U12246 ( .A1(n15615), .A2(n17143), .ZN(n17147) );
  INV_X1 U12247 ( .A(n17138), .ZN(n17146) );
  NAND2_X1 U12248 ( .A1(n17190), .A2(n17152), .ZN(n17188) );
  NOR2_X1 U12249 ( .A1(n17192), .A2(n17234), .ZN(n17231) );
  BUF_X1 U12250 ( .A(n17231), .Z(n20800) );
  NAND2_X1 U12251 ( .A1(n16198), .A2(n9984), .ZN(n16178) );
  OAI22_X1 U12252 ( .A1(n17636), .A2(n17628), .B1(n17637), .B2(n17482), .ZN(
        n17292) );
  NAND2_X1 U12253 ( .A1(n17619), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n17460) );
  NOR2_X1 U12254 ( .A1(n17440), .A2(n17435), .ZN(n17688) );
  NOR2_X1 U12255 ( .A1(n17415), .A2(n17414), .ZN(n17400) );
  NAND2_X1 U12256 ( .A1(n17733), .A2(n17498), .ZN(n17424) );
  INV_X1 U12257 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17442) );
  INV_X1 U12258 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17497) );
  INV_X1 U12259 ( .A(n17516), .ZN(n17529) );
  INV_X1 U12260 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17534) );
  INV_X1 U12261 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17546) );
  INV_X1 U12262 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17555) );
  INV_X1 U12263 ( .A(n17619), .ZN(n17554) );
  INV_X1 U12264 ( .A(n17614), .ZN(n17607) );
  NOR2_X1 U12265 ( .A1(n17582), .A2(n17584), .ZN(n17619) );
  NOR2_X1 U12266 ( .A1(n16314), .A2(n17192), .ZN(n17615) );
  NAND2_X1 U12267 ( .A1(n17460), .A2(n17399), .ZN(n17614) );
  NAND2_X1 U12268 ( .A1(n9937), .A2(n11310), .ZN(n17274) );
  NAND2_X1 U12269 ( .A1(n17493), .A2(n9955), .ZN(n17432) );
  NOR2_X1 U12270 ( .A1(n17430), .A2(n11498), .ZN(n17866) );
  NOR2_X1 U12271 ( .A1(n17541), .A2(n9949), .ZN(n11498) );
  OR2_X1 U12272 ( .A1(n11297), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9949) );
  INV_X1 U12273 ( .A(n17850), .ZN(n17870) );
  NAND2_X1 U12274 ( .A1(n9945), .A2(n9946), .ZN(n17578) );
  NOR2_X1 U12275 ( .A1(n18590), .A2(n9563), .ZN(n17932) );
  INV_X1 U12276 ( .A(n18403), .ZN(n17942) );
  INV_X1 U12277 ( .A(n17939), .ZN(n17945) );
  INV_X1 U12278 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20820) );
  INV_X1 U12279 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15525) );
  OAI211_X1 U12280 ( .C1(n18450), .C2(n18433), .A(n17959), .B(n15521), .ZN(
        n18573) );
  INV_X1 U12281 ( .A(n16659), .ZN(n18452) );
  INV_X1 U12282 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18543) );
  INV_X1 U12283 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18475) );
  INV_X2 U12284 ( .A(n19966), .ZN(n19965) );
  NOR2_X1 U12285 ( .A1(n13021), .A2(n12167), .ZN(n16225) );
  INV_X1 U12287 ( .A(n14721), .ZN(n14454) );
  NAND2_X1 U12288 ( .A1(n14533), .A2(n9863), .ZN(n14535) );
  AND2_X1 U12289 ( .A1(n15730), .A2(n14532), .ZN(n9863) );
  AOI211_X1 U12290 ( .C1(n19916), .C2(n13919), .A(n13906), .B(n13905), .ZN(
        n13907) );
  INV_X1 U12291 ( .A(n9763), .ZN(n9762) );
  OAI21_X1 U12292 ( .B1(n14453), .B2(n19955), .A(n9764), .ZN(n9763) );
  NOR3_X1 U12293 ( .A1(n12131), .A2(n13955), .A3(n12130), .ZN(n9764) );
  OAI211_X1 U12294 ( .C1(n14722), .C2(n19925), .A(n9783), .B(n9781), .ZN(
        P1_U3001) );
  NAND2_X1 U12295 ( .A1(n14721), .A2(n19936), .ZN(n9781) );
  NOR2_X1 U12296 ( .A1(n9784), .A2(n14720), .ZN(n9783) );
  AOI21_X1 U12297 ( .B1(n14718), .B2(n14719), .A(n14717), .ZN(n9784) );
  NAND2_X1 U12298 ( .A1(n14034), .A2(n14033), .ZN(n14035) );
  OAI21_X1 U12299 ( .B1(n15155), .B2(n18984), .A(n10066), .ZN(n14004) );
  NOR2_X1 U12300 ( .A1(n14002), .A2(n10067), .ZN(n10066) );
  NAND2_X1 U12301 ( .A1(n15088), .A2(n9687), .ZN(P2_U2994) );
  NAND2_X1 U12302 ( .A1(n9688), .A2(n16102), .ZN(n9687) );
  OAI21_X1 U12303 ( .B1(n16052), .B2(n18984), .A(n9919), .ZN(P2_U2999) );
  AOI21_X1 U12304 ( .B1(n16054), .B2(n16102), .A(n9920), .ZN(n9919) );
  INV_X1 U12305 ( .A(n9921), .ZN(n9920) );
  AOI21_X1 U12306 ( .B1(n16053), .B2(n18988), .A(n9922), .ZN(n9921) );
  NOR2_X1 U12307 ( .A1(n9874), .A2(n15153), .ZN(n9873) );
  OAI21_X1 U12308 ( .B1(n10008), .B2(n16365), .A(n10002), .ZN(P3_U2642) );
  NOR2_X1 U12309 ( .A1(n16368), .A2(n10003), .ZN(n10002) );
  INV_X1 U12310 ( .A(n10009), .ZN(n10008) );
  NAND2_X1 U12311 ( .A1(n10005), .A2(n10004), .ZN(n10003) );
  AOI21_X1 U12312 ( .B1(n9934), .B2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n9928), .ZN(n9927) );
  AND2_X1 U12313 ( .A1(n11515), .A2(n11514), .ZN(n11516) );
  AOI21_X1 U12314 ( .B1(n12138), .B2(n17865), .A(n11513), .ZN(n11514) );
  INV_X1 U12315 ( .A(n10670), .ZN(n10063) );
  NOR2_X2 U12316 ( .A1(n11185), .A2(n11186), .ZN(n11269) );
  AND2_X1 U12317 ( .A1(n14091), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10384) );
  AND4_X1 U12318 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n9926), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U12319 ( .A1(n12198), .A2(n9615), .ZN(n12194) );
  INV_X1 U12320 ( .A(n13307), .ZN(n9693) );
  AND2_X1 U12321 ( .A1(n15362), .A2(n10057), .ZN(n9603) );
  NOR2_X1 U12322 ( .A1(n13561), .A2(n9853), .ZN(n14413) );
  AND2_X1 U12323 ( .A1(n9834), .A2(n9661), .ZN(n9604) );
  AOI22_X1 U12324 ( .A1(n9640), .A2(n14231), .B1(n14253), .B2(n14867), .ZN(
        n14862) );
  NOR2_X1 U12325 ( .A1(n14891), .A2(n14892), .ZN(n9605) );
  AOI21_X1 U12326 ( .B1(n15994), .B2(n15933), .A(n18830), .ZN(n9906) );
  AND2_X1 U12327 ( .A1(n19999), .A2(n19972), .ZN(n9606) );
  AND2_X1 U12328 ( .A1(n11310), .A2(n17454), .ZN(n9607) );
  AND2_X1 U12329 ( .A1(n12447), .A2(n12349), .ZN(n9608) );
  AND2_X1 U12330 ( .A1(n10557), .A2(n9666), .ZN(n9610) );
  AND2_X1 U12331 ( .A1(n11047), .A2(n11043), .ZN(n9611) );
  AND2_X1 U12332 ( .A1(n9603), .A2(n10088), .ZN(n9612) );
  NAND4_X2 U12333 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10858) );
  NAND2_X1 U12334 ( .A1(n10073), .A2(n10762), .ZN(n10774) );
  NAND2_X1 U12335 ( .A1(n12190), .A2(n12189), .ZN(n15543) );
  OR2_X1 U12336 ( .A1(n13270), .A2(n9885), .ZN(n13323) );
  NOR2_X1 U12337 ( .A1(n15351), .A2(n9664), .ZN(n13207) );
  OR2_X1 U12338 ( .A1(n10012), .A2(n17310), .ZN(n9613) );
  AND2_X1 U12339 ( .A1(n13008), .A2(n13010), .ZN(n9614) );
  AND2_X1 U12340 ( .A1(n9912), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9615) );
  AND2_X1 U12341 ( .A1(n11834), .A2(n11833), .ZN(n9616) );
  NAND2_X1 U12342 ( .A1(n15041), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15042) );
  NAND2_X1 U12343 ( .A1(n10035), .A2(n9614), .ZN(n10036) );
  AND2_X1 U12344 ( .A1(n10581), .A2(n9672), .ZN(n9617) );
  AND2_X1 U12345 ( .A1(n9902), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9618) );
  NAND2_X1 U12346 ( .A1(n14156), .A2(n14155), .ZN(n9619) );
  OR2_X1 U12347 ( .A1(n9857), .A2(n9856), .ZN(n9620) );
  AND2_X1 U12348 ( .A1(n15209), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9621) );
  NOR2_X1 U12349 ( .A1(n12772), .A2(n11990), .ZN(n11994) );
  INV_X1 U12350 ( .A(n11994), .ZN(n9707) );
  OR2_X1 U12351 ( .A1(n13337), .A2(n13359), .ZN(n9622) );
  AND2_X2 U12352 ( .A1(n14282), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10349) );
  INV_X1 U12353 ( .A(n9570), .ZN(n9937) );
  NAND2_X1 U12354 ( .A1(n10659), .A2(n10565), .ZN(n10567) );
  NAND2_X1 U12355 ( .A1(n17330), .A2(n17358), .ZN(n17359) );
  NAND2_X1 U12356 ( .A1(n10558), .A2(n10557), .ZN(n13259) );
  INV_X1 U12357 ( .A(n10247), .ZN(n10268) );
  NAND2_X1 U12358 ( .A1(n10336), .A2(n14093), .ZN(n9623) );
  AND2_X1 U12359 ( .A1(n14391), .A2(n13776), .ZN(n9624) );
  NOR2_X1 U12360 ( .A1(n18551), .A2(n18420), .ZN(n11264) );
  NOR2_X1 U12361 ( .A1(n13561), .A2(n13498), .ZN(n9625) );
  NOR2_X1 U12362 ( .A1(n15327), .A2(n15326), .ZN(n9626) );
  NAND2_X1 U12363 ( .A1(n9970), .A2(n9969), .ZN(n9627) );
  NAND2_X1 U12364 ( .A1(n9992), .A2(n9991), .ZN(n9628) );
  OR2_X1 U12365 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9629) );
  AND2_X1 U12366 ( .A1(n16041), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15039) );
  NOR2_X1 U12367 ( .A1(n14897), .A2(n14887), .ZN(n14879) );
  AND2_X2 U12368 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10337) );
  INV_X1 U12369 ( .A(n9934), .ZN(n16176) );
  OAI21_X1 U12370 ( .B1(n16177), .B2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n9935), .ZN(n9934) );
  AND2_X1 U12371 ( .A1(n10059), .A2(n10057), .ZN(n15359) );
  AND2_X1 U12372 ( .A1(n11686), .A2(n9849), .ZN(n9630) );
  AND3_X1 U12373 ( .A1(n12039), .A2(n12884), .A3(n9771), .ZN(n9631) );
  AND2_X1 U12374 ( .A1(n15175), .A2(n9811), .ZN(n9632) );
  NAND2_X1 U12375 ( .A1(n10308), .A2(n9636), .ZN(n10412) );
  AND2_X1 U12376 ( .A1(n14879), .A2(n14880), .ZN(n13533) );
  AND2_X1 U12377 ( .A1(n11168), .A2(n10551), .ZN(n9633) );
  NAND2_X1 U12378 ( .A1(n14327), .A2(n13904), .ZN(n13908) );
  INV_X1 U12379 ( .A(n10314), .ZN(n9734) );
  AND2_X1 U12380 ( .A1(n14667), .A2(n12128), .ZN(n9634) );
  AND2_X1 U12381 ( .A1(n9978), .A2(n9977), .ZN(n9635) );
  NOR2_X1 U12382 ( .A1(n14873), .A2(n14872), .ZN(n14871) );
  AND2_X1 U12383 ( .A1(n9598), .A2(n12349), .ZN(n9636) );
  AND3_X1 U12384 ( .A1(n9930), .A2(n12141), .A3(n9929), .ZN(n9637) );
  NOR2_X1 U12385 ( .A1(n10656), .A2(n10658), .ZN(n9638) );
  AND2_X1 U12386 ( .A1(n10069), .A2(n10239), .ZN(n9639) );
  AND2_X1 U12387 ( .A1(n14234), .A2(n10027), .ZN(n9640) );
  OR2_X1 U12388 ( .A1(n11130), .A2(n10269), .ZN(n9641) );
  AND3_X1 U12389 ( .A1(n10170), .A2(n10168), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9642) );
  AND2_X1 U12390 ( .A1(n9808), .A2(n15209), .ZN(n9643) );
  OAI21_X1 U12391 ( .B1(n15146), .B2(n16117), .A(n14001), .ZN(n14002) );
  INV_X1 U12392 ( .A(n12998), .ZN(n12043) );
  OR2_X1 U12393 ( .A1(n9632), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9644) );
  AND2_X1 U12394 ( .A1(n9607), .A2(n9937), .ZN(n9645) );
  AND2_X1 U12395 ( .A1(n12481), .A2(n12482), .ZN(n9646) );
  AND2_X1 U12396 ( .A1(n10081), .A2(n17269), .ZN(n9647) );
  NOR2_X1 U12397 ( .A1(n11168), .A2(n11173), .ZN(n9648) );
  AND2_X1 U12398 ( .A1(n14391), .A2(n9871), .ZN(n9649) );
  INV_X2 U12399 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10141) );
  AND2_X1 U12400 ( .A1(n9711), .A2(n14630), .ZN(n9650) );
  AND2_X1 U12401 ( .A1(n10422), .A2(n10420), .ZN(n9651) );
  NOR2_X1 U12402 ( .A1(n10653), .A2(n9749), .ZN(n9652) );
  INV_X1 U12403 ( .A(n10675), .ZN(n9744) );
  AND2_X1 U12404 ( .A1(n11525), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n9653) );
  AND2_X1 U12405 ( .A1(n9743), .A2(n9744), .ZN(n9654) );
  INV_X1 U12406 ( .A(n10827), .ZN(n10835) );
  INV_X1 U12407 ( .A(n9776), .ZN(n18439) );
  OR2_X1 U12408 ( .A1(n17859), .A2(n18598), .ZN(n9776) );
  NAND2_X1 U12409 ( .A1(n9988), .A2(n9992), .ZN(n12168) );
  OR2_X1 U12410 ( .A1(n12744), .A2(n9962), .ZN(n9655) );
  NAND2_X1 U12411 ( .A1(n20024), .A2(n11759), .ZN(n12955) );
  NOR2_X1 U12412 ( .A1(n13119), .A2(n13118), .ZN(n13106) );
  NAND2_X1 U12413 ( .A1(n9852), .A2(n9855), .ZN(n14432) );
  NAND2_X1 U12414 ( .A1(n14488), .A2(n14474), .ZN(n14405) );
  NOR2_X1 U12415 ( .A1(n12197), .A2(n16067), .ZN(n12198) );
  NOR2_X1 U12416 ( .A1(n12210), .A2(n15098), .ZN(n12212) );
  NOR2_X1 U12417 ( .A1(n12203), .A2(n16106), .ZN(n12204) );
  NOR2_X1 U12418 ( .A1(n12199), .A2(n18743), .ZN(n12200) );
  NOR2_X1 U12419 ( .A1(n12201), .A2(n16094), .ZN(n12202) );
  AND2_X1 U12420 ( .A1(n12198), .A2(n9911), .ZN(n12195) );
  AND2_X1 U12421 ( .A1(n12198), .A2(n9912), .ZN(n12196) );
  NAND2_X1 U12422 ( .A1(n9961), .A2(n9958), .ZN(n13028) );
  NOR2_X1 U12423 ( .A1(n13028), .A2(n13203), .ZN(n13202) );
  INV_X1 U12424 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15559) );
  AND2_X1 U12425 ( .A1(n13106), .A2(n13105), .ZN(n13227) );
  NOR2_X1 U12426 ( .A1(n11954), .A2(n11963), .ZN(n11957) );
  INV_X1 U12427 ( .A(n11957), .ZN(n9789) );
  NOR2_X1 U12428 ( .A1(n16134), .A2(n16135), .ZN(n15349) );
  AND2_X1 U12429 ( .A1(n15154), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9656) );
  NAND2_X1 U12430 ( .A1(n11690), .A2(n12814), .ZN(n12770) );
  INV_X1 U12431 ( .A(n10506), .ZN(n9836) );
  OR2_X1 U12432 ( .A1(n15328), .A2(n9887), .ZN(n9657) );
  NOR3_X1 U12433 ( .A1(n12628), .A2(n9655), .A3(n13004), .ZN(n13003) );
  OR2_X1 U12434 ( .A1(n9657), .A2(n15293), .ZN(n9658) );
  NAND2_X1 U12435 ( .A1(n10048), .A2(n10047), .ZN(n13445) );
  NAND2_X1 U12436 ( .A1(n9815), .A2(n11884), .ZN(n15777) );
  OR2_X1 U12437 ( .A1(n15351), .A2(n9657), .ZN(n15292) );
  NAND2_X1 U12438 ( .A1(n17405), .A2(n17528), .ZN(n17330) );
  NAND2_X1 U12439 ( .A1(n13409), .A2(n13410), .ZN(n13561) );
  INV_X1 U12440 ( .A(n13561), .ZN(n9852) );
  AND2_X1 U12441 ( .A1(n13558), .A2(n11921), .ZN(n9659) );
  NOR2_X1 U12442 ( .A1(n14905), .A2(n10033), .ZN(n14891) );
  NAND2_X1 U12443 ( .A1(n14884), .A2(n14886), .ZN(n14885) );
  INV_X1 U12444 ( .A(n10222), .ZN(n12345) );
  AND2_X1 U12445 ( .A1(n17493), .A2(n9953), .ZN(n17447) );
  NOR2_X1 U12446 ( .A1(n20053), .A2(n19970), .ZN(n9660) );
  AND2_X1 U12447 ( .A1(n10507), .A2(n9833), .ZN(n9661) );
  AND2_X1 U12448 ( .A1(n12234), .A2(n12235), .ZN(n12233) );
  NOR2_X1 U12449 ( .A1(n15351), .A2(n9658), .ZN(n9662) );
  AND2_X1 U12450 ( .A1(n15000), .A2(n15001), .ZN(n12234) );
  AND2_X1 U12451 ( .A1(n9984), .A2(n9983), .ZN(n9663) );
  AND2_X1 U12452 ( .A1(n12212), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12190) );
  NOR2_X1 U12453 ( .A1(n15351), .A2(n15328), .ZN(n15314) );
  INV_X1 U12454 ( .A(n14392), .ZN(n13776) );
  INV_X1 U12455 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20571) );
  INV_X1 U12456 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17618) );
  INV_X1 U12457 ( .A(n9758), .ZN(n9757) );
  OR2_X1 U12458 ( .A1(n14407), .A2(n9759), .ZN(n9758) );
  OR2_X1 U12459 ( .A1(n9658), .A2(n9888), .ZN(n9664) );
  INV_X1 U12460 ( .A(n9985), .ZN(n9984) );
  NAND2_X1 U12461 ( .A1(n9986), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9985) );
  AND2_X1 U12462 ( .A1(n10507), .A2(n10506), .ZN(n9665) );
  AND2_X1 U12463 ( .A1(n13312), .A2(n13310), .ZN(n9666) );
  AND2_X1 U12464 ( .A1(n10368), .A2(n10395), .ZN(n9667) );
  AND2_X1 U12465 ( .A1(n9973), .A2(n9972), .ZN(n9668) );
  AOI21_X1 U12466 ( .B1(n16412), .B2(n10001), .A(n9999), .ZN(n9996) );
  AND2_X1 U12467 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9669) );
  AND2_X1 U12468 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9670) );
  INV_X1 U12469 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16122) );
  INV_X1 U12470 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9990) );
  AND2_X1 U12471 ( .A1(n10038), .A2(n10037), .ZN(n12597) );
  NAND2_X1 U12472 ( .A1(n12981), .A2(n12980), .ZN(n12982) );
  AND2_X1 U12473 ( .A1(n16121), .A2(n19652), .ZN(n18988) );
  INV_X1 U12474 ( .A(n18988), .ZN(n16117) );
  NAND2_X1 U12475 ( .A1(n9966), .A2(n9970), .ZN(n12551) );
  NAND2_X1 U12476 ( .A1(n13232), .A2(n13231), .ZN(n13230) );
  NOR2_X1 U12477 ( .A1(n15543), .A2(n20721), .ZN(n15041) );
  OR2_X1 U12478 ( .A1(n14526), .A2(n14525), .ZN(n9671) );
  NAND2_X1 U12479 ( .A1(n10718), .A2(n10217), .ZN(n12220) );
  NAND2_X1 U12480 ( .A1(n13232), .A2(n9754), .ZN(n9751) );
  AND2_X1 U12481 ( .A1(n16121), .A2(n12336), .ZN(n16107) );
  INV_X1 U12482 ( .A(n16107), .ZN(n18992) );
  NOR2_X1 U12483 ( .A1(n12864), .A2(n12863), .ZN(n12627) );
  NOR2_X1 U12484 ( .A1(n12628), .A2(n12744), .ZN(n12745) );
  NOR2_X1 U12485 ( .A1(n13270), .A2(n9882), .ZN(n15370) );
  AOI21_X1 U12486 ( .B1(n11424), .B2(n11423), .A(n11426), .ZN(n18591) );
  INV_X1 U12487 ( .A(n10858), .ZN(n9804) );
  NAND2_X1 U12488 ( .A1(n11262), .A2(n12137), .ZN(n17528) );
  INV_X1 U12489 ( .A(n17528), .ZN(n17454) );
  OR2_X1 U12490 ( .A1(n10468), .A2(n12963), .ZN(n9672) );
  AND2_X1 U12491 ( .A1(n10188), .A2(n10187), .ZN(n11018) );
  OR2_X1 U12492 ( .A1(n10468), .A2(n10590), .ZN(n9673) );
  AOI21_X1 U12493 ( .B1(n18644), .B2(n9917), .A(n18830), .ZN(n9914) );
  AND2_X1 U12494 ( .A1(n10636), .A2(n9841), .ZN(n9674) );
  OR2_X1 U12495 ( .A1(n14785), .A2(n14781), .ZN(n9675) );
  INV_X1 U12496 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9993) );
  OR2_X1 U12497 ( .A1(n12845), .A2(n13962), .ZN(n13964) );
  OR2_X1 U12498 ( .A1(n10961), .A2(n10960), .ZN(n13010) );
  AND2_X1 U12499 ( .A1(n10035), .A2(n13008), .ZN(n9676) );
  OR2_X1 U12500 ( .A1(n12628), .A2(n9655), .ZN(n9677) );
  AND2_X1 U12501 ( .A1(n15041), .A2(n9902), .ZN(n9678) );
  NOR2_X1 U12502 ( .A1(n14863), .A2(n10026), .ZN(n9679) );
  AND2_X1 U12503 ( .A1(n9838), .A2(n18744), .ZN(n9680) );
  AOI21_X1 U12504 ( .B1(n12178), .B2(n10001), .A(n10014), .ZN(n10010) );
  AND2_X1 U12505 ( .A1(n9866), .A2(n13295), .ZN(n9681) );
  AND2_X1 U12506 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18396) );
  INV_X1 U12507 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10103) );
  AND2_X1 U12508 ( .A1(n12323), .A2(n19683), .ZN(n16114) );
  INV_X1 U12509 ( .A(n16114), .ZN(n18984) );
  BUF_X1 U12510 ( .A(n12456), .Z(n19005) );
  OR2_X1 U12511 ( .A1(n12324), .A2(n19683), .ZN(n18982) );
  INV_X1 U12512 ( .A(n18982), .ZN(n16102) );
  INV_X1 U12513 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9710) );
  AND2_X1 U12514 ( .A1(n16198), .A2(n9986), .ZN(n9682) );
  NAND3_X1 U12515 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .A3(n18553), .ZN(n18450) );
  AND2_X1 U12516 ( .A1(n12273), .A2(n12228), .ZN(n18852) );
  AND2_X1 U12517 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n9683) );
  INV_X1 U12518 ( .A(n14429), .ZN(n9856) );
  AND2_X1 U12519 ( .A1(n13523), .A2(n12191), .ZN(n13988) );
  OR2_X1 U12520 ( .A1(n16056), .A2(n16121), .ZN(n9684) );
  INV_X1 U12521 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n9839) );
  AND2_X1 U12522 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9685) );
  INV_X1 U12523 ( .A(n15781), .ZN(n19967) );
  AND2_X1 U12524 ( .A1(n12260), .A2(n20518), .ZN(n15781) );
  NAND2_X1 U12525 ( .A1(n17560), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16599) );
  INV_X1 U12526 ( .A(n14614), .ZN(n9715) );
  INV_X1 U12527 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18553) );
  INV_X1 U12528 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9987) );
  INV_X1 U12529 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n9954) );
  INV_X1 U12530 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9983) );
  INV_X1 U12531 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9814) );
  INV_X1 U12532 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9904) );
  AOI22_X2 U12533 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20014), .B1(DATAI_26_), 
        .B2(n20013), .ZN(n20534) );
  AOI22_X2 U12534 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20014), .B1(DATAI_28_), 
        .B2(n20013), .ZN(n20546) );
  AOI22_X2 U12535 ( .A1(DATAI_21_), .A2(n20013), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20014), .ZN(n20458) );
  NAND3_X1 U12536 ( .A1(n9686), .A2(n9667), .A3(n9803), .ZN(n11153) );
  NAND4_X1 U12537 ( .A1(n10383), .A2(n10380), .A3(n10381), .A4(n10382), .ZN(
        n9686) );
  NOR2_X2 U12538 ( .A1(n15108), .A2(n15096), .ZN(n15095) );
  OR2_X2 U12539 ( .A1(n15122), .A2(n15247), .ZN(n15108) );
  NAND2_X2 U12540 ( .A1(n15302), .A2(n15084), .ZN(n15122) );
  AND2_X2 U12541 ( .A1(n15327), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15302) );
  NAND2_X2 U12542 ( .A1(n10253), .A2(n9691), .ZN(n10274) );
  AND2_X2 U12543 ( .A1(n10210), .A2(n10211), .ZN(n10253) );
  XNOR2_X1 U12544 ( .A(n11140), .B(n9692), .ZN(n12741) );
  NAND2_X1 U12545 ( .A1(n10056), .A2(n13265), .ZN(n9694) );
  NAND2_X1 U12546 ( .A1(n10114), .A2(n10141), .ZN(n9695) );
  NAND2_X1 U12547 ( .A1(n10109), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9696) );
  AND2_X2 U12548 ( .A1(n9697), .A2(n12813), .ZN(n11612) );
  OAI21_X1 U12549 ( .B1(n14754), .B2(n19925), .A(n9698), .ZN(P1_U3004) );
  AND2_X1 U12550 ( .A1(n14752), .A2(n14753), .ZN(n9698) );
  NAND3_X2 U12551 ( .A1(n11915), .A2(n11916), .A3(n11914), .ZN(n14666) );
  AND2_X1 U12552 ( .A1(n14666), .A2(n14667), .ZN(n14778) );
  XNOR2_X2 U12553 ( .A(n9700), .B(n11670), .ZN(n20094) );
  NAND2_X2 U12554 ( .A1(n15737), .A2(n11920), .ZN(n14613) );
  NOR2_X2 U12555 ( .A1(n11815), .A2(n12854), .ZN(n11841) );
  AND2_X1 U12556 ( .A1(n9707), .A2(n11668), .ZN(n9709) );
  NAND2_X1 U12557 ( .A1(n11672), .A2(n11668), .ZN(n9848) );
  NAND4_X1 U12558 ( .A1(n11672), .A2(n9602), .A3(n9709), .A4(n9708), .ZN(n9845) );
  INV_X1 U12559 ( .A(n11666), .ZN(n11672) );
  NAND2_X1 U12560 ( .A1(n14631), .A2(n9650), .ZN(P1_U2972) );
  NOR2_X1 U12561 ( .A1(n9712), .A2(n9714), .ZN(n9713) );
  NAND3_X1 U12562 ( .A1(n14641), .A2(n9713), .A3(n9609), .ZN(n14625) );
  NAND2_X1 U12563 ( .A1(n11662), .A2(n9717), .ZN(n9716) );
  NAND2_X4 U12564 ( .A1(n11897), .A2(n11896), .ZN(n14777) );
  OAI21_X1 U12565 ( .B1(n13960), .B2(n19925), .A(n9762), .ZN(P1_U3000) );
  OAI21_X1 U12566 ( .B1(n12013), .B2(n19972), .A(n9720), .ZN(n11666) );
  NAND3_X1 U12567 ( .A1(n12927), .A2(n9723), .A3(n11665), .ZN(n9722) );
  NAND2_X1 U12568 ( .A1(n15779), .A2(n9724), .ZN(n9726) );
  NAND2_X1 U12569 ( .A1(n11884), .A2(n9725), .ZN(n9724) );
  NAND2_X1 U12570 ( .A1(n9727), .A2(n11882), .ZN(n9725) );
  NAND2_X1 U12571 ( .A1(n11894), .A2(n15901), .ZN(n15779) );
  NAND2_X1 U12572 ( .A1(n15787), .A2(n11864), .ZN(n13062) );
  INV_X1 U12573 ( .A(n11864), .ZN(n9727) );
  NAND2_X1 U12574 ( .A1(n15779), .A2(n11882), .ZN(n9728) );
  INV_X1 U12575 ( .A(n11894), .ZN(n9729) );
  NAND2_X1 U12576 ( .A1(n15785), .A2(n15784), .ZN(n15787) );
  OAI21_X1 U12577 ( .B1(n14730), .B2(n19925), .A(n14729), .ZN(P1_U3002) );
  NAND2_X1 U12578 ( .A1(n9732), .A2(n14777), .ZN(n9731) );
  NAND2_X1 U12579 ( .A1(n14626), .A2(n11921), .ZN(n9732) );
  AND2_X2 U12580 ( .A1(n10710), .A2(n9733), .ZN(n10170) );
  NAND2_X2 U12581 ( .A1(n10019), .A2(n10017), .ZN(n10704) );
  AND2_X2 U12582 ( .A1(n10214), .A2(n10202), .ZN(n10710) );
  NAND3_X1 U12583 ( .A1(n10431), .A2(n10430), .A3(n9736), .ZN(n10445) );
  XNOR2_X2 U12584 ( .A(n9738), .B(n10446), .ZN(n11158) );
  INV_X1 U12585 ( .A(n10447), .ZN(n9738) );
  NAND2_X1 U12586 ( .A1(n10447), .A2(n10446), .ZN(n10550) );
  NAND3_X1 U12587 ( .A1(n9741), .A2(n9742), .A3(n9739), .ZN(n13531) );
  NAND3_X1 U12588 ( .A1(n9740), .A2(n10675), .A3(n9745), .ZN(n9739) );
  NAND2_X1 U12589 ( .A1(n9831), .A2(n9743), .ZN(n9745) );
  NAND2_X1 U12590 ( .A1(n10671), .A2(n9744), .ZN(n9741) );
  NAND2_X1 U12591 ( .A1(n9831), .A2(n9654), .ZN(n9742) );
  INV_X1 U12592 ( .A(n9745), .ZN(n13557) );
  AND2_X2 U12593 ( .A1(n9748), .A2(n9746), .ZN(n15173) );
  NAND2_X1 U12594 ( .A1(n10647), .A2(n10646), .ZN(n15036) );
  INV_X1 U12595 ( .A(n10646), .ZN(n9749) );
  NAND2_X1 U12596 ( .A1(n10059), .A2(n9612), .ZN(n15052) );
  NOR2_X2 U12597 ( .A1(n19972), .A2(n19985), .ZN(n12477) );
  INV_X1 U12598 ( .A(n9761), .ZN(n14465) );
  NAND3_X1 U12599 ( .A1(n12929), .A2(n14331), .A3(n12529), .ZN(n9769) );
  NAND3_X1 U12600 ( .A1(n12039), .A2(n12884), .A3(n12043), .ZN(n13122) );
  NOR2_X2 U12601 ( .A1(n17981), .A2(n11390), .ZN(n11485) );
  NAND3_X1 U12602 ( .A1(n9778), .A2(n11349), .A3(n11348), .ZN(n9777) );
  INV_X1 U12603 ( .A(n11936), .ZN(n11952) );
  NAND2_X1 U12604 ( .A1(n9788), .A2(n11942), .ZN(n11945) );
  NAND2_X1 U12605 ( .A1(n9790), .A2(n9789), .ZN(n9788) );
  NAND2_X2 U12606 ( .A1(n19985), .A2(n12926), .ZN(n12927) );
  NAND2_X2 U12608 ( .A1(n9896), .A2(n9894), .ZN(n9798) );
  NAND2_X1 U12609 ( .A1(n9798), .A2(n11035), .ZN(n11036) );
  OAI21_X1 U12610 ( .B1(n9798), .B2(n11035), .A(n11034), .ZN(n11037) );
  NAND2_X1 U12611 ( .A1(n10277), .A2(n9798), .ZN(n9796) );
  OR2_X2 U12612 ( .A1(n9798), .A2(n10285), .ZN(n9797) );
  NAND2_X1 U12613 ( .A1(n14036), .A2(n9799), .ZN(P2_U2983) );
  OR2_X2 U12614 ( .A1(n14058), .A2(n18982), .ZN(n9799) );
  NAND2_X1 U12615 ( .A1(n14057), .A2(n9800), .ZN(P2_U3015) );
  OR2_X2 U12616 ( .A1(n14058), .A2(n16152), .ZN(n9800) );
  AND2_X4 U12617 ( .A1(n10337), .A2(n12581), .ZN(n14104) );
  NAND4_X1 U12618 ( .A1(n10328), .A2(n10326), .A3(n10325), .A4(n10327), .ZN(
        n9803) );
  NOR2_X4 U12619 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12813) );
  NAND2_X1 U12620 ( .A1(n14626), .A2(n9659), .ZN(n9826) );
  OAI21_X1 U12621 ( .B1(n14626), .B2(n9820), .A(n9817), .ZN(n14606) );
  NAND2_X1 U12622 ( .A1(n14626), .A2(n9818), .ZN(n9817) );
  AND2_X1 U12623 ( .A1(n9659), .A2(n14719), .ZN(n9818) );
  INV_X1 U12624 ( .A(n14626), .ZN(n9823) );
  AND2_X1 U12625 ( .A1(n9826), .A2(n9819), .ZN(n14607) );
  NAND2_X1 U12626 ( .A1(n9821), .A2(n14719), .ZN(n9820) );
  AOI21_X1 U12627 ( .B1(n14606), .B2(n15769), .A(n9824), .ZN(n11922) );
  NAND3_X1 U12628 ( .A1(n11759), .A2(n20571), .A3(n20024), .ZN(n9847) );
  NAND2_X1 U12629 ( .A1(n14015), .A2(n9827), .ZN(n10666) );
  OAI21_X1 U12630 ( .B1(n9830), .B2(n18810), .A(n9829), .ZN(n9828) );
  NAND2_X1 U12631 ( .A1(n18838), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9829) );
  XNOR2_X1 U12632 ( .A(n13981), .B(n10063), .ZN(n9831) );
  NAND3_X1 U12633 ( .A1(n9834), .A2(n10507), .A3(n9832), .ZN(n10564) );
  NAND2_X1 U12634 ( .A1(n10567), .A2(n9680), .ZN(n10579) );
  NAND2_X1 U12635 ( .A1(n10578), .A2(n9617), .ZN(n10605) );
  AND2_X1 U12636 ( .A1(n10582), .A2(n9840), .ZN(n18736) );
  XNOR2_X1 U12637 ( .A(n9840), .B(n9672), .ZN(n18725) );
  NAND2_X1 U12638 ( .A1(n9842), .A2(n10642), .ZN(n10643) );
  NAND2_X1 U12639 ( .A1(n10635), .A2(n10636), .ZN(n9842) );
  NAND2_X1 U12640 ( .A1(n9842), .A2(n10639), .ZN(n15549) );
  NAND2_X1 U12641 ( .A1(n9845), .A2(n9669), .ZN(n9846) );
  AND2_X2 U12642 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14844) );
  INV_X2 U12643 ( .A(n14777), .ZN(n15769) );
  OR2_X2 U12644 ( .A1(n20094), .A2(n11758), .ZN(n11759) );
  NAND2_X1 U12645 ( .A1(n9848), .A2(n9670), .ZN(n10044) );
  NAND2_X1 U12646 ( .A1(n11758), .A2(n11688), .ZN(n9849) );
  OAI21_X1 U12647 ( .B1(n12824), .B2(n12634), .A(n9858), .ZN(n12635) );
  XNOR2_X2 U12648 ( .A(n11766), .B(n11793), .ZN(n12824) );
  INV_X1 U12649 ( .A(n12634), .ZN(n9860) );
  NAND2_X1 U12650 ( .A1(n14346), .A2(n9861), .ZN(n9865) );
  INV_X1 U12651 ( .A(n13954), .ZN(n9864) );
  NAND3_X1 U12652 ( .A1(n13227), .A2(n13228), .A3(n13295), .ZN(n13379) );
  NAND2_X1 U12653 ( .A1(n9867), .A2(n12882), .ZN(n13119) );
  OAI21_X1 U12654 ( .B1(n12984), .B2(n9872), .A(n10821), .ZN(n12985) );
  OAI21_X1 U12655 ( .B1(n9565), .B2(n16152), .A(n9873), .ZN(P2_U3017) );
  OAI21_X1 U12656 ( .B1(n15155), .B2(n18994), .A(n9875), .ZN(n9874) );
  NAND2_X1 U12657 ( .A1(n11015), .A2(n9876), .ZN(n14306) );
  INV_X1 U12658 ( .A(n14306), .ZN(n14935) );
  NAND3_X1 U12659 ( .A1(n9878), .A2(n12839), .A3(n12982), .ZN(n12840) );
  NAND2_X2 U12660 ( .A1(n10761), .A2(n9566), .ZN(n12268) );
  NAND2_X1 U12661 ( .A1(n9596), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9893) );
  NAND3_X1 U12662 ( .A1(n10260), .A2(n10258), .A3(n10259), .ZN(n10287) );
  NAND2_X1 U12663 ( .A1(n10294), .A2(n10293), .ZN(n9896) );
  NAND3_X1 U12664 ( .A1(n12836), .A2(n11157), .A3(n9899), .ZN(n11165) );
  NAND2_X1 U12665 ( .A1(n11165), .A2(n10086), .ZN(n11163) );
  NAND2_X1 U12666 ( .A1(n9900), .A2(n18814), .ZN(n15941) );
  INV_X1 U12667 ( .A(n9918), .ZN(n15935) );
  OR2_X1 U12668 ( .A1(n15302), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9923) );
  NAND3_X1 U12669 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n9926), .A3(
        n9924), .ZN(n12203) );
  NOR2_X1 U12670 ( .A1(n16122), .A2(n9925), .ZN(n9924) );
  NAND3_X1 U12671 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n9926), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12206) );
  INV_X2 U12672 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18560) );
  NAND3_X1 U12673 ( .A1(n12142), .A2(n12140), .A3(n9927), .ZN(P3_U2799) );
  AND2_X2 U12674 ( .A1(n9933), .A2(n9932), .ZN(n18415) );
  NOR2_X1 U12675 ( .A1(n9570), .A2(n9607), .ZN(n16204) );
  INV_X2 U12676 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18575) );
  NAND2_X1 U12677 ( .A1(n9939), .A2(n9943), .ZN(n9938) );
  NAND2_X1 U12678 ( .A1(n9940), .A2(n17580), .ZN(n9943) );
  INV_X1 U12679 ( .A(n9947), .ZN(n9939) );
  INV_X1 U12680 ( .A(n17590), .ZN(n9945) );
  INV_X1 U12681 ( .A(n17580), .ZN(n9948) );
  INV_X1 U12682 ( .A(n9943), .ZN(n9946) );
  INV_X1 U12683 ( .A(n11286), .ZN(n9940) );
  NAND2_X1 U12684 ( .A1(n9942), .A2(n9944), .ZN(n17564) );
  INV_X1 U12685 ( .A(n17566), .ZN(n9941) );
  NOR2_X1 U12686 ( .A1(n17590), .A2(n11286), .ZN(n17579) );
  NAND2_X1 U12687 ( .A1(n9950), .A2(n9952), .ZN(n17513) );
  NOR2_X1 U12688 ( .A1(n11294), .A2(n11293), .ZN(n11297) );
  INV_X1 U12689 ( .A(n12628), .ZN(n9961) );
  NAND2_X1 U12690 ( .A1(n9965), .A2(n9611), .ZN(n12845) );
  INV_X1 U12691 ( .A(n13964), .ZN(n9966) );
  NAND2_X1 U12692 ( .A1(n9966), .A2(n9967), .ZN(n12864) );
  INV_X1 U12693 ( .A(n9979), .ZN(n16381) );
  INV_X1 U12694 ( .A(n9978), .ZN(n16374) );
  OR2_X1 U12695 ( .A1(n16392), .A2(n10012), .ZN(n9979) );
  NAND3_X1 U12696 ( .A1(n9982), .A2(n9981), .A3(n9980), .ZN(n12176) );
  INV_X1 U12697 ( .A(n17415), .ZN(n9988) );
  NAND2_X1 U12698 ( .A1(n9988), .A2(n9989), .ZN(n17345) );
  NOR2_X2 U12699 ( .A1(n9995), .A2(n9994), .ZN(n16393) );
  INV_X1 U12700 ( .A(n12178), .ZN(n10013) );
  OAI21_X2 U12701 ( .B1(n10013), .B2(n10012), .A(n10011), .ZN(n16434) );
  NAND2_X1 U12702 ( .A1(n10018), .A2(n10141), .ZN(n10017) );
  NAND4_X1 U12703 ( .A1(n10155), .A2(n10154), .A3(n10152), .A4(n10153), .ZN(
        n10018) );
  NAND2_X1 U12704 ( .A1(n10020), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10019) );
  NAND4_X1 U12705 ( .A1(n10159), .A2(n10158), .A3(n10156), .A4(n10157), .ZN(
        n10020) );
  OAI21_X1 U12706 ( .B1(n11130), .B2(n10240), .A(n9639), .ZN(n10241) );
  NAND2_X1 U12707 ( .A1(n14253), .A2(n9679), .ZN(n10021) );
  NAND2_X1 U12708 ( .A1(n14231), .A2(n14234), .ZN(n14873) );
  NAND3_X1 U12709 ( .A1(n10031), .A2(n10032), .A3(n9619), .ZN(n10029) );
  NAND2_X1 U12710 ( .A1(n14132), .A2(n14156), .ZN(n10031) );
  INV_X1 U12711 ( .A(n10036), .ZN(n13190) );
  NAND2_X1 U12712 ( .A1(n12555), .A2(n12546), .ZN(n12979) );
  AND3_X2 U12713 ( .A1(n10762), .A2(n10071), .A3(n10767), .ZN(n10247) );
  AND2_X4 U12714 ( .A1(n11526), .A2(n11525), .ZN(n13731) );
  NAND2_X1 U12715 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11639) );
  AOI22_X1 U12716 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13731), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U12717 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13731), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11533) );
  AOI21_X1 U12718 ( .B1(n11806), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n10041), .ZN(n11569) );
  NAND2_X1 U12719 ( .A1(n11774), .A2(n11772), .ZN(n10042) );
  AND2_X2 U12720 ( .A1(n11633), .A2(n19972), .ZN(n11659) );
  NAND2_X1 U12721 ( .A1(n13330), .A2(n11903), .ZN(n10048) );
  NAND2_X2 U12722 ( .A1(n14708), .A2(n13446), .ZN(n13481) );
  NAND2_X1 U12723 ( .A1(n10050), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10049) );
  NAND4_X1 U12724 ( .A1(n10163), .A2(n10162), .A3(n10160), .A4(n10161), .ZN(
        n10050) );
  NAND2_X1 U12725 ( .A1(n10052), .A2(n10141), .ZN(n10051) );
  NAND4_X1 U12726 ( .A1(n10167), .A2(n10165), .A3(n10166), .A4(n10164), .ZN(
        n10052) );
  NAND2_X1 U12727 ( .A1(n10558), .A2(n9610), .ZN(n10059) );
  NAND2_X1 U12728 ( .A1(n13982), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10065) );
  INV_X1 U12729 ( .A(n10238), .ZN(n10762) );
  NAND3_X1 U12730 ( .A1(n10767), .A2(n10070), .A3(n10762), .ZN(n10069) );
  NAND3_X1 U12731 ( .A1(n11168), .A2(n10551), .A3(n9804), .ZN(n10074) );
  NAND2_X1 U12732 ( .A1(n10074), .A2(n18802), .ZN(n10556) );
  NAND2_X1 U12733 ( .A1(n11659), .A2(n19824), .ZN(n19828) );
  NAND2_X1 U12734 ( .A1(n14876), .A2(n14878), .ZN(n14877) );
  XNOR2_X1 U12735 ( .A(n14204), .B(n14205), .ZN(n14876) );
  NAND2_X1 U12736 ( .A1(n12470), .A2(n12469), .ZN(n12545) );
  OAI21_X1 U12737 ( .B1(n12511), .B2(n19827), .A(n11785), .ZN(n11787) );
  NAND2_X1 U12738 ( .A1(n12545), .A2(n12544), .ZN(n12557) );
  INV_X1 U12739 ( .A(n12547), .ZN(n12541) );
  AND2_X1 U12740 ( .A1(n12468), .A2(n12419), .ZN(n19654) );
  INV_X1 U12741 ( .A(n11022), .ZN(n14026) );
  NAND2_X1 U12742 ( .A1(n11022), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10259) );
  OAI22_X4 U12743 ( .A1(n14031), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12317), 
        .B2(n14025), .ZN(n18814) );
  NAND2_X1 U12744 ( .A1(n10283), .A2(n10282), .ZN(n10284) );
  AOI21_X1 U12745 ( .B1(n9598), .B2(n12455), .A(n12416), .ZN(n12417) );
  XNOR2_X1 U12746 ( .A(n11786), .B(n11787), .ZN(n12889) );
  NOR2_X1 U12747 ( .A1(n10255), .A2(n10254), .ZN(n10260) );
  AOI22_X1 U12748 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10123) );
  AND2_X1 U12749 ( .A1(n10279), .A2(n10280), .ZN(n10277) );
  AOI22_X1 U12750 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U12751 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U12752 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10110) );
  OR2_X1 U12753 ( .A1(n15596), .A2(n16183), .ZN(n10075) );
  AND2_X1 U12754 ( .A1(n15596), .A2(n11311), .ZN(n10076) );
  OR2_X1 U12755 ( .A1(n17528), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10077) );
  AND2_X2 U12756 ( .A1(n18968), .A2(n19679), .ZN(n18966) );
  NOR2_X1 U12757 ( .A1(n20379), .A2(n20348), .ZN(n10078) );
  NOR2_X1 U12758 ( .A1(n11501), .A2(n11282), .ZN(n10079) );
  NOR2_X1 U12759 ( .A1(n17264), .A2(n17263), .ZN(n10081) );
  OR2_X1 U12760 ( .A1(n15599), .A2(n16191), .ZN(n10084) );
  AND2_X1 U12761 ( .A1(n12176), .A2(n10089), .ZN(n10085) );
  AND2_X1 U12762 ( .A1(n9633), .A2(n11164), .ZN(n10086) );
  NAND2_X1 U12763 ( .A1(n17454), .A2(n17630), .ZN(n10087) );
  INV_X2 U12764 ( .A(n18612), .ZN(n18532) );
  INV_X1 U12765 ( .A(n14290), .ZN(n14263) );
  NAND2_X1 U12766 ( .A1(n10575), .A2(n11075), .ZN(n10088) );
  INV_X1 U12767 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14437) );
  INV_X1 U12768 ( .A(n12166), .ZN(n13211) );
  INV_X1 U12769 ( .A(n10295), .ZN(n12447) );
  INV_X1 U12770 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19633) );
  OR2_X1 U12771 ( .A1(n16491), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10089) );
  AND2_X1 U12772 ( .A1(n15016), .A2(n15014), .ZN(n10090) );
  INV_X1 U12773 ( .A(n13607), .ZN(n13706) );
  INV_X1 U12774 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15917) );
  INV_X1 U12775 ( .A(n20140), .ZN(n20001) );
  NAND2_X1 U12776 ( .A1(n20571), .A2(n19971), .ZN(n20140) );
  AND2_X1 U12777 ( .A1(n19824), .A2(n19823), .ZN(n19899) );
  OR2_X1 U12778 ( .A1(n19802), .A2(n20667), .ZN(n19801) );
  INV_X2 U12779 ( .A(n19801), .ZN(n19820) );
  INV_X1 U12780 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11288) );
  INV_X1 U12781 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14425) );
  AND2_X1 U12782 ( .A1(n17192), .A2(n17238), .ZN(n17246) );
  INV_X2 U12783 ( .A(n17246), .ZN(n17244) );
  OR2_X1 U12784 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10091) );
  NOR2_X1 U12785 ( .A1(n20379), .A2(n20187), .ZN(n10092) );
  AND2_X1 U12786 ( .A1(n10257), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10094) );
  INV_X1 U12787 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U12788 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15608), .ZN(n19555) );
  INV_X1 U12789 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12670) );
  INV_X1 U12790 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12648) );
  INV_X1 U12791 ( .A(n10812), .ZN(n11004) );
  AND2_X1 U12792 ( .A1(n16995), .A2(n17991), .ZN(n16993) );
  INV_X2 U12793 ( .A(n16993), .ZN(n16984) );
  NOR2_X1 U12794 ( .A1(n11183), .A2(n11185), .ZN(n11267) );
  INV_X1 U12795 ( .A(n10279), .ZN(n10281) );
  AND2_X1 U12796 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10096) );
  AND3_X1 U12797 ( .A1(n11571), .A2(n11570), .A3(n11569), .ZN(n10097) );
  OR2_X1 U12798 ( .A1(n12246), .A2(n19972), .ZN(n10098) );
  AND2_X1 U12799 ( .A1(n11702), .A2(n20015), .ZN(n10099) );
  AND4_X1 U12800 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n10101) );
  OR2_X1 U12801 ( .A1(n11832), .A2(n11831), .ZN(n11855) );
  NAND2_X1 U12802 ( .A1(n10238), .A2(n10221), .ZN(n10215) );
  INV_X1 U12803 ( .A(n11899), .ZN(n11723) );
  AND2_X1 U12804 ( .A1(n15584), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11681) );
  XNOR2_X1 U12805 ( .A(n11518), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11929) );
  OAI22_X1 U12806 ( .A1(n10310), .A2(n10426), .B1(n10412), .B2(n10309), .ZN(
        n10311) );
  OR2_X1 U12807 ( .A1(n10467), .A2(n10219), .ZN(n10228) );
  INV_X1 U12808 ( .A(n11939), .ZN(n11934) );
  NOR2_X1 U12809 ( .A1(n11723), .A2(n11800), .ZN(n11740) );
  AOI22_X1 U12810 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10329), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10181) );
  INV_X1 U12811 ( .A(n10228), .ZN(n10220) );
  INV_X1 U12812 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U12813 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10157) );
  AOI21_X1 U12814 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20820), .A(
        n11405), .ZN(n11406) );
  INV_X1 U12815 ( .A(n15632), .ZN(n13745) );
  INV_X1 U12816 ( .A(n13953), .ZN(n13670) );
  OR2_X1 U12817 ( .A1(n11701), .A2(n11700), .ZN(n11703) );
  OR2_X1 U12818 ( .A1(n11874), .A2(n11873), .ZN(n11888) );
  NAND3_X1 U12819 ( .A1(n19999), .A2(n19972), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11954) );
  INV_X1 U12820 ( .A(n10662), .ZN(n10663) );
  OR2_X1 U12821 ( .A1(n14129), .A2(n14128), .ZN(n14151) );
  INV_X1 U12822 ( .A(n10350), .ZN(n13418) );
  OAI21_X1 U12823 ( .B1(n16121), .B2(n13999), .A(n15151), .ZN(n14000) );
  AND2_X1 U12824 ( .A1(n10632), .A2(n15078), .ZN(n10633) );
  INV_X1 U12825 ( .A(n12542), .ZN(n12540) );
  NAND2_X1 U12826 ( .A1(n10119), .A2(n10141), .ZN(n10126) );
  INV_X1 U12827 ( .A(n12512), .ZN(n13793) );
  NAND2_X1 U12828 ( .A1(n13746), .A2(n13745), .ZN(n13747) );
  INV_X1 U12829 ( .A(n13289), .ZN(n12916) );
  INV_X1 U12830 ( .A(n13096), .ZN(n13097) );
  INV_X1 U12831 ( .A(n11703), .ZN(n11817) );
  INV_X1 U12832 ( .A(n11954), .ZN(n11958) );
  NAND2_X1 U12833 ( .A1(n10184), .A2(n10141), .ZN(n10185) );
  OR2_X1 U12834 ( .A1(n10443), .A2(n10442), .ZN(n10481) );
  OR2_X1 U12835 ( .A1(n14181), .A2(n14180), .ZN(n14182) );
  INV_X1 U12836 ( .A(n10291), .ZN(n11034) );
  INV_X1 U12837 ( .A(n10828), .ZN(n11003) );
  AOI22_X1 U12838 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18405), .B2(n18568), .ZN(
        n11420) );
  OAI22_X1 U12839 ( .A1(n11416), .A2(n18425), .B1(n11415), .B2(n11414), .ZN(
        n11422) );
  AND2_X1 U12840 ( .A1(n17372), .A2(n17262), .ZN(n17263) );
  AND2_X1 U12841 ( .A1(n17454), .A2(n18552), .ZN(n11313) );
  NOR2_X1 U12842 ( .A1(n17144), .A2(n11484), .ZN(n11497) );
  NOR2_X1 U12843 ( .A1(n17128), .A2(n11287), .ZN(n11263) );
  INV_X1 U12844 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15452) );
  INV_X1 U12845 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n20729) );
  INV_X1 U12846 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20819) );
  AND2_X1 U12847 ( .A1(n12086), .A2(n12085), .ZN(n14493) );
  OR2_X1 U12848 ( .A1(n13674), .A2(n14482), .ZN(n13693) );
  INV_X1 U12849 ( .A(n13793), .ZN(n13900) );
  INV_X1 U12850 ( .A(n13797), .ZN(n13952) );
  INV_X1 U12851 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19727) );
  NAND2_X1 U12852 ( .A1(n11654), .A2(n10099), .ZN(n11667) );
  INV_X1 U12853 ( .A(n20190), .ZN(n20225) );
  AND2_X1 U12854 ( .A1(n20379), .A2(n20503), .ZN(n20312) );
  INV_X1 U12855 ( .A(n13007), .ZN(n13008) );
  NAND3_X1 U12856 ( .A1(n12345), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n9573), 
        .ZN(n14227) );
  INV_X1 U12857 ( .A(n13010), .ZN(n13009) );
  XNOR2_X1 U12858 ( .A(n11034), .B(n11033), .ZN(n10292) );
  AND2_X1 U12859 ( .A1(n10668), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15169) );
  NAND2_X1 U12860 ( .A1(n12340), .A2(n12455), .ZN(n12344) );
  CLKBUF_X3 U12861 ( .A(n11330), .Z(n15501) );
  OR2_X1 U12862 ( .A1(n11490), .A2(n15419), .ZN(n17189) );
  NOR2_X1 U12863 ( .A1(n11314), .A2(n11313), .ZN(n11315) );
  NOR2_X1 U12864 ( .A1(n18590), .A2(n17118), .ZN(n16208) );
  NAND2_X1 U12865 ( .A1(n11263), .A2(n17124), .ZN(n11290) );
  NOR2_X1 U12866 ( .A1(n11479), .A2(n17969), .ZN(n11477) );
  AND2_X1 U12867 ( .A1(n12485), .A2(n11975), .ZN(n12375) );
  INV_X1 U12868 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15699) );
  INV_X1 U12869 ( .A(n19779), .ZN(n19728) );
  OR3_X1 U12870 ( .A1(n12934), .A2(n12931), .A3(n12930), .ZN(n15629) );
  AND3_X1 U12871 ( .A1(n12065), .A2(n12090), .A3(n12064), .ZN(n14525) );
  OR2_X1 U12872 ( .A1(n14346), .A2(n13903), .ZN(n13904) );
  NAND2_X1 U12873 ( .A1(n11675), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13607) );
  NOR2_X1 U12874 ( .A1(n12247), .A2(n12246), .ZN(n15572) );
  AND2_X1 U12875 ( .A1(n12072), .A2(n12071), .ZN(n14513) );
  NAND2_X1 U12876 ( .A1(n12794), .A2(n12793), .ZN(n15561) );
  AND2_X1 U12877 ( .A1(n11814), .A2(n11813), .ZN(n12854) );
  NOR2_X1 U12878 ( .A1(n20141), .A2(n20140), .ZN(n20480) );
  AOI21_X1 U12879 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20428), .A(n20140), 
        .ZN(n20516) );
  NOR2_X1 U12880 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12706) );
  INV_X1 U12881 ( .A(n13202), .ZN(n13339) );
  AND2_X1 U12882 ( .A1(n10951), .A2(n10950), .ZN(n15328) );
  NAND2_X1 U12883 ( .A1(n18892), .A2(n12994), .ZN(n13212) );
  INV_X1 U12884 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15117) );
  INV_X1 U12885 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12760) );
  INV_X1 U12886 ( .A(n16150), .ZN(n18995) );
  NOR2_X1 U12887 ( .A1(n10739), .A2(n12239), .ZN(n19669) );
  OR2_X1 U12888 ( .A1(n12557), .A2(n12556), .ZN(n12558) );
  NOR2_X1 U12889 ( .A1(n19636), .A2(n19633), .ZN(n19225) );
  INV_X1 U12890 ( .A(n19632), .ZN(n19303) );
  OR2_X1 U12891 ( .A1(n19389), .A2(n19384), .ZN(n19438) );
  INV_X1 U12892 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19493) );
  NOR2_X1 U12893 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16444), .ZN(n16435) );
  NOR2_X1 U12894 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16476), .ZN(n16466) );
  INV_X1 U12895 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16857) );
  INV_X1 U12896 ( .A(n17136), .ZN(n17058) );
  NAND2_X1 U12897 ( .A1(n11426), .A2(n11425), .ZN(n18430) );
  NOR2_X1 U12898 ( .A1(n18600), .A2(n17189), .ZN(n17191) );
  INV_X1 U12899 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17483) );
  INV_X1 U12900 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17585) );
  INV_X1 U12901 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16215) );
  NOR2_X1 U12902 ( .A1(n17630), .A2(n17298), .ZN(n17637) );
  NOR2_X1 U12903 ( .A1(n11303), .A2(n11302), .ZN(n17340) );
  INV_X1 U12904 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17435) );
  INV_X1 U12905 ( .A(n18411), .ZN(n18429) );
  INV_X1 U12906 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18405) );
  AOI21_X1 U12907 ( .B1(n17950), .B2(n18602), .A(n18569), .ZN(n17958) );
  NOR2_X1 U12908 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18543), .ZN(n18329) );
  NAND2_X1 U12909 ( .A1(n19828), .A2(n12426), .ZN(n20664) );
  OR3_X1 U12910 ( .A1(n12934), .A2(n12926), .A3(n12928), .ZN(n19747) );
  OR3_X1 U12911 ( .A1(n19725), .A2(n15697), .A3(n14402), .ZN(n14419) );
  AND2_X1 U12912 ( .A1(n13915), .A2(n12922), .ZN(n19755) );
  AND2_X1 U12913 ( .A1(n13915), .A2(n12936), .ZN(n19778) );
  INV_X1 U12914 ( .A(n19761), .ZN(n19773) );
  INV_X1 U12915 ( .A(n20015), .ZN(n14532) );
  AND2_X1 U12916 ( .A1(n15730), .A2(n12494), .ZN(n13909) );
  INV_X2 U12917 ( .A(n19901), .ZN(n19894) );
  NAND2_X1 U12918 ( .A1(n13711), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13773) );
  AND2_X1 U12919 ( .A1(n13405), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13494) );
  NAND2_X1 U12920 ( .A1(n13221), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13289) );
  INV_X2 U12921 ( .A(n14677), .ZN(n19914) );
  INV_X1 U12922 ( .A(n12895), .ZN(n15889) );
  NOR2_X1 U12923 ( .A1(n14823), .A2(n12894), .ZN(n19945) );
  INV_X1 U12924 ( .A(n19925), .ZN(n19952) );
  NOR2_X1 U12925 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19700) );
  OAI22_X1 U12926 ( .A1(n19982), .A2(n19981), .B1(n20318), .B2(n20136), .ZN(
        n20020) );
  OAI22_X1 U12927 ( .A1(n20062), .A2(n20061), .B1(n20194), .B2(n20318), .ZN(
        n20086) );
  AND2_X1 U12928 ( .A1(n19969), .A2(n19968), .ZN(n20100) );
  OAI221_X1 U12929 ( .B1(n10092), .B2(n20386), .C1(n10092), .C2(n20142), .A(
        n20480), .ZN(n20159) );
  OAI22_X1 U12930 ( .A1(n20196), .A2(n20195), .B1(n20194), .B2(n20473), .ZN(
        n20220) );
  INV_X1 U12931 ( .A(n20355), .ZN(n20231) );
  INV_X1 U12932 ( .A(n20342), .ZN(n20310) );
  OR2_X1 U12933 ( .A1(n20053), .A2(n20052), .ZN(n20287) );
  OAI211_X1 U12934 ( .C1(n20320), .C2(n20317), .A(n20316), .B(n20315), .ZN(
        n20345) );
  OAI22_X1 U12935 ( .A1(n20391), .A2(n20390), .B1(n20473), .B2(n20389), .ZN(
        n20421) );
  AND2_X1 U12936 ( .A1(n20475), .A2(n9660), .ZN(n20466) );
  INV_X1 U12937 ( .A(n20398), .ZN(n20529) );
  INV_X1 U12938 ( .A(n20410), .ZN(n20547) );
  AND2_X1 U12939 ( .A1(n15581), .A2(n15580), .ZN(n15586) );
  INV_X1 U12940 ( .A(n20666), .ZN(n20585) );
  INV_X1 U12941 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20592) );
  NAND2_X1 U12942 ( .A1(n12679), .A2(n12989), .ZN(n12272) );
  INV_X1 U12943 ( .A(n18852), .ZN(n18810) );
  AND2_X1 U12944 ( .A1(n10991), .A2(n10990), .ZN(n13437) );
  NOR2_X1 U12945 ( .A1(n18853), .A2(n19639), .ZN(n18838) );
  INV_X1 U12946 ( .A(n19555), .ZN(n18818) );
  AND2_X1 U12947 ( .A1(n18973), .A2(n19633), .ZN(n18854) );
  OR2_X1 U12948 ( .A1(n10974), .A2(n10973), .ZN(n13189) );
  OR2_X1 U12949 ( .A1(n10917), .A2(n10916), .ZN(n12748) );
  INV_X1 U12950 ( .A(n14929), .ZN(n14907) );
  OR2_X1 U12951 ( .A1(n13201), .A2(n13200), .ZN(n13465) );
  AND2_X1 U12952 ( .A1(n10863), .A2(n10862), .ZN(n13269) );
  INV_X1 U12953 ( .A(n18892), .ZN(n18920) );
  INV_X1 U12954 ( .A(n13211), .ZN(n13021) );
  INV_X1 U12955 ( .A(n15369), .ZN(n18764) );
  OR2_X1 U12956 ( .A1(n15186), .A2(n10793), .ZN(n13542) );
  XNOR2_X1 U12957 ( .A(n11171), .B(n13317), .ZN(n13307) );
  AND2_X1 U12958 ( .A1(n11174), .A2(n11021), .ZN(n16150) );
  NOR2_X2 U12959 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19642) );
  INV_X1 U12960 ( .A(n19548), .ZN(n19052) );
  NOR2_X2 U12961 ( .A1(n19066), .A2(n19229), .ZN(n19112) );
  NAND2_X1 U12962 ( .A1(n13017), .A2(n13016), .ZN(n19392) );
  NOR2_X2 U12963 ( .A1(n19229), .A2(n19394), .ZN(n19216) );
  NOR2_X1 U12964 ( .A1(n19147), .A2(n19445), .ZN(n19220) );
  NOR2_X2 U12965 ( .A1(n19445), .A2(n19229), .ZN(n19279) );
  NOR2_X2 U12966 ( .A1(n19446), .A2(n19066), .ZN(n19297) );
  NOR2_X1 U12967 ( .A1(n19446), .A2(n19303), .ZN(n19307) );
  NOR2_X1 U12968 ( .A1(n19446), .A2(n19394), .ZN(n19380) );
  INV_X1 U12969 ( .A(n19515), .ZN(n19464) );
  INV_X1 U12970 ( .A(n19392), .ZN(n19496) );
  AND2_X1 U12971 ( .A1(n19043), .A2(n19049), .ZN(n19533) );
  INV_X1 U12972 ( .A(n19558), .ZN(n10754) );
  NOR2_X1 U12973 ( .A1(n19493), .A2(n13184), .ZN(n13014) );
  INV_X1 U12974 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19578) );
  NAND2_X1 U12975 ( .A1(n12179), .A2(n18598), .ZN(n11488) );
  NAND2_X1 U12976 ( .A1(n12181), .A2(n18444), .ZN(n16664) );
  OR4_X1 U12977 ( .A1(n18512), .A2(n16452), .A3(n18510), .A4(n18508), .ZN(
        n16432) );
  INV_X1 U12978 ( .A(n16672), .ZN(n16663) );
  NOR3_X1 U12979 ( .A1(n16664), .A2(n16507), .A3(n12182), .ZN(n16473) );
  INV_X1 U12980 ( .A(n16658), .ZN(n16603) );
  NOR2_X1 U12981 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16572), .ZN(n16553) );
  INV_X1 U12982 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16595) );
  INV_X1 U12983 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16616) );
  OAI211_X1 U12984 ( .C1(n18603), .C2(n18446), .A(n16632), .B(n18616), .ZN(
        n16674) );
  NOR2_X1 U12985 ( .A1(n16771), .A2(n16772), .ZN(n16744) );
  NOR2_X1 U12986 ( .A1(n16974), .A2(n16810), .ZN(n16797) );
  INV_X1 U12987 ( .A(n16995), .ZN(n16974) );
  NOR3_X1 U12988 ( .A1(n17991), .A2(n17076), .A3(n17196), .ZN(n17068) );
  NAND3_X1 U12989 ( .A1(n11261), .A2(n11260), .A3(n11259), .ZN(n12137) );
  NOR2_X1 U12990 ( .A1(n15418), .A2(n15417), .ZN(n15614) );
  INV_X1 U12991 ( .A(n17188), .ZN(n17177) );
  INV_X1 U12992 ( .A(n17424), .ZN(n17372) );
  NAND2_X1 U12993 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17446), .ZN(
        n17767) );
  INV_X1 U12994 ( .A(n17520), .ZN(n17498) );
  NOR2_X1 U12995 ( .A1(n9578), .A2(n16215), .ZN(n16216) );
  NOR2_X1 U12996 ( .A1(n17668), .A2(n17673), .ZN(n17299) );
  NAND2_X1 U12997 ( .A1(n17852), .A2(n9563), .ZN(n17900) );
  INV_X1 U12998 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17713) );
  NOR2_X1 U12999 ( .A1(n17435), .A2(n17755), .ZN(n17733) );
  NOR2_X1 U13000 ( .A1(n17821), .A2(n17807), .ZN(n17800) );
  NOR2_X1 U13001 ( .A1(n17812), .A2(n9563), .ZN(n17848) );
  INV_X1 U13002 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17874) );
  INV_X1 U13003 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17897) );
  INV_X1 U13004 ( .A(n17900), .ZN(n17936) );
  NOR3_X1 U13005 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n20687), .ZN(n18298) );
  NOR2_X1 U13006 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18543), .ZN(
        n18569) );
  INV_X1 U13007 ( .A(n18041), .ZN(n18059) );
  INV_X1 U13008 ( .A(n18084), .ZN(n18105) );
  INV_X1 U13009 ( .A(n18117), .ZN(n18151) );
  INV_X1 U13010 ( .A(n18143), .ZN(n18172) );
  INV_X1 U13011 ( .A(n18176), .ZN(n18195) );
  INV_X1 U13012 ( .A(n18199), .ZN(n18219) );
  INV_X1 U13013 ( .A(n18358), .ZN(n18280) );
  INV_X1 U13014 ( .A(n18346), .ZN(n18304) );
  AND2_X1 U13015 ( .A1(n18273), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18348) );
  INV_X1 U13016 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18478) );
  INV_X1 U13017 ( .A(U212), .ZN(n16257) );
  INV_X1 U13018 ( .A(n20664), .ZN(n12934) );
  INV_X1 U13019 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20055) );
  OR3_X1 U13020 ( .A1(n12934), .A2(n12933), .A3(n12932), .ZN(n19761) );
  INV_X1 U13021 ( .A(n19755), .ZN(n15657) );
  INV_X1 U13022 ( .A(n15745), .ZN(n14577) );
  INV_X1 U13023 ( .A(n19802), .ZN(n19822) );
  OAI21_X1 U13024 ( .B1(n14416), .B2(n14415), .A(n14491), .ZN(n14682) );
  INV_X1 U13025 ( .A(n19916), .ZN(n19912) );
  INV_X1 U13026 ( .A(n19917), .ZN(n19708) );
  NAND2_X1 U13027 ( .A1(n20100), .A2(n9660), .ZN(n20041) );
  NAND2_X1 U13028 ( .A1(n20100), .A2(n20426), .ZN(n20084) );
  NAND2_X1 U13029 ( .A1(n20100), .A2(n20231), .ZN(n20137) );
  NAND2_X1 U13030 ( .A1(n20232), .A2(n9660), .ZN(n20186) );
  NAND2_X1 U13031 ( .A1(n20232), .A2(n20426), .ZN(n20218) );
  NAND2_X1 U13032 ( .A1(n20232), .A2(n20474), .ZN(n20243) );
  NAND2_X1 U13033 ( .A1(n20283), .A2(n9660), .ZN(n20307) );
  OR2_X1 U13034 ( .A1(n20356), .A2(n20287), .ZN(n20342) );
  OR2_X1 U13035 ( .A1(n20356), .A2(n20308), .ZN(n20378) );
  OR2_X1 U13036 ( .A1(n20356), .A2(n20355), .ZN(n20425) );
  NAND2_X1 U13037 ( .A1(n20475), .A2(n20426), .ZN(n20502) );
  NAND2_X1 U13038 ( .A1(n20475), .A2(n20474), .ZN(n20568) );
  NOR2_X1 U13039 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20670) );
  NAND2_X1 U13040 ( .A1(n20590), .A2(n20675), .ZN(n20649) );
  INV_X1 U13041 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20595) );
  NAND2_X1 U13042 ( .A1(n20663), .A2(n20592), .ZN(n20639) );
  OR2_X1 U13043 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n19698), .ZN(n20675) );
  AND2_X1 U13044 ( .A1(n12681), .A2(n12223), .ZN(n18623) );
  NAND2_X1 U13045 ( .A1(n12267), .A2(n12266), .ZN(n12324) );
  INV_X1 U13046 ( .A(n18838), .ZN(n18742) );
  INV_X1 U13047 ( .A(n18855), .ZN(n18842) );
  INV_X1 U13048 ( .A(n18854), .ZN(n18822) );
  INV_X1 U13049 ( .A(n19636), .ZN(n13034) );
  AND2_X1 U13050 ( .A1(n18869), .A2(n18868), .ZN(n18890) );
  INV_X1 U13051 ( .A(n18874), .ZN(n18927) );
  OR2_X1 U13052 ( .A1(n18968), .A2(n12367), .ZN(n18930) );
  NAND2_X1 U13053 ( .A1(n12366), .A2(n19688), .ZN(n18968) );
  INV_X1 U13054 ( .A(n18973), .ZN(n12430) );
  INV_X1 U13055 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16035) );
  INV_X1 U13056 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16056) );
  INV_X1 U13057 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18743) );
  INV_X1 U13058 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16106) );
  INV_X1 U13059 ( .A(n12340), .ZN(n12349) );
  INV_X1 U13060 ( .A(n16154), .ZN(n18994) );
  INV_X1 U13061 ( .A(n18999), .ZN(n16152) );
  INV_X1 U13062 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19666) );
  NAND2_X1 U13063 ( .A1(n19064), .A2(n19087), .ZN(n19086) );
  INV_X1 U13064 ( .A(n19142), .ZN(n19116) );
  INV_X1 U13065 ( .A(n19197), .ZN(n19175) );
  AOI21_X1 U13066 ( .B1(n19177), .B2(n19180), .A(n19176), .ZN(n19201) );
  AOI211_X2 U13067 ( .C1(n13020), .C2(n13019), .A(n19496), .B(n13018), .ZN(
        n19219) );
  INV_X1 U13068 ( .A(n19220), .ZN(n19248) );
  AOI211_X2 U13069 ( .C1(n19253), .C2(n19254), .A(n19496), .B(n19252), .ZN(
        n19284) );
  AOI211_X2 U13070 ( .C1(n13039), .C2(n13044), .A(n19496), .B(n13038), .ZN(
        n19302) );
  INV_X1 U13071 ( .A(n19307), .ZN(n19361) );
  AOI211_X2 U13072 ( .C1(n13130), .C2(n13129), .A(n19496), .B(n13128), .ZN(
        n19379) );
  INV_X1 U13073 ( .A(n19380), .ZN(n19443) );
  AOI211_X2 U13074 ( .C1(n19454), .C2(n19456), .A(n19496), .B(n19452), .ZN(
        n19488) );
  NAND2_X1 U13075 ( .A1(n19017), .A2(n19500), .ZN(n19548) );
  NAND2_X1 U13076 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10754), .ZN(n16174) );
  INV_X1 U13077 ( .A(n19631), .ZN(n19559) );
  NAND2_X1 U13078 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19560), .ZN(n19695) );
  NOR2_X1 U13079 ( .A1(n18431), .A2(n17151), .ZN(n18620) );
  INV_X1 U13080 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n20687) );
  INV_X1 U13081 ( .A(n16473), .ZN(n16500) );
  INV_X1 U13082 ( .A(n16673), .ZN(n16638) );
  NAND2_X1 U13083 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16674), .ZN(n16658) );
  NOR2_X1 U13084 ( .A1(n16678), .A2(n16738), .ZN(n16743) );
  INV_X1 U13085 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16966) );
  NOR2_X1 U13086 ( .A1(n20684), .A2(n16971), .ZN(n16970) );
  INV_X1 U13087 ( .A(n17074), .ZN(n17049) );
  NOR3_X1 U13088 ( .A1(n17111), .A2(n17240), .A3(n17142), .ZN(n17114) );
  NOR2_X1 U13089 ( .A1(n11204), .A2(n11203), .ZN(n17128) );
  NAND2_X1 U13090 ( .A1(n17177), .A2(n17960), .ZN(n17168) );
  OR2_X1 U13091 ( .A1(n18553), .A2(n17624), .ZN(n17179) );
  INV_X1 U13092 ( .A(n17234), .ZN(n17238) );
  INV_X1 U13093 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17492) );
  NAND2_X1 U13094 ( .A1(n18247), .A2(n18298), .ZN(n17995) );
  OAI21_X1 U13095 ( .B1(n16218), .B2(n16217), .A(n16216), .ZN(n16219) );
  INV_X1 U13096 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18404) );
  INV_X1 U13097 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18425) );
  INV_X2 U13098 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18551) );
  INV_X1 U13099 ( .A(n18321), .ZN(n18318) );
  INV_X1 U13100 ( .A(n18341), .ZN(n18386) );
  INV_X1 U13101 ( .A(n18541), .ZN(n18459) );
  INV_X1 U13102 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18487) );
  NOR2_X1 U13103 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12167), .ZN(n16300)
         );
  INV_X1 U13104 ( .A(n16268), .ZN(n16259) );
  INV_X1 U13105 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19581) );
  OR4_X1 U13106 ( .A1(n12244), .A2(n12243), .A3(n12242), .A4(n12241), .ZN(
        P2_U2834) );
  OR4_X1 U13107 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        P3_U2651) );
  NAND2_X1 U13108 ( .A1(n11517), .A2(n11516), .ZN(P3_U2831) );
  INV_X1 U13109 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10102) );
  AND2_X2 U13110 ( .A1(n10102), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10336) );
  AND2_X4 U13111 ( .A1(n10336), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14278) );
  AOI22_X1 U13112 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10108) );
  AND2_X2 U13113 ( .A1(n10103), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12657) );
  AND2_X4 U13114 ( .A1(n12657), .A2(n12581), .ZN(n14091) );
  NAND2_X1 U13115 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10104) );
  NOR2_X2 U13116 ( .A1(n10104), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10128) );
  AOI22_X1 U13117 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10107) );
  AND2_X4 U13118 ( .A1(n12650), .A2(n10493), .ZN(n10329) );
  NOR2_X2 U13119 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10334) );
  AND2_X4 U13120 ( .A1(n10334), .A2(n12581), .ZN(n14282) );
  AOI22_X1 U13121 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U13122 ( .A1(n9568), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10105) );
  NAND4_X1 U13123 ( .A1(n10108), .A2(n10107), .A3(n10106), .A4(n10105), .ZN(
        n10109) );
  AOI22_X1 U13124 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10113) );
  AOI22_X1 U13125 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U13126 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10111) );
  NAND4_X1 U13127 ( .A1(n10113), .A2(n10112), .A3(n10111), .A4(n10110), .ZN(
        n10114) );
  AOI22_X1 U13128 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U13129 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U13130 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U13131 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10115) );
  NAND4_X1 U13132 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10119) );
  AOI22_X1 U13133 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U13134 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10121) );
  NAND4_X1 U13135 ( .A1(n10123), .A2(n10122), .A3(n10121), .A4(n10120), .ZN(
        n10124) );
  NAND2_X1 U13136 ( .A1(n10124), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10125) );
  AOI22_X1 U13137 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10132) );
  INV_X2 U13138 ( .A(n12645), .ZN(n14214) );
  AOI22_X1 U13139 ( .A1(n9568), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U13140 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U13141 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10128), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10129) );
  NAND4_X1 U13142 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .ZN(
        n10133) );
  NAND2_X1 U13143 ( .A1(n10133), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10140) );
  AOI22_X1 U13144 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U13145 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U13146 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U13147 ( .A1(n9568), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10134) );
  NAND4_X1 U13148 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10138) );
  NAND2_X1 U13149 ( .A1(n10138), .A2(n10141), .ZN(n10139) );
  AOI22_X1 U13150 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10144) );
  AOI22_X1 U13151 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U13152 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10142) );
  NAND4_X1 U13153 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10151) );
  AOI22_X1 U13154 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U13155 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U13156 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10146) );
  NAND4_X1 U13157 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10150) );
  AOI22_X1 U13158 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U13159 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13160 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U13161 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U13162 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13163 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U13164 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U13165 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14214), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U13166 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U13167 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13168 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13169 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U13170 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10164) );
  INV_X1 U13171 ( .A(n10718), .ZN(n10188) );
  INV_X1 U13172 ( .A(n10212), .ZN(n10169) );
  NAND2_X1 U13173 ( .A1(n10170), .A2(n10169), .ZN(n10739) );
  NAND2_X1 U13174 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10172) );
  AOI22_X1 U13175 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10329), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13176 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10174) );
  NAND4_X1 U13177 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  NAND2_X1 U13178 ( .A1(n10177), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10186) );
  NAND2_X1 U13179 ( .A1(n14278), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10178) );
  AOI22_X1 U13180 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13181 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10180) );
  NAND4_X1 U13182 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n10184) );
  NAND3_X1 U13183 ( .A1(n10739), .A2(n10712), .A3(n10219), .ZN(n10187) );
  AOI22_X1 U13184 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U13185 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13186 ( .A1(n10329), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13187 ( .A1(n14214), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10189) );
  NAND4_X1 U13188 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10193) );
  AOI22_X1 U13189 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U13190 ( .A1(n14091), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10329), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13191 ( .A1(n9568), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14104), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U13192 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14282), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10194) );
  NAND4_X1 U13193 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10198) );
  NAND2_X1 U13194 ( .A1(n10217), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12367) );
  NAND2_X1 U13195 ( .A1(n11018), .A2(n19690), .ZN(n10211) );
  NAND4_X1 U13196 ( .A1(n10127), .A2(n10222), .A3(n10705), .A4(n12991), .ZN(
        n10238) );
  NAND2_X1 U13197 ( .A1(n10766), .A2(n10238), .ZN(n10257) );
  NAND2_X1 U13198 ( .A1(n10257), .A2(n12691), .ZN(n10208) );
  NAND4_X1 U13199 ( .A1(n10705), .A2(n10221), .A3(n10214), .A4(n10704), .ZN(
        n10200) );
  INV_X1 U13200 ( .A(n10218), .ZN(n10207) );
  MUX2_X1 U13201 ( .A(n10222), .B(n10214), .S(n10201), .Z(n10205) );
  AND2_X1 U13202 ( .A1(n10212), .A2(n10712), .ZN(n10204) );
  NAND2_X1 U13203 ( .A1(n10229), .A2(n10759), .ZN(n10203) );
  NAND3_X1 U13204 ( .A1(n10205), .A2(n10204), .A3(n10203), .ZN(n10206) );
  NAND3_X1 U13205 ( .A1(n10207), .A2(n10206), .A3(n12691), .ZN(n10771) );
  NAND2_X1 U13206 ( .A1(n10208), .A2(n10771), .ZN(n10209) );
  NAND2_X1 U13207 ( .A1(n10209), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U13208 ( .A1(n10213), .A2(n10212), .ZN(n10716) );
  NAND2_X1 U13209 ( .A1(n10229), .A2(n13054), .ZN(n10708) );
  OAI211_X1 U13210 ( .C1(n10716), .C2(n13054), .A(n10708), .B(n19050), .ZN(
        n10757) );
  NAND2_X1 U13211 ( .A1(n10757), .A2(n10759), .ZN(n10216) );
  NAND2_X1 U13212 ( .A1(n10216), .A2(n10215), .ZN(n10256) );
  INV_X1 U13213 ( .A(n11017), .ZN(n10224) );
  NAND4_X1 U13214 ( .A1(n10803), .A2(n12691), .A3(n10767), .A4(n19043), .ZN(
        n10223) );
  NAND2_X2 U13215 ( .A1(n10224), .A2(n10223), .ZN(n11133) );
  AOI22_X1 U13216 ( .A1(n11133), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12706), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U13217 ( .A1(n10228), .A2(n19043), .ZN(n10230) );
  INV_X1 U13218 ( .A(n10229), .ZN(n10811) );
  NAND2_X2 U13219 ( .A1(n10232), .A2(n10231), .ZN(n11019) );
  NOR2_X1 U13220 ( .A1(n10219), .A2(n12317), .ZN(n10233) );
  NAND4_X1 U13221 ( .A1(n10803), .A2(n12691), .A3(n10767), .A4(n12341), .ZN(
        n10234) );
  INV_X1 U13222 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12421) );
  NAND2_X1 U13223 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10239) );
  INV_X1 U13224 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10240) );
  INV_X1 U13225 ( .A(n10242), .ZN(n10243) );
  NOR2_X1 U13226 ( .A1(n10243), .A2(n10237), .ZN(n10244) );
  AOI22_X1 U13227 ( .A1(n12585), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12706), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U13228 ( .A1(n10247), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10252) );
  INV_X1 U13229 ( .A(n12706), .ZN(n10251) );
  NAND2_X1 U13230 ( .A1(n10248), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U13231 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10249) );
  NAND4_X1 U13232 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .ZN(
        n10255) );
  INV_X1 U13233 ( .A(n10253), .ZN(n10254) );
  NAND2_X1 U13234 ( .A1(n10256), .A2(n10094), .ZN(n10258) );
  NAND2_X1 U13235 ( .A1(n10274), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10263) );
  NAND2_X1 U13236 ( .A1(n12706), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10262) );
  NAND2_X1 U13237 ( .A1(n10263), .A2(n10262), .ZN(n11039) );
  NAND2_X1 U13238 ( .A1(n11022), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10267) );
  INV_X1 U13239 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12737) );
  OAI21_X1 U13240 ( .B1(n11130), .B2(n12737), .A(n10264), .ZN(n10265) );
  INV_X1 U13241 ( .A(n10265), .ZN(n10266) );
  INV_X1 U13242 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10469) );
  INV_X1 U13243 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U13244 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10270) );
  OAI211_X1 U13245 ( .C1(n10268), .C2(n10469), .A(n9641), .B(n10270), .ZN(
        n10271) );
  INV_X1 U13246 ( .A(n10271), .ZN(n10273) );
  NAND2_X1 U13247 ( .A1(n11022), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10272) );
  NAND2_X1 U13248 ( .A1(n10274), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10276) );
  AOI21_X1 U13249 ( .B1(n12317), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U13250 ( .A1(n10281), .A2(n10278), .ZN(n10285) );
  NAND2_X1 U13251 ( .A1(n11033), .A2(n10291), .ZN(n10280) );
  NAND2_X1 U13252 ( .A1(n10279), .A2(n10278), .ZN(n10283) );
  INV_X1 U13253 ( .A(n10286), .ZN(n10289) );
  INV_X1 U13254 ( .A(n10287), .ZN(n10288) );
  NAND2_X1 U13255 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  INV_X2 U13256 ( .A(n12456), .ZN(n10318) );
  INV_X1 U13257 ( .A(n10411), .ZN(n13132) );
  AOI22_X1 U13258 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10524), .B1(
        n13132), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10328) );
  INV_X1 U13259 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10299) );
  NAND2_X1 U13260 ( .A1(n12340), .A2(n10297), .ZN(n10314) );
  INV_X1 U13261 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10298) );
  INV_X1 U13262 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10300) );
  INV_X1 U13263 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14133) );
  NOR2_X1 U13264 ( .A1(n10302), .A2(n10301), .ZN(n10327) );
  INV_X1 U13265 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10307) );
  INV_X1 U13266 ( .A(n10297), .ZN(n10304) );
  NAND2_X1 U13267 ( .A1(n12340), .A2(n10304), .ZN(n10316) );
  INV_X1 U13268 ( .A(n10316), .ZN(n10305) );
  INV_X1 U13269 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10306) );
  OAI22_X1 U13270 ( .A1(n10307), .A2(n10514), .B1(n10516), .B2(n10306), .ZN(
        n10312) );
  INV_X1 U13271 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10310) );
  INV_X1 U13272 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10309) );
  NOR2_X1 U13273 ( .A1(n10312), .A2(n10311), .ZN(n10326) );
  NOR2_X2 U13274 ( .A1(n10320), .A2(n10313), .ZN(n10407) );
  NOR2_X2 U13275 ( .A1(n10315), .A2(n19005), .ZN(n10415) );
  AOI22_X1 U13276 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10415), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10324) );
  NOR2_X2 U13277 ( .A1(n10315), .A2(n10318), .ZN(n19491) );
  NOR2_X1 U13278 ( .A1(n10317), .A2(n19005), .ZN(n10416) );
  AOI22_X1 U13279 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19491), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10323) );
  NOR2_X2 U13280 ( .A1(n10317), .A2(n10318), .ZN(n19382) );
  AOI21_X1 U13281 ( .B1(n19382), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n19683), .ZN(n10322) );
  NAND2_X1 U13282 ( .A1(n10318), .A2(n9598), .ZN(n10319) );
  NAND2_X1 U13283 ( .A1(n19308), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10321) );
  AND4_X1 U13284 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10325) );
  AOI22_X1 U13285 ( .A1(n10344), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13286 ( .A1(n10432), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13287 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10331) );
  AND2_X2 U13288 ( .A1(n14295), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10400) );
  AOI22_X1 U13289 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10330) );
  NAND4_X1 U13290 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10343) );
  AOI22_X1 U13291 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13292 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10340) );
  AND2_X2 U13293 ( .A1(n12657), .A2(n14093), .ZN(n14123) );
  NAND3_X1 U13294 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10743) );
  INV_X1 U13295 ( .A(n10743), .ZN(n10335) );
  AOI22_X1 U13296 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14122), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10339) );
  AND2_X1 U13297 ( .A1(n14093), .A2(n10337), .ZN(n10350) );
  AOI22_X1 U13298 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10338) );
  NAND4_X1 U13299 ( .A1(n10341), .A2(n10340), .A3(n10339), .A4(n10338), .ZN(
        n10342) );
  AND2_X1 U13300 ( .A1(n19683), .A2(n10492), .ZN(n12320) );
  AOI22_X1 U13301 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13302 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10384), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13303 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13304 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10345) );
  NAND4_X1 U13305 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10356) );
  AOI22_X1 U13306 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10437), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13307 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n10350), .ZN(n10353) );
  AOI22_X1 U13308 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n14122), .ZN(n10352) );
  AOI22_X1 U13309 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14123), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10351) );
  NAND4_X1 U13310 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10355) );
  AND2_X1 U13311 ( .A1(n12320), .A2(n11141), .ZN(n11146) );
  AOI22_X1 U13312 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14114), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13313 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10344), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13314 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14120), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13315 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10357) );
  NAND4_X1 U13316 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10367) );
  AOI22_X1 U13317 ( .A1(n10437), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13318 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n14121), .ZN(n10364) );
  AOI22_X1 U13319 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n14122), .ZN(n10363) );
  AOI22_X1 U13320 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10362) );
  NAND4_X1 U13321 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10366) );
  OR2_X1 U13322 ( .A1(n11146), .A2(n10824), .ZN(n10368) );
  INV_X1 U13323 ( .A(n10418), .ZN(n19222) );
  AOI22_X1 U13324 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19222), .B1(
        n19149), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10373) );
  INV_X1 U13325 ( .A(n10417), .ZN(n10369) );
  NAND2_X1 U13326 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10372) );
  AOI22_X1 U13327 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19382), .B1(
        n10415), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13328 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19491), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10370) );
  INV_X1 U13329 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14191) );
  NAND2_X1 U13330 ( .A1(n19308), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10375) );
  NAND2_X1 U13331 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10374) );
  OAI211_X1 U13332 ( .C1(n10411), .C2(n14191), .A(n10375), .B(n10374), .ZN(
        n10376) );
  INV_X1 U13333 ( .A(n10376), .ZN(n10382) );
  INV_X1 U13334 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12539) );
  INV_X1 U13335 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10377) );
  OAI22_X1 U13336 ( .A1(n12539), .A2(n10514), .B1(n10516), .B2(n10377), .ZN(
        n10379) );
  INV_X1 U13337 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13419) );
  INV_X1 U13338 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14185) );
  OAI22_X1 U13339 ( .A1(n13419), .A2(n10426), .B1(n10412), .B2(n14185), .ZN(
        n10378) );
  NOR2_X1 U13340 ( .A1(n10379), .A2(n10378), .ZN(n10381) );
  INV_X1 U13341 ( .A(n10423), .ZN(n19088) );
  AOI22_X1 U13342 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10344), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13343 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10864), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13344 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13345 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10385) );
  NAND4_X1 U13346 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10394) );
  AOI22_X1 U13347 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14120), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U13348 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14121), .ZN(n10391) );
  AOI22_X1 U13349 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n14122), .ZN(n10390) );
  AOI22_X1 U13350 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10389) );
  NAND4_X1 U13351 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10393) );
  NOR2_X1 U13352 ( .A1(n10394), .A2(n10393), .ZN(n10838) );
  NAND2_X1 U13353 ( .A1(n10838), .A2(n19683), .ZN(n10395) );
  AOI22_X1 U13354 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14114), .B1(
        n10344), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13355 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10864), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13356 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10384), .B1(
        n14120), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13357 ( .A1(n10437), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10396) );
  NAND4_X1 U13358 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10406) );
  AOI22_X1 U13359 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U13360 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n14121), .ZN(n10403) );
  AOI22_X1 U13361 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n14122), .ZN(n10402) );
  AOI22_X1 U13362 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10401) );
  NAND4_X1 U13363 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10405) );
  INV_X1 U13364 ( .A(n10480), .ZN(n11152) );
  INV_X1 U13365 ( .A(n10524), .ZN(n10410) );
  INV_X1 U13366 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U13367 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10409) );
  NAND2_X1 U13368 ( .A1(n19308), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10408) );
  OAI211_X1 U13369 ( .C1(n10410), .C2(n14245), .A(n10409), .B(n10408), .ZN(
        n10414) );
  INV_X1 U13370 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14243) );
  INV_X1 U13371 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14237) );
  OAI22_X1 U13372 ( .A1(n10411), .A2(n14243), .B1(n14237), .B2(n10412), .ZN(
        n10413) );
  NOR2_X1 U13373 ( .A1(n10414), .A2(n10413), .ZN(n10431) );
  AOI22_X1 U13374 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19382), .B1(
        n19491), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U13376 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n10415), .B1(
        n13042), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10421) );
  INV_X1 U13377 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10419) );
  NAND2_X1 U13378 ( .A1(n19022), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10420) );
  INV_X1 U13379 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10425) );
  INV_X1 U13380 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10424) );
  OAI22_X1 U13381 ( .A1(n10425), .A2(n10516), .B1(n10423), .B2(n10424), .ZN(
        n10429) );
  INV_X1 U13382 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10427) );
  INV_X1 U13383 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14235) );
  OAI22_X1 U13384 ( .A1(n10427), .A2(n10426), .B1(n10526), .B2(n14235), .ZN(
        n10428) );
  NOR2_X1 U13385 ( .A1(n10429), .A2(n10428), .ZN(n10430) );
  AOI22_X1 U13386 ( .A1(n10344), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13387 ( .A1(n10432), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13388 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13389 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10433) );
  NAND4_X1 U13390 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n10443) );
  AOI22_X1 U13391 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13392 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13393 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14122), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13394 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10438) );
  NAND4_X1 U13395 ( .A1(n10441), .A2(n10440), .A3(n10439), .A4(n10438), .ZN(
        n10442) );
  INV_X1 U13396 ( .A(n10481), .ZN(n10848) );
  NAND2_X1 U13397 ( .A1(n10848), .A2(n19683), .ZN(n10444) );
  NAND2_X1 U13398 ( .A1(n10344), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10451) );
  NAND2_X1 U13399 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10450) );
  NAND2_X1 U13400 ( .A1(n10432), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10449) );
  NAND2_X1 U13401 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10448) );
  AOI22_X1 U13402 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14120), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U13403 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10455) );
  NAND2_X1 U13404 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10454) );
  NAND2_X1 U13405 ( .A1(n14115), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10453) );
  NAND2_X1 U13406 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10452) );
  AOI22_X1 U13407 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10459) );
  NAND2_X1 U13408 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10458) );
  AOI22_X1 U13409 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n14122), .ZN(n10457) );
  NAND2_X1 U13410 ( .A1(n14121), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10456) );
  MUX2_X1 U13411 ( .A(n10817), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10678) );
  NAND2_X1 U13412 ( .A1(n10678), .A2(n10679), .ZN(n10465) );
  NAND2_X1 U13413 ( .A1(n10817), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13414 ( .A1(n10465), .A2(n10464), .ZN(n10472) );
  XNOR2_X1 U13415 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10471) );
  INV_X1 U13416 ( .A(n10471), .ZN(n10466) );
  XNOR2_X1 U13417 ( .A(n10472), .B(n10466), .ZN(n10719) );
  MUX2_X1 U13418 ( .A(n10824), .B(n10719), .S(n9567), .Z(n10729) );
  MUX2_X1 U13419 ( .A(n10729), .B(n10469), .S(n13985), .Z(n10491) );
  NOR2_X1 U13420 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10470) );
  MUX2_X1 U13421 ( .A(n10470), .B(n11141), .S(n10468), .Z(n10490) );
  NAND2_X1 U13422 ( .A1(n10491), .A2(n10490), .ZN(n10487) );
  NAND2_X1 U13423 ( .A1(n10472), .A2(n10471), .ZN(n10474) );
  NAND2_X1 U13424 ( .A1(n19651), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10473) );
  MUX2_X1 U13425 ( .A(n12670), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10477) );
  INV_X1 U13426 ( .A(n10477), .ZN(n10475) );
  INV_X1 U13427 ( .A(n10720), .ZN(n10691) );
  MUX2_X1 U13428 ( .A(n10838), .B(n10691), .S(n9567), .Z(n10733) );
  NOR2_X4 U13429 ( .A1(n10487), .A2(n10486), .ZN(n10507) );
  NOR2_X1 U13430 ( .A1(n10141), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10476) );
  INV_X1 U13431 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15610) );
  NOR2_X1 U13432 ( .A1(n15610), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10479) );
  NAND2_X1 U13433 ( .A1(n10694), .A2(n10479), .ZN(n10721) );
  MUX2_X1 U13434 ( .A(n10480), .B(n10721), .S(n9567), .Z(n10734) );
  INV_X1 U13435 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18825) );
  MUX2_X1 U13436 ( .A(n10734), .B(n18825), .S(n13985), .Z(n10506) );
  INV_X1 U13437 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11050) );
  MUX2_X1 U13438 ( .A(n11050), .B(n10481), .S(n10468), .Z(n10482) );
  OAI21_X1 U13439 ( .B1(n9665), .B2(n10482), .A(n10554), .ZN(n18811) );
  INV_X1 U13440 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11159) );
  INV_X1 U13441 ( .A(n10507), .ZN(n10489) );
  NAND2_X1 U13442 ( .A1(n10487), .A2(n10486), .ZN(n10488) );
  NAND2_X1 U13443 ( .A1(n10489), .A2(n10488), .ZN(n12759) );
  OAI21_X2 U13444 ( .B1(n11140), .B2(n10858), .A(n12759), .ZN(n10502) );
  NAND2_X1 U13445 ( .A1(n10502), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12723) );
  INV_X1 U13446 ( .A(n10490), .ZN(n10498) );
  XNOR2_X1 U13447 ( .A(n10491), .B(n10498), .ZN(n13076) );
  INV_X1 U13448 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19007) );
  XNOR2_X1 U13449 ( .A(n13076), .B(n19007), .ZN(n13971) );
  INV_X1 U13450 ( .A(n10492), .ZN(n11142) );
  AND2_X1 U13451 ( .A1(n10493), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10494) );
  NOR2_X1 U13452 ( .A1(n10679), .A2(n10494), .ZN(n10682) );
  INV_X1 U13453 ( .A(n10682), .ZN(n10741) );
  MUX2_X1 U13454 ( .A(n11142), .B(n10741), .S(n9567), .Z(n10732) );
  INV_X1 U13455 ( .A(n10732), .ZN(n10495) );
  MUX2_X1 U13456 ( .A(n10495), .B(P2_EBX_REG_0__SCAN_IN), .S(n13985), .Z(
        n18851) );
  NAND2_X1 U13457 ( .A1(n18851), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12331) );
  AND2_X1 U13458 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10496) );
  NAND2_X1 U13459 ( .A1(n13985), .A2(n10496), .ZN(n10497) );
  NAND2_X1 U13460 ( .A1(n10498), .A2(n10497), .ZN(n12329) );
  INV_X1 U13461 ( .A(n12329), .ZN(n18839) );
  NAND2_X1 U13462 ( .A1(n18839), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10500) );
  INV_X1 U13463 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13182) );
  AND2_X1 U13464 ( .A1(n12329), .A2(n13182), .ZN(n10499) );
  AOI21_X1 U13465 ( .B1(n12331), .B2(n10500), .A(n10499), .ZN(n13970) );
  NAND2_X1 U13466 ( .A1(n13971), .A2(n13970), .ZN(n13969) );
  NAND2_X1 U13467 ( .A1(n13076), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10501) );
  AND2_X1 U13468 ( .A1(n13969), .A2(n10501), .ZN(n12725) );
  NAND2_X1 U13469 ( .A1(n12723), .A2(n12725), .ZN(n10505) );
  INV_X1 U13470 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10503) );
  XNOR2_X1 U13471 ( .A(n10507), .B(n9836), .ZN(n18823) );
  XNOR2_X1 U13472 ( .A(n18823), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12834) );
  INV_X1 U13473 ( .A(n18823), .ZN(n10508) );
  INV_X1 U13474 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12844) );
  NAND2_X1 U13475 ( .A1(n16108), .A2(n16109), .ZN(n10511) );
  NAND2_X1 U13476 ( .A1(n10509), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10510) );
  NAND2_X1 U13477 ( .A1(n10511), .A2(n10510), .ZN(n13163) );
  INV_X1 U13478 ( .A(n10550), .ZN(n10549) );
  AOI22_X1 U13479 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19382), .B1(
        n13042), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13480 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19491), .B1(
        n10415), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10519) );
  INV_X1 U13481 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10513) );
  INV_X1 U13482 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10512) );
  OAI22_X1 U13483 ( .A1(n10514), .A2(n10513), .B1(n10412), .B2(n10512), .ZN(
        n10515) );
  INV_X1 U13484 ( .A(n10515), .ZN(n10518) );
  NAND2_X1 U13485 ( .A1(n19058), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10517) );
  INV_X1 U13486 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14266) );
  NAND2_X1 U13487 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10522) );
  NAND2_X1 U13488 ( .A1(n19308), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10521) );
  OAI211_X1 U13489 ( .C1(n10411), .C2(n14266), .A(n10522), .B(n10521), .ZN(
        n10523) );
  INV_X1 U13490 ( .A(n10523), .ZN(n10534) );
  INV_X1 U13491 ( .A(n10426), .ZN(n10525) );
  AOI22_X1 U13492 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n10525), .ZN(n10533) );
  INV_X1 U13493 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10527) );
  INV_X1 U13494 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14256) );
  OAI22_X1 U13495 ( .A1(n19123), .A2(n10527), .B1(n10526), .B2(n14256), .ZN(
        n10531) );
  INV_X1 U13496 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10529) );
  INV_X1 U13497 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10528) );
  OAI22_X1 U13498 ( .A1(n10423), .A2(n10529), .B1(n10418), .B2(n10528), .ZN(
        n10530) );
  NOR2_X1 U13499 ( .A1(n10531), .A2(n10530), .ZN(n10532) );
  NAND4_X1 U13500 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10547) );
  AOI22_X1 U13501 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13502 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10384), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13503 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13504 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10536) );
  NAND4_X1 U13505 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10545) );
  AOI22_X1 U13506 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10437), .B1(
        n14120), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13507 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n14121), .ZN(n10542) );
  AOI22_X1 U13508 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n14122), .ZN(n10541) );
  AOI22_X1 U13509 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10540) );
  NAND4_X1 U13510 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10544) );
  NAND2_X1 U13511 ( .A1(n10552), .A2(n19683), .ZN(n10546) );
  NAND2_X1 U13512 ( .A1(n10550), .A2(n11161), .ZN(n10551) );
  MUX2_X1 U13513 ( .A(n10552), .B(P2_EBX_REG_6__SCAN_IN), .S(n13985), .Z(
        n10553) );
  AND2_X1 U13514 ( .A1(n10554), .A2(n10553), .ZN(n10555) );
  OR2_X1 U13515 ( .A1(n10555), .A2(n9604), .ZN(n18802) );
  INV_X1 U13516 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13166) );
  XNOR2_X1 U13517 ( .A(n10556), .B(n13166), .ZN(n13162) );
  NAND2_X1 U13518 ( .A1(n13163), .A2(n13162), .ZN(n10558) );
  NAND2_X1 U13519 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10557) );
  INV_X1 U13520 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11057) );
  MUX2_X1 U13521 ( .A(n11057), .B(n10858), .S(n10468), .Z(n10560) );
  NAND2_X1 U13522 ( .A1(n13985), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10559) );
  XNOR2_X1 U13523 ( .A(n10564), .B(n10559), .ZN(n18777) );
  AND2_X1 U13524 ( .A1(n10858), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11172) );
  NAND2_X1 U13525 ( .A1(n18777), .A2(n11172), .ZN(n13312) );
  INV_X1 U13526 ( .A(n10560), .ZN(n10561) );
  XNOR2_X1 U13527 ( .A(n9604), .B(n10561), .ZN(n18790) );
  NAND2_X1 U13528 ( .A1(n18790), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13310) );
  NAND2_X1 U13529 ( .A1(n18777), .A2(n10858), .ZN(n10562) );
  INV_X1 U13530 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13317) );
  NAND2_X1 U13531 ( .A1(n10562), .A2(n13317), .ZN(n13313) );
  OR2_X1 U13532 ( .A1(n18790), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13309) );
  AND2_X1 U13533 ( .A1(n13313), .A2(n13309), .ZN(n10563) );
  OR2_X2 U13534 ( .A1(n10564), .A2(n13985), .ZN(n10659) );
  INV_X1 U13535 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11066) );
  NOR2_X1 U13536 ( .A1(n10468), .A2(n11066), .ZN(n10566) );
  XNOR2_X1 U13537 ( .A(n10567), .B(n10566), .ZN(n18767) );
  NAND2_X1 U13538 ( .A1(n18767), .A2(n10858), .ZN(n10576) );
  INV_X1 U13539 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15380) );
  AND2_X1 U13540 ( .A1(n10576), .A2(n15380), .ZN(n15392) );
  NAND2_X1 U13541 ( .A1(n13985), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10568) );
  MUX2_X1 U13542 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n10568), .S(n10570), .Z(
        n10569) );
  AND2_X1 U13543 ( .A1(n10569), .A2(n10659), .ZN(n18757) );
  NAND2_X1 U13544 ( .A1(n18757), .A2(n10858), .ZN(n10577) );
  INV_X1 U13545 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15368) );
  NAND2_X1 U13546 ( .A1(n10577), .A2(n15368), .ZN(n15362) );
  NAND2_X1 U13547 ( .A1(n13985), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10571) );
  OR2_X1 U13548 ( .A1(n10572), .A2(n10571), .ZN(n10574) );
  INV_X1 U13549 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18744) );
  NAND2_X1 U13550 ( .A1(n10659), .A2(n10579), .ZN(n10578) );
  INV_X1 U13551 ( .A(n10578), .ZN(n10573) );
  NAND2_X1 U13552 ( .A1(n10574), .A2(n10573), .ZN(n18747) );
  OR2_X1 U13553 ( .A1(n18747), .A2(n9804), .ZN(n10575) );
  INV_X1 U13554 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11075) );
  OR2_X1 U13555 ( .A1(n10575), .A2(n11075), .ZN(n16075) );
  NOR2_X1 U13556 ( .A1(n10576), .A2(n15380), .ZN(n15391) );
  NOR2_X1 U13557 ( .A1(n15368), .A2(n10577), .ZN(n15360) );
  NOR2_X1 U13558 ( .A1(n15391), .A2(n15360), .ZN(n16073) );
  AND2_X1 U13559 ( .A1(n16075), .A2(n16073), .ZN(n15051) );
  NAND2_X1 U13560 ( .A1(n13985), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10581) );
  INV_X1 U13561 ( .A(n10579), .ZN(n10580) );
  OR2_X1 U13562 ( .A1(n10581), .A2(n10580), .ZN(n10582) );
  NAND2_X1 U13563 ( .A1(n18736), .A2(n10858), .ZN(n10583) );
  INV_X1 U13564 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15332) );
  NOR2_X1 U13565 ( .A1(n10583), .A2(n15332), .ZN(n15344) );
  NAND2_X1 U13566 ( .A1(n10583), .A2(n15332), .ZN(n15048) );
  NAND2_X1 U13567 ( .A1(n13985), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10586) );
  INV_X1 U13568 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12963) );
  INV_X1 U13569 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11087) );
  NOR2_X1 U13570 ( .A1(n10468), .A2(n11087), .ZN(n10603) );
  NAND2_X1 U13571 ( .A1(n13985), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U13572 ( .A1(n10608), .A2(n10607), .ZN(n10610) );
  NOR2_X1 U13573 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(P2_EBX_REG_17__SCAN_IN), 
        .ZN(n10584) );
  NOR2_X1 U13574 ( .A1(n10468), .A2(n10584), .ZN(n10585) );
  MUX2_X1 U13575 ( .A(n13985), .B(n10586), .S(n10600), .Z(n10587) );
  OR2_X1 U13576 ( .A1(n10600), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U13577 ( .A1(n10587), .A2(n10589), .ZN(n18666) );
  INV_X1 U13578 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15247) );
  OAI21_X1 U13579 ( .B1(n18666), .B2(n9804), .A(n15247), .ZN(n15104) );
  INV_X1 U13580 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11106) );
  NOR2_X1 U13581 ( .A1(n10468), .A2(n11106), .ZN(n10588) );
  NAND2_X1 U13582 ( .A1(n10589), .A2(n10588), .ZN(n10591) );
  INV_X1 U13583 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n18667) );
  AND2_X1 U13584 ( .A1(n18667), .A2(n11106), .ZN(n10590) );
  NAND2_X1 U13585 ( .A1(n10591), .A2(n10612), .ZN(n18660) );
  INV_X1 U13586 ( .A(n18660), .ZN(n10592) );
  NAND2_X1 U13587 ( .A1(n10592), .A2(n10858), .ZN(n10625) );
  INV_X1 U13588 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15096) );
  NAND2_X1 U13589 ( .A1(n10625), .A2(n15096), .ZN(n15089) );
  AND2_X1 U13590 ( .A1(n15104), .A2(n15089), .ZN(n15075) );
  NAND2_X1 U13591 ( .A1(n13985), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10593) );
  XNOR2_X1 U13592 ( .A(n10612), .B(n10593), .ZN(n18647) );
  NAND2_X1 U13593 ( .A1(n18647), .A2(n10858), .ZN(n10630) );
  INV_X1 U13594 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10594) );
  NAND2_X1 U13595 ( .A1(n10630), .A2(n10594), .ZN(n15077) );
  AND2_X1 U13596 ( .A1(n15075), .A2(n15077), .ZN(n15063) );
  INV_X1 U13597 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11094) );
  NOR2_X1 U13598 ( .A1(n10468), .A2(n11094), .ZN(n10596) );
  INV_X1 U13599 ( .A(n10659), .ZN(n10595) );
  AOI21_X1 U13600 ( .B1(n10610), .B2(n10596), .A(n10595), .ZN(n10597) );
  OR2_X1 U13601 ( .A1(n10610), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10599) );
  AND2_X1 U13602 ( .A1(n10597), .A2(n10599), .ZN(n18689) );
  NAND2_X1 U13603 ( .A1(n18689), .A2(n10858), .ZN(n10621) );
  XNOR2_X1 U13604 ( .A(n10621), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15129) );
  INV_X1 U13605 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11098) );
  NOR2_X1 U13606 ( .A1(n10468), .A2(n11098), .ZN(n10598) );
  NAND2_X1 U13607 ( .A1(n10599), .A2(n10598), .ZN(n10601) );
  NAND2_X1 U13608 ( .A1(n10601), .A2(n10600), .ZN(n18678) );
  OR2_X1 U13609 ( .A1(n18678), .A2(n9804), .ZN(n10602) );
  INV_X1 U13610 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15275) );
  NAND2_X1 U13611 ( .A1(n10602), .A2(n15275), .ZN(n15059) );
  INV_X1 U13612 ( .A(n10603), .ZN(n10604) );
  XNOR2_X1 U13613 ( .A(n10605), .B(n10604), .ZN(n18712) );
  NAND2_X1 U13614 ( .A1(n18712), .A2(n10858), .ZN(n10606) );
  INV_X1 U13615 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15311) );
  NAND2_X1 U13616 ( .A1(n10606), .A2(n15311), .ZN(n15305) );
  OR2_X1 U13617 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  AND2_X1 U13618 ( .A1(n10610), .A2(n10609), .ZN(n18705) );
  NAND2_X1 U13619 ( .A1(n18705), .A2(n10858), .ZN(n10618) );
  INV_X1 U13620 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15298) );
  NAND2_X1 U13621 ( .A1(n10618), .A2(n15298), .ZN(n15287) );
  NAND2_X1 U13622 ( .A1(n18725), .A2(n10858), .ZN(n10611) );
  INV_X1 U13623 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15333) );
  NAND2_X1 U13624 ( .A1(n10611), .A2(n15333), .ZN(n15323) );
  AND4_X1 U13625 ( .A1(n15059), .A2(n15305), .A3(n15287), .A4(n15323), .ZN(
        n10616) );
  NAND2_X1 U13626 ( .A1(n13985), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10613) );
  INV_X1 U13627 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11112) );
  OAI211_X1 U13628 ( .C1(n10614), .C2(n10613), .A(n10659), .B(n10638), .ZN(
        n12229) );
  OR2_X1 U13629 ( .A1(n12229), .A2(n9804), .ZN(n10615) );
  INV_X1 U13630 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15068) );
  NAND2_X1 U13631 ( .A1(n10615), .A2(n15068), .ZN(n15065) );
  NAND4_X1 U13632 ( .A1(n15063), .A2(n15129), .A3(n10616), .A4(n15065), .ZN(
        n10634) );
  NAND2_X1 U13633 ( .A1(n10858), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10617) );
  OR2_X1 U13634 ( .A1(n12229), .A2(n10617), .ZN(n15064) );
  INV_X1 U13635 ( .A(n10618), .ZN(n10619) );
  NAND2_X1 U13636 ( .A1(n10619), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15288) );
  AND2_X1 U13637 ( .A1(n10858), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10620) );
  NAND2_X1 U13638 ( .A1(n18725), .A2(n10620), .ZN(n15322) );
  AND2_X1 U13639 ( .A1(n15288), .A2(n15322), .ZN(n10624) );
  INV_X1 U13640 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n20764) );
  OR2_X1 U13641 ( .A1(n10621), .A2(n20764), .ZN(n15056) );
  NAND2_X1 U13642 ( .A1(n10858), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10622) );
  OR2_X1 U13643 ( .A1(n18678), .A2(n10622), .ZN(n15058) );
  AND2_X1 U13644 ( .A1(n10858), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10623) );
  NAND2_X1 U13645 ( .A1(n18712), .A2(n10623), .ZN(n15304) );
  AND4_X1 U13646 ( .A1(n10624), .A2(n15056), .A3(n15058), .A4(n15304), .ZN(
        n10629) );
  INV_X1 U13647 ( .A(n10625), .ZN(n10626) );
  NAND2_X1 U13648 ( .A1(n10626), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15090) );
  INV_X1 U13649 ( .A(n18666), .ZN(n10628) );
  AND2_X1 U13650 ( .A1(n10858), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10627) );
  NAND2_X1 U13651 ( .A1(n10628), .A2(n10627), .ZN(n15103) );
  AND4_X1 U13652 ( .A1(n15064), .A2(n10629), .A3(n15090), .A4(n15103), .ZN(
        n10632) );
  INV_X1 U13653 ( .A(n10630), .ZN(n10631) );
  NAND2_X1 U13654 ( .A1(n10631), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15078) );
  NAND2_X1 U13655 ( .A1(n10638), .A2(n10659), .ZN(n10635) );
  NAND2_X1 U13656 ( .A1(n13985), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10636) );
  INV_X1 U13657 ( .A(n10636), .ZN(n10637) );
  NAND2_X1 U13658 ( .A1(n10638), .A2(n10637), .ZN(n10639) );
  OR2_X1 U13659 ( .A1(n15549), .A2(n9804), .ZN(n10640) );
  INV_X1 U13660 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U13661 ( .A1(n10640), .A2(n15197), .ZN(n15200) );
  NAND2_X1 U13662 ( .A1(n15201), .A2(n15200), .ZN(n10641) );
  OR3_X1 U13663 ( .A1(n15549), .A2(n9804), .A3(n15197), .ZN(n15199) );
  NAND2_X1 U13664 ( .A1(n10641), .A2(n15199), .ZN(n16037) );
  INV_X1 U13665 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11029) );
  NOR2_X1 U13666 ( .A1(n10468), .A2(n11029), .ZN(n10642) );
  NAND2_X1 U13667 ( .A1(n10649), .A2(n10643), .ZN(n16019) );
  OR2_X1 U13668 ( .A1(n16019), .A2(n9804), .ZN(n10644) );
  XNOR2_X1 U13669 ( .A(n10644), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16038) );
  NAND2_X1 U13670 ( .A1(n16037), .A2(n16038), .ZN(n10647) );
  NAND2_X1 U13671 ( .A1(n10858), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10645) );
  OR2_X1 U13672 ( .A1(n16019), .A2(n10645), .ZN(n10646) );
  INV_X1 U13673 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14898) );
  NOR2_X1 U13674 ( .A1(n10468), .A2(n14898), .ZN(n10648) );
  NAND2_X1 U13675 ( .A1(n10649), .A2(n10648), .ZN(n10650) );
  NAND2_X1 U13676 ( .A1(n10650), .A2(n10659), .ZN(n10651) );
  NOR2_X1 U13677 ( .A1(n10655), .A2(n10651), .ZN(n16003) );
  NAND2_X1 U13678 ( .A1(n16003), .A2(n10858), .ZN(n15037) );
  INV_X1 U13679 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15192) );
  NOR2_X1 U13680 ( .A1(n15037), .A2(n15192), .ZN(n10653) );
  NAND2_X1 U13681 ( .A1(n15037), .A2(n15192), .ZN(n10652) );
  NAND2_X1 U13682 ( .A1(n13985), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10654) );
  OAI21_X1 U13683 ( .B1(n10655), .B2(n10654), .A(n10659), .ZN(n10656) );
  INV_X1 U13684 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14889) );
  NAND2_X1 U13685 ( .A1(n9638), .A2(n10858), .ZN(n10667) );
  INV_X1 U13686 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15159) );
  AND2_X1 U13687 ( .A1(n10667), .A2(n15159), .ZN(n15168) );
  NAND2_X1 U13688 ( .A1(n13985), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10657) );
  OR2_X1 U13689 ( .A1(n10658), .A2(n10657), .ZN(n10660) );
  INV_X1 U13690 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11124) );
  NAND2_X1 U13691 ( .A1(n10659), .A2(n10662), .ZN(n10661) );
  INV_X1 U13692 ( .A(n10661), .ZN(n14015) );
  XNOR2_X1 U13693 ( .A(n10666), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15029) );
  NAND2_X1 U13694 ( .A1(n13985), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10664) );
  NAND2_X1 U13695 ( .A1(n10661), .A2(n10664), .ZN(n10672) );
  OR2_X1 U13696 ( .A1(n10664), .A2(n10663), .ZN(n10665) );
  AND2_X1 U13697 ( .A1(n10672), .A2(n10665), .ZN(n15970) );
  NAND2_X1 U13698 ( .A1(n15970), .A2(n10858), .ZN(n10670) );
  INV_X1 U13699 ( .A(n10666), .ZN(n10669) );
  INV_X1 U13700 ( .A(n10667), .ZN(n10668) );
  AOI21_X1 U13701 ( .B1(n10669), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15169), .ZN(n13983) );
  INV_X1 U13702 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13543) );
  AOI21_X1 U13703 ( .B1(n13981), .B2(n13983), .A(n10670), .ZN(n10671) );
  INV_X1 U13704 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11025) );
  NOR2_X1 U13705 ( .A1(n10468), .A2(n11025), .ZN(n10673) );
  AOI21_X1 U13706 ( .B1(n10673), .B2(n10672), .A(n14009), .ZN(n10674) );
  INV_X1 U13707 ( .A(n10674), .ZN(n15965) );
  XNOR2_X1 U13708 ( .A(n13982), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10675) );
  NAND2_X1 U13709 ( .A1(n10734), .A2(n10720), .ZN(n10676) );
  NAND2_X1 U13710 ( .A1(n10676), .A2(n9567), .ZN(n10692) );
  NAND2_X1 U13711 ( .A1(n12367), .A2(n9573), .ZN(n10677) );
  MUX2_X1 U13712 ( .A(n10677), .B(n9567), .S(n10719), .Z(n10690) );
  INV_X1 U13713 ( .A(n10678), .ZN(n10731) );
  INV_X1 U13714 ( .A(n10679), .ZN(n10680) );
  XNOR2_X1 U13715 ( .A(n10731), .B(n10680), .ZN(n10722) );
  INV_X1 U13716 ( .A(n10722), .ZN(n10681) );
  OAI21_X1 U13717 ( .B1(n9573), .B2(n10682), .A(n10681), .ZN(n10684) );
  NAND2_X1 U13718 ( .A1(n19683), .A2(n10719), .ZN(n10683) );
  NAND2_X1 U13719 ( .A1(n10684), .A2(n10683), .ZN(n10685) );
  NAND2_X1 U13720 ( .A1(n10685), .A2(n12691), .ZN(n10688) );
  OAI21_X1 U13721 ( .B1(n10731), .B2(n10741), .A(n10686), .ZN(n10687) );
  NAND2_X1 U13722 ( .A1(n10688), .A2(n10687), .ZN(n10689) );
  NAND3_X1 U13723 ( .A1(n10692), .A2(n10690), .A3(n10689), .ZN(n10700) );
  NAND2_X1 U13724 ( .A1(n10692), .A2(n10691), .ZN(n10699) );
  NAND2_X1 U13725 ( .A1(n15610), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10693) );
  NAND2_X1 U13726 ( .A1(n10694), .A2(n10693), .ZN(n10696) );
  INV_X1 U13727 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15531) );
  NAND2_X1 U13728 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15531), .ZN(
        n10695) );
  OAI21_X1 U13729 ( .B1(n9567), .B2(n10721), .A(n10737), .ZN(n10697) );
  INV_X1 U13730 ( .A(n10697), .ZN(n10698) );
  NAND3_X1 U13731 ( .A1(n10700), .A2(n10699), .A3(n10698), .ZN(n10701) );
  MUX2_X1 U13732 ( .A(n10701), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n12317), .Z(n10706) );
  INV_X1 U13733 ( .A(n10737), .ZN(n10702) );
  NAND2_X1 U13734 ( .A1(n10702), .A2(n19690), .ZN(n10703) );
  NAND2_X1 U13735 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19685) );
  INV_X1 U13736 ( .A(n19685), .ZN(n19680) );
  INV_X1 U13737 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20696) );
  NOR2_X1 U13738 ( .A1(n20696), .A2(n19578), .ZN(n19570) );
  NOR2_X1 U13739 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19572) );
  NOR3_X1 U13740 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19570), .A3(n19572), 
        .ZN(n19688) );
  INV_X1 U13741 ( .A(n19688), .ZN(n19566) );
  NOR2_X1 U13742 ( .A1(n19680), .A2(n19566), .ZN(n12575) );
  NAND2_X1 U13743 ( .A1(n12575), .A2(n10704), .ZN(n10753) );
  AOI21_X1 U13744 ( .B1(n10706), .B2(n12691), .A(n10705), .ZN(n10707) );
  NAND2_X1 U13745 ( .A1(n12574), .A2(n10707), .ZN(n10752) );
  NAND2_X1 U13746 ( .A1(n10708), .A2(n10712), .ZN(n10709) );
  NAND2_X1 U13747 ( .A1(n12693), .A2(n10709), .ZN(n10715) );
  NAND2_X1 U13748 ( .A1(n19683), .A2(n13054), .ZN(n10776) );
  NAND2_X1 U13749 ( .A1(n10776), .A2(n12691), .ZN(n10711) );
  NAND2_X1 U13750 ( .A1(n10711), .A2(n10710), .ZN(n10713) );
  NAND2_X1 U13751 ( .A1(n10713), .A2(n10712), .ZN(n10714) );
  NAND2_X1 U13752 ( .A1(n10715), .A2(n10714), .ZN(n10778) );
  INV_X1 U13753 ( .A(n10778), .ZN(n10726) );
  NAND2_X1 U13754 ( .A1(n19683), .A2(n10217), .ZN(n12239) );
  AOI21_X1 U13755 ( .B1(n10716), .B2(n19050), .A(n12239), .ZN(n10777) );
  NOR2_X1 U13756 ( .A1(n10716), .A2(n13054), .ZN(n10717) );
  NOR2_X1 U13757 ( .A1(n10777), .A2(n10717), .ZN(n10725) );
  NAND3_X1 U13758 ( .A1(n10721), .A2(n10720), .A3(n10719), .ZN(n10742) );
  OR2_X1 U13759 ( .A1(n10742), .A2(n10722), .ZN(n10723) );
  NAND3_X1 U13760 ( .A1(n10718), .A2(n12679), .A3(n12575), .ZN(n10724) );
  AND3_X1 U13761 ( .A1(n10726), .A2(n10725), .A3(n10724), .ZN(n12572) );
  MUX2_X1 U13762 ( .A(n10718), .B(n10704), .S(n19683), .Z(n10727) );
  NAND3_X1 U13763 ( .A1(n10727), .A2(n12679), .A3(n19685), .ZN(n10728) );
  NAND2_X1 U13764 ( .A1(n12572), .A2(n10728), .ZN(n10750) );
  INV_X1 U13765 ( .A(n10729), .ZN(n10730) );
  OAI21_X1 U13766 ( .B1(n10732), .B2(n10731), .A(n10730), .ZN(n10736) );
  INV_X1 U13767 ( .A(n10733), .ZN(n10735) );
  NAND3_X1 U13768 ( .A1(n10736), .A2(n10735), .A3(n10734), .ZN(n10738) );
  AND2_X1 U13769 ( .A1(n10738), .A2(n10737), .ZN(n19675) );
  NAND2_X1 U13770 ( .A1(n19675), .A2(n19669), .ZN(n10749) );
  AND2_X1 U13771 ( .A1(n12679), .A2(n13184), .ZN(n10740) );
  OAI21_X1 U13772 ( .B1(n10742), .B2(n10741), .A(n10740), .ZN(n10745) );
  AND2_X1 U13773 ( .A1(n15531), .A2(n10743), .ZN(n15527) );
  INV_X1 U13774 ( .A(n15527), .ZN(n12690) );
  INV_X1 U13775 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12689) );
  OAI21_X1 U13776 ( .B1(n10432), .B2(n12690), .A(n12689), .ZN(n16171) );
  NAND2_X1 U13777 ( .A1(n16171), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10744) );
  INV_X1 U13778 ( .A(n19670), .ZN(n10747) );
  INV_X1 U13779 ( .A(n10739), .ZN(n10746) );
  NAND3_X1 U13780 ( .A1(n10747), .A2(n10746), .A3(n9573), .ZN(n10748) );
  NAND2_X1 U13781 ( .A1(n10749), .A2(n10748), .ZN(n12267) );
  NOR2_X1 U13782 ( .A1(n10750), .A2(n12267), .ZN(n10751) );
  OAI211_X1 U13783 ( .C1(n12574), .C2(n10753), .A(n10752), .B(n10751), .ZN(
        n10755) );
  NAND2_X1 U13784 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13184), .ZN(n19558) );
  NOR2_X1 U13785 ( .A1(n10739), .A2(n9567), .ZN(n19671) );
  INV_X1 U13786 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12319) );
  NOR2_X1 U13787 ( .A1(n13182), .A2(n12319), .ZN(n19008) );
  AND2_X1 U13788 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19008), .ZN(
        n10781) );
  NAND2_X1 U13789 ( .A1(n10757), .A2(n9573), .ZN(n12656) );
  INV_X1 U13790 ( .A(n10777), .ZN(n10758) );
  NAND2_X1 U13791 ( .A1(n12656), .A2(n10758), .ZN(n10760) );
  NAND2_X1 U13792 ( .A1(n10760), .A2(n10759), .ZN(n10773) );
  NOR2_X1 U13793 ( .A1(n10237), .A2(n10761), .ZN(n10763) );
  NAND2_X1 U13794 ( .A1(n10763), .A2(n10762), .ZN(n12987) );
  NAND2_X1 U13795 ( .A1(n10217), .A2(n10704), .ZN(n10764) );
  OAI211_X1 U13796 ( .C1(n10705), .C2(n12268), .A(n12987), .B(n10764), .ZN(
        n10765) );
  INV_X1 U13797 ( .A(n10765), .ZN(n10770) );
  OAI21_X1 U13798 ( .B1(n10762), .B2(n10766), .A(n12268), .ZN(n10768) );
  NAND2_X1 U13799 ( .A1(n10768), .A2(n10767), .ZN(n10769) );
  AND3_X1 U13800 ( .A1(n10771), .A2(n10770), .A3(n10769), .ZN(n10772) );
  AND2_X1 U13801 ( .A1(n10773), .A2(n10772), .ZN(n12644) );
  NAND2_X1 U13802 ( .A1(n12644), .A2(n10774), .ZN(n10775) );
  NAND2_X1 U13803 ( .A1(n11174), .A2(n10775), .ZN(n19006) );
  NAND2_X1 U13804 ( .A1(n11174), .A2(n12684), .ZN(n15258) );
  OR2_X1 U13805 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19008), .ZN(
        n10795) );
  OR2_X1 U13806 ( .A1(n15258), .A2(n10795), .ZN(n19012) );
  INV_X1 U13807 ( .A(n11174), .ZN(n10780) );
  NOR2_X1 U13808 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19634) );
  NOR2_X1 U13809 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n10779) );
  AND2_X2 U13810 ( .A1(n19634), .A2(n10779), .ZN(n18980) );
  INV_X2 U13811 ( .A(n18980), .ZN(n19016) );
  NAND2_X1 U13812 ( .A1(n10780), .A2(n19016), .ZN(n19001) );
  OAI211_X1 U13813 ( .C1(n10781), .C2(n19006), .A(n19012), .B(n19001), .ZN(
        n12728) );
  INV_X1 U13814 ( .A(n12728), .ZN(n10788) );
  OR2_X1 U13815 ( .A1(n15400), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10782) );
  NAND2_X1 U13816 ( .A1(n10788), .A2(n10782), .ZN(n16151) );
  NOR2_X1 U13817 ( .A1(n12844), .A2(n11159), .ZN(n13268) );
  NAND4_X1 U13818 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n13268), .ZN(n10798) );
  INV_X1 U13819 ( .A(n10798), .ZN(n10783) );
  NOR2_X1 U13820 ( .A1(n15400), .A2(n10783), .ZN(n10784) );
  NOR2_X1 U13821 ( .A1(n16151), .A2(n10784), .ZN(n15366) );
  AND2_X1 U13822 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15269) );
  NAND3_X1 U13823 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15270) );
  INV_X1 U13824 ( .A(n15270), .ZN(n10785) );
  AND2_X1 U13825 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n10785), .ZN(
        n10786) );
  AND2_X1 U13826 ( .A1(n15269), .A2(n10786), .ZN(n15260) );
  AND3_X1 U13827 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15084) );
  NAND2_X1 U13828 ( .A1(n15260), .A2(n15084), .ZN(n15223) );
  INV_X1 U13829 ( .A(n15223), .ZN(n15222) );
  AND3_X1 U13830 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13831 ( .A1(n15222), .A2(n10787), .ZN(n15214) );
  NOR2_X1 U13832 ( .A1(n15068), .A2(n15214), .ZN(n10789) );
  AOI21_X1 U13833 ( .B1(n15366), .B2(n10789), .A(n15365), .ZN(n16124) );
  NAND2_X1 U13834 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16128) );
  INV_X1 U13835 ( .A(n16128), .ZN(n10790) );
  NOR2_X1 U13836 ( .A1(n15365), .A2(n10790), .ZN(n10791) );
  OR2_X1 U13837 ( .A1(n16124), .A2(n10791), .ZN(n15186) );
  AND2_X1 U13838 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15158) );
  AND2_X1 U13839 ( .A1(n15158), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10792) );
  NOR2_X1 U13840 ( .A1(n15365), .A2(n10792), .ZN(n10793) );
  INV_X1 U13841 ( .A(n13542), .ZN(n10802) );
  NAND2_X1 U13842 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19008), .ZN(
        n10794) );
  NAND2_X1 U13843 ( .A1(n15258), .A2(n10794), .ZN(n10796) );
  NAND2_X1 U13844 ( .A1(n10796), .A2(n10795), .ZN(n10797) );
  NOR2_X1 U13845 ( .A1(n15400), .A2(n10797), .ZN(n12729) );
  NAND2_X1 U13846 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12729), .ZN(
        n12842) );
  NOR3_X1 U13847 ( .A1(n15068), .A2(n15214), .A3(n15385), .ZN(n16129) );
  INV_X1 U13848 ( .A(n16129), .ZN(n10799) );
  NOR2_X1 U13849 ( .A1(n16128), .A2(n10799), .ZN(n15193) );
  NAND2_X1 U13850 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15193), .ZN(
        n15176) );
  INV_X1 U13851 ( .A(n15176), .ZN(n10800) );
  NAND2_X1 U13852 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14043) );
  NAND2_X1 U13853 ( .A1(n15149), .A2(n14043), .ZN(n10801) );
  NAND2_X1 U13854 ( .A1(n10802), .A2(n10801), .ZN(n15154) );
  INV_X1 U13855 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10804) );
  OR2_X1 U13856 ( .A1(n10827), .A2(n10804), .ZN(n10809) );
  INV_X1 U13857 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n10806) );
  NAND2_X1 U13858 ( .A1(n9573), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10805) );
  OAI211_X1 U13859 ( .C1(n19050), .C2(n10806), .A(n10805), .B(n19639), .ZN(
        n10807) );
  INV_X1 U13860 ( .A(n10807), .ZN(n10808) );
  NAND2_X1 U13861 ( .A1(n10809), .A2(n10808), .ZN(n12984) );
  AND2_X1 U13862 ( .A1(n10468), .A2(n19639), .ZN(n10810) );
  AND2_X1 U13863 ( .A1(n9573), .A2(n19639), .ZN(n10828) );
  NAND2_X1 U13864 ( .A1(n10811), .A2(n10828), .ZN(n10826) );
  NOR2_X1 U13865 ( .A1(n19050), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10812) );
  AND2_X1 U13866 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10813) );
  NOR2_X1 U13867 ( .A1(n10812), .A2(n10813), .ZN(n10814) );
  OR2_X1 U13868 ( .A1(n10827), .A2(n10240), .ZN(n10816) );
  AOI22_X1 U13869 ( .A1(n10812), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10828), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10815) );
  AND2_X1 U13870 ( .A1(n10816), .A2(n10815), .ZN(n10822) );
  XNOR2_X1 U13871 ( .A(n10821), .B(n10822), .ZN(n12434) );
  NAND2_X1 U13872 ( .A1(n10229), .A2(n19050), .ZN(n10818) );
  MUX2_X1 U13873 ( .A(n10818), .B(n10817), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10820) );
  INV_X1 U13874 ( .A(n10978), .ZN(n10859) );
  NAND2_X1 U13875 ( .A1(n10859), .A2(n11141), .ZN(n10819) );
  NAND2_X1 U13876 ( .A1(n10820), .A2(n10819), .ZN(n12433) );
  NAND2_X1 U13877 ( .A1(n10822), .A2(n10821), .ZN(n10823) );
  NAND2_X1 U13878 ( .A1(n12436), .A2(n10823), .ZN(n10832) );
  INV_X1 U13879 ( .A(n10824), .ZN(n11147) );
  NAND2_X1 U13880 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10825) );
  OAI211_X1 U13881 ( .C1(n11147), .C2(n10978), .A(n10826), .B(n10825), .ZN(
        n10831) );
  XNOR2_X1 U13882 ( .A(n10832), .B(n10831), .ZN(n12981) );
  OR2_X1 U13883 ( .A1(n10827), .A2(n10269), .ZN(n10830) );
  INV_X2 U13884 ( .A(n11004), .ZN(n10987) );
  INV_X2 U13885 ( .A(n11003), .ZN(n14040) );
  AOI22_X1 U13886 ( .A1(n10987), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n14040), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10829) );
  AND2_X1 U13887 ( .A1(n10830), .A2(n10829), .ZN(n12980) );
  INV_X1 U13888 ( .A(n10831), .ZN(n10833) );
  NAND2_X1 U13889 ( .A1(n10833), .A2(n10832), .ZN(n10834) );
  OR2_X1 U13890 ( .A1(n10827), .A2(n12737), .ZN(n10841) );
  AOI22_X1 U13891 ( .A1(n14040), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10837) );
  NAND2_X1 U13892 ( .A1(n10987), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10836) );
  OAI211_X1 U13893 ( .C1(n10838), .C2(n10978), .A(n10837), .B(n10836), .ZN(
        n10839) );
  INV_X1 U13894 ( .A(n10839), .ZN(n10840) );
  AND2_X1 U13895 ( .A1(n10841), .A2(n10840), .ZN(n12730) );
  INV_X1 U13896 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10842) );
  OR2_X1 U13897 ( .A1(n10827), .A2(n10842), .ZN(n10844) );
  AOI22_X1 U13898 ( .A1(n10987), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n14040), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10843) );
  OAI211_X1 U13899 ( .C1(n11152), .C2(n10978), .A(n10844), .B(n10843), .ZN(
        n12839) );
  INV_X1 U13900 ( .A(n12840), .ZN(n10852) );
  INV_X1 U13901 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10845) );
  OR2_X1 U13902 ( .A1(n10827), .A2(n10845), .ZN(n10851) );
  NAND2_X1 U13903 ( .A1(n10987), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U13904 ( .A1(n14040), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10846) );
  OAI211_X1 U13905 ( .C1(n10978), .C2(n10848), .A(n10847), .B(n10846), .ZN(
        n10849) );
  INV_X1 U13906 ( .A(n10849), .ZN(n10850) );
  NAND2_X1 U13907 ( .A1(n10851), .A2(n10850), .ZN(n16146) );
  NAND2_X1 U13908 ( .A1(n10852), .A2(n16146), .ZN(n16147) );
  NAND2_X1 U13909 ( .A1(n10859), .A2(n10853), .ZN(n10854) );
  INV_X1 U13910 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10855) );
  OR2_X1 U13911 ( .A1(n10827), .A2(n10855), .ZN(n10857) );
  AOI22_X1 U13912 ( .A1(n10987), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n14040), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10856) );
  NAND2_X1 U13913 ( .A1(n10857), .A2(n10856), .ZN(n13168) );
  NAND2_X1 U13914 ( .A1(n13169), .A2(n13168), .ZN(n13167) );
  NAND2_X1 U13915 ( .A1(n10859), .A2(n10858), .ZN(n10860) );
  INV_X1 U13916 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10861) );
  OR2_X1 U13917 ( .A1(n10827), .A2(n10861), .ZN(n10863) );
  AOI22_X1 U13918 ( .A1(n10987), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n14040), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13919 ( .A1(n10432), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13920 ( .A1(n10344), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13921 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13922 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10865) );
  NAND4_X1 U13923 ( .A1(n10868), .A2(n10867), .A3(n10866), .A4(n10865), .ZN(
        n10874) );
  AOI22_X1 U13924 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U13925 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13926 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14122), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13927 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10869) );
  NAND4_X1 U13928 ( .A1(n10872), .A2(n10871), .A3(n10870), .A4(n10869), .ZN(
        n10873) );
  INV_X1 U13929 ( .A(n12602), .ZN(n10878) );
  INV_X1 U13930 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10875) );
  OR2_X1 U13931 ( .A1(n10827), .A2(n10875), .ZN(n10877) );
  AOI22_X1 U13932 ( .A1(n10987), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n14040), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10876) );
  OAI211_X1 U13933 ( .C1(n10878), .C2(n10978), .A(n10877), .B(n10876), .ZN(
        n13322) );
  INV_X1 U13934 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n10879) );
  OR2_X1 U13935 ( .A1(n10827), .A2(n10879), .ZN(n10894) );
  AOI22_X1 U13936 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U13937 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10384), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U13938 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13939 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10880) );
  NAND4_X1 U13940 ( .A1(n10883), .A2(n10882), .A3(n10881), .A4(n10880), .ZN(
        n10889) );
  AOI22_X1 U13941 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14120), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13942 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14121), .ZN(n10886) );
  AOI22_X1 U13943 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n14122), .ZN(n10885) );
  AOI22_X1 U13944 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10884) );
  NAND4_X1 U13945 ( .A1(n10887), .A2(n10886), .A3(n10885), .A4(n10884), .ZN(
        n10888) );
  NOR2_X1 U13946 ( .A1(n10889), .A2(n10888), .ZN(n12624) );
  NAND2_X1 U13947 ( .A1(n10987), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n10891) );
  NAND2_X1 U13948 ( .A1(n14040), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10890) );
  OAI211_X1 U13949 ( .C1(n10978), .C2(n12624), .A(n10891), .B(n10890), .ZN(
        n10892) );
  INV_X1 U13950 ( .A(n10892), .ZN(n10893) );
  AOI22_X1 U13951 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13952 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10384), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13953 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10400), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13954 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10895) );
  NAND4_X1 U13955 ( .A1(n10898), .A2(n10897), .A3(n10896), .A4(n10895), .ZN(
        n10904) );
  AOI22_X1 U13956 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13957 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__2__SCAN_IN), .B2(n10350), .ZN(n10901) );
  AOI22_X1 U13958 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n14122), .ZN(n10900) );
  AOI22_X1 U13959 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14123), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10899) );
  NAND4_X1 U13960 ( .A1(n10902), .A2(n10901), .A3(n10900), .A4(n10899), .ZN(
        n10903) );
  INV_X1 U13961 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10905) );
  OR2_X1 U13962 ( .A1(n10827), .A2(n10905), .ZN(n10907) );
  AOI22_X1 U13963 ( .A1(n10987), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10906) );
  OAI211_X1 U13964 ( .C1(n12867), .C2(n10978), .A(n10907), .B(n10906), .ZN(
        n15371) );
  AOI22_X1 U13965 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10911) );
  INV_X1 U13966 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20810) );
  AOI22_X1 U13967 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10384), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13968 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13969 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10908) );
  NAND4_X1 U13970 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n10917) );
  AOI22_X1 U13971 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14120), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13972 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n14121), .ZN(n10914) );
  AOI22_X1 U13973 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14122), .ZN(n10913) );
  AOI22_X1 U13974 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10912) );
  NAND4_X1 U13975 ( .A1(n10915), .A2(n10914), .A3(n10913), .A4(n10912), .ZN(
        n10916) );
  INV_X1 U13976 ( .A(n12748), .ZN(n10918) );
  NOR2_X1 U13977 ( .A1(n10978), .A2(n10918), .ZN(n10921) );
  NAND2_X1 U13978 ( .A1(n10987), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n10919) );
  OAI21_X1 U13979 ( .B1(n11003), .B2(n11075), .A(n10919), .ZN(n10920) );
  AOI211_X1 U13980 ( .C1(n10835), .C2(P2_REIP_REG_11__SCAN_IN), .A(n10921), 
        .B(n10920), .ZN(n16135) );
  AOI22_X1 U13981 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10384), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13982 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U13983 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10400), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13984 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10922) );
  NAND4_X1 U13985 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n10931) );
  AOI22_X1 U13986 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13987 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__4__SCAN_IN), .B2(n10350), .ZN(n10928) );
  AOI22_X1 U13988 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n14122), .ZN(n10927) );
  AOI22_X1 U13989 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14123), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10926) );
  NAND4_X1 U13990 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n10930) );
  INV_X1 U13991 ( .A(n12751), .ZN(n10935) );
  INV_X1 U13992 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10932) );
  OR2_X1 U13993 ( .A1(n10827), .A2(n10932), .ZN(n10934) );
  AOI22_X1 U13994 ( .A1(n10987), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10933) );
  OAI211_X1 U13995 ( .C1(n10935), .C2(n10978), .A(n10934), .B(n10933), .ZN(
        n15350) );
  INV_X1 U13996 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n10936) );
  OR2_X1 U13997 ( .A1(n10827), .A2(n10936), .ZN(n10951) );
  AOI22_X1 U13998 ( .A1(n10344), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U13999 ( .A1(n10432), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U14000 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U14001 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10937) );
  NAND4_X1 U14002 ( .A1(n10940), .A2(n10939), .A3(n10938), .A4(n10937), .ZN(
        n10946) );
  AOI22_X1 U14003 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U14004 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U14005 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14122), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U14006 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10941) );
  NAND4_X1 U14007 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n10945) );
  NOR2_X1 U14008 ( .A1(n10946), .A2(n10945), .ZN(n13007) );
  NAND2_X1 U14009 ( .A1(n10987), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n10948) );
  NAND2_X1 U14010 ( .A1(n14040), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10947) );
  OAI211_X1 U14011 ( .C1(n10978), .C2(n13007), .A(n10948), .B(n10947), .ZN(
        n10949) );
  INV_X1 U14012 ( .A(n10949), .ZN(n10950) );
  AOI22_X1 U14013 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10432), .B1(
        n10344), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U14014 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10384), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U14015 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U14016 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10952) );
  NAND4_X1 U14017 ( .A1(n10955), .A2(n10954), .A3(n10953), .A4(n10952), .ZN(
        n10961) );
  AOI22_X1 U14018 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10437), .B1(
        n14120), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U14019 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n10350), .ZN(n10958) );
  AOI22_X1 U14020 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n14122), .ZN(n10957) );
  AOI22_X1 U14021 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14123), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10956) );
  NAND4_X1 U14022 ( .A1(n10959), .A2(n10958), .A3(n10957), .A4(n10956), .ZN(
        n10960) );
  INV_X1 U14023 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10962) );
  OR2_X1 U14024 ( .A1(n10827), .A2(n10962), .ZN(n10964) );
  AOI22_X1 U14025 ( .A1(n10987), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10963) );
  OAI211_X1 U14026 ( .C1(n13009), .C2(n10978), .A(n10964), .B(n10963), .ZN(
        n15315) );
  INV_X1 U14027 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n11091) );
  OR2_X1 U14028 ( .A1(n10827), .A2(n11091), .ZN(n10981) );
  AOI22_X1 U14029 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U14030 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n10432), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U14031 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10966) );
  AOI22_X1 U14032 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10965) );
  NAND4_X1 U14033 ( .A1(n10968), .A2(n10967), .A3(n10966), .A4(n10965), .ZN(
        n10974) );
  AOI22_X1 U14034 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n14120), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U14035 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14121), .ZN(n10971) );
  AOI22_X1 U14036 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n14122), .ZN(n10970) );
  AOI22_X1 U14037 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10969) );
  NAND4_X1 U14038 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10973) );
  INV_X1 U14039 ( .A(n13189), .ZN(n10977) );
  NAND2_X1 U14040 ( .A1(n10987), .A2(P2_EAX_REG_15__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U14041 ( .A1(n14040), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10975) );
  OAI211_X1 U14042 ( .C1(n10978), .C2(n10977), .A(n10976), .B(n10975), .ZN(
        n10979) );
  INV_X1 U14043 ( .A(n10979), .ZN(n10980) );
  INV_X1 U14044 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19595) );
  OR2_X1 U14045 ( .A1(n10827), .A2(n19595), .ZN(n10983) );
  AOI22_X1 U14046 ( .A1(n10987), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U14047 ( .A1(n10983), .A2(n10982), .ZN(n13208) );
  INV_X1 U14048 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n10984) );
  OR2_X1 U14049 ( .A1(n10827), .A2(n10984), .ZN(n10986) );
  AOI22_X1 U14050 ( .A1(n10987), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U14051 ( .A1(n10986), .A2(n10985), .ZN(n13248) );
  INV_X1 U14052 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19598) );
  OR2_X1 U14053 ( .A1(n10827), .A2(n19598), .ZN(n10989) );
  AOI22_X1 U14054 ( .A1(n10987), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U14055 ( .A1(n10989), .A2(n10988), .ZN(n13384) );
  INV_X1 U14056 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n15097) );
  OR2_X1 U14057 ( .A1(n10827), .A2(n15097), .ZN(n10991) );
  AOI22_X1 U14058 ( .A1(n10987), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10990) );
  INV_X1 U14059 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19601) );
  OR2_X1 U14060 ( .A1(n10827), .A2(n19601), .ZN(n10993) );
  AOI22_X1 U14061 ( .A1(n10987), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U14062 ( .A1(n10993), .A2(n10992), .ZN(n15001) );
  INV_X1 U14063 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19602) );
  OR2_X1 U14064 ( .A1(n10827), .A2(n19602), .ZN(n10995) );
  AOI22_X1 U14065 ( .A1(n10987), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10994) );
  NAND2_X1 U14066 ( .A1(n10995), .A2(n10994), .ZN(n12235) );
  INV_X1 U14067 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19604) );
  OR2_X1 U14068 ( .A1(n10827), .A2(n19604), .ZN(n10997) );
  AOI22_X1 U14069 ( .A1(n10987), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10996) );
  NAND2_X1 U14070 ( .A1(n10997), .A2(n10996), .ZN(n14983) );
  INV_X1 U14071 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n10998) );
  OR2_X1 U14072 ( .A1(n10827), .A2(n10998), .ZN(n11000) );
  AOI22_X1 U14073 ( .A1(n10987), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10999) );
  NAND2_X1 U14074 ( .A1(n11000), .A2(n10999), .ZN(n16012) );
  INV_X1 U14075 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19607) );
  OR2_X1 U14076 ( .A1(n10827), .A2(n19607), .ZN(n11002) );
  AOI22_X1 U14077 ( .A1(n10987), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11001) );
  AND2_X1 U14078 ( .A1(n11002), .A2(n11001), .ZN(n14975) );
  INV_X1 U14079 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14967) );
  OAI22_X1 U14080 ( .A1(n11004), .A2(n14967), .B1(n15159), .B2(n11003), .ZN(
        n11005) );
  AOI21_X1 U14081 ( .B1(n10835), .B2(P2_REIP_REG_25__SCAN_IN), .A(n11005), 
        .ZN(n14964) );
  INV_X1 U14082 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19611) );
  OR2_X1 U14083 ( .A1(n10827), .A2(n19611), .ZN(n11007) );
  AOI22_X1 U14084 ( .A1(n10987), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U14085 ( .A1(n11007), .A2(n11006), .ZN(n14955) );
  NAND2_X1 U14086 ( .A1(n14965), .A2(n14955), .ZN(n14957) );
  INV_X1 U14087 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19615) );
  OR2_X1 U14088 ( .A1(n10827), .A2(n19615), .ZN(n11009) );
  AOI22_X1 U14089 ( .A1(n10987), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11008) );
  INV_X1 U14090 ( .A(n11015), .ZN(n11012) );
  INV_X1 U14091 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19616) );
  OR2_X1 U14092 ( .A1(n10827), .A2(n19616), .ZN(n11011) );
  AOI22_X1 U14093 ( .A1(n10987), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11010) );
  AND2_X1 U14094 ( .A1(n11011), .A2(n11010), .ZN(n11013) );
  AND2_X1 U14095 ( .A1(n11012), .A2(n11013), .ZN(n11016) );
  INV_X1 U14096 ( .A(n11013), .ZN(n11014) );
  AND2_X1 U14097 ( .A1(n12681), .A2(n9573), .ZN(n11020) );
  NOR2_X1 U14098 ( .A1(n11018), .A2(n11019), .ZN(n12682) );
  OR2_X1 U14099 ( .A1(n11020), .A2(n12682), .ZN(n11021) );
  NAND2_X1 U14100 ( .A1(n14022), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U14101 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11023) );
  OAI211_X1 U14102 ( .C1(n13993), .C2(n11025), .A(n11024), .B(n11023), .ZN(
        n11026) );
  AOI21_X1 U14103 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11026), .ZN(n11132) );
  NAND2_X1 U14104 ( .A1(n13995), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11032) );
  NAND2_X1 U14105 ( .A1(n14022), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U14106 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11027) );
  OAI211_X1 U14107 ( .C1(n13993), .C2(n11029), .A(n11028), .B(n11027), .ZN(
        n11030) );
  INV_X1 U14108 ( .A(n11030), .ZN(n11031) );
  NAND2_X1 U14109 ( .A1(n11032), .A2(n11031), .ZN(n14902) );
  INV_X1 U14110 ( .A(n11033), .ZN(n11035) );
  NAND2_X1 U14111 ( .A1(n11037), .A2(n11036), .ZN(n11038) );
  INV_X1 U14112 ( .A(n11039), .ZN(n11042) );
  INV_X1 U14113 ( .A(n11040), .ZN(n11041) );
  NAND2_X1 U14114 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  NAND2_X1 U14115 ( .A1(n14022), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11045) );
  NAND2_X1 U14116 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11044) );
  OAI211_X1 U14117 ( .C1(n13993), .C2(n18825), .A(n11045), .B(n11044), .ZN(
        n11046) );
  AOI21_X1 U14118 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11046), .ZN(n12848) );
  NAND2_X1 U14119 ( .A1(n14022), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11049) );
  NAND2_X1 U14120 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11048) );
  OAI211_X1 U14121 ( .C1(n11050), .C2(n13993), .A(n11049), .B(n11048), .ZN(
        n11051) );
  AOI21_X1 U14122 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11051), .ZN(n13962) );
  INV_X1 U14123 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12569) );
  NAND2_X1 U14124 ( .A1(n14022), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U14125 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11052) );
  OAI211_X1 U14126 ( .C1(n12569), .C2(n13993), .A(n11053), .B(n11052), .ZN(
        n11054) );
  AOI21_X1 U14127 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11054), .ZN(n12564) );
  NAND2_X1 U14128 ( .A1(n13995), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11060) );
  NAND2_X1 U14129 ( .A1(n14022), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11056) );
  NAND2_X1 U14130 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11055) );
  OAI211_X1 U14131 ( .C1(n11057), .C2(n13993), .A(n11056), .B(n11055), .ZN(
        n11058) );
  INV_X1 U14132 ( .A(n11058), .ZN(n11059) );
  NAND2_X1 U14133 ( .A1(n11060), .A2(n11059), .ZN(n12550) );
  INV_X1 U14134 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12610) );
  NAND2_X1 U14135 ( .A1(n14022), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U14136 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11061) );
  OAI211_X1 U14137 ( .C1(n12610), .C2(n13993), .A(n11062), .B(n11061), .ZN(
        n11063) );
  AOI21_X1 U14138 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11063), .ZN(n12604) );
  NAND2_X1 U14139 ( .A1(n13995), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11069) );
  NAND2_X1 U14140 ( .A1(n14022), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11065) );
  NAND2_X1 U14141 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11064) );
  OAI211_X1 U14142 ( .C1(n11066), .C2(n13993), .A(n11065), .B(n11064), .ZN(
        n11067) );
  INV_X1 U14143 ( .A(n11067), .ZN(n11068) );
  NAND2_X1 U14144 ( .A1(n11069), .A2(n11068), .ZN(n12598) );
  NAND2_X1 U14145 ( .A1(n14022), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11071) );
  NAND2_X1 U14146 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11070) );
  OAI211_X1 U14147 ( .C1(n9839), .C2(n13993), .A(n11071), .B(n11070), .ZN(
        n11072) );
  AOI21_X1 U14148 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11072), .ZN(n12863) );
  AOI22_X1 U14149 ( .A1(n10247), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11074) );
  NAND2_X1 U14150 ( .A1(n14022), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11073) );
  OAI211_X1 U14151 ( .C1(n14026), .C2(n11075), .A(n11074), .B(n11073), .ZN(
        n12629) );
  NAND2_X1 U14152 ( .A1(n12627), .A2(n12629), .ZN(n12628) );
  INV_X1 U14153 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U14154 ( .A1(n14022), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11077) );
  NAND2_X1 U14155 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11076) );
  OAI211_X1 U14156 ( .C1(n11078), .C2(n13993), .A(n11077), .B(n11076), .ZN(
        n11079) );
  AOI21_X1 U14157 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11079), .ZN(n12744) );
  NAND2_X1 U14158 ( .A1(n13995), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11084) );
  NAND2_X1 U14159 ( .A1(n14022), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U14160 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11080) );
  OAI211_X1 U14161 ( .C1(n12963), .C2(n13993), .A(n11081), .B(n11080), .ZN(
        n11082) );
  INV_X1 U14162 ( .A(n11082), .ZN(n11083) );
  NAND2_X1 U14163 ( .A1(n11084), .A2(n11083), .ZN(n12961) );
  NAND2_X1 U14164 ( .A1(n14022), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11086) );
  NAND2_X1 U14165 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11085) );
  OAI211_X1 U14166 ( .C1(n11087), .C2(n13993), .A(n11086), .B(n11085), .ZN(
        n11088) );
  AOI21_X1 U14167 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11088), .ZN(n13004) );
  NAND2_X1 U14168 ( .A1(n13995), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11090) );
  AOI22_X1 U14169 ( .A1(n10247), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11089) );
  OAI211_X1 U14170 ( .C1(n11130), .C2(n11091), .A(n11090), .B(n11089), .ZN(
        n13029) );
  NAND2_X1 U14171 ( .A1(n14022), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11093) );
  NAND2_X1 U14172 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11092) );
  OAI211_X1 U14173 ( .C1(n11094), .C2(n13993), .A(n11093), .B(n11092), .ZN(
        n11095) );
  AOI21_X1 U14174 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11095), .ZN(n13203) );
  NAND2_X1 U14175 ( .A1(n14022), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U14176 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11096) );
  OAI211_X1 U14177 ( .C1(n11098), .C2(n13993), .A(n11097), .B(n11096), .ZN(
        n11099) );
  AOI21_X1 U14178 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11099), .ZN(n13338) );
  NAND2_X1 U14179 ( .A1(n13202), .A2(n11100), .ZN(n13337) );
  NAND2_X1 U14180 ( .A1(n14022), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U14181 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11101) );
  OAI211_X1 U14182 ( .C1(n13993), .C2(n18667), .A(n11102), .B(n11101), .ZN(
        n11103) );
  AOI21_X1 U14183 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11103), .ZN(n13359) );
  NAND2_X1 U14184 ( .A1(n14022), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14185 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11104) );
  OAI211_X1 U14186 ( .C1(n11106), .C2(n13993), .A(n11105), .B(n11104), .ZN(
        n11107) );
  AOI21_X1 U14187 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11107), .ZN(n14924) );
  NAND2_X1 U14188 ( .A1(n13995), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11109) );
  AOI22_X1 U14189 ( .A1(n10247), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11108) );
  OAI211_X1 U14190 ( .C1(n11130), .C2(n19601), .A(n11109), .B(n11108), .ZN(
        n13472) );
  NAND2_X1 U14191 ( .A1(n14022), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U14192 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11110) );
  OAI211_X1 U14193 ( .C1(n11112), .C2(n13993), .A(n11111), .B(n11110), .ZN(
        n11113) );
  AOI21_X1 U14194 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11113), .ZN(n12230) );
  AOI22_X1 U14195 ( .A1(n10247), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11114) );
  OAI21_X1 U14196 ( .B1(n11130), .B2(n19604), .A(n11114), .ZN(n11115) );
  AOI21_X1 U14197 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11115), .ZN(n14914) );
  NAND2_X1 U14198 ( .A1(n14902), .A2(n14913), .ZN(n14901) );
  NAND2_X1 U14199 ( .A1(n14022), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11117) );
  NAND2_X1 U14200 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11116) );
  OAI211_X1 U14201 ( .C1(n13993), .C2(n14898), .A(n11117), .B(n11116), .ZN(
        n11118) );
  AOI21_X1 U14202 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11118), .ZN(n14895) );
  NAND2_X1 U14203 ( .A1(n14022), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11120) );
  NAND2_X1 U14204 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11119) );
  OAI211_X1 U14205 ( .C1(n13993), .C2(n14889), .A(n11120), .B(n11119), .ZN(
        n11121) );
  AOI21_X1 U14206 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11121), .ZN(n14887) );
  NAND2_X1 U14207 ( .A1(n13995), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11127) );
  NAND2_X1 U14208 ( .A1(n14022), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11123) );
  NAND2_X1 U14209 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11122) );
  OAI211_X1 U14210 ( .C1(n13993), .C2(n11124), .A(n11123), .B(n11122), .ZN(
        n11125) );
  INV_X1 U14211 ( .A(n11125), .ZN(n11126) );
  NAND2_X1 U14212 ( .A1(n11127), .A2(n11126), .ZN(n14880) );
  NAND2_X1 U14213 ( .A1(n13995), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11129) );
  AOI22_X1 U14214 ( .A1(n10247), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11128) );
  OAI211_X1 U14215 ( .C1(n11130), .C2(n19615), .A(n11129), .B(n11128), .ZN(
        n13534) );
  INV_X1 U14216 ( .A(n13997), .ZN(n11131) );
  AOI21_X1 U14217 ( .B1(n11132), .B2(n13536), .A(n11131), .ZN(n13525) );
  NAND2_X1 U14218 ( .A1(n11133), .A2(n19683), .ZN(n11135) );
  INV_X1 U14219 ( .A(n12585), .ZN(n11134) );
  NAND2_X1 U14220 ( .A1(n11135), .A2(n11134), .ZN(n11136) );
  NAND2_X1 U14221 ( .A1(n11174), .A2(n11136), .ZN(n16158) );
  AND2_X1 U14222 ( .A1(n18980), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n13524) );
  AOI21_X1 U14223 ( .B1(n13525), .B2(n19004), .A(n13524), .ZN(n11137) );
  OAI21_X1 U14224 ( .B1(n15969), .B2(n18995), .A(n11137), .ZN(n11139) );
  NOR2_X1 U14225 ( .A1(n13542), .A2(n14043), .ZN(n14045) );
  INV_X1 U14226 ( .A(n15149), .ZN(n13538) );
  NOR3_X1 U14227 ( .A1(n14045), .A2(n13538), .A3(n13543), .ZN(n11138) );
  AOI211_X1 U14228 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15154), .A(
        n11139), .B(n11138), .ZN(n11176) );
  INV_X1 U14229 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13984) );
  OR2_X1 U14230 ( .A1(n12320), .A2(n12319), .ZN(n12322) );
  INV_X1 U14231 ( .A(n12322), .ZN(n11143) );
  XNOR2_X1 U14232 ( .A(n11142), .B(n11141), .ZN(n11144) );
  NAND2_X1 U14233 ( .A1(n11143), .A2(n11144), .ZN(n11145) );
  XNOR2_X1 U14234 ( .A(n11144), .B(n12322), .ZN(n12333) );
  NAND2_X1 U14235 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12333), .ZN(
        n12332) );
  NAND2_X1 U14236 ( .A1(n11145), .A2(n12332), .ZN(n11148) );
  XNOR2_X1 U14237 ( .A(n19007), .B(n11148), .ZN(n13977) );
  XOR2_X1 U14238 ( .A(n11147), .B(n11146), .Z(n13976) );
  NAND2_X1 U14239 ( .A1(n13977), .A2(n13976), .ZN(n13975) );
  NAND2_X1 U14240 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11148), .ZN(
        n11149) );
  NAND2_X1 U14241 ( .A1(n13975), .A2(n11149), .ZN(n11150) );
  XNOR2_X1 U14242 ( .A(n11150), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12727) );
  NAND2_X1 U14243 ( .A1(n11150), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11151) );
  XNOR2_X1 U14244 ( .A(n11153), .B(n11152), .ZN(n11154) );
  XNOR2_X1 U14245 ( .A(n11156), .B(n11154), .ZN(n12837) );
  INV_X1 U14246 ( .A(n11154), .ZN(n11155) );
  OR2_X1 U14247 ( .A1(n11156), .A2(n11155), .ZN(n11157) );
  INV_X1 U14248 ( .A(n11158), .ZN(n11160) );
  INV_X1 U14249 ( .A(n11164), .ZN(n16111) );
  NAND2_X1 U14250 ( .A1(n16111), .A2(n11161), .ZN(n11162) );
  OAI211_X1 U14251 ( .C1(n11165), .C2(n9633), .A(n11163), .B(n11162), .ZN(
        n13161) );
  NAND2_X1 U14252 ( .A1(n13161), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13160) );
  NAND2_X1 U14253 ( .A1(n11165), .A2(n11164), .ZN(n11166) );
  NAND2_X1 U14254 ( .A1(n11166), .A2(n9633), .ZN(n11167) );
  INV_X1 U14255 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11169) );
  NAND2_X1 U14256 ( .A1(n11170), .A2(n11169), .ZN(n13262) );
  INV_X1 U14257 ( .A(n11172), .ZN(n11173) );
  INV_X1 U14258 ( .A(n15214), .ZN(n15209) );
  AOI21_X1 U14259 ( .B1(n13984), .B2(n13553), .A(n9632), .ZN(n13529) );
  NAND2_X1 U14260 ( .A1(n13529), .A2(n16154), .ZN(n11175) );
  AND2_X1 U14261 ( .A1(n11176), .A2(n11175), .ZN(n11177) );
  OAI21_X1 U14262 ( .B1(n13531), .B2(n16152), .A(n11177), .ZN(P2_U3018) );
  AOI22_X1 U14263 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14264 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11180) );
  AOI22_X1 U14265 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11179) );
  INV_X2 U14266 ( .A(n11264), .ZN(n11194) );
  AOI22_X1 U14267 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11178) );
  NAND4_X1 U14268 ( .A1(n11181), .A2(n11180), .A3(n11179), .A4(n11178), .ZN(
        n11193) );
  INV_X2 U14269 ( .A(n11271), .ZN(n16864) );
  INV_X2 U14270 ( .A(n10095), .ZN(n16862) );
  AOI22_X1 U14271 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14272 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11190) );
  INV_X4 U14273 ( .A(n15484), .ZN(n16881) );
  AOI22_X1 U14274 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14275 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11188) );
  NAND4_X1 U14276 ( .A1(n11191), .A2(n11190), .A3(n11189), .A4(n11188), .ZN(
        n11192) );
  AOI22_X1 U14277 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14278 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14279 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14280 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11195) );
  NAND4_X1 U14281 ( .A1(n11198), .A2(n11197), .A3(n11196), .A4(n11195), .ZN(
        n11204) );
  AOI22_X1 U14282 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14283 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14284 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11200) );
  AOI22_X1 U14285 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11199) );
  NAND4_X1 U14286 ( .A1(n11202), .A2(n11201), .A3(n11200), .A4(n11199), .ZN(
        n11203) );
  INV_X2 U14287 ( .A(n16696), .ZN(n16943) );
  AOI22_X1 U14288 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14289 ( .A1(n11267), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14290 ( .A1(n11268), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11264), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11206) );
  INV_X2 U14291 ( .A(n10095), .ZN(n16927) );
  AOI22_X1 U14292 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11265), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11205) );
  NAND4_X1 U14293 ( .A1(n11208), .A2(n11207), .A3(n11206), .A4(n11205), .ZN(
        n11214) );
  INV_X1 U14294 ( .A(n11269), .ZN(n15484) );
  AOI22_X1 U14295 ( .A1(n11269), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11212) );
  INV_X2 U14296 ( .A(n11251), .ZN(n16950) );
  AOI22_X1 U14297 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14298 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14299 ( .A1(n11323), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11209) );
  NAND4_X1 U14300 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11213) );
  NOR2_X2 U14301 ( .A1(n11214), .A2(n11213), .ZN(n17137) );
  INV_X1 U14302 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n20711) );
  AOI22_X1 U14303 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11330), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n11216), .ZN(n11217) );
  OAI21_X1 U14304 ( .B1(n20711), .B2(n11251), .A(n11217), .ZN(n11223) );
  AOI22_X1 U14305 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11264), .B1(
        n16845), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14306 ( .A1(n11270), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n11268), .ZN(n11220) );
  AOI22_X1 U14307 ( .A1(n11241), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11265), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14308 ( .A1(n11267), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11271), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11218) );
  NAND4_X1 U14309 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11222) );
  AOI22_X1 U14310 ( .A1(n11269), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11224) );
  INV_X1 U14311 ( .A(n11224), .ZN(n11227) );
  AOI22_X1 U14312 ( .A1(n11323), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n16933), .ZN(n11225) );
  INV_X1 U14313 ( .A(n11225), .ZN(n11226) );
  AOI22_X1 U14314 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U14315 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11238) );
  AOI22_X1 U14316 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11230) );
  OAI21_X1 U14317 ( .B1(n15484), .B2(n20729), .A(n11230), .ZN(n11236) );
  AOI22_X1 U14318 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14319 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U14320 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11232) );
  AOI22_X1 U14321 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11231) );
  NAND4_X1 U14322 ( .A1(n11234), .A2(n11233), .A3(n11232), .A4(n11231), .ZN(
        n11235) );
  AOI211_X1 U14323 ( .C1(n16899), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n11236), .B(n11235), .ZN(n11237) );
  NAND3_X1 U14324 ( .A1(n11239), .A2(n11238), .A3(n11237), .ZN(n17131) );
  NAND2_X1 U14325 ( .A1(n11450), .A2(n17131), .ZN(n11287) );
  AOI22_X1 U14326 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14327 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14328 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11240) );
  OAI21_X1 U14329 ( .B1(n11194), .B2(n20785), .A(n11240), .ZN(n11247) );
  AOI22_X1 U14330 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14331 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14332 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14333 ( .A1(n11268), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11242) );
  NAND4_X1 U14334 ( .A1(n11245), .A2(n11244), .A3(n11243), .A4(n11242), .ZN(
        n11246) );
  AOI211_X1 U14335 ( .C1(n9574), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n11247), .B(n11246), .ZN(n11248) );
  NAND3_X1 U14336 ( .A1(n11250), .A2(n11249), .A3(n11248), .ZN(n17124) );
  AOI22_X1 U14337 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14338 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11260) );
  BUF_X4 U14339 ( .A(n11268), .Z(n16951) );
  AOI22_X1 U14340 ( .A1(n15502), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11252) );
  OAI21_X1 U14341 ( .B1(n11194), .B2(n16966), .A(n11252), .ZN(n11258) );
  AOI22_X1 U14342 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14343 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14344 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14345 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11253) );
  NAND4_X1 U14346 ( .A1(n11256), .A2(n11255), .A3(n11254), .A4(n11253), .ZN(
        n11257) );
  AOI211_X1 U14347 ( .C1(n16951), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n11258), .B(n11257), .ZN(n11259) );
  OAI21_X1 U14348 ( .B1(n11262), .B2(n12137), .A(n17528), .ZN(n11293) );
  XNOR2_X1 U14349 ( .A(n17124), .B(n11263), .ZN(n17566) );
  INV_X1 U14350 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11501) );
  XNOR2_X1 U14351 ( .A(n11501), .B(n11282), .ZN(n17605) );
  INV_X1 U14352 ( .A(n17605), .ZN(n11284) );
  AOI22_X1 U14353 ( .A1(n11330), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11265), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11266) );
  OAI21_X1 U14354 ( .B1(n11194), .B2(n15452), .A(n11266), .ZN(n11277) );
  AOI22_X1 U14355 ( .A1(n11267), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11268), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U14356 ( .A1(n11270), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11269), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14357 ( .A1(n16845), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14358 ( .A1(n11323), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11271), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11272) );
  NAND4_X1 U14359 ( .A1(n11275), .A2(n11274), .A3(n11273), .A4(n11272), .ZN(
        n11276) );
  AOI211_X1 U14360 ( .C1(n11215), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n11277), .B(n11276), .ZN(n11280) );
  AOI22_X1 U14361 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U14362 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11278) );
  NAND3_X1 U14363 ( .A1(n11280), .A2(n11279), .A3(n11278), .ZN(n15617) );
  NAND2_X1 U14364 ( .A1(n15617), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17620) );
  NOR2_X1 U14365 ( .A1(n11452), .A2(n17620), .ZN(n17613) );
  INV_X1 U14366 ( .A(n17604), .ZN(n11283) );
  AOI21_X2 U14367 ( .B1(n11284), .B2(n11283), .A(n10079), .ZN(n11285) );
  NOR2_X1 U14368 ( .A1(n11285), .A2(n17897), .ZN(n11286) );
  XNOR2_X1 U14369 ( .A(n17131), .B(n11450), .ZN(n17592) );
  XNOR2_X1 U14370 ( .A(n11285), .B(n17897), .ZN(n17591) );
  NOR2_X1 U14371 ( .A1(n17592), .A2(n17591), .ZN(n17590) );
  XNOR2_X1 U14372 ( .A(n17128), .B(n11287), .ZN(n17580) );
  NAND2_X1 U14373 ( .A1(n17566), .A2(n17564), .ZN(n11289) );
  AOI21_X1 U14374 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n11289), .A(
        n17565), .ZN(n17553) );
  XOR2_X1 U14375 ( .A(n17121), .B(n11290), .Z(n11291) );
  XNOR2_X1 U14376 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n11291), .ZN(
        n17552) );
  NOR2_X1 U14377 ( .A1(n17553), .A2(n17552), .ZN(n17551) );
  NOR2_X2 U14378 ( .A1(n17551), .A2(n11292), .ZN(n11294) );
  INV_X1 U14379 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17838) );
  INV_X1 U14380 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17455) );
  AND2_X1 U14381 ( .A1(n17492), .A2(n17455), .ZN(n11295) );
  NOR2_X1 U14382 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11296) );
  OR2_X1 U14383 ( .A1(n17541), .A2(n11297), .ZN(n11298) );
  NAND2_X1 U14384 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17827) );
  NOR2_X1 U14385 ( .A1(n17827), .A2(n17492), .ZN(n17810) );
  NAND2_X1 U14386 ( .A1(n17810), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17807) );
  INV_X1 U14387 ( .A(n17807), .ZN(n17781) );
  NAND3_X1 U14388 ( .A1(n17781), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17755) );
  INV_X1 U14389 ( .A(n17733), .ZN(n17410) );
  NOR2_X2 U14390 ( .A1(n17452), .A2(n17410), .ZN(n11302) );
  INV_X1 U14391 ( .A(n11302), .ZN(n11299) );
  INV_X1 U14392 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17423) );
  NOR3_X2 U14393 ( .A1(n11303), .A2(n11301), .A3(n11300), .ZN(n17406) );
  INV_X1 U14394 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17745) );
  NAND2_X1 U14395 ( .A1(n17406), .A2(n17745), .ZN(n17405) );
  INV_X1 U14396 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17672) );
  NAND2_X1 U14397 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17669) );
  INV_X1 U14398 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17695) );
  NOR2_X1 U14399 ( .A1(n17713), .A2(n17695), .ZN(n17708) );
  NAND3_X1 U14400 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17708), .ZN(n11306) );
  NOR2_X1 U14401 ( .A1(n17669), .A2(n11306), .ZN(n17693) );
  NAND2_X1 U14402 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17693), .ZN(
        n17664) );
  NOR2_X1 U14403 ( .A1(n17672), .A2(n17664), .ZN(n11474) );
  INV_X1 U14404 ( .A(n11474), .ZN(n17315) );
  NOR2_X1 U14405 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17454), .ZN(
        n17395) );
  NAND2_X1 U14406 ( .A1(n17395), .A2(n17713), .ZN(n11304) );
  NOR2_X1 U14407 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11304), .ZN(
        n17360) );
  INV_X1 U14408 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17352) );
  NAND2_X1 U14409 ( .A1(n17360), .A2(n17352), .ZN(n17339) );
  INV_X1 U14410 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n20760) );
  NAND2_X1 U14411 ( .A1(n17672), .A2(n20760), .ZN(n17682) );
  OAI22_X1 U14412 ( .A1(n17340), .A2(n17315), .B1(n17339), .B2(n17682), .ZN(
        n11305) );
  NOR2_X2 U14413 ( .A1(n17309), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17308) );
  NOR2_X1 U14414 ( .A1(n20760), .A2(n11306), .ZN(n17670) );
  INV_X1 U14415 ( .A(n17669), .ZN(n17737) );
  INV_X1 U14416 ( .A(n17340), .ZN(n17411) );
  NAND2_X1 U14417 ( .A1(n17737), .A2(n17411), .ZN(n17358) );
  NAND2_X1 U14418 ( .A1(n17670), .A2(n17359), .ZN(n17331) );
  INV_X1 U14419 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17653) );
  INV_X1 U14420 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17634) );
  NOR2_X1 U14421 ( .A1(n17653), .A2(n17634), .ZN(n11506) );
  INV_X1 U14422 ( .A(n11506), .ZN(n17630) );
  NOR2_X1 U14423 ( .A1(n16204), .A2(n10091), .ZN(n11312) );
  NAND2_X1 U14424 ( .A1(n11312), .A2(n17528), .ZN(n15597) );
  INV_X1 U14425 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16183) );
  NAND2_X1 U14426 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16183), .ZN(
        n11509) );
  OAI22_X1 U14427 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17528), .B1(
        n15597), .B2(n11509), .ZN(n11318) );
  NAND3_X1 U14428 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11507) );
  INV_X1 U14429 ( .A(n11507), .ZN(n16184) );
  NAND2_X1 U14430 ( .A1(n16184), .A2(n16207), .ZN(n15596) );
  INV_X1 U14431 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18552) );
  NAND2_X1 U14432 ( .A1(n18552), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11311) );
  OAI21_X1 U14433 ( .B1(n11312), .B2(n17454), .A(n10076), .ZN(n11316) );
  AOI21_X1 U14434 ( .B1(n17454), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n18552), .ZN(n11314) );
  AND2_X1 U14435 ( .A1(n11316), .A2(n11315), .ZN(n11317) );
  AOI22_X1 U14436 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11322) );
  AOI22_X1 U14437 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14438 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14439 ( .A1(n11393), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11319) );
  NAND4_X1 U14440 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(
        n11329) );
  AOI22_X1 U14441 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14442 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14443 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14444 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11324) );
  NAND4_X1 U14445 ( .A1(n11327), .A2(n11326), .A3(n11325), .A4(n11324), .ZN(
        n11328) );
  AOI22_X1 U14446 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14447 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11339) );
  INV_X1 U14448 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U14449 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11331) );
  OAI21_X1 U14450 ( .B1(n11392), .B2(n16985), .A(n11331), .ZN(n11337) );
  AOI22_X1 U14451 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14452 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14453 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14454 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11332) );
  NAND4_X1 U14455 ( .A1(n11335), .A2(n11334), .A3(n11333), .A4(n11332), .ZN(
        n11336) );
  NOR2_X1 U14456 ( .A1(n17192), .A2(n17969), .ZN(n11428) );
  AOI22_X1 U14457 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14458 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14459 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11341) );
  OAI21_X1 U14460 ( .B1(n11194), .B2(n20819), .A(n11341), .ZN(n11347) );
  AOI22_X1 U14461 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14462 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14463 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14464 ( .A1(n16862), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11393), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11342) );
  NAND4_X1 U14465 ( .A1(n11345), .A2(n11344), .A3(n11343), .A4(n11342), .ZN(
        n11346) );
  NAND2_X1 U14466 ( .A1(n11428), .A2(n17985), .ZN(n11443) );
  AOI22_X1 U14467 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14468 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14469 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14470 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11350) );
  NAND4_X1 U14471 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n11359) );
  AOI22_X1 U14472 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14473 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14474 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14475 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11354) );
  NAND4_X1 U14476 ( .A1(n11357), .A2(n11356), .A3(n11355), .A4(n11354), .ZN(
        n11358) );
  AOI22_X1 U14477 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14478 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11393), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14479 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11360) );
  OAI21_X1 U14480 ( .B1(n11392), .B2(n20785), .A(n11360), .ZN(n11366) );
  AOI22_X1 U14481 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14482 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14483 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14484 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11361) );
  NAND4_X1 U14485 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11365) );
  NAND2_X1 U14486 ( .A1(n11390), .A2(n17981), .ZN(n18399) );
  AOI22_X1 U14487 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11393), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11370) );
  OAI21_X1 U14488 ( .B1(n11392), .B2(n16966), .A(n11370), .ZN(n11376) );
  AOI22_X1 U14489 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14490 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14491 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14492 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11371) );
  NAND4_X1 U14493 ( .A1(n11374), .A2(n11373), .A3(n11372), .A4(n11371), .ZN(
        n11375) );
  AOI22_X1 U14494 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14495 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14496 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11380) );
  OAI21_X1 U14497 ( .B1(n10095), .B2(n20729), .A(n11380), .ZN(n11386) );
  AOI22_X1 U14498 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14499 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14500 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14501 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11381) );
  NAND4_X1 U14502 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .ZN(
        n11385) );
  AOI211_X1 U14503 ( .C1(n9574), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n11386), .B(n11385), .ZN(n11387) );
  NAND3_X1 U14504 ( .A1(n11389), .A2(n11388), .A3(n11387), .ZN(n17973) );
  AOI22_X1 U14505 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14506 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14507 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11391) );
  OAI21_X1 U14508 ( .B1(n11392), .B2(n15452), .A(n11391), .ZN(n11399) );
  AOI22_X1 U14509 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14510 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14511 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11393), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14512 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11394) );
  NAND4_X1 U14513 ( .A1(n11397), .A2(n11396), .A3(n11395), .A4(n11394), .ZN(
        n11398) );
  AOI211_X1 U14514 ( .C1(n16899), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n11399), .B(n11398), .ZN(n11400) );
  INV_X1 U14515 ( .A(n17969), .ZN(n11429) );
  NAND2_X1 U14516 ( .A1(n11488), .A2(n11429), .ZN(n11434) );
  NOR2_X1 U14517 ( .A1(n11485), .A2(n11434), .ZN(n11403) );
  OAI211_X1 U14518 ( .C1(n11435), .C2(n15616), .A(n11497), .B(n11403), .ZN(
        n11430) );
  INV_X1 U14519 ( .A(n18427), .ZN(n18590) );
  OAI21_X1 U14520 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18404), .A(
        n11410), .ZN(n11421) );
  INV_X1 U14521 ( .A(n11421), .ZN(n11419) );
  INV_X1 U14522 ( .A(n11420), .ZN(n11411) );
  INV_X1 U14523 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18426) );
  NOR2_X1 U14524 ( .A1(n11420), .A2(n11410), .ZN(n11404) );
  OAI22_X1 U14525 ( .A1(n18560), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n20820), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11412) );
  NOR2_X1 U14526 ( .A1(n11413), .A2(n11412), .ZN(n11405) );
  OAI21_X1 U14527 ( .B1(n18425), .B2(n11415), .A(n11416), .ZN(n11407) );
  INV_X1 U14528 ( .A(n11407), .ZN(n11408) );
  NAND2_X1 U14529 ( .A1(n11411), .A2(n11410), .ZN(n11409) );
  XNOR2_X1 U14530 ( .A(n11413), .B(n11412), .ZN(n11418) );
  NAND2_X1 U14531 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15525), .ZN(
        n11414) );
  OAI21_X1 U14532 ( .B1(n11419), .B2(n11425), .A(n11426), .ZN(n18589) );
  INV_X1 U14533 ( .A(n18589), .ZN(n11445) );
  NOR2_X1 U14534 ( .A1(n11421), .A2(n11420), .ZN(n11424) );
  INV_X1 U14535 ( .A(n11422), .ZN(n11423) );
  INV_X1 U14536 ( .A(n18430), .ZN(n16312) );
  NAND2_X2 U14537 ( .A1(n18532), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18537) );
  OAI211_X1 U14538 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18475), .B(n18537), .ZN(n18468) );
  OAI21_X1 U14539 ( .B1(n11429), .B2(n18598), .A(n18468), .ZN(n11427) );
  OAI21_X1 U14540 ( .B1(n11428), .B2(n11427), .A(n18608), .ZN(n16310) );
  NOR3_X1 U14541 ( .A1(n11477), .A2(n16312), .A3(n16310), .ZN(n11442) );
  NOR2_X1 U14542 ( .A1(n17144), .A2(n17960), .ZN(n11431) );
  NOR2_X1 U14543 ( .A1(n11390), .A2(n11479), .ZN(n11437) );
  NAND4_X1 U14544 ( .A1(n11435), .A2(n11484), .A3(n11431), .A4(n11437), .ZN(
        n18414) );
  INV_X1 U14545 ( .A(n11430), .ZN(n11441) );
  INV_X1 U14546 ( .A(n11431), .ZN(n11439) );
  NOR2_X1 U14547 ( .A1(n17144), .A2(n11437), .ZN(n11433) );
  NOR2_X1 U14548 ( .A1(n11435), .A2(n17985), .ZN(n18390) );
  INV_X1 U14549 ( .A(n11478), .ZN(n11432) );
  OAI22_X1 U14550 ( .A1(n11435), .A2(n11433), .B1(n17960), .B2(n11432), .ZN(
        n11486) );
  INV_X1 U14551 ( .A(n11434), .ZN(n11436) );
  INV_X1 U14552 ( .A(n11435), .ZN(n17976) );
  OAI22_X1 U14553 ( .A1(n11437), .A2(n11436), .B1(n17976), .B2(n18399), .ZN(
        n11438) );
  AOI211_X1 U14554 ( .C1(n11484), .C2(n11439), .A(n11486), .B(n11438), .ZN(
        n11481) );
  NAND2_X1 U14555 ( .A1(n17192), .A2(n17960), .ZN(n11491) );
  INV_X1 U14556 ( .A(n11491), .ZN(n11440) );
  NAND2_X1 U14557 ( .A1(n17991), .A2(n18399), .ZN(n15615) );
  NAND2_X1 U14558 ( .A1(n11440), .A2(n15615), .ZN(n11482) );
  OAI211_X1 U14559 ( .C1(n11487), .C2(n11441), .A(n11481), .B(n11482), .ZN(
        n15515) );
  AOI211_X1 U14560 ( .C1(n11477), .C2(n18591), .A(n11442), .B(n15515), .ZN(
        n11444) );
  NAND2_X1 U14561 ( .A1(n12132), .A2(n17850), .ZN(n11517) );
  INV_X1 U14562 ( .A(n11451), .ZN(n17145) );
  NAND2_X1 U14563 ( .A1(n15617), .A2(n17145), .ZN(n11454) );
  NAND2_X1 U14564 ( .A1(n17137), .A2(n11454), .ZN(n11448) );
  NAND2_X1 U14565 ( .A1(n11448), .A2(n17131), .ZN(n11459) );
  NOR2_X1 U14566 ( .A1(n17128), .A2(n11459), .ZN(n11446) );
  NAND2_X1 U14567 ( .A1(n11446), .A2(n17124), .ZN(n11462) );
  NOR2_X1 U14568 ( .A1(n17121), .A2(n11462), .ZN(n11466) );
  NAND2_X1 U14569 ( .A1(n11466), .A2(n12137), .ZN(n11467) );
  XOR2_X1 U14570 ( .A(n11446), .B(n17124), .Z(n11447) );
  AND2_X1 U14571 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11447), .ZN(
        n11461) );
  XNOR2_X1 U14572 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11447), .ZN(
        n17563) );
  XOR2_X1 U14573 ( .A(n17131), .B(n11448), .Z(n11457) );
  AND2_X1 U14574 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11457), .ZN(
        n11458) );
  INV_X1 U14575 ( .A(n11448), .ZN(n11449) );
  AOI21_X1 U14576 ( .B1(n11450), .B2(n15617), .A(n11449), .ZN(n11455) );
  NOR2_X1 U14577 ( .A1(n11455), .A2(n11501), .ZN(n11456) );
  INV_X1 U14578 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20679) );
  NAND2_X1 U14579 ( .A1(n11451), .A2(n20679), .ZN(n11453) );
  NOR2_X1 U14580 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15617), .ZN(
        n17622) );
  NAND2_X1 U14581 ( .A1(n17622), .A2(n11452), .ZN(n17611) );
  NAND3_X1 U14582 ( .A1(n11454), .A2(n11453), .A3(n17611), .ZN(n17603) );
  XNOR2_X1 U14583 ( .A(n11501), .B(n11455), .ZN(n17602) );
  NOR2_X1 U14584 ( .A1(n17603), .A2(n17602), .ZN(n17601) );
  NOR2_X1 U14585 ( .A1(n11456), .A2(n17601), .ZN(n17595) );
  XNOR2_X1 U14586 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11457), .ZN(
        n17594) );
  NOR2_X1 U14587 ( .A1(n17595), .A2(n17594), .ZN(n17593) );
  NOR2_X1 U14588 ( .A1(n11458), .A2(n17593), .ZN(n17574) );
  XNOR2_X1 U14589 ( .A(n11459), .B(n17128), .ZN(n17575) );
  NOR2_X1 U14590 ( .A1(n17574), .A2(n17575), .ZN(n11460) );
  NAND2_X1 U14591 ( .A1(n17574), .A2(n17575), .ZN(n17573) );
  OAI21_X1 U14592 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n11460), .A(
        n17573), .ZN(n17562) );
  NOR2_X1 U14593 ( .A1(n17563), .A2(n17562), .ZN(n17561) );
  NOR2_X1 U14594 ( .A1(n11461), .A2(n17561), .ZN(n11463) );
  XNOR2_X1 U14595 ( .A(n11462), .B(n17121), .ZN(n11464) );
  NOR2_X1 U14596 ( .A1(n11463), .A2(n11464), .ZN(n11465) );
  INV_X1 U14597 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17858) );
  XNOR2_X1 U14598 ( .A(n11464), .B(n11463), .ZN(n17549) );
  NOR2_X1 U14599 ( .A1(n17858), .A2(n17549), .ZN(n17548) );
  NOR2_X1 U14600 ( .A1(n11465), .A2(n17548), .ZN(n11468) );
  XNOR2_X1 U14601 ( .A(n11466), .B(n12137), .ZN(n11469) );
  NAND2_X1 U14602 ( .A1(n11468), .A2(n11469), .ZN(n17536) );
  NAND2_X1 U14603 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17536), .ZN(
        n11471) );
  NOR2_X1 U14604 ( .A1(n11467), .A2(n11471), .ZN(n11473) );
  INV_X1 U14605 ( .A(n11467), .ZN(n11472) );
  OR2_X1 U14606 ( .A1(n11469), .A2(n11468), .ZN(n17537) );
  OAI21_X1 U14607 ( .B1(n11472), .B2(n11471), .A(n17537), .ZN(n11470) );
  AOI21_X1 U14608 ( .B1(n11472), .B2(n11471), .A(n11470), .ZN(n17526) );
  INV_X1 U14609 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17862) );
  NAND3_X1 U14610 ( .A1(n17800), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17440) );
  NAND2_X1 U14611 ( .A1(n17688), .A2(n11474), .ZN(n17668) );
  INV_X1 U14612 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17673) );
  NAND2_X1 U14613 ( .A1(n17299), .A2(n11506), .ZN(n17260) );
  NAND2_X1 U14614 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11475) );
  NOR2_X1 U14615 ( .A1(n17260), .A2(n11475), .ZN(n16189) );
  INV_X1 U14616 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16191) );
  NOR3_X1 U14617 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16191), .A3(
        n16183), .ZN(n11499) );
  NOR2_X1 U14618 ( .A1(n17260), .A2(n11507), .ZN(n16190) );
  NAND2_X1 U14619 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16190), .ZN(
        n11476) );
  AOI22_X1 U14620 ( .A1(n16189), .A2(n11499), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11476), .ZN(n12139) );
  NAND2_X1 U14621 ( .A1(n11491), .A2(n11488), .ZN(n18615) );
  OR2_X1 U14622 ( .A1(n11478), .A2(n11477), .ZN(n11483) );
  NAND2_X1 U14623 ( .A1(n18390), .A2(n11480), .ZN(n15519) );
  OAI211_X1 U14624 ( .C1(n11484), .C2(n11483), .A(n11482), .B(n11481), .ZN(
        n11494) );
  NOR2_X1 U14625 ( .A1(n18414), .A2(n11494), .ZN(n18394) );
  NOR2_X1 U14626 ( .A1(n17969), .A2(n17973), .ZN(n18389) );
  NAND2_X1 U14627 ( .A1(n11485), .A2(n18389), .ZN(n15416) );
  NAND2_X1 U14628 ( .A1(n17192), .A2(n12179), .ZN(n15612) );
  NAND2_X1 U14629 ( .A1(n17189), .A2(n15522), .ZN(n15611) );
  NAND2_X1 U14630 ( .A1(n18598), .A2(n18415), .ZN(n11496) );
  INV_X1 U14631 ( .A(n11494), .ZN(n11495) );
  OAI21_X1 U14632 ( .B1(n11497), .B2(n11496), .A(n11495), .ZN(n18388) );
  NAND2_X1 U14633 ( .A1(n18439), .A2(n9564), .ZN(n17939) );
  OR2_X1 U14634 ( .A1(n12139), .A2(n17939), .ZN(n11515) );
  NAND2_X1 U14635 ( .A1(n17866), .A2(n17528), .ZN(n17527) );
  NAND2_X1 U14636 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17665), .ZN(
        n17298) );
  NAND3_X1 U14637 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n17637), .ZN(n16211) );
  INV_X1 U14638 ( .A(n11499), .ZN(n11510) );
  NAND2_X1 U14639 ( .A1(n16184), .A2(n17637), .ZN(n15535) );
  OAI21_X1 U14640 ( .B1(n16183), .B2(n15535), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11500) );
  OAI21_X1 U14641 ( .B1(n16211), .B2(n11510), .A(n11500), .ZN(n12138) );
  NAND2_X1 U14642 ( .A1(n18427), .A2(n17118), .ZN(n17823) );
  NOR2_X1 U14643 ( .A1(n9563), .A2(n17823), .ZN(n17865) );
  NOR2_X1 U14644 ( .A1(n11501), .A2(n20679), .ZN(n17730) );
  INV_X1 U14645 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17890) );
  NOR3_X1 U14646 ( .A1(n17890), .A2(n17897), .A3(n11288), .ZN(n17871) );
  NAND2_X1 U14647 ( .A1(n17730), .A2(n17871), .ZN(n17856) );
  NAND2_X1 U14648 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17855) );
  NOR2_X1 U14649 ( .A1(n17856), .A2(n17855), .ZN(n17843) );
  NAND2_X1 U14650 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17843), .ZN(
        n17783) );
  NOR2_X1 U14651 ( .A1(n17410), .A2(n17783), .ZN(n17689) );
  NOR2_X1 U14652 ( .A1(n17315), .A2(n17673), .ZN(n11502) );
  NAND2_X1 U14653 ( .A1(n17689), .A2(n11502), .ZN(n17631) );
  INV_X1 U14654 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17638) );
  INV_X1 U14655 ( .A(n11502), .ZN(n17652) );
  NOR3_X1 U14656 ( .A1(n17630), .A2(n17638), .A3(n17652), .ZN(n16203) );
  INV_X1 U14657 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18572) );
  NOR2_X1 U14658 ( .A1(n18572), .A2(n17783), .ZN(n17819) );
  INV_X1 U14659 ( .A(n17819), .ZN(n17842) );
  NOR2_X1 U14660 ( .A1(n17410), .A2(n17842), .ZN(n17753) );
  AOI21_X1 U14661 ( .B1(n16203), .B2(n17753), .A(n9569), .ZN(n11503) );
  AOI21_X1 U14662 ( .B1(n18403), .B2(n17631), .A(n11503), .ZN(n11505) );
  AOI21_X1 U14663 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17913) );
  INV_X1 U14664 ( .A(n17855), .ZN(n11504) );
  NAND3_X1 U14665 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17871), .A3(
        n11504), .ZN(n17731) );
  NOR2_X1 U14666 ( .A1(n17913), .A2(n17731), .ZN(n17780) );
  NAND2_X1 U14667 ( .A1(n17733), .A2(n17780), .ZN(n17692) );
  OAI21_X1 U14668 ( .B1(n17692), .B2(n17652), .A(n18411), .ZN(n17632) );
  OAI211_X1 U14669 ( .C1(n17836), .C2(n11506), .A(n11505), .B(n17632), .ZN(
        n15537) );
  AOI21_X1 U14670 ( .B1(n17859), .B2(n11507), .A(n15537), .ZN(n11508) );
  NAND2_X1 U14671 ( .A1(n18553), .A2(n18543), .ZN(n18556) );
  NOR2_X1 U14672 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18556), .ZN(n18617) );
  NAND2_X2 U14673 ( .A1(n18617), .A2(n18603), .ZN(n17852) );
  AOI21_X1 U14674 ( .B1(n9564), .B2(n11508), .A(n9578), .ZN(n15601) );
  INV_X1 U14675 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18534) );
  NOR2_X1 U14676 ( .A1(n18534), .A2(n17852), .ZN(n12136) );
  INV_X1 U14677 ( .A(n9569), .ZN(n18395) );
  AOI21_X1 U14678 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18395), .A(
        n18403), .ZN(n17914) );
  INV_X1 U14679 ( .A(n17689), .ZN(n17734) );
  OAI22_X1 U14680 ( .A1(n18429), .A2(n17692), .B1(n17914), .B2(n17734), .ZN(
        n17651) );
  NAND4_X1 U14681 ( .A1(n9564), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16203), .A4(n17651), .ZN(n15533) );
  NAND2_X1 U14682 ( .A1(n9564), .A2(n17859), .ZN(n17929) );
  OAI22_X1 U14683 ( .A1(n11510), .A2(n15533), .B1(n11509), .B2(n17929), .ZN(
        n11511) );
  AOI211_X1 U14684 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n15601), .A(
        n12136), .B(n11511), .ZN(n11512) );
  INV_X1 U14685 ( .A(n11512), .ZN(n11513) );
  NOR2_X1 U14686 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11906) );
  INV_X1 U14687 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11518) );
  AND2_X2 U14688 ( .A1(n11518), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11528) );
  INV_X1 U14689 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11519) );
  AND2_X2 U14690 ( .A1(n11528), .A2(n11527), .ZN(n11575) );
  AOI22_X1 U14691 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11709), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11524) );
  INV_X1 U14692 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14693 ( .A1(n13682), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11574), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11523) );
  AND2_X2 U14694 ( .A1(n12813), .A2(n11525), .ZN(n11716) );
  AOI22_X1 U14695 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11522) );
  AND2_X2 U14696 ( .A1(n11527), .A2(n11529), .ZN(n11581) );
  AND2_X2 U14697 ( .A1(n12813), .A2(n11529), .ZN(n11597) );
  AOI22_X1 U14698 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11521) );
  NAND4_X1 U14699 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11535) );
  AND2_X2 U14700 ( .A1(n11526), .A2(n11528), .ZN(n11710) );
  AOI22_X1 U14701 ( .A1(n11826), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11532) );
  AND2_X2 U14702 ( .A1(n11529), .A2(n14844), .ZN(n11602) );
  AOI22_X1 U14703 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14704 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11582), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U14705 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11534) );
  OR2_X2 U14706 ( .A1(n11535), .A2(n11534), .ZN(n11974) );
  AOI22_X1 U14707 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11709), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14708 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14709 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13682), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14710 ( .A1(n11574), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14711 ( .A1(n11826), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14712 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11542) );
  BUF_X4 U14713 ( .A(n11582), .Z(n13932) );
  AOI22_X1 U14714 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14715 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11540) );
  NAND2_X1 U14716 ( .A1(n12003), .A2(n19994), .ZN(n11979) );
  NAND2_X1 U14717 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11548) );
  NAND2_X1 U14718 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14719 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11546) );
  NAND2_X1 U14720 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11545) );
  NAND2_X1 U14721 ( .A1(n13682), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11552) );
  NAND2_X1 U14722 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11551) );
  NAND2_X1 U14723 ( .A1(n11574), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11550) );
  NAND2_X1 U14724 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11549) );
  NAND2_X1 U14725 ( .A1(n11826), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11556) );
  NAND2_X1 U14726 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11555) );
  NAND2_X1 U14727 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11554) );
  NAND2_X1 U14728 ( .A1(n11716), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11553) );
  NAND2_X1 U14729 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11560) );
  NAND2_X1 U14730 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11559) );
  NAND2_X1 U14731 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11558) );
  NAND2_X1 U14732 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11557) );
  NOR2_X1 U14733 ( .A1(n11979), .A2(n14532), .ZN(n11611) );
  AOI22_X1 U14734 ( .A1(n11574), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14735 ( .A1(n11716), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14736 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11582), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14737 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11709), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14738 ( .A1(n11826), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14739 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11572) );
  NAND3_X2 U14740 ( .A1(n11573), .A2(n10097), .A3(n11572), .ZN(n11655) );
  AOI22_X1 U14741 ( .A1(n11826), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14742 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11574), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14743 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11709), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14744 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14745 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14746 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14747 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11582), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11583) );
  NAND2_X1 U14748 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11591) );
  NAND2_X1 U14749 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11590) );
  NAND2_X1 U14750 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11589) );
  NAND2_X1 U14751 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11588) );
  INV_X1 U14752 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11592) );
  NAND2_X1 U14753 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11595) );
  NAND2_X1 U14754 ( .A1(n11574), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11594) );
  NAND2_X1 U14755 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11593) );
  NAND2_X1 U14756 ( .A1(n11826), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U14757 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U14758 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11599) );
  NAND2_X1 U14759 ( .A1(n11716), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11598) );
  NAND2_X1 U14760 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U14761 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14762 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11604) );
  NAND2_X1 U14763 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11603) );
  NAND2_X1 U14764 ( .A1(n11611), .A2(n12381), .ZN(n11988) );
  INV_X1 U14765 ( .A(n11988), .ZN(n11633) );
  NAND2_X1 U14766 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11616) );
  NAND2_X1 U14767 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11615) );
  NAND2_X1 U14768 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11614) );
  NAND2_X1 U14769 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11613) );
  NAND2_X1 U14770 ( .A1(n13682), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11620) );
  NAND2_X1 U14771 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11619) );
  NAND2_X1 U14772 ( .A1(n11574), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11618) );
  NAND2_X1 U14773 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11617) );
  NAND2_X1 U14774 ( .A1(n11826), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11624) );
  NAND2_X1 U14775 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11623) );
  NAND2_X1 U14776 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11622) );
  NAND2_X1 U14777 ( .A1(n11716), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11621) );
  NAND2_X1 U14778 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11628) );
  NAND2_X1 U14779 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11627) );
  NAND2_X1 U14780 ( .A1(n13932), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11626) );
  NAND2_X1 U14781 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11625) );
  NAND4_X4 U14782 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n19972) );
  NAND2_X1 U14783 ( .A1(n11709), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11637) );
  NAND2_X1 U14784 ( .A1(n11576), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11636) );
  NAND2_X1 U14785 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11635) );
  NAND2_X1 U14786 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11634) );
  NAND2_X1 U14787 ( .A1(n11826), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11641) );
  NAND2_X1 U14788 ( .A1(n11574), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11640) );
  NAND2_X1 U14789 ( .A1(n11716), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11638) );
  NAND2_X1 U14790 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11645) );
  NAND2_X1 U14791 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11644) );
  NAND2_X1 U14792 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11643) );
  NAND2_X1 U14793 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11642) );
  NAND2_X1 U14794 ( .A1(n11806), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11649) );
  NAND2_X1 U14795 ( .A1(n11695), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11648) );
  NAND2_X1 U14796 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11647) );
  NAND2_X1 U14797 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11646) );
  NAND2_X1 U14798 ( .A1(n11659), .A2(n19985), .ZN(n12479) );
  NAND2_X1 U14799 ( .A1(n11675), .A2(n11767), .ZN(n11673) );
  INV_X1 U14800 ( .A(n11673), .ZN(n11654) );
  NAND2_X1 U14801 ( .A1(n11667), .A2(n19994), .ZN(n11658) );
  NAND2_X1 U14802 ( .A1(n12003), .A2(n11767), .ZN(n11781) );
  NAND2_X1 U14803 ( .A1(n11781), .A2(n12494), .ZN(n11656) );
  NAND2_X1 U14804 ( .A1(n10099), .A2(n11675), .ZN(n11964) );
  NAND2_X1 U14805 ( .A1(n11656), .A2(n11964), .ZN(n11657) );
  NAND2_X1 U14806 ( .A1(n11658), .A2(n11657), .ZN(n11664) );
  NAND2_X2 U14807 ( .A1(n12482), .A2(n11767), .ZN(n12246) );
  NAND2_X1 U14808 ( .A1(n20592), .A2(n19698), .ZN(n20577) );
  NAND2_X1 U14809 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_1__SCAN_IN), 
        .ZN(n11660) );
  NOR2_X2 U14810 ( .A1(n11974), .A2(n19994), .ZN(n12801) );
  NAND3_X1 U14811 ( .A1(n12801), .A2(n12477), .A3(n11937), .ZN(n12772) );
  AND2_X1 U14812 ( .A1(n12246), .A2(n11974), .ZN(n11663) );
  NAND2_X1 U14813 ( .A1(n11974), .A2(n19972), .ZN(n11665) );
  NAND2_X1 U14814 ( .A1(n11937), .A2(n20015), .ZN(n12495) );
  NAND2_X1 U14815 ( .A1(n12495), .A2(n11990), .ZN(n12490) );
  NAND2_X1 U14816 ( .A1(n9646), .A2(n12490), .ZN(n11983) );
  AOI21_X1 U14817 ( .B1(n11983), .B2(n14061), .A(n12801), .ZN(n11668) );
  NAND2_X1 U14818 ( .A1(n19700), .A2(n20571), .ZN(n12248) );
  INV_X1 U14819 ( .A(n12248), .ZN(n11797) );
  NAND2_X1 U14820 ( .A1(n20507), .A2(n20428), .ZN(n20379) );
  NAND2_X1 U14821 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20503) );
  AOI21_X1 U14822 ( .B1(n11797), .B2(n20312), .A(n11681), .ZN(n11669) );
  INV_X1 U14823 ( .A(n11684), .ZN(n11670) );
  INV_X1 U14824 ( .A(n15584), .ZN(n15591) );
  MUX2_X1 U14825 ( .A(n15591), .B(n12248), .S(n20428), .Z(n11671) );
  INV_X1 U14826 ( .A(n12477), .ZN(n12923) );
  AND2_X1 U14827 ( .A1(n12923), .A2(n12025), .ZN(n12429) );
  NAND2_X1 U14828 ( .A1(n11999), .A2(n19994), .ZN(n11674) );
  NAND2_X1 U14829 ( .A1(n12481), .A2(n20015), .ZN(n11976) );
  AOI22_X1 U14830 ( .A1(n12429), .A2(n11674), .B1(n11976), .B2(n19826), .ZN(
        n11678) );
  NAND3_X1 U14831 ( .A1(n11983), .A2(n19985), .A3(n14061), .ZN(n11677) );
  AND2_X1 U14832 ( .A1(n19700), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11676) );
  NAND2_X1 U14833 ( .A1(n12801), .A2(n11675), .ZN(n12016) );
  NAND4_X1 U14834 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n12016), .ZN(
        n11679) );
  INV_X1 U14836 ( .A(n11707), .ZN(n11680) );
  NAND2_X1 U14837 ( .A1(n11708), .A2(n11680), .ZN(n11758) );
  INV_X1 U14838 ( .A(n11681), .ZN(n11682) );
  AND2_X1 U14839 ( .A1(n11682), .A2(n11520), .ZN(n11683) );
  AND2_X1 U14840 ( .A1(n15584), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11685) );
  XNOR2_X1 U14841 ( .A(n20503), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19980) );
  NAND2_X1 U14842 ( .A1(n11797), .A2(n19980), .ZN(n11687) );
  NAND2_X1 U14843 ( .A1(n11689), .A2(n11687), .ZN(n11686) );
  NAND4_X1 U14844 ( .A1(n11759), .A2(n11689), .A3(n11688), .A4(n11687), .ZN(
        n11690) );
  AOI22_X1 U14845 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14846 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14847 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11692) );
  INV_X1 U14848 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n20697) );
  AOI22_X1 U14849 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11691) );
  NAND4_X1 U14850 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11701) );
  AOI22_X1 U14851 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14852 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14853 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14854 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11696) );
  NAND4_X1 U14855 ( .A1(n11699), .A2(n11698), .A3(n11697), .A4(n11696), .ZN(
        n11700) );
  INV_X1 U14856 ( .A(n11801), .ZN(n11704) );
  AOI22_X1 U14857 ( .A1(n11704), .A2(n11703), .B1(n11958), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11705) );
  XNOR2_X1 U14858 ( .A(n11706), .B(n11705), .ZN(n11792) );
  INV_X1 U14859 ( .A(n11792), .ZN(n11766) );
  NAND2_X1 U14860 ( .A1(n12253), .A2(n20571), .ZN(n11736) );
  AOI22_X1 U14861 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14862 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14863 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11574), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14864 ( .A1(n13887), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11711) );
  NAND4_X1 U14865 ( .A1(n11714), .A2(n11713), .A3(n11712), .A4(n11711), .ZN(
        n11722) );
  AOI22_X1 U14866 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14867 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13889), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14868 ( .A1(n13879), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14869 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11717) );
  NAND4_X1 U14870 ( .A1(n11720), .A2(n11719), .A3(n11718), .A4(n11717), .ZN(
        n11721) );
  NOR2_X1 U14871 ( .A1(n11800), .A2(n11899), .ZN(n11751) );
  AOI22_X1 U14872 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14873 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14874 ( .A1(n13879), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14875 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11724) );
  NAND4_X1 U14876 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n11733) );
  AOI22_X1 U14877 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14878 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11574), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14879 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14880 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11728) );
  NAND4_X1 U14881 ( .A1(n11731), .A2(n11730), .A3(n11729), .A4(n11728), .ZN(
        n11732) );
  MUX2_X1 U14882 ( .A(n11740), .B(n11751), .S(n11780), .Z(n11734) );
  INV_X1 U14883 ( .A(n11734), .ZN(n11735) );
  INV_X1 U14884 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11739) );
  AOI21_X1 U14885 ( .B1(n12926), .B2(n11780), .A(n20571), .ZN(n11738) );
  NAND2_X1 U14886 ( .A1(n12482), .A2(n11899), .ZN(n11737) );
  OAI211_X1 U14887 ( .C1(n11954), .C2(n11739), .A(n11738), .B(n11737), .ZN(
        n11772) );
  INV_X1 U14888 ( .A(n11740), .ZN(n11895) );
  AOI22_X1 U14889 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14890 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14891 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14892 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11741) );
  NAND4_X1 U14893 ( .A1(n11744), .A2(n11743), .A3(n11742), .A4(n11741), .ZN(
        n11750) );
  AOI22_X1 U14894 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U14895 ( .A1(n13879), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U14896 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U14897 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11745) );
  NAND4_X1 U14898 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n11749) );
  INV_X1 U14899 ( .A(n11779), .ZN(n11754) );
  INV_X1 U14900 ( .A(n11751), .ZN(n11753) );
  NAND2_X1 U14901 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11752) );
  OAI211_X1 U14902 ( .C1(n11801), .C2(n11754), .A(n11753), .B(n11752), .ZN(
        n11755) );
  NAND2_X1 U14903 ( .A1(n11756), .A2(n11755), .ZN(n11757) );
  INV_X1 U14904 ( .A(n11800), .ZN(n11760) );
  NAND2_X1 U14905 ( .A1(n11760), .A2(n11779), .ZN(n11761) );
  INV_X1 U14906 ( .A(n12511), .ZN(n11762) );
  NAND2_X1 U14907 ( .A1(n11763), .A2(n11762), .ZN(n11765) );
  AND2_X2 U14908 ( .A1(n11765), .A2(n11764), .ZN(n11793) );
  INV_X1 U14909 ( .A(n11963), .ZN(n11893) );
  NAND2_X1 U14910 ( .A1(n12824), .A2(n11893), .ZN(n11771) );
  NAND2_X1 U14911 ( .A1(n11779), .A2(n11780), .ZN(n11818) );
  XNOR2_X1 U14912 ( .A(n11818), .B(n11817), .ZN(n11769) );
  NAND2_X1 U14913 ( .A1(n12926), .A2(n19994), .ZN(n11775) );
  INV_X1 U14914 ( .A(n11775), .ZN(n11768) );
  AOI21_X1 U14915 ( .B1(n11769), .B2(n19826), .A(n11768), .ZN(n11770) );
  NAND2_X1 U14916 ( .A1(n11771), .A2(n11770), .ZN(n12718) );
  INV_X1 U14917 ( .A(n11772), .ZN(n11773) );
  XNOR2_X1 U14918 ( .A(n11774), .B(n11773), .ZN(n12251) );
  NAND2_X1 U14919 ( .A1(n12251), .A2(n11893), .ZN(n11778) );
  OAI21_X1 U14920 ( .B1(n9590), .B2(n11780), .A(n11775), .ZN(n11776) );
  INV_X1 U14921 ( .A(n11776), .ZN(n11777) );
  OAI21_X1 U14922 ( .B1(n11780), .B2(n11779), .A(n11818), .ZN(n11783) );
  INV_X1 U14923 ( .A(n11781), .ZN(n11782) );
  OAI21_X1 U14924 ( .B1(n11783), .B2(n9590), .A(n11782), .ZN(n11784) );
  INV_X1 U14925 ( .A(n11784), .ZN(n11785) );
  NAND2_X1 U14926 ( .A1(n12889), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12891) );
  INV_X1 U14927 ( .A(n11786), .ZN(n11788) );
  NAND2_X1 U14928 ( .A1(n11788), .A2(n11787), .ZN(n11789) );
  NAND2_X1 U14929 ( .A1(n12891), .A2(n11789), .ZN(n11790) );
  INV_X1 U14930 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19961) );
  XNOR2_X1 U14931 ( .A(n11790), .B(n19961), .ZN(n12719) );
  NAND2_X1 U14932 ( .A1(n12718), .A2(n12719), .ZN(n12720) );
  NAND2_X1 U14933 ( .A1(n11790), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11791) );
  INV_X1 U14934 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19943) );
  NAND2_X1 U14935 ( .A1(n11793), .A2(n11792), .ZN(n11815) );
  NAND2_X1 U14936 ( .A1(n11794), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11799) );
  OAI21_X1 U14937 ( .B1(n20503), .B2(n20256), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11796) );
  INV_X1 U14938 ( .A(n20503), .ZN(n20091) );
  NAND2_X1 U14939 ( .A1(n20058), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20187) );
  INV_X1 U14940 ( .A(n20187), .ZN(n11795) );
  NAND2_X1 U14941 ( .A1(n20091), .A2(n11795), .ZN(n20224) );
  NAND2_X1 U14942 ( .A1(n11796), .A2(n20224), .ZN(n20257) );
  AOI22_X1 U14943 ( .A1(n11797), .A2(n20257), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15584), .ZN(n11798) );
  AOI22_X1 U14944 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U14945 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U14946 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14947 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11802) );
  NAND4_X1 U14948 ( .A1(n11805), .A2(n11804), .A3(n11803), .A4(n11802), .ZN(
        n11812) );
  AOI22_X1 U14949 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14950 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U14951 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U14952 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11807) );
  NAND4_X1 U14953 ( .A1(n11810), .A2(n11809), .A3(n11808), .A4(n11807), .ZN(
        n11811) );
  AOI22_X1 U14954 ( .A1(n11936), .A2(n11856), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n11958), .ZN(n11813) );
  AND2_X1 U14955 ( .A1(n11815), .A2(n12854), .ZN(n11816) );
  NAND2_X1 U14956 ( .A1(n11818), .A2(n11817), .ZN(n11858) );
  XNOR2_X1 U14957 ( .A(n11858), .B(n11856), .ZN(n11819) );
  OAI22_X1 U14958 ( .A1(n19969), .A2(n11963), .B1(n9590), .B2(n11819), .ZN(
        n12903) );
  NAND2_X1 U14959 ( .A1(n12904), .A2(n12903), .ZN(n12902) );
  NAND2_X1 U14960 ( .A1(n11820), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11821) );
  NAND2_X1 U14961 ( .A1(n12902), .A2(n11821), .ZN(n19904) );
  AOI22_X1 U14962 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14963 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14964 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13806), .B1(
        n13889), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14965 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n13932), .B1(
        n13881), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11822) );
  NAND4_X1 U14966 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n11832) );
  AOI22_X1 U14967 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13821), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14968 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13880), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14969 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n13887), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14970 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9594), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11827) );
  NAND4_X1 U14971 ( .A1(n11830), .A2(n11829), .A3(n11828), .A4(n11827), .ZN(
        n11831) );
  NAND2_X1 U14972 ( .A1(n11936), .A2(n11855), .ZN(n11834) );
  NAND2_X1 U14973 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11833) );
  XNOR2_X1 U14974 ( .A(n11841), .B(n9616), .ZN(n12951) );
  NAND2_X1 U14975 ( .A1(n12951), .A2(n11893), .ZN(n11838) );
  NAND2_X1 U14976 ( .A1(n11858), .A2(n11856), .ZN(n11835) );
  XNOR2_X1 U14977 ( .A(n11835), .B(n11855), .ZN(n11836) );
  NAND2_X1 U14978 ( .A1(n11836), .A2(n19826), .ZN(n11837) );
  NAND2_X1 U14979 ( .A1(n11838), .A2(n11837), .ZN(n11839) );
  INV_X1 U14980 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19933) );
  XNOR2_X1 U14981 ( .A(n11839), .B(n19933), .ZN(n19903) );
  NAND2_X1 U14982 ( .A1(n19904), .A2(n19903), .ZN(n19906) );
  NAND2_X1 U14983 ( .A1(n11839), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11840) );
  AOI22_X1 U14984 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U14985 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14986 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U14987 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11842) );
  NAND4_X1 U14988 ( .A1(n11845), .A2(n11844), .A3(n11843), .A4(n11842), .ZN(
        n11851) );
  AOI22_X1 U14989 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14990 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14991 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14992 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11846) );
  NAND4_X1 U14993 ( .A1(n11849), .A2(n11848), .A3(n11847), .A4(n11846), .ZN(
        n11850) );
  AOI22_X1 U14994 ( .A1(n11936), .A2(n11877), .B1(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n11958), .ZN(n11852) );
  NAND2_X1 U14995 ( .A1(n11853), .A2(n11852), .ZN(n11854) );
  NAND2_X1 U14996 ( .A1(n11876), .A2(n11854), .ZN(n13098) );
  OR2_X1 U14997 ( .A1(n13098), .A2(n11963), .ZN(n11862) );
  AND2_X1 U14998 ( .A1(n11856), .A2(n11855), .ZN(n11857) );
  AND2_X1 U14999 ( .A1(n11858), .A2(n11857), .ZN(n11878) );
  INV_X1 U15000 ( .A(n11877), .ZN(n11859) );
  XNOR2_X1 U15001 ( .A(n11878), .B(n11859), .ZN(n11860) );
  NAND2_X1 U15002 ( .A1(n11860), .A2(n19826), .ZN(n11861) );
  NAND2_X1 U15003 ( .A1(n11862), .A2(n11861), .ZN(n11863) );
  INV_X1 U15004 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13065) );
  XNOR2_X1 U15005 ( .A(n11863), .B(n13065), .ZN(n15784) );
  NAND2_X1 U15006 ( .A1(n11863), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11864) );
  AOI22_X1 U15007 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U15008 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11574), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U15009 ( .A1(n13879), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U15010 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11865) );
  NAND4_X1 U15011 ( .A1(n11868), .A2(n11867), .A3(n11866), .A4(n11865), .ZN(
        n11874) );
  AOI22_X1 U15012 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13821), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U15013 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U15014 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U15015 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11869) );
  NAND4_X1 U15016 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11873) );
  AOI22_X1 U15017 ( .A1(n11936), .A2(n11888), .B1(n11958), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U15018 ( .A1(n11876), .A2(n11875), .ZN(n13088) );
  NAND3_X1 U15019 ( .A1(n11897), .A2(n11893), .A3(n13088), .ZN(n11881) );
  NAND2_X1 U15020 ( .A1(n11878), .A2(n11877), .ZN(n11889) );
  XNOR2_X1 U15021 ( .A(n11888), .B(n11889), .ZN(n11879) );
  NAND2_X1 U15022 ( .A1(n19826), .A2(n11879), .ZN(n11880) );
  NAND2_X1 U15023 ( .A1(n13063), .A2(n15890), .ZN(n11882) );
  INV_X1 U15024 ( .A(n13063), .ZN(n11883) );
  NAND2_X1 U15025 ( .A1(n11883), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11884) );
  NAND2_X1 U15026 ( .A1(n11936), .A2(n11899), .ZN(n11886) );
  NAND2_X1 U15027 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11885) );
  NAND2_X1 U15028 ( .A1(n11886), .A2(n11885), .ZN(n11887) );
  XNOR2_X1 U15029 ( .A(n11897), .B(n11887), .ZN(n13220) );
  INV_X1 U15030 ( .A(n11888), .ZN(n11890) );
  NOR2_X1 U15031 ( .A1(n11890), .A2(n11889), .ZN(n11898) );
  XNOR2_X1 U15032 ( .A(n11899), .B(n11898), .ZN(n11891) );
  NOR2_X1 U15033 ( .A1(n11891), .A2(n9590), .ZN(n11892) );
  AOI21_X1 U15034 ( .B1(n13220), .B2(n11893), .A(n11892), .ZN(n11894) );
  INV_X1 U15035 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15901) );
  NOR2_X1 U15036 ( .A1(n11895), .A2(n11963), .ZN(n11896) );
  NAND2_X1 U15037 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  NOR2_X1 U15038 ( .A1(n9590), .A2(n11900), .ZN(n11901) );
  INV_X1 U15039 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11902) );
  NAND2_X1 U15040 ( .A1(n13331), .A2(n11902), .ZN(n11903) );
  INV_X1 U15041 ( .A(n13331), .ZN(n11904) );
  INV_X1 U15042 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11905) );
  NAND2_X1 U15043 ( .A1(n14777), .A2(n11905), .ZN(n13446) );
  NAND2_X1 U15044 ( .A1(n11906), .A2(n13481), .ZN(n11907) );
  NAND2_X1 U15045 ( .A1(n11907), .A2(n15769), .ZN(n11916) );
  NOR2_X1 U15046 ( .A1(n15769), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14683) );
  NAND2_X1 U15047 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11908) );
  NAND2_X1 U15048 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11909) );
  NAND2_X1 U15049 ( .A1(n14685), .A2(n11909), .ZN(n14809) );
  NOR2_X1 U15050 ( .A1(n15769), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14807) );
  XNOR2_X1 U15051 ( .A(n15769), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14812) );
  NOR2_X1 U15052 ( .A1(n14807), .A2(n14812), .ZN(n11910) );
  INV_X1 U15053 ( .A(n13481), .ZN(n11911) );
  NAND3_X1 U15054 ( .A1(n14671), .A2(n11911), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11915) );
  NAND2_X1 U15055 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14697) );
  INV_X1 U15056 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12057) );
  INV_X1 U15057 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U15058 ( .A1(n12057), .A2(n11912), .ZN(n11913) );
  NAND2_X1 U15059 ( .A1(n15769), .A2(n11913), .ZN(n14694) );
  NAND2_X1 U15060 ( .A1(n14697), .A2(n14694), .ZN(n13482) );
  NOR2_X1 U15061 ( .A1(n14809), .A2(n13482), .ZN(n11914) );
  INV_X1 U15062 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15834) );
  XNOR2_X1 U15063 ( .A(n15769), .B(n15834), .ZN(n14667) );
  NAND2_X1 U15064 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14787) );
  INV_X1 U15065 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20808) );
  NOR2_X1 U15066 ( .A1(n14787), .A2(n20808), .ZN(n12128) );
  NAND2_X1 U15067 ( .A1(n11917), .A2(n14777), .ZN(n15738) );
  INV_X1 U15068 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14798) );
  INV_X1 U15069 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14796) );
  NAND4_X1 U15070 ( .A1(n15834), .A2(n20808), .A3(n14798), .A4(n14796), .ZN(
        n11918) );
  NOR2_X1 U15071 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11919) );
  INV_X1 U15072 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15808) );
  NAND2_X1 U15073 ( .A1(n11919), .A2(n15808), .ZN(n14615) );
  NAND3_X1 U15074 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14614) );
  NAND2_X1 U15075 ( .A1(n11920), .A2(n14777), .ZN(n14641) );
  NAND2_X1 U15076 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14734) );
  INV_X1 U15077 ( .A(n14734), .ZN(n11921) );
  INV_X1 U15078 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14723) );
  NOR2_X1 U15079 ( .A1(n15769), .A2(n14723), .ZN(n13558) );
  INV_X1 U15080 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14750) );
  INV_X1 U15081 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14731) );
  NAND2_X1 U15082 ( .A1(n14750), .A2(n14731), .ZN(n14733) );
  NOR2_X1 U15083 ( .A1(n14777), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13559) );
  INV_X1 U15084 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14719) );
  XNOR2_X1 U15085 ( .A(n11922), .B(n12023), .ZN(n13960) );
  XNOR2_X1 U15086 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11935) );
  NAND2_X1 U15087 ( .A1(n20428), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U15088 ( .A1(n11935), .A2(n11934), .ZN(n11924) );
  NAND2_X1 U15089 ( .A1(n20507), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11923) );
  NOR2_X1 U15090 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19964), .ZN(
        n11925) );
  NAND2_X1 U15091 ( .A1(n11970), .A2(n11957), .ZN(n11962) );
  NAND2_X1 U15092 ( .A1(n11970), .A2(n11936), .ZN(n11961) );
  NAND3_X1 U15093 ( .A1(n15917), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n11926), .ZN(n11968) );
  AOI21_X1 U15094 ( .B1(n11929), .B2(n11928), .A(n11927), .ZN(n11930) );
  INV_X1 U15095 ( .A(n11930), .ZN(n11967) );
  NAND2_X1 U15096 ( .A1(n11937), .A2(n19972), .ZN(n11931) );
  NAND2_X1 U15097 ( .A1(n11931), .A2(n19827), .ZN(n11953) );
  XNOR2_X1 U15098 ( .A(n11933), .B(n11932), .ZN(n11966) );
  XNOR2_X1 U15099 ( .A(n11935), .B(n11934), .ZN(n11965) );
  INV_X1 U15100 ( .A(n11948), .ZN(n11938) );
  NOR2_X1 U15101 ( .A1(n11965), .A2(n11938), .ZN(n11943) );
  OAI21_X1 U15102 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20428), .A(
        n11939), .ZN(n11940) );
  INV_X1 U15103 ( .A(n11940), .ZN(n11941) );
  OAI211_X1 U15104 ( .C1(n12926), .C2(n12246), .A(n11953), .B(n11941), .ZN(
        n11942) );
  AND2_X1 U15105 ( .A1(n11943), .A2(n11945), .ZN(n11951) );
  OAI21_X1 U15106 ( .B1(n11952), .B2(n11966), .A(n11953), .ZN(n11944) );
  AOI21_X1 U15107 ( .B1(n11958), .B2(n11966), .A(n11944), .ZN(n11950) );
  INV_X1 U15108 ( .A(n11965), .ZN(n11947) );
  AOI211_X1 U15109 ( .C1(n11948), .C2(n19985), .A(n11947), .B(n11946), .ZN(
        n11949) );
  OAI33_X1 U15110 ( .A1(n11953), .A2(n11952), .A3(n11966), .B1(n11951), .B2(
        n11950), .B3(n11949), .ZN(n11956) );
  NAND2_X1 U15111 ( .A1(n11954), .A2(n11967), .ZN(n11955) );
  AOI22_X1 U15112 ( .A1(n11957), .A2(n11967), .B1(n11956), .B2(n11955), .ZN(
        n11960) );
  NOR2_X1 U15113 ( .A1(n11958), .A2(n11968), .ZN(n11959) );
  OR3_X1 U15114 ( .A1(n12822), .A2(n11964), .A3(n11963), .ZN(n11986) );
  NOR3_X1 U15115 ( .A1(n11967), .A2(n11966), .A3(n11965), .ZN(n11969) );
  OAI21_X1 U15116 ( .B1(n11970), .B2(n11969), .A(n11968), .ZN(n12485) );
  INV_X1 U15117 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n11971) );
  NAND2_X1 U15118 ( .A1(n11972), .A2(n11971), .ZN(n15605) );
  NAND2_X1 U15119 ( .A1(n19985), .A2(n15605), .ZN(n11973) );
  NAND4_X1 U15120 ( .A1(n11974), .A2(n12485), .A3(n20666), .A4(n11973), .ZN(
        n11985) );
  INV_X1 U15121 ( .A(n11975), .ZN(n12385) );
  INV_X1 U15122 ( .A(n11976), .ZN(n11978) );
  OR2_X1 U15123 ( .A1(n11999), .A2(n19999), .ZN(n11977) );
  AOI21_X1 U15124 ( .B1(n14061), .B2(n12926), .A(n11979), .ZN(n11980) );
  NAND2_X1 U15125 ( .A1(n12011), .A2(n11980), .ZN(n12247) );
  INV_X1 U15126 ( .A(n12247), .ZN(n12478) );
  NAND2_X1 U15127 ( .A1(n11999), .A2(n19972), .ZN(n11981) );
  NAND2_X1 U15128 ( .A1(n11981), .A2(n9590), .ZN(n11982) );
  NAND2_X1 U15129 ( .A1(n11983), .A2(n11982), .ZN(n12009) );
  NAND2_X1 U15130 ( .A1(n12478), .A2(n12009), .ZN(n11984) );
  NAND2_X1 U15131 ( .A1(n12385), .A2(n11984), .ZN(n12788) );
  NAND3_X1 U15132 ( .A1(n11986), .A2(n11985), .A3(n12788), .ZN(n11987) );
  NAND2_X1 U15133 ( .A1(n11987), .A2(n19701), .ZN(n11993) );
  INV_X1 U15134 ( .A(n15605), .ZN(n11989) );
  OAI21_X1 U15135 ( .B1(n19985), .B2(n11989), .A(n20666), .ZN(n12925) );
  OAI211_X1 U15136 ( .C1(n12784), .C2(n12925), .A(n19972), .B(n11990), .ZN(
        n11991) );
  NAND3_X1 U15137 ( .A1(n19824), .A2(n12003), .A3(n11991), .ZN(n11992) );
  INV_X1 U15138 ( .A(n12246), .ZN(n11995) );
  OR2_X1 U15139 ( .A1(n11995), .A2(n12477), .ZN(n11996) );
  NAND2_X1 U15140 ( .A1(n12478), .A2(n11996), .ZN(n12383) );
  OAI211_X1 U15141 ( .C1(n12482), .C2(n9707), .A(n9602), .B(n12383), .ZN(
        n11997) );
  INV_X1 U15142 ( .A(n11997), .ZN(n11998) );
  NOR2_X1 U15143 ( .A1(n11999), .A2(n19827), .ZN(n12000) );
  NAND2_X1 U15144 ( .A1(n12001), .A2(n12000), .ZN(n12776) );
  NAND2_X1 U15145 ( .A1(n11975), .A2(n19985), .ZN(n15558) );
  INV_X1 U15146 ( .A(n12927), .ZN(n12002) );
  AOI22_X1 U15147 ( .A1(n12002), .A2(n12246), .B1(n19972), .B2(n11974), .ZN(
        n12008) );
  OAI21_X1 U15148 ( .B1(n12003), .B2(n11655), .A(n20015), .ZN(n12004) );
  OAI21_X1 U15149 ( .B1(n12004), .B2(n12801), .A(n19985), .ZN(n12007) );
  INV_X1 U15150 ( .A(n19994), .ZN(n12005) );
  NAND2_X1 U15151 ( .A1(n12005), .A2(n19972), .ZN(n12040) );
  NAND2_X1 U15152 ( .A1(n12121), .A2(n11979), .ZN(n12006) );
  AND3_X1 U15153 ( .A1(n12008), .A2(n12007), .A3(n12006), .ZN(n12010) );
  OAI211_X1 U15154 ( .C1(n12011), .C2(n12114), .A(n12010), .B(n12009), .ZN(
        n12012) );
  INV_X1 U15155 ( .A(n12012), .ZN(n12015) );
  OR2_X1 U15156 ( .A1(n12013), .A2(n12923), .ZN(n12014) );
  AND2_X1 U15157 ( .A1(n12015), .A2(n12014), .ZN(n12774) );
  OAI211_X1 U15158 ( .C1(n12771), .C2(n19972), .A(n12774), .B(n12016), .ZN(
        n12017) );
  NAND2_X1 U15159 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15813) );
  INV_X1 U15160 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15890) );
  NOR3_X1 U15161 ( .A1(n11902), .A2(n15901), .A3(n15890), .ZN(n15871) );
  NAND3_X1 U15162 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15871), .ZN(n15860) );
  NOR2_X1 U15163 ( .A1(n11912), .A2(n15860), .ZN(n14826) );
  NAND2_X1 U15164 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14826), .ZN(
        n12020) );
  INV_X1 U15165 ( .A(n12020), .ZN(n12019) );
  NOR2_X1 U15166 ( .A1(n19933), .A2(n19943), .ZN(n19924) );
  INV_X1 U15167 ( .A(n19924), .ZN(n13069) );
  NAND2_X1 U15168 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13066) );
  NOR3_X1 U15169 ( .A1(n13065), .A2(n13069), .A3(n13066), .ZN(n14824) );
  NAND2_X1 U15170 ( .A1(n12019), .A2(n14824), .ZN(n14785) );
  INV_X1 U15171 ( .A(n14823), .ZN(n19950) );
  INV_X1 U15172 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15848) );
  INV_X1 U15173 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14815) );
  NOR2_X1 U15174 ( .A1(n15848), .A2(n14815), .ZN(n15835) );
  NAND3_X1 U15175 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n15835), .ZN(n15827) );
  NOR2_X1 U15176 ( .A1(n15834), .A2(n15827), .ZN(n12127) );
  NAND2_X1 U15177 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12127), .ZN(
        n14781) );
  INV_X1 U15178 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19947) );
  INV_X1 U15179 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19951) );
  OAI21_X1 U15180 ( .B1(n19947), .B2(n19951), .A(n19961), .ZN(n19922) );
  NAND3_X1 U15181 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n19924), .A3(
        n19922), .ZN(n13072) );
  NOR2_X1 U15182 ( .A1(n13072), .A2(n12020), .ZN(n14783) );
  NAND2_X1 U15183 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14783), .ZN(
        n13488) );
  INV_X1 U15184 ( .A(n13488), .ZN(n12021) );
  OR2_X2 U15185 ( .A1(n12248), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19927) );
  AOI22_X1 U15186 ( .A1(n12126), .A2(n19927), .B1(n10093), .B2(n19947), .ZN(
        n13067) );
  OAI221_X1 U15187 ( .B1(n19946), .B2(n12021), .C1(n19946), .C2(n12127), .A(
        n13067), .ZN(n12022) );
  NAND2_X1 U15188 ( .A1(n12895), .A2(n13067), .ZN(n15866) );
  OAI21_X1 U15189 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n19946), .A(
        n15809), .ZN(n14769) );
  AOI21_X1 U15190 ( .B1(n15889), .B2(n14614), .A(n14769), .ZN(n15801) );
  AND2_X1 U15191 ( .A1(n15809), .A2(n12895), .ZN(n14751) );
  AOI21_X1 U15192 ( .B1(n11921), .B2(n14756), .A(n14751), .ZN(n14728) );
  INV_X1 U15193 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12023) );
  NOR3_X1 U15194 ( .A1(n14717), .A2(n14751), .A3(n12023), .ZN(n12131) );
  AND2_X1 U15195 ( .A1(n12528), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12024) );
  AOI21_X1 U15196 ( .B1(n12121), .B2(P1_EBX_REG_30__SCAN_IN), .A(n12024), .ZN(
        n14332) );
  INV_X1 U15197 ( .A(n12025), .ZN(n14331) );
  NAND2_X1 U15198 ( .A1(n12040), .A2(n19951), .ZN(n12027) );
  INV_X1 U15199 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12529) );
  NAND2_X1 U15200 ( .A1(n12929), .A2(n12529), .ZN(n12026) );
  NAND3_X1 U15201 ( .A1(n12027), .A2(n12114), .A3(n12026), .ZN(n12028) );
  NAND2_X1 U15202 ( .A1(n12040), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12030) );
  INV_X1 U15203 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12622) );
  NAND2_X1 U15204 ( .A1(n12114), .A2(n12622), .ZN(n12029) );
  NAND2_X1 U15205 ( .A1(n12030), .A2(n12029), .ZN(n12614) );
  INV_X1 U15206 ( .A(n12031), .ZN(n12032) );
  AOI21_X1 U15207 ( .B1(n12958), .B2(n12929), .A(n12032), .ZN(n12639) );
  OR2_X1 U15208 ( .A1(n12120), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12037) );
  NAND2_X1 U15209 ( .A1(n12040), .A2(n19961), .ZN(n12035) );
  INV_X1 U15210 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U15211 ( .A1(n12929), .A2(n12033), .ZN(n12034) );
  NAND3_X1 U15212 ( .A1(n12035), .A2(n12114), .A3(n12034), .ZN(n12036) );
  NAND2_X1 U15213 ( .A1(n12037), .A2(n12036), .ZN(n12640) );
  MUX2_X1 U15214 ( .A(n12113), .B(n12114), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12038) );
  OAI21_X1 U15215 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n12121), .A(
        n12038), .ZN(n12886) );
  INV_X1 U15216 ( .A(n12886), .ZN(n12039) );
  MUX2_X1 U15217 ( .A(n12120), .B(n12040), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12042) );
  INV_X1 U15218 ( .A(n12040), .ZN(n12074) );
  NAND2_X1 U15219 ( .A1(n12074), .A2(n12528), .ZN(n12090) );
  NAND2_X1 U15220 ( .A1(n12528), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12041) );
  AND3_X1 U15221 ( .A1(n12042), .A2(n12090), .A3(n12041), .ZN(n12998) );
  NAND2_X1 U15222 ( .A1(n12114), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12044) );
  OAI211_X1 U15223 ( .C1(P1_EBX_REG_5__SCAN_IN), .C2(n12528), .A(n12040), .B(
        n12044), .ZN(n12045) );
  OAI21_X1 U15224 ( .B1(n12113), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12045), .ZN(
        n13121) );
  NAND2_X1 U15225 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12528), .ZN(
        n12046) );
  AND2_X1 U15226 ( .A1(n12090), .A2(n12046), .ZN(n12048) );
  MUX2_X1 U15227 ( .A(n12120), .B(n12040), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12047) );
  NAND2_X1 U15228 ( .A1(n12048), .A2(n12047), .ZN(n13073) );
  INV_X1 U15229 ( .A(n12113), .ZN(n12049) );
  INV_X1 U15230 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13234) );
  NAND2_X1 U15231 ( .A1(n12049), .A2(n13234), .ZN(n12052) );
  NAND2_X1 U15232 ( .A1(n12114), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12050) );
  OAI211_X1 U15233 ( .C1(n12528), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12040), .B(
        n12050), .ZN(n12051) );
  AND2_X1 U15234 ( .A1(n12052), .A2(n12051), .ZN(n13231) );
  MUX2_X1 U15235 ( .A(n12120), .B(n12040), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12054) );
  NAND2_X1 U15236 ( .A1(n12528), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12053) );
  NAND2_X1 U15237 ( .A1(n12114), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12055) );
  OAI211_X1 U15238 ( .C1(n12528), .C2(P1_EBX_REG_9__SCAN_IN), .A(n12040), .B(
        n12055), .ZN(n12056) );
  OAI21_X1 U15239 ( .B1(n12113), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12056), .ZN(
        n15879) );
  INV_X1 U15240 ( .A(n12120), .ZN(n12082) );
  INV_X1 U15241 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13478) );
  NAND2_X1 U15242 ( .A1(n12082), .A2(n13478), .ZN(n12061) );
  NAND2_X1 U15243 ( .A1(n12040), .A2(n12057), .ZN(n12059) );
  NAND2_X1 U15244 ( .A1(n12929), .A2(n13478), .ZN(n12058) );
  NAND3_X1 U15245 ( .A1(n12059), .A2(n12114), .A3(n12058), .ZN(n12060) );
  MUX2_X1 U15246 ( .A(n12113), .B(n12114), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12062) );
  OAI21_X1 U15247 ( .B1(n12121), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12062), .ZN(n13513) );
  INV_X1 U15248 ( .A(n13513), .ZN(n12063) );
  NAND2_X1 U15249 ( .A1(n13510), .A2(n12063), .ZN(n14526) );
  MUX2_X1 U15250 ( .A(n12120), .B(n12040), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12065) );
  NAND2_X1 U15251 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n12528), .ZN(
        n12064) );
  MUX2_X1 U15252 ( .A(n12113), .B(n12114), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12066) );
  OAI21_X1 U15253 ( .B1(n12121), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12066), .ZN(n14435) );
  INV_X1 U15254 ( .A(n14435), .ZN(n12067) );
  MUX2_X1 U15255 ( .A(n12113), .B(n12114), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12068) );
  OAI21_X1 U15256 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n12121), .A(
        n12068), .ZN(n14514) );
  OR2_X1 U15257 ( .A1(n12120), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n12072) );
  INV_X1 U15258 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14814) );
  NAND2_X1 U15259 ( .A1(n12040), .A2(n14814), .ZN(n12070) );
  INV_X1 U15260 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15716) );
  NAND2_X1 U15261 ( .A1(n12929), .A2(n15716), .ZN(n12069) );
  NAND3_X1 U15262 ( .A1(n12070), .A2(n12114), .A3(n12069), .ZN(n12071) );
  NOR2_X1 U15263 ( .A1(n14514), .A2(n14513), .ZN(n12073) );
  OR2_X1 U15264 ( .A1(n12120), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n12078) );
  NAND2_X1 U15265 ( .A1(n12040), .A2(n14815), .ZN(n12076) );
  INV_X1 U15266 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14507) );
  NAND2_X1 U15267 ( .A1(n12929), .A2(n14507), .ZN(n12075) );
  NAND3_X1 U15268 ( .A1(n12076), .A2(n12114), .A3(n12075), .ZN(n12077) );
  NAND2_X1 U15269 ( .A1(n12078), .A2(n12077), .ZN(n14504) );
  MUX2_X1 U15270 ( .A(n12113), .B(n12114), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12081) );
  INV_X1 U15271 ( .A(n12121), .ZN(n12616) );
  INV_X1 U15272 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12079) );
  NAND2_X1 U15273 ( .A1(n12616), .A2(n12079), .ZN(n12080) );
  NAND2_X1 U15274 ( .A1(n12081), .A2(n12080), .ZN(n14422) );
  INV_X1 U15275 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14497) );
  NAND2_X1 U15276 ( .A1(n12082), .A2(n14497), .ZN(n12086) );
  NAND2_X1 U15277 ( .A1(n12040), .A2(n15834), .ZN(n12084) );
  NAND2_X1 U15278 ( .A1(n12929), .A2(n14497), .ZN(n12083) );
  NAND3_X1 U15279 ( .A1(n12084), .A2(n12114), .A3(n12083), .ZN(n12085) );
  MUX2_X1 U15280 ( .A(n12113), .B(n12114), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12088) );
  OR2_X1 U15281 ( .A1(n12121), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12087) );
  NAND2_X1 U15282 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12528), .ZN(
        n12089) );
  AND2_X1 U15283 ( .A1(n12090), .A2(n12089), .ZN(n12092) );
  MUX2_X1 U15284 ( .A(n12120), .B(n12040), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12091) );
  NAND2_X1 U15285 ( .A1(n12092), .A2(n12091), .ZN(n14474) );
  MUX2_X1 U15286 ( .A(n12113), .B(n12114), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12093) );
  OAI21_X1 U15287 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n12121), .A(
        n12093), .ZN(n14407) );
  MUX2_X1 U15288 ( .A(n12113), .B(n12114), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12095) );
  OR2_X1 U15289 ( .A1(n12121), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12094) );
  AND2_X1 U15290 ( .A1(n12095), .A2(n12094), .ZN(n14393) );
  OR2_X1 U15291 ( .A1(n12120), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n12100) );
  INV_X1 U15292 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12096) );
  NAND2_X1 U15293 ( .A1(n12040), .A2(n12096), .ZN(n12098) );
  INV_X1 U15294 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15713) );
  NAND2_X1 U15295 ( .A1(n12929), .A2(n15713), .ZN(n12097) );
  NAND3_X1 U15296 ( .A1(n12098), .A2(n12114), .A3(n12097), .ZN(n12099) );
  NAND2_X1 U15297 ( .A1(n12100), .A2(n12099), .ZN(n15635) );
  NAND2_X1 U15298 ( .A1(n14393), .A2(n15635), .ZN(n12101) );
  OR2_X1 U15299 ( .A1(n12120), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n12105) );
  INV_X1 U15300 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15793) );
  NAND2_X1 U15301 ( .A1(n12040), .A2(n15793), .ZN(n12103) );
  INV_X1 U15302 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14468) );
  NAND2_X1 U15303 ( .A1(n12929), .A2(n14468), .ZN(n12102) );
  NAND3_X1 U15304 ( .A1(n12103), .A2(n12114), .A3(n12102), .ZN(n12104) );
  NAND2_X1 U15305 ( .A1(n12105), .A2(n12104), .ZN(n14464) );
  NAND2_X1 U15306 ( .A1(n12114), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12106) );
  OAI211_X1 U15307 ( .C1(n12528), .C2(P1_EBX_REG_25__SCAN_IN), .A(n12040), .B(
        n12106), .ZN(n12107) );
  OAI21_X1 U15308 ( .B1(n12113), .B2(P1_EBX_REG_25__SCAN_IN), .A(n12107), .ZN(
        n14381) );
  MUX2_X1 U15309 ( .A(n12120), .B(n12040), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12110) );
  NAND2_X1 U15310 ( .A1(n12528), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12109) );
  AND2_X1 U15311 ( .A1(n12110), .A2(n12109), .ZN(n14367) );
  NAND2_X1 U15312 ( .A1(n12114), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12111) );
  OAI211_X1 U15313 ( .C1(n12528), .C2(P1_EBX_REG_27__SCAN_IN), .A(n12040), .B(
        n12111), .ZN(n12112) );
  OAI21_X1 U15314 ( .B1(n12113), .B2(P1_EBX_REG_27__SCAN_IN), .A(n12112), .ZN(
        n14358) );
  NAND2_X1 U15315 ( .A1(n12040), .A2(n14731), .ZN(n12115) );
  OAI211_X1 U15316 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n12528), .A(n12115), .B(
        n12114), .ZN(n12117) );
  OR2_X1 U15317 ( .A1(n12120), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n12116) );
  NAND2_X1 U15318 ( .A1(n12117), .A2(n12116), .ZN(n14342) );
  OR2_X1 U15319 ( .A1(n12121), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12119) );
  INV_X1 U15320 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n13928) );
  NAND2_X1 U15321 ( .A1(n12929), .A2(n13928), .ZN(n12118) );
  NAND2_X1 U15322 ( .A1(n12119), .A2(n12118), .ZN(n14329) );
  OAI22_X1 U15323 ( .A1(n14329), .A2(n14331), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12120), .ZN(n13923) );
  NAND2_X1 U15324 ( .A1(n14344), .A2(n13923), .ZN(n13922) );
  MUX2_X1 U15325 ( .A(n14332), .B(n12114), .S(n13922), .Z(n12123) );
  AOI22_X1 U15326 ( .A1(n12121), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12528), .ZN(n12122) );
  NOR2_X1 U15327 ( .A1(n12784), .A2(n9590), .ZN(n19823) );
  AND2_X1 U15328 ( .A1(n11994), .A2(n12482), .ZN(n12124) );
  NOR2_X1 U15329 ( .A1(n19823), .A2(n12124), .ZN(n12125) );
  INV_X1 U15330 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20640) );
  NOR2_X1 U15331 ( .A1(n19927), .A2(n20640), .ZN(n13955) );
  NOR2_X1 U15332 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12611), .ZN(
        n12894) );
  INV_X1 U15333 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15857) );
  NOR2_X1 U15334 ( .A1(n15857), .A2(n14785), .ZN(n13490) );
  NAND2_X1 U15335 ( .A1(n19945), .A2(n13490), .ZN(n14768) );
  OAI21_X1 U15336 ( .B1(n13488), .B2(n19946), .A(n14768), .ZN(n14813) );
  NAND4_X1 U15337 ( .A1(n12128), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n12127), .A4(n14813), .ZN(n15792) );
  NAND2_X1 U15338 ( .A1(n9715), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12129) );
  NOR2_X1 U15339 ( .A1(n15792), .A2(n12129), .ZN(n14745) );
  NAND3_X1 U15340 ( .A1(n14745), .A2(n11921), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14718) );
  NOR3_X1 U15341 ( .A1(n14718), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14719), .ZN(n12130) );
  NAND2_X1 U15342 ( .A1(n12132), .A2(n17516), .ZN(n12142) );
  NAND2_X1 U15343 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17950) );
  NAND2_X1 U15344 ( .A1(n18543), .A2(n17950), .ZN(n18605) );
  NOR2_X1 U15345 ( .A1(n18553), .A2(n20687), .ZN(n17584) );
  NAND2_X1 U15346 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17583) );
  NAND2_X1 U15347 ( .A1(n16551), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16549) );
  NOR2_X1 U15348 ( .A1(n16549), .A2(n17497), .ZN(n16501) );
  NAND2_X1 U15349 ( .A1(n17535), .A2(n16501), .ZN(n16539) );
  NAND2_X1 U15350 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17443) );
  NOR2_X1 U15351 ( .A1(n17443), .A2(n17442), .ZN(n17413) );
  NAND2_X1 U15352 ( .A1(n16492), .A2(n17413), .ZN(n17415) );
  NAND2_X1 U15353 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17414) );
  NAND2_X1 U15354 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17384) );
  NAND2_X1 U15355 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17346) );
  NAND2_X1 U15356 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17328), .ZN(
        n16337) );
  NAND2_X1 U15357 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17304) );
  NAND2_X1 U15358 ( .A1(n17285), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16333) );
  NAND2_X1 U15359 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17270) );
  INV_X1 U15360 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16371) );
  NAND2_X1 U15361 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16198), .ZN(
        n12133) );
  INV_X1 U15362 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18599) );
  NOR2_X1 U15363 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18599), .ZN(n17296) );
  NAND2_X1 U15364 ( .A1(n18553), .A2(n18599), .ZN(n18602) );
  NOR2_X1 U15365 ( .A1(n9987), .A2(n16177), .ZN(n12135) );
  NOR2_X1 U15366 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17399), .ZN(
        n16196) );
  INV_X1 U15367 ( .A(n16195), .ZN(n16334) );
  INV_X1 U15368 ( .A(n17296), .ZN(n17624) );
  INV_X2 U15369 ( .A(n17995), .ZN(n18273) );
  NAND2_X1 U15370 ( .A1(n18273), .A2(n12133), .ZN(n12134) );
  OAI211_X1 U15371 ( .C1(n16334), .C2(n17624), .A(n12134), .B(n9597), .ZN(
        n16197) );
  NAND2_X1 U15372 ( .A1(n12138), .A2(n9600), .ZN(n12141) );
  OR2_X1 U15373 ( .A1(n12139), .A2(n17628), .ZN(n12140) );
  NOR2_X1 U15374 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12144) );
  NOR4_X1 U15375 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12143) );
  NAND4_X1 U15376 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12144), .A4(n12143), .ZN(n12167) );
  NOR4_X1 U15377 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12148) );
  NOR4_X1 U15378 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12147) );
  NOR4_X1 U15379 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12146) );
  NOR4_X1 U15380 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12145) );
  AND4_X1 U15381 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12153) );
  NOR4_X1 U15382 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12151) );
  NOR4_X1 U15383 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12150) );
  NOR4_X1 U15384 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12149) );
  AND4_X1 U15385 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n20595), .ZN(
        n12152) );
  NAND2_X1 U15386 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  INV_X1 U15387 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20662) );
  NOR3_X1 U15388 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20662), .ZN(n12156) );
  NOR4_X1 U15389 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12155) );
  NAND4_X1 U15390 ( .A1(n19965), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12156), .A4(
        n12155), .ZN(U214) );
  NOR4_X1 U15391 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12160) );
  NOR4_X1 U15392 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12159) );
  NOR4_X1 U15393 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12158) );
  NOR4_X1 U15394 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12157) );
  NAND4_X1 U15395 ( .A1(n12160), .A2(n12159), .A3(n12158), .A4(n12157), .ZN(
        n12165) );
  NOR4_X1 U15396 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12163) );
  NOR4_X1 U15397 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12162) );
  NOR4_X1 U15398 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12161) );
  NAND4_X1 U15399 ( .A1(n12163), .A2(n12162), .A3(n12161), .A4(n19581), .ZN(
        n12164) );
  NAND2_X1 U15400 ( .A1(n16225), .A2(U214), .ZN(U212) );
  NAND2_X1 U15401 ( .A1(n17366), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12169) );
  NOR2_X1 U15402 ( .A1(n9990), .A2(n12169), .ZN(n16347) );
  AOI21_X1 U15403 ( .B1(n9990), .B2(n12169), .A(n16347), .ZN(n17370) );
  INV_X1 U15404 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12171) );
  NOR2_X1 U15405 ( .A1(n12168), .A2(n17618), .ZN(n17375) );
  NAND2_X1 U15406 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17375), .ZN(
        n12170) );
  INV_X1 U15407 ( .A(n12169), .ZN(n17342) );
  AOI21_X1 U15408 ( .B1(n12171), .B2(n12170), .A(n17342), .ZN(n17376) );
  XOR2_X1 U15409 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B(n17375), .Z(
        n17389) );
  NOR2_X1 U15410 ( .A1(n17415), .A2(n17618), .ZN(n17416) );
  INV_X1 U15411 ( .A(n17416), .ZN(n12172) );
  NOR2_X1 U15412 ( .A1(n17414), .A2(n12172), .ZN(n12174) );
  INV_X1 U15413 ( .A(n12174), .ZN(n12173) );
  AOI21_X1 U15414 ( .B1(n9993), .B2(n12173), .A(n17375), .ZN(n17404) );
  INV_X1 U15415 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12175) );
  NAND2_X1 U15416 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17416), .ZN(
        n16491) );
  AOI21_X1 U15417 ( .B1(n12175), .B2(n16491), .A(n12174), .ZN(n17417) );
  NOR2_X1 U15418 ( .A1(n17376), .A2(n16454), .ZN(n16453) );
  NOR2_X1 U15419 ( .A1(n16453), .A2(n10012), .ZN(n12178) );
  NOR3_X1 U15420 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18457) );
  AOI211_X1 U15421 ( .C1(n17370), .C2(n12178), .A(n16348), .B(n16659), .ZN(
        n12188) );
  NOR3_X1 U15422 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16650) );
  INV_X1 U15423 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20694) );
  NAND2_X1 U15424 ( .A1(n16650), .A2(n20694), .ZN(n16635) );
  NOR2_X1 U15425 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16635), .ZN(n16624) );
  NAND2_X1 U15426 ( .A1(n16624), .A2(n16616), .ZN(n16615) );
  NOR2_X1 U15427 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16615), .ZN(n16598) );
  NAND2_X1 U15428 ( .A1(n16598), .A2(n16595), .ZN(n16594) );
  INV_X1 U15429 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16923) );
  NAND2_X1 U15430 ( .A1(n16577), .A2(n16923), .ZN(n16572) );
  INV_X1 U15431 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16906) );
  NAND2_X1 U15432 ( .A1(n16553), .A2(n16906), .ZN(n16546) );
  INV_X1 U15433 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16876) );
  NAND2_X1 U15434 ( .A1(n16525), .A2(n16876), .ZN(n16515) );
  NAND2_X1 U15435 ( .A1(n16505), .A2(n16857), .ZN(n16494) );
  INV_X1 U15436 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16825) );
  NAND2_X1 U15437 ( .A1(n16486), .A2(n16825), .ZN(n16476) );
  INV_X1 U15438 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16457) );
  NAND2_X1 U15439 ( .A1(n16466), .A2(n16457), .ZN(n16455) );
  INV_X1 U15440 ( .A(n18450), .ZN(n18606) );
  INV_X1 U15441 ( .A(n12181), .ZN(n18618) );
  NAND2_X1 U15442 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18598), .ZN(n12180) );
  AOI211_X4 U15443 ( .C1(n20687), .C2(n18608), .A(n18618), .B(n12180), .ZN(
        n16672) );
  AOI211_X1 U15444 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16455), .A(n16445), .B(
        n16663), .ZN(n12187) );
  NAND2_X1 U15445 ( .A1(n18329), .A2(n18553), .ZN(n18446) );
  NOR2_X1 U15446 ( .A1(n9578), .A2(n18452), .ZN(n16632) );
  INV_X1 U15447 ( .A(n18608), .ZN(n18600) );
  AOI211_X1 U15448 ( .C1(n18468), .C2(n17192), .A(n18600), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18444) );
  AOI211_X4 U15449 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18598), .A(n18444), .B(
        n18618), .ZN(n16673) );
  INV_X1 U15450 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16759) );
  OAI22_X1 U15451 ( .A1(n9990), .A2(n16658), .B1(n16638), .B2(n16759), .ZN(
        n12186) );
  NAND2_X1 U15452 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16460) );
  INV_X1 U15453 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18504) );
  INV_X1 U15454 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18502) );
  NOR2_X1 U15455 ( .A1(n18504), .A2(n18502), .ZN(n16485) );
  NAND2_X1 U15456 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16485), .ZN(n16452) );
  INV_X1 U15457 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18497) );
  INV_X1 U15458 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18493) );
  INV_X1 U15459 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18489) );
  INV_X1 U15460 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18482) );
  NAND2_X1 U15461 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16644) );
  NOR2_X1 U15462 ( .A1(n18482), .A2(n16644), .ZN(n16626) );
  NAND3_X1 U15463 ( .A1(n16626), .A2(P3_REIP_REG_5__SCAN_IN), .A3(
        P3_REIP_REG_4__SCAN_IN), .ZN(n16589) );
  NOR3_X1 U15464 ( .A1(n18489), .A2(n18487), .A3(n16589), .ZN(n16578) );
  NAND2_X1 U15465 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16578), .ZN(n16554) );
  NOR2_X1 U15466 ( .A1(n18493), .A2(n16554), .ZN(n16556) );
  NAND2_X1 U15467 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16556), .ZN(n16536) );
  NOR2_X1 U15468 ( .A1(n18497), .A2(n16536), .ZN(n16532) );
  NAND2_X1 U15469 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16532), .ZN(n16507) );
  NAND2_X1 U15470 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n12182) );
  NOR2_X1 U15471 ( .A1(n16452), .A2(n16500), .ZN(n16461) );
  INV_X1 U15472 ( .A(n16461), .ZN(n16472) );
  NOR2_X1 U15473 ( .A1(n16460), .A2(n16472), .ZN(n12184) );
  INV_X1 U15474 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18512) );
  INV_X1 U15475 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18510) );
  INV_X1 U15476 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18508) );
  NOR2_X1 U15477 ( .A1(n16507), .A2(n12182), .ZN(n16327) );
  NAND2_X1 U15478 ( .A1(n16327), .A2(n16674), .ZN(n16508) );
  NAND2_X1 U15479 ( .A1(n16664), .A2(n16674), .ZN(n16671) );
  OAI21_X1 U15480 ( .B1(n16432), .B2(n16508), .A(n16671), .ZN(n16451) );
  INV_X1 U15481 ( .A(n16451), .ZN(n12183) );
  MUX2_X1 U15482 ( .A(n12184), .B(n12183), .S(P3_REIP_REG_20__SCAN_IN), .Z(
        n12185) );
  INV_X1 U15483 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15069) );
  NAND2_X1 U15484 ( .A1(n12204), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12201) );
  NAND2_X1 U15485 ( .A1(n12202), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12199) );
  NAND2_X1 U15486 ( .A1(n12200), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12197) );
  NAND2_X1 U15487 ( .A1(n12195), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12210) );
  INV_X1 U15488 ( .A(n12190), .ZN(n12214) );
  AND2_X1 U15489 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12190), .ZN(
        n15544) );
  AOI21_X1 U15490 ( .B1(n15069), .B2(n12214), .A(n15544), .ZN(n15071) );
  AND2_X1 U15491 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12189) );
  INV_X1 U15492 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13548) );
  AND2_X1 U15493 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12191) );
  NAND2_X1 U15494 ( .A1(n13988), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12193) );
  INV_X1 U15495 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12192) );
  INV_X1 U15496 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14025) );
  AOI21_X1 U15497 ( .B1(n15117), .B2(n12194), .A(n12195), .ZN(n15118) );
  AOI21_X1 U15498 ( .B1(n16056), .B2(n12209), .A(n12196), .ZN(n18703) );
  AOI21_X1 U15499 ( .B1(n16067), .B2(n12208), .A(n12198), .ZN(n18724) );
  AOI21_X1 U15500 ( .B1(n18743), .B2(n12199), .A(n12200), .ZN(n18753) );
  AOI21_X1 U15501 ( .B1(n16094), .B2(n12201), .A(n12202), .ZN(n18772) );
  AOI21_X1 U15502 ( .B1(n16106), .B2(n12203), .A(n12204), .ZN(n18788) );
  AOI21_X1 U15503 ( .B1(n16122), .B2(n12206), .A(n9601), .ZN(n18816) );
  AOI21_X1 U15504 ( .B1(n12760), .B2(n12205), .A(n12207), .ZN(n12758) );
  OAI22_X1 U15505 ( .A1(n12317), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n13183) );
  INV_X1 U15506 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18846) );
  OAI22_X1 U15507 ( .A1(n12317), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n18846), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13181) );
  AND2_X1 U15508 ( .A1(n13183), .A2(n13181), .ZN(n13081) );
  OAI21_X1 U15509 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12205), .ZN(n13974) );
  NAND2_X1 U15510 ( .A1(n13081), .A2(n13974), .ZN(n12756) );
  NOR2_X1 U15511 ( .A1(n12758), .A2(n12756), .ZN(n18829) );
  OAI21_X1 U15512 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12207), .A(
        n12206), .ZN(n18991) );
  NAND2_X1 U15513 ( .A1(n18829), .A2(n18991), .ZN(n18813) );
  NOR2_X1 U15514 ( .A1(n18816), .A2(n18813), .ZN(n18798) );
  OAI21_X1 U15515 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9601), .A(
        n12203), .ZN(n18799) );
  NAND2_X1 U15516 ( .A1(n18798), .A2(n18799), .ZN(n18787) );
  NOR2_X1 U15517 ( .A1(n18788), .A2(n18787), .ZN(n18780) );
  OAI21_X1 U15518 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12204), .A(
        n12201), .ZN(n18781) );
  NAND2_X1 U15519 ( .A1(n18780), .A2(n18781), .ZN(n18770) );
  NOR2_X1 U15520 ( .A1(n18772), .A2(n18770), .ZN(n18760) );
  OAI21_X1 U15521 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12202), .A(
        n12199), .ZN(n18761) );
  NAND2_X1 U15522 ( .A1(n18760), .A2(n18761), .ZN(n18750) );
  NOR2_X1 U15523 ( .A1(n18753), .A2(n18750), .ZN(n18737) );
  OAI21_X1 U15524 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12200), .A(
        n12208), .ZN(n18738) );
  NAND2_X1 U15525 ( .A1(n18737), .A2(n18738), .ZN(n18722) );
  NOR2_X1 U15526 ( .A1(n18724), .A2(n18722), .ZN(n18715) );
  OAI21_X1 U15527 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12198), .A(
        n12209), .ZN(n18716) );
  NAND2_X1 U15528 ( .A1(n18715), .A2(n18716), .ZN(n18702) );
  NOR2_X1 U15529 ( .A1(n18703), .A2(n18702), .ZN(n18692) );
  OAI21_X1 U15530 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12196), .A(
        n12194), .ZN(n18694) );
  NAND2_X1 U15531 ( .A1(n18692), .A2(n18694), .ZN(n18682) );
  NOR2_X1 U15532 ( .A1(n15118), .A2(n18682), .ZN(n18670) );
  OAI21_X1 U15533 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12195), .A(
        n12213), .ZN(n18671) );
  NAND2_X1 U15534 ( .A1(n18670), .A2(n18671), .ZN(n12211) );
  AOI21_X1 U15535 ( .B1(n12213), .B2(n15098), .A(n12212), .ZN(n18657) );
  OAI21_X1 U15536 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12212), .A(
        n12214), .ZN(n15083) );
  INV_X1 U15537 ( .A(n15083), .ZN(n18646) );
  OR2_X1 U15538 ( .A1(n18657), .A2(n18646), .ZN(n12215) );
  NOR2_X1 U15539 ( .A1(n18656), .A2(n12215), .ZN(n12218) );
  AND2_X1 U15540 ( .A1(n15083), .A2(n12216), .ZN(n12217) );
  OR2_X1 U15541 ( .A1(n12218), .A2(n12217), .ZN(n18644) );
  NOR3_X1 U15542 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15608) );
  AOI211_X1 U15543 ( .C1(n15071), .C2(n12219), .A(n15545), .B(n19555), .ZN(
        n12244) );
  AND2_X1 U15544 ( .A1(n12575), .A2(n19633), .ZN(n12237) );
  NOR2_X1 U15545 ( .A1(n12432), .A2(n12237), .ZN(n15929) );
  AOI21_X1 U15546 ( .B1(n19685), .B2(n19633), .A(P2_EBX_REG_31__SCAN_IN), .ZN(
        n12221) );
  AND2_X1 U15547 ( .A1(n12273), .A2(n12221), .ZN(n12222) );
  OR2_X2 U15548 ( .A1(n15929), .A2(n12222), .ZN(n18856) );
  INV_X1 U15549 ( .A(n18856), .ZN(n18826) );
  INV_X1 U15550 ( .A(n12272), .ZN(n12223) );
  NAND2_X1 U15551 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19493), .ZN(n19551) );
  NOR2_X1 U15552 ( .A1(n19558), .A2(n19551), .ZN(n16168) );
  NOR2_X1 U15553 ( .A1(n18980), .A2(n16168), .ZN(n12224) );
  NAND2_X1 U15554 ( .A1(n19555), .A2(n12224), .ZN(n12225) );
  OAI22_X1 U15555 ( .A1(n18826), .A2(n11112), .B1(n19602), .B2(n18792), .ZN(
        n12243) );
  OAI21_X1 U15556 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19680), .A(
        P2_EBX_REG_31__SCAN_IN), .ZN(n12226) );
  INV_X1 U15557 ( .A(n12226), .ZN(n12227) );
  AND2_X1 U15558 ( .A1(n9573), .A2(n12227), .ZN(n12228) );
  OAI22_X1 U15559 ( .A1(n15069), .A2(n18742), .B1(n12229), .B2(n18810), .ZN(
        n12242) );
  NAND2_X1 U15560 ( .A1(n13471), .A2(n12230), .ZN(n12231) );
  NAND2_X1 U15561 ( .A1(n14915), .A2(n12231), .ZN(n15213) );
  AND2_X1 U15562 ( .A1(n9573), .A2(n19685), .ZN(n12232) );
  NOR2_X1 U15563 ( .A1(n12234), .A2(n12235), .ZN(n12236) );
  NOR2_X1 U15564 ( .A1(n12233), .A2(n12236), .ZN(n15210) );
  INV_X1 U15565 ( .A(n15210), .ZN(n12240) );
  INV_X1 U15566 ( .A(n12237), .ZN(n12238) );
  NOR2_X1 U15567 ( .A1(n12239), .A2(n12238), .ZN(n12707) );
  OAI22_X1 U15568 ( .A1(n15213), .A2(n18822), .B1(n12240), .B2(n18842), .ZN(
        n12241) );
  NAND2_X1 U15569 ( .A1(n20571), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15585) );
  NAND2_X1 U15570 ( .A1(n20055), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12245) );
  AND2_X1 U15571 ( .A1(n15585), .A2(n12245), .ZN(n12713) );
  NAND2_X1 U15572 ( .A1(n20509), .A2(n12248), .ZN(n20665) );
  AND2_X1 U15573 ( .A1(n20665), .A2(n20571), .ZN(n12249) );
  INV_X1 U15574 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12250) );
  AOI21_X1 U15575 ( .B1(n12713), .B2(n14677), .A(n12250), .ZN(n12264) );
  INV_X1 U15576 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20659) );
  NOR2_X1 U15577 ( .A1(n19927), .A2(n20659), .ZN(n12617) );
  NAND2_X1 U15578 ( .A1(n20052), .A2(n11675), .ZN(n12252) );
  NAND2_X1 U15579 ( .A1(n12252), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12258) );
  INV_X1 U15580 ( .A(n12258), .ZN(n12259) );
  NAND2_X1 U15581 ( .A1(n12494), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12944) );
  NAND2_X1 U15582 ( .A1(n20573), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12255) );
  NAND2_X1 U15583 ( .A1(n12512), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12254) );
  OAI211_X1 U15584 ( .C1(n12944), .C2(n15559), .A(n12255), .B(n12254), .ZN(
        n12256) );
  AOI21_X1 U15585 ( .B1(n12253), .B2(n13706), .A(n12256), .ZN(n12257) );
  INV_X1 U15586 ( .A(n12257), .ZN(n12518) );
  OR2_X1 U15587 ( .A1(n12258), .A2(n12257), .ZN(n12520) );
  OAI21_X1 U15588 ( .B1(n12259), .B2(n12518), .A(n12520), .ZN(n12941) );
  NAND3_X1 U15589 ( .A1(n20571), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15920) );
  INV_X1 U15590 ( .A(n15920), .ZN(n12260) );
  NOR2_X1 U15591 ( .A1(n12941), .A2(n19967), .ZN(n12263) );
  OAI21_X1 U15592 ( .B1(n12261), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11786), .ZN(n12620) );
  NOR2_X1 U15593 ( .A1(n12620), .A2(n19708), .ZN(n12262) );
  OR4_X1 U15594 ( .A1(n12264), .A2(n12617), .A3(n12263), .A4(n12262), .ZN(
        P1_U2999) );
  AND2_X1 U15595 ( .A1(n12268), .A2(n19685), .ZN(n12570) );
  NOR2_X1 U15596 ( .A1(n12570), .A2(n12575), .ZN(n12265) );
  AND3_X1 U15597 ( .A1(n12681), .A2(n12679), .A3(n12265), .ZN(n12696) );
  NOR2_X1 U15598 ( .A1(n12696), .A2(n16174), .ZN(n19676) );
  AND2_X1 U15599 ( .A1(n10217), .A2(n12989), .ZN(n12266) );
  OAI21_X1 U15600 ( .B1(n19676), .B2(n12689), .A(n12324), .ZN(P2_U2819) );
  INV_X1 U15601 ( .A(n12268), .ZN(n12271) );
  INV_X1 U15602 ( .A(n18623), .ZN(n19678) );
  NAND2_X1 U15603 ( .A1(n19642), .A2(n13184), .ZN(n18622) );
  INV_X1 U15604 ( .A(n18622), .ZN(n12269) );
  OAI21_X1 U15605 ( .B1(n12269), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19678), 
        .ZN(n12270) );
  OAI21_X1 U15606 ( .B1(n12271), .B2(n19678), .A(n12270), .ZN(P2_U3612) );
  INV_X1 U15607 ( .A(n12693), .ZN(n12576) );
  INV_X1 U15608 ( .A(n12576), .ZN(n15528) );
  NOR2_X1 U15609 ( .A1(n12272), .A2(n15528), .ZN(n18857) );
  INV_X1 U15610 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19697) );
  INV_X1 U15611 ( .A(n12273), .ZN(n12274) );
  OAI211_X1 U15612 ( .C1(n18857), .C2(n19697), .A(n12274), .B(n18622), .ZN(
        P2_U2814) );
  INV_X2 U15613 ( .A(n12432), .ZN(n18975) );
  INV_X1 U15614 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15615 ( .A1(n13211), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13021), .ZN(n18928) );
  NOR2_X1 U15616 ( .A1(n12430), .A2(n18928), .ZN(n12279) );
  AOI21_X1 U15617 ( .B1(n18975), .B2(P2_EAX_REG_16__SCAN_IN), .A(n12279), .ZN(
        n12275) );
  OAI21_X1 U15618 ( .B1(n12392), .B2(n12276), .A(n12275), .ZN(P2_U2952) );
  INV_X1 U15619 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15620 ( .A1(n13211), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13021), .ZN(n19029) );
  NOR2_X1 U15621 ( .A1(n12430), .A2(n19029), .ZN(n12287) );
  AOI21_X1 U15622 ( .B1(n18975), .B2(P2_EAX_REG_18__SCAN_IN), .A(n12287), .ZN(
        n12277) );
  OAI21_X1 U15623 ( .B1(n12392), .B2(n12278), .A(n12277), .ZN(P2_U2954) );
  INV_X1 U15624 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12281) );
  AOI21_X1 U15625 ( .B1(n18975), .B2(P2_EAX_REG_0__SCAN_IN), .A(n12279), .ZN(
        n12280) );
  OAI21_X1 U15626 ( .B1(n12392), .B2(n12281), .A(n12280), .ZN(P2_U2967) );
  INV_X1 U15627 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15628 ( .A1(n13211), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13021), .ZN(n19040) );
  NOR2_X1 U15629 ( .A1(n12430), .A2(n19040), .ZN(n12284) );
  AOI21_X1 U15630 ( .B1(n18975), .B2(P2_EAX_REG_5__SCAN_IN), .A(n12284), .ZN(
        n12282) );
  OAI21_X1 U15631 ( .B1(n12392), .B2(n12283), .A(n12282), .ZN(P2_U2972) );
  INV_X1 U15632 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n12286) );
  AOI21_X1 U15633 ( .B1(n18975), .B2(P2_EAX_REG_21__SCAN_IN), .A(n12284), .ZN(
        n12285) );
  OAI21_X1 U15634 ( .B1(n12392), .B2(n12286), .A(n12285), .ZN(P2_U2957) );
  INV_X1 U15635 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n12289) );
  AOI21_X1 U15636 ( .B1(n18975), .B2(P2_EAX_REG_2__SCAN_IN), .A(n12287), .ZN(
        n12288) );
  OAI21_X1 U15637 ( .B1(n12392), .B2(n12289), .A(n12288), .ZN(P2_U2969) );
  INV_X1 U15638 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15639 ( .A1(n13211), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13021), .ZN(n15004) );
  NOR2_X1 U15640 ( .A1(n12430), .A2(n15004), .ZN(n12396) );
  AOI21_X1 U15641 ( .B1(n18975), .B2(P2_EAX_REG_4__SCAN_IN), .A(n12396), .ZN(
        n12290) );
  OAI21_X1 U15642 ( .B1(n12392), .B2(n12291), .A(n12290), .ZN(P2_U2971) );
  INV_X1 U15643 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15644 ( .A1(n13211), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13021), .ZN(n19034) );
  NOR2_X1 U15645 ( .A1(n12430), .A2(n19034), .ZN(n12393) );
  AOI21_X1 U15646 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n18975), .A(n12393), .ZN(
        n12292) );
  OAI21_X1 U15647 ( .B1(n12392), .B2(n12293), .A(n12292), .ZN(P2_U2970) );
  INV_X1 U15648 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15649 ( .A1(n13211), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13021), .ZN(n18919) );
  NOR2_X1 U15650 ( .A1(n12430), .A2(n18919), .ZN(n12296) );
  AOI21_X1 U15651 ( .B1(n18975), .B2(P2_EAX_REG_1__SCAN_IN), .A(n12296), .ZN(
        n12294) );
  OAI21_X1 U15652 ( .B1(n12392), .B2(n12295), .A(n12294), .ZN(P2_U2968) );
  INV_X1 U15653 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n12298) );
  AOI21_X1 U15654 ( .B1(n18975), .B2(P2_EAX_REG_17__SCAN_IN), .A(n12296), .ZN(
        n12297) );
  OAI21_X1 U15655 ( .B1(n12392), .B2(n12298), .A(n12297), .ZN(P2_U2953) );
  INV_X1 U15656 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n12304) );
  INV_X1 U15657 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12299) );
  OR2_X1 U15658 ( .A1(n12166), .A2(n12299), .ZN(n12301) );
  NAND2_X1 U15659 ( .A1(n12166), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12300) );
  AND2_X1 U15660 ( .A1(n12301), .A2(n12300), .ZN(n18882) );
  INV_X1 U15661 ( .A(n18882), .ZN(n12302) );
  NAND2_X1 U15662 ( .A1(n18973), .A2(n12302), .ZN(n12354) );
  NAND2_X1 U15663 ( .A1(n18975), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n12303) );
  OAI211_X1 U15664 ( .C1(n12392), .C2(n12304), .A(n12354), .B(n12303), .ZN(
        P2_U2978) );
  INV_X1 U15665 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n12310) );
  INV_X1 U15666 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12305) );
  OR2_X1 U15667 ( .A1(n12166), .A2(n12305), .ZN(n12307) );
  NAND2_X1 U15668 ( .A1(n12166), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12306) );
  AND2_X1 U15669 ( .A1(n12307), .A2(n12306), .ZN(n18887) );
  INV_X1 U15670 ( .A(n18887), .ZN(n12308) );
  NAND2_X1 U15671 ( .A1(n18973), .A2(n12308), .ZN(n12352) );
  NAND2_X1 U15672 ( .A1(n18975), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n12309) );
  OAI211_X1 U15673 ( .C1(n12392), .C2(n12310), .A(n12352), .B(n12309), .ZN(
        P2_U2976) );
  INV_X1 U15674 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n12316) );
  INV_X1 U15675 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n12311) );
  OR2_X1 U15676 ( .A1(n12166), .A2(n12311), .ZN(n12313) );
  NAND2_X1 U15677 ( .A1(n12166), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12312) );
  AND2_X1 U15678 ( .A1(n12313), .A2(n12312), .ZN(n18883) );
  INV_X1 U15679 ( .A(n18883), .ZN(n12314) );
  NAND2_X1 U15680 ( .A1(n18973), .A2(n12314), .ZN(n12357) );
  NAND2_X1 U15681 ( .A1(n18975), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n12315) );
  OAI211_X1 U15682 ( .C1(n12392), .C2(n12316), .A(n12357), .B(n12315), .ZN(
        P2_U2977) );
  OR2_X1 U15683 ( .A1(n19642), .A2(n19634), .ZN(n19662) );
  NAND2_X1 U15684 ( .A1(n19662), .A2(n12317), .ZN(n12318) );
  AND2_X1 U15685 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19652) );
  NAND2_X1 U15686 ( .A1(n12320), .A2(n12319), .ZN(n12321) );
  AND2_X1 U15687 ( .A1(n12322), .A2(n12321), .ZN(n15399) );
  INV_X1 U15688 ( .A(n12324), .ZN(n12323) );
  NOR2_X1 U15689 ( .A1(n19016), .A2(n10804), .ZN(n15398) );
  OAI21_X1 U15690 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18851), .A(
        n12331), .ZN(n15396) );
  NOR2_X1 U15691 ( .A1(n18982), .A2(n15396), .ZN(n12325) );
  AOI211_X1 U15692 ( .C1(n15399), .C2(n16114), .A(n15398), .B(n12325), .ZN(
        n12328) );
  INV_X1 U15693 ( .A(n12455), .ZN(n12538) );
  NAND2_X1 U15694 ( .A1(n19633), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U15695 ( .A1(n12538), .A2(n12326), .ZN(n12336) );
  OAI21_X1 U15696 ( .B1(n18979), .B2(n12336), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12327) );
  OAI211_X1 U15697 ( .C1(n16117), .C2(n12349), .A(n12328), .B(n12327), .ZN(
        P2_U3014) );
  XNOR2_X1 U15698 ( .A(n12329), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12330) );
  XNOR2_X1 U15699 ( .A(n12331), .B(n12330), .ZN(n12445) );
  OAI21_X1 U15700 ( .B1(n12333), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n12332), .ZN(n12442) );
  INV_X1 U15701 ( .A(n12442), .ZN(n12334) );
  NAND2_X1 U15702 ( .A1(n16114), .A2(n12334), .ZN(n12335) );
  NAND2_X1 U15703 ( .A1(n18980), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12437) );
  OAI211_X1 U15704 ( .C1(n18846), .C2(n16121), .A(n12335), .B(n12437), .ZN(
        n12338) );
  NOR2_X1 U15705 ( .A1(n18992), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12337) );
  AOI211_X1 U15706 ( .C1(n16102), .C2(n12445), .A(n12338), .B(n12337), .ZN(
        n12339) );
  OAI21_X1 U15707 ( .B1(n12447), .B2(n16117), .A(n12339), .ZN(P2_U3013) );
  INV_X1 U15708 ( .A(n12341), .ZN(n12342) );
  AOI22_X1 U15709 ( .A1(n12536), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19642), .B2(n19666), .ZN(n12343) );
  NAND2_X1 U15710 ( .A1(n12344), .A2(n12343), .ZN(n12414) );
  NAND2_X1 U15711 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12346) );
  INV_X1 U15712 ( .A(n19663), .ZN(n13040) );
  INV_X1 U15713 ( .A(n12683), .ZN(n12685) );
  NAND2_X1 U15714 ( .A1(n12685), .A2(n12682), .ZN(n12573) );
  NAND2_X1 U15715 ( .A1(n12573), .A2(n10774), .ZN(n12348) );
  INV_X2 U15716 ( .A(n14918), .ZN(n12420) );
  INV_X1 U15717 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12350) );
  MUX2_X1 U15718 ( .A(n12350), .B(n12349), .S(n14918), .Z(n12351) );
  OAI21_X1 U15719 ( .B1(n13040), .B2(n14929), .A(n12351), .ZN(P2_U2887) );
  INV_X1 U15720 ( .A(n12392), .ZN(n18976) );
  NAND2_X1 U15721 ( .A1(n18976), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12353) );
  OAI211_X1 U15722 ( .C1(n12432), .C2(n14967), .A(n12353), .B(n12352), .ZN(
        P2_U2961) );
  INV_X1 U15723 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14947) );
  NAND2_X1 U15724 ( .A1(n18976), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12355) );
  OAI211_X1 U15725 ( .C1(n12432), .C2(n14947), .A(n12355), .B(n12354), .ZN(
        P2_U2963) );
  INV_X1 U15726 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18941) );
  NAND2_X1 U15727 ( .A1(n18976), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n12356) );
  MUX2_X1 U15728 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n12166), .Z(n18875) );
  NAND2_X1 U15729 ( .A1(n18973), .A2(n18875), .ZN(n18969) );
  OAI211_X1 U15730 ( .C1(n18941), .C2(n12432), .A(n12356), .B(n18969), .ZN(
        P2_U2980) );
  INV_X1 U15731 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U15732 ( .A1(n18976), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12358) );
  OAI211_X1 U15733 ( .C1(n12432), .C2(n14958), .A(n12358), .B(n12357), .ZN(
        P2_U2962) );
  INV_X1 U15734 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14940) );
  NAND2_X1 U15735 ( .A1(n18976), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12363) );
  INV_X1 U15736 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n12359) );
  OR2_X1 U15737 ( .A1(n12166), .A2(n12359), .ZN(n12361) );
  NAND2_X1 U15738 ( .A1(n12166), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12360) );
  AND2_X1 U15739 ( .A1(n12361), .A2(n12360), .ZN(n18878) );
  INV_X1 U15740 ( .A(n18878), .ZN(n12362) );
  NAND2_X1 U15741 ( .A1(n18973), .A2(n12362), .ZN(n12424) );
  OAI211_X1 U15742 ( .C1(n12432), .C2(n14940), .A(n12363), .B(n12424), .ZN(
        P2_U2964) );
  NAND2_X1 U15743 ( .A1(n12375), .A2(n19701), .ZN(n12426) );
  NOR2_X1 U15744 ( .A1(n20509), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12427) );
  INV_X1 U15745 ( .A(n19828), .ZN(n19825) );
  AOI211_X1 U15746 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n12426), .A(n12427), 
        .B(n19825), .ZN(n12364) );
  INV_X1 U15747 ( .A(n12364), .ZN(P1_U2801) );
  INV_X1 U15748 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13210) );
  OR2_X1 U15749 ( .A1(n15528), .A2(n16174), .ZN(n12365) );
  NAND2_X1 U15750 ( .A1(n13014), .A2(n12317), .ZN(n19679) );
  INV_X2 U15751 ( .A(n19679), .ZN(n18963) );
  AOI22_X1 U15752 ( .A1(n18963), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12368) );
  OAI21_X1 U15753 ( .B1(n13210), .B2(n18930), .A(n12368), .ZN(P2_U2935) );
  INV_X1 U15754 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14986) );
  AOI22_X1 U15755 ( .A1(n18963), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12369) );
  OAI21_X1 U15756 ( .B1(n14986), .B2(n18930), .A(n12369), .ZN(P2_U2929) );
  INV_X1 U15757 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U15758 ( .A1(n18963), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12370) );
  OAI21_X1 U15759 ( .B1(n14978), .B2(n18930), .A(n12370), .ZN(P2_U2927) );
  INV_X1 U15760 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14993) );
  AOI22_X1 U15761 ( .A1(n18963), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12371) );
  OAI21_X1 U15762 ( .B1(n14993), .B2(n18930), .A(n12371), .ZN(P2_U2930) );
  AOI22_X1 U15763 ( .A1(n18963), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12372) );
  OAI21_X1 U15764 ( .B1(n14967), .B2(n18930), .A(n12372), .ZN(P2_U2926) );
  AOI22_X1 U15765 ( .A1(n18963), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12373) );
  OAI21_X1 U15766 ( .B1(n14947), .B2(n18930), .A(n12373), .ZN(P2_U2924) );
  INV_X1 U15767 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n15003) );
  AOI22_X1 U15768 ( .A1(n18963), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12374) );
  OAI21_X1 U15769 ( .B1(n15003), .B2(n18930), .A(n12374), .ZN(P2_U2931) );
  OR2_X1 U15770 ( .A1(n12822), .A2(n12477), .ZN(n12378) );
  INV_X1 U15771 ( .A(n12375), .ZN(n12376) );
  NAND2_X1 U15772 ( .A1(n12378), .A2(n12377), .ZN(n19703) );
  NAND3_X1 U15773 ( .A1(n12923), .A2(n15605), .A3(n12528), .ZN(n12379) );
  AND2_X1 U15774 ( .A1(n12379), .A2(n20666), .ZN(n20668) );
  OR2_X1 U15775 ( .A1(n19703), .A2(n20668), .ZN(n15576) );
  AND2_X1 U15776 ( .A1(n15576), .A2(n19701), .ZN(n19710) );
  INV_X1 U15777 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12391) );
  INV_X1 U15778 ( .A(n12822), .ZN(n15554) );
  INV_X1 U15779 ( .A(n11979), .ZN(n12380) );
  NAND3_X1 U15780 ( .A1(n12381), .A2(n12380), .A3(n19972), .ZN(n12382) );
  AND2_X1 U15781 ( .A1(n12383), .A2(n12382), .ZN(n12384) );
  OR2_X1 U15782 ( .A1(n12822), .A2(n12384), .ZN(n12387) );
  OR2_X1 U15783 ( .A1(n12485), .A2(n12385), .ZN(n12386) );
  OAI211_X1 U15784 ( .C1(n15554), .C2(n12776), .A(n12387), .B(n12386), .ZN(
        n12388) );
  NAND2_X1 U15785 ( .A1(n12388), .A2(n20015), .ZN(n15574) );
  INV_X1 U15786 ( .A(n15574), .ZN(n12389) );
  NAND2_X1 U15787 ( .A1(n12389), .A2(n19710), .ZN(n12390) );
  OAI21_X1 U15788 ( .B1(n19710), .B2(n12391), .A(n12390), .ZN(P1_U3484) );
  INV_X1 U15789 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n12395) );
  AOI21_X1 U15790 ( .B1(n18975), .B2(P2_EAX_REG_19__SCAN_IN), .A(n12393), .ZN(
        n12394) );
  OAI21_X1 U15791 ( .B1(n12392), .B2(n12395), .A(n12394), .ZN(P2_U2955) );
  INV_X1 U15792 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n12398) );
  AOI21_X1 U15793 ( .B1(n18975), .B2(P2_EAX_REG_20__SCAN_IN), .A(n12396), .ZN(
        n12397) );
  OAI21_X1 U15794 ( .B1(n12392), .B2(n12398), .A(n12397), .ZN(P2_U2956) );
  INV_X1 U15795 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15796 ( .A1(n13211), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13021), .ZN(n18888) );
  NOR2_X1 U15797 ( .A1(n12430), .A2(n18888), .ZN(n12408) );
  AOI21_X1 U15798 ( .B1(n18975), .B2(P2_EAX_REG_24__SCAN_IN), .A(n12408), .ZN(
        n12399) );
  OAI21_X1 U15799 ( .B1(n12392), .B2(n12400), .A(n12399), .ZN(P2_U2960) );
  INV_X1 U15800 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15801 ( .A1(n13211), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13021), .ZN(n19044) );
  NOR2_X1 U15802 ( .A1(n12430), .A2(n19044), .ZN(n12411) );
  AOI21_X1 U15803 ( .B1(n18975), .B2(P2_EAX_REG_6__SCAN_IN), .A(n12411), .ZN(
        n12401) );
  OAI21_X1 U15804 ( .B1(n12392), .B2(n12402), .A(n12401), .ZN(P2_U2973) );
  INV_X1 U15805 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n12404) );
  INV_X1 U15806 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16260) );
  INV_X1 U15807 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n17992) );
  AOI22_X1 U15808 ( .A1(n13211), .A2(n16260), .B1(n17992), .B2(n13021), .ZN(
        n16023) );
  INV_X1 U15809 ( .A(n16023), .ZN(n19053) );
  NOR2_X1 U15810 ( .A1(n12430), .A2(n19053), .ZN(n12405) );
  AOI21_X1 U15811 ( .B1(n18975), .B2(P2_EAX_REG_23__SCAN_IN), .A(n12405), .ZN(
        n12403) );
  OAI21_X1 U15812 ( .B1(n12392), .B2(n12404), .A(n12403), .ZN(P2_U2959) );
  INV_X1 U15813 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n12407) );
  AOI21_X1 U15814 ( .B1(n18975), .B2(P2_EAX_REG_7__SCAN_IN), .A(n12405), .ZN(
        n12406) );
  OAI21_X1 U15815 ( .B1(n12392), .B2(n12407), .A(n12406), .ZN(P2_U2974) );
  INV_X1 U15816 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n12410) );
  AOI21_X1 U15817 ( .B1(n18975), .B2(P2_EAX_REG_8__SCAN_IN), .A(n12408), .ZN(
        n12409) );
  OAI21_X1 U15818 ( .B1(n12392), .B2(n12410), .A(n12409), .ZN(P2_U2975) );
  INV_X1 U15819 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n12413) );
  AOI21_X1 U15820 ( .B1(n18975), .B2(P2_EAX_REG_22__SCAN_IN), .A(n12411), .ZN(
        n12412) );
  OAI21_X1 U15821 ( .B1(n12392), .B2(n12413), .A(n12412), .ZN(P2_U2958) );
  NAND2_X1 U15822 ( .A1(n14201), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12465) );
  XNOR2_X1 U15823 ( .A(n12414), .B(n12465), .ZN(n12418) );
  NAND2_X1 U15824 ( .A1(n12536), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12415) );
  NAND2_X1 U15825 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19335) );
  NAND2_X1 U15826 ( .A1(n10817), .A2(n19666), .ZN(n19250) );
  AND2_X1 U15827 ( .A1(n19335), .A2(n19250), .ZN(n13125) );
  NAND2_X1 U15828 ( .A1(n13125), .A2(n19642), .ZN(n19305) );
  NAND2_X1 U15829 ( .A1(n12415), .A2(n19305), .ZN(n12416) );
  NAND2_X1 U15830 ( .A1(n12418), .A2(n12417), .ZN(n12468) );
  OR2_X1 U15831 ( .A1(n12418), .A2(n12417), .ZN(n12419) );
  MUX2_X1 U15832 ( .A(n12447), .B(n12421), .S(n12420), .Z(n12422) );
  OAI21_X1 U15833 ( .B1(n19654), .B2(n14929), .A(n12422), .ZN(P2_U2886) );
  INV_X1 U15834 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n12425) );
  NAND2_X1 U15835 ( .A1(n18975), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n12423) );
  OAI211_X1 U15836 ( .C1(n12392), .C2(n12425), .A(n12424), .B(n12423), .ZN(
        P2_U2979) );
  OAI21_X1 U15837 ( .B1(n12427), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n12934), 
        .ZN(n12428) );
  OAI21_X1 U15838 ( .B1(n12429), .B2(n12934), .A(n12428), .ZN(P1_U3487) );
  INV_X1 U15839 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n18937) );
  INV_X1 U15840 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15841 ( .A1(n13211), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13021), .ZN(n18870) );
  OAI222_X1 U15842 ( .A1(n12432), .A2(n18937), .B1(n12392), .B2(n12431), .C1(
        n12430), .C2(n18870), .ZN(P2_U2982) );
  NAND2_X1 U15843 ( .A1(n12434), .A2(n12433), .ZN(n12435) );
  NAND2_X1 U15844 ( .A1(n12436), .A2(n12435), .ZN(n19658) );
  NAND2_X1 U15845 ( .A1(n16150), .A2(n19658), .ZN(n12438) );
  NAND2_X1 U15846 ( .A1(n12438), .A2(n12437), .ZN(n12444) );
  INV_X1 U15847 ( .A(n15400), .ZN(n15263) );
  INV_X1 U15848 ( .A(n19008), .ZN(n12439) );
  OAI211_X1 U15849 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15263), .B(n12439), .ZN(n12441) );
  OR2_X1 U15850 ( .A1(n19001), .A2(n13182), .ZN(n12440) );
  OAI211_X1 U15851 ( .C1(n12442), .C2(n18994), .A(n12441), .B(n12440), .ZN(
        n12443) );
  AOI211_X1 U15852 ( .C1(n18999), .C2(n12445), .A(n12444), .B(n12443), .ZN(
        n12446) );
  OAI21_X1 U15853 ( .B1(n12447), .B2(n16158), .A(n12446), .ZN(P2_U3045) );
  INV_X1 U15854 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15855 ( .A1(n18963), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12448) );
  OAI21_X1 U15856 ( .B1(n12449), .B2(n18930), .A(n12448), .ZN(P2_U2928) );
  AOI22_X1 U15857 ( .A1(n18963), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12450) );
  OAI21_X1 U15858 ( .B1(n14958), .B2(n18930), .A(n12450), .ZN(P2_U2925) );
  INV_X1 U15859 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U15860 ( .A1(n18963), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12451) );
  OAI21_X1 U15861 ( .B1(n13250), .B2(n18930), .A(n12451), .ZN(P2_U2934) );
  INV_X1 U15862 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U15863 ( .A1(n18963), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12452) );
  OAI21_X1 U15864 ( .B1(n13438), .B2(n18930), .A(n12452), .ZN(P2_U2932) );
  AOI22_X1 U15865 ( .A1(n18963), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12453) );
  OAI21_X1 U15866 ( .B1(n14940), .B2(n18930), .A(n12453), .ZN(P2_U2923) );
  INV_X1 U15867 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13387) );
  AOI22_X1 U15868 ( .A1(n18963), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12454) );
  OAI21_X1 U15869 ( .B1(n13387), .B2(n18930), .A(n12454), .ZN(P2_U2933) );
  NAND2_X1 U15870 ( .A1(n12456), .A2(n12455), .ZN(n12460) );
  NAND2_X1 U15871 ( .A1(n19335), .A2(n19651), .ZN(n12458) );
  NAND2_X1 U15872 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19489) );
  INV_X1 U15873 ( .A(n19489), .ZN(n12457) );
  NAND2_X1 U15874 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12457), .ZN(
        n12534) );
  AND2_X1 U15875 ( .A1(n12458), .A2(n12534), .ZN(n13126) );
  AOI22_X1 U15876 ( .A1(n12536), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19642), .B2(n13126), .ZN(n12459) );
  NAND2_X1 U15877 ( .A1(n12460), .A2(n12459), .ZN(n12463) );
  INV_X1 U15878 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12461) );
  NOR2_X1 U15879 ( .A1(n14227), .A2(n12461), .ZN(n12462) );
  OR2_X1 U15880 ( .A1(n12463), .A2(n12462), .ZN(n12464) );
  NAND2_X1 U15881 ( .A1(n12463), .A2(n12462), .ZN(n12544) );
  INV_X1 U15882 ( .A(n12414), .ZN(n12466) );
  NAND2_X1 U15883 ( .A1(n12466), .A2(n12465), .ZN(n12467) );
  NOR2_X1 U15884 ( .A1(n10318), .A2(n12420), .ZN(n12471) );
  AOI21_X1 U15885 ( .B1(P2_EBX_REG_2__SCAN_IN), .B2(n12420), .A(n12471), .ZN(
        n12472) );
  OAI21_X1 U15886 ( .B1(n19647), .B2(n14929), .A(n12472), .ZN(P2_U2885) );
  INV_X1 U15887 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n19831) );
  INV_X1 U15888 ( .A(n19823), .ZN(n12473) );
  AOI21_X1 U15889 ( .B1(n12473), .B2(n15558), .A(n15605), .ZN(n12474) );
  NAND2_X1 U15890 ( .A1(n19802), .A2(n19972), .ZN(n19798) );
  INV_X1 U15891 ( .A(n12829), .ZN(n15922) );
  AOI22_X1 U15892 ( .A1(n20667), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12475) );
  OAI21_X1 U15893 ( .B1(n19831), .B2(n19798), .A(n12475), .ZN(P1_U2919) );
  INV_X1 U15894 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n20815) );
  AOI22_X1 U15895 ( .A1(n20667), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12476) );
  OAI21_X1 U15896 ( .B1(n20815), .B2(n19798), .A(n12476), .ZN(P1_U2920) );
  NAND2_X1 U15897 ( .A1(n12478), .A2(n12477), .ZN(n12785) );
  OAI21_X1 U15898 ( .B1(n12479), .B2(n20585), .A(n12785), .ZN(n12480) );
  NAND2_X1 U15899 ( .A1(n12822), .A2(n12480), .ZN(n12782) );
  INV_X1 U15900 ( .A(n12481), .ZN(n12483) );
  NAND4_X1 U15901 ( .A1(n12483), .A2(n12482), .A3(n14532), .A4(n12801), .ZN(
        n12526) );
  NOR2_X1 U15902 ( .A1(n12484), .A2(n20585), .ZN(n12486) );
  NAND2_X1 U15903 ( .A1(n12486), .A2(n12485), .ZN(n12789) );
  OAI21_X1 U15904 ( .B1(n12526), .B2(n12923), .A(n12789), .ZN(n12487) );
  INV_X1 U15905 ( .A(n12487), .ZN(n12488) );
  NAND2_X1 U15906 ( .A1(n12782), .A2(n12488), .ZN(n12489) );
  INV_X1 U15907 ( .A(n12490), .ZN(n12491) );
  INV_X1 U15908 ( .A(DATAI_0_), .ZN(n12493) );
  NAND2_X1 U15909 ( .A1(n19965), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12492) );
  OAI21_X1 U15910 ( .B1(n19965), .B2(n12493), .A(n12492), .ZN(n19856) );
  INV_X1 U15911 ( .A(n19856), .ZN(n19978) );
  INV_X1 U15912 ( .A(n13909), .ZN(n12497) );
  INV_X1 U15913 ( .A(n12495), .ZN(n12496) );
  INV_X1 U15914 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19858) );
  OAI222_X1 U15915 ( .A1(n9576), .A2(n12941), .B1(n19978), .B2(n14601), .C1(
        n15730), .C2(n19858), .ZN(P1_U2904) );
  INV_X1 U15916 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n19841) );
  AOI22_X1 U15917 ( .A1(n20667), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12498) );
  OAI21_X1 U15918 ( .B1(n19841), .B2(n19798), .A(n12498), .ZN(P1_U2914) );
  INV_X1 U15919 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n19837) );
  AOI22_X1 U15920 ( .A1(n20667), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12499) );
  OAI21_X1 U15921 ( .B1(n19837), .B2(n19798), .A(n12499), .ZN(P1_U2916) );
  INV_X1 U15922 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n19835) );
  AOI22_X1 U15923 ( .A1(n20667), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12500) );
  OAI21_X1 U15924 ( .B1(n19835), .B2(n19798), .A(n12500), .ZN(P1_U2917) );
  INV_X1 U15925 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n19833) );
  AOI22_X1 U15926 ( .A1(n20667), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12501) );
  OAI21_X1 U15927 ( .B1(n19833), .B2(n19798), .A(n12501), .ZN(P1_U2918) );
  INV_X1 U15928 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n19843) );
  AOI22_X1 U15929 ( .A1(n20667), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12502) );
  OAI21_X1 U15930 ( .B1(n19843), .B2(n19798), .A(n12502), .ZN(P1_U2913) );
  AOI22_X1 U15931 ( .A1(n20667), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12503) );
  OAI21_X1 U15932 ( .B1(n14563), .B2(n19798), .A(n12503), .ZN(P1_U2912) );
  INV_X1 U15933 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n19850) );
  AOI22_X1 U15934 ( .A1(n20667), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12504) );
  OAI21_X1 U15935 ( .B1(n19850), .B2(n19798), .A(n12504), .ZN(P1_U2909) );
  INV_X1 U15936 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n19852) );
  AOI22_X1 U15937 ( .A1(n20667), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12505) );
  OAI21_X1 U15938 ( .B1(n19852), .B2(n19798), .A(n12505), .ZN(P1_U2908) );
  INV_X1 U15939 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n19839) );
  AOI22_X1 U15940 ( .A1(n20667), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12506) );
  OAI21_X1 U15941 ( .B1(n19839), .B2(n19798), .A(n12506), .ZN(P1_U2915) );
  INV_X1 U15942 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n19846) );
  AOI22_X1 U15943 ( .A1(n20667), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12507) );
  OAI21_X1 U15944 ( .B1(n19846), .B2(n19798), .A(n12507), .ZN(P1_U2911) );
  INV_X1 U15945 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n19848) );
  AOI22_X1 U15946 ( .A1(n20667), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12508) );
  OAI21_X1 U15947 ( .B1(n19848), .B2(n19798), .A(n12508), .ZN(P1_U2910) );
  INV_X1 U15948 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n19854) );
  AOI22_X1 U15949 ( .A1(n20667), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12509) );
  OAI21_X1 U15950 ( .B1(n19854), .B2(n19798), .A(n12509), .ZN(P1_U2907) );
  NAND2_X1 U15951 ( .A1(n20053), .A2(n13706), .ZN(n12517) );
  AOI22_X1 U15952 ( .A1(n12512), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20573), .ZN(n12515) );
  INV_X1 U15953 ( .A(n12944), .ZN(n12513) );
  NAND2_X1 U15954 ( .A1(n12513), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12514) );
  AND2_X1 U15955 ( .A1(n12515), .A2(n12514), .ZN(n12516) );
  NAND2_X1 U15956 ( .A1(n12517), .A2(n12516), .ZN(n12522) );
  OR2_X1 U15957 ( .A1(n12518), .A2(n13952), .ZN(n12519) );
  NAND2_X1 U15958 ( .A1(n12520), .A2(n12519), .ZN(n12521) );
  NAND2_X1 U15959 ( .A1(n12522), .A2(n12521), .ZN(n12636) );
  OR2_X1 U15960 ( .A1(n12522), .A2(n12521), .ZN(n12523) );
  NAND2_X1 U15961 ( .A1(n12636), .A2(n12523), .ZN(n19921) );
  INV_X1 U15962 ( .A(DATAI_1_), .ZN(n12525) );
  NAND2_X1 U15963 ( .A1(n19965), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12524) );
  OAI21_X1 U15964 ( .B1(n19965), .B2(n12525), .A(n12524), .ZN(n19859) );
  INV_X1 U15965 ( .A(n19859), .ZN(n19987) );
  INV_X1 U15966 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19861) );
  OAI222_X1 U15967 ( .A1(n9576), .A2(n19921), .B1(n19987), .B2(n14601), .C1(
        n15730), .C2(n19861), .ZN(P1_U2903) );
  OR2_X1 U15968 ( .A1(n12776), .A2(n12822), .ZN(n12792) );
  NAND2_X1 U15969 ( .A1(n19797), .A2(n14532), .ZN(n14528) );
  XNOR2_X1 U15970 ( .A(n12958), .B(n12528), .ZN(n12893) );
  OAI22_X1 U15971 ( .A1(n14528), .A2(n12893), .B1(n12529), .B2(n19797), .ZN(
        n12530) );
  INV_X1 U15972 ( .A(n12530), .ZN(n12531) );
  OAI21_X1 U15973 ( .B1(n19921), .B2(n14530), .A(n12531), .ZN(P1_U2871) );
  INV_X1 U15974 ( .A(n12534), .ZN(n12533) );
  NAND2_X1 U15975 ( .A1(n12533), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19497) );
  NAND2_X1 U15976 ( .A1(n12670), .A2(n12534), .ZN(n12535) );
  AND3_X1 U15977 ( .A1(n19497), .A2(n19642), .A3(n12535), .ZN(n13131) );
  AOI21_X1 U15978 ( .B1(n12536), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13131), .ZN(n12537) );
  NOR2_X1 U15979 ( .A1(n14227), .A2(n12539), .ZN(n12542) );
  NAND2_X1 U15980 ( .A1(n12541), .A2(n12540), .ZN(n12543) );
  NAND2_X1 U15981 ( .A1(n12547), .A2(n12542), .ZN(n12977) );
  NAND2_X1 U15982 ( .A1(n12556), .A2(n12557), .ZN(n12555) );
  NAND2_X1 U15983 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19043), .ZN(
        n12546) );
  AND2_X1 U15984 ( .A1(n12547), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12548) );
  INV_X1 U15985 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12549) );
  NOR2_X1 U15986 ( .A1(n14227), .A2(n12549), .ZN(n12975) );
  XNOR2_X1 U15987 ( .A(n12597), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12554) );
  OR2_X1 U15988 ( .A1(n12565), .A2(n12550), .ZN(n12552) );
  NAND2_X1 U15989 ( .A1(n12552), .A2(n12551), .ZN(n18793) );
  MUX2_X1 U15990 ( .A(n18793), .B(n11057), .S(n12420), .Z(n12553) );
  OAI21_X1 U15991 ( .B1(n12554), .B2(n14929), .A(n12553), .ZN(P2_U2880) );
  NOR2_X1 U15992 ( .A1(n12532), .A2(n12420), .ZN(n12559) );
  AOI21_X1 U15993 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n12420), .A(n12559), .ZN(
        n12560) );
  OAI21_X1 U15994 ( .B1(n13034), .B2(n14929), .A(n12560), .ZN(P2_U2884) );
  INV_X1 U15995 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12561) );
  NOR2_X1 U15996 ( .A1(n13961), .A2(n12561), .ZN(n12563) );
  INV_X1 U15997 ( .A(n12597), .ZN(n12562) );
  OAI211_X1 U15998 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n12563), .A(
        n12562), .B(n14907), .ZN(n12568) );
  AND2_X1 U15999 ( .A1(n13964), .A2(n12564), .ZN(n12566) );
  OR2_X1 U16000 ( .A1(n12566), .A2(n12565), .ZN(n13175) );
  INV_X1 U16001 ( .A(n13175), .ZN(n18805) );
  NAND2_X1 U16002 ( .A1(n18805), .A2(n14918), .ZN(n12567) );
  OAI211_X1 U16003 ( .C1(n14918), .C2(n12569), .A(n12568), .B(n12567), .ZN(
        P2_U2881) );
  NAND2_X1 U16004 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13014), .ZN(n12710) );
  INV_X1 U16005 ( .A(n12710), .ZN(n15609) );
  AND3_X1 U16006 ( .A1(n12681), .A2(n12679), .A3(n12570), .ZN(n12571) );
  AOI21_X1 U16007 ( .B1(n12683), .B2(n12684), .A(n12571), .ZN(n12988) );
  AND3_X1 U16008 ( .A1(n12988), .A2(n12573), .A3(n12572), .ZN(n12579) );
  INV_X1 U16009 ( .A(n12574), .ZN(n12577) );
  NAND3_X1 U16010 ( .A1(n12577), .A2(n12576), .A3(n12575), .ZN(n12578) );
  OAI22_X1 U16011 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19639), .B1(n12702), 
        .B2(n16174), .ZN(n12580) );
  AOI21_X1 U16012 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15609), .A(n12580), .ZN(
        n15414) );
  OR2_X1 U16013 ( .A1(n12532), .A2(n12644), .ZN(n12593) );
  INV_X1 U16014 ( .A(n11133), .ZN(n12663) );
  NAND2_X1 U16015 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12587) );
  OR2_X1 U16016 ( .A1(n12684), .A2(n12682), .ZN(n12647) );
  INV_X1 U16017 ( .A(n10337), .ZN(n12582) );
  NAND2_X1 U16018 ( .A1(n12582), .A2(n12581), .ZN(n12646) );
  NAND2_X1 U16019 ( .A1(n12647), .A2(n12646), .ZN(n12583) );
  OAI21_X1 U16020 ( .B1(n12663), .B2(n12587), .A(n12583), .ZN(n12590) );
  INV_X1 U16021 ( .A(n10774), .ZN(n12584) );
  NOR2_X1 U16022 ( .A1(n12585), .A2(n12584), .ZN(n12654) );
  INV_X1 U16023 ( .A(n12646), .ZN(n12586) );
  AOI21_X1 U16024 ( .B1(n11133), .B2(n12587), .A(n12586), .ZN(n12588) );
  OAI21_X1 U16025 ( .B1(n12654), .B2(n14296), .A(n12588), .ZN(n12589) );
  MUX2_X1 U16026 ( .A(n12590), .B(n12589), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12591) );
  NOR2_X1 U16027 ( .A1(n12591), .A2(n14115), .ZN(n12592) );
  NAND2_X1 U16028 ( .A1(n12593), .A2(n12592), .ZN(n12678) );
  AOI22_X1 U16029 ( .A1(n19636), .A2(n16167), .B1(n19634), .B2(n12678), .ZN(
        n12595) );
  NAND2_X1 U16030 ( .A1(n15414), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12594) );
  OAI21_X1 U16031 ( .B1(n15414), .B2(n12595), .A(n12594), .ZN(P2_U3596) );
  NAND2_X1 U16032 ( .A1(n12597), .A2(n12596), .ZN(n12623) );
  XNOR2_X1 U16033 ( .A(n12623), .B(n12624), .ZN(n12601) );
  OR2_X1 U16034 ( .A1(n12598), .A2(n12605), .ZN(n12599) );
  NAND2_X1 U16035 ( .A1(n12864), .A2(n12599), .ZN(n18776) );
  MUX2_X1 U16036 ( .A(n11066), .B(n18776), .S(n14918), .Z(n12600) );
  OAI21_X1 U16037 ( .B1(n12601), .B2(n14929), .A(n12600), .ZN(P2_U2878) );
  AND2_X1 U16038 ( .A1(n12597), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12603) );
  OAI211_X1 U16039 ( .C1(n12603), .C2(n12602), .A(n14907), .B(n12623), .ZN(
        n12609) );
  NAND2_X1 U16040 ( .A1(n12604), .A2(n12551), .ZN(n12607) );
  INV_X1 U16041 ( .A(n12605), .ZN(n12606) );
  AND2_X1 U16042 ( .A1(n12607), .A2(n12606), .ZN(n18783) );
  NAND2_X1 U16043 ( .A1(n14918), .A2(n18783), .ZN(n12608) );
  OAI211_X1 U16044 ( .C1(n14918), .C2(n12610), .A(n12609), .B(n12608), .ZN(
        P2_U2879) );
  INV_X1 U16045 ( .A(n13067), .ZN(n19948) );
  AOI21_X1 U16046 ( .B1(n14784), .B2(n19947), .A(n19948), .ZN(n12896) );
  INV_X1 U16047 ( .A(n12611), .ZN(n14801) );
  NOR3_X1 U16048 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14784), .A3(
        n10093), .ZN(n12612) );
  AOI21_X1 U16049 ( .B1(n12896), .B2(n14801), .A(n12612), .ZN(n12613) );
  INV_X1 U16050 ( .A(n12613), .ZN(n12619) );
  INV_X1 U16051 ( .A(n12614), .ZN(n12615) );
  AOI21_X1 U16052 ( .B1(n12616), .B2(n19947), .A(n12615), .ZN(n12935) );
  AOI21_X1 U16053 ( .B1(n19936), .B2(n12935), .A(n12617), .ZN(n12618) );
  OAI211_X1 U16054 ( .C1(n19925), .C2(n12620), .A(n12619), .B(n12618), .ZN(
        P1_U3031) );
  INV_X1 U16055 ( .A(n12935), .ZN(n12621) );
  OAI222_X1 U16056 ( .A1(n12941), .A2(n14530), .B1(n12622), .B2(n19797), .C1(
        n12621), .C2(n14528), .ZN(P1_U2872) );
  INV_X1 U16057 ( .A(n12623), .ZN(n12626) );
  INV_X1 U16058 ( .A(n12624), .ZN(n12625) );
  NAND2_X1 U16059 ( .A1(n12626), .A2(n12625), .ZN(n12866) );
  XNOR2_X1 U16060 ( .A(n12750), .B(n12748), .ZN(n12631) );
  OAI21_X1 U16061 ( .B1(n12627), .B2(n12629), .A(n12628), .ZN(n18756) );
  MUX2_X1 U16062 ( .A(n18744), .B(n18756), .S(n14918), .Z(n12630) );
  OAI21_X1 U16063 ( .B1(n12631), .B2(n14929), .A(n12630), .ZN(P2_U2876) );
  XNOR2_X1 U16064 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12712) );
  AOI21_X1 U16065 ( .B1(n13946), .B2(n12712), .A(n13953), .ZN(n12633) );
  NAND2_X1 U16066 ( .A1(n12512), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12632) );
  OAI211_X1 U16067 ( .C1(n12944), .C2(n9710), .A(n12633), .B(n12632), .ZN(
        n12634) );
  NAND2_X1 U16068 ( .A1(n13953), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12871) );
  INV_X1 U16069 ( .A(n12636), .ZN(n12638) );
  INV_X1 U16070 ( .A(n12635), .ZN(n12637) );
  NAND2_X1 U16071 ( .A1(n12637), .A2(n12638), .ZN(n12872) );
  OAI21_X1 U16072 ( .B1(n12637), .B2(n12638), .A(n12872), .ZN(n12974) );
  NOR2_X1 U16073 ( .A1(n12639), .A2(n12640), .ZN(n12641) );
  OR2_X1 U16074 ( .A1(n12884), .A2(n12641), .ZN(n19954) );
  INV_X1 U16075 ( .A(n19954), .ZN(n12642) );
  AOI22_X1 U16076 ( .A1(n19792), .A2(n12642), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14520), .ZN(n12643) );
  OAI21_X1 U16077 ( .B1(n12974), .B2(n14530), .A(n12643), .ZN(P1_U2870) );
  INV_X1 U16078 ( .A(n12644), .ZN(n12661) );
  NAND2_X1 U16079 ( .A1(n12645), .A2(n12646), .ZN(n12653) );
  NAND2_X1 U16080 ( .A1(n12647), .A2(n12653), .ZN(n12652) );
  NOR2_X1 U16081 ( .A1(n12648), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12649) );
  OAI21_X1 U16082 ( .B1(n12650), .B2(n12649), .A(n11133), .ZN(n12651) );
  OAI211_X1 U16083 ( .C1(n12654), .C2(n12653), .A(n12652), .B(n12651), .ZN(
        n12655) );
  AOI21_X1 U16084 ( .B1(n19005), .B2(n12661), .A(n12655), .ZN(n13185) );
  INV_X1 U16085 ( .A(n12702), .ZN(n12677) );
  MUX2_X1 U16086 ( .A(n12581), .B(n13185), .S(n12677), .Z(n12699) );
  NOR2_X1 U16087 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12699), .ZN(
        n12673) );
  NAND2_X1 U16088 ( .A1(n11133), .A2(n10103), .ZN(n12659) );
  NAND2_X1 U16089 ( .A1(n12656), .A2(n11019), .ZN(n12662) );
  OAI21_X1 U16090 ( .B1(n12657), .B2(n10336), .A(n12662), .ZN(n12658) );
  NAND2_X1 U16091 ( .A1(n12659), .A2(n12658), .ZN(n12660) );
  AOI21_X1 U16092 ( .B1(n9598), .B2(n12661), .A(n12660), .ZN(n15410) );
  AOI21_X1 U16093 ( .B1(n15410), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n12702), .ZN(n12669) );
  NAND2_X1 U16094 ( .A1(n12340), .A2(n12661), .ZN(n12666) );
  INV_X1 U16095 ( .A(n12662), .ZN(n12664) );
  MUX2_X1 U16096 ( .A(n12664), .B(n12663), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n12665) );
  NAND2_X1 U16097 ( .A1(n12666), .A2(n12665), .ZN(n15405) );
  NOR2_X1 U16098 ( .A1(n15405), .A2(n19666), .ZN(n12667) );
  OAI21_X1 U16099 ( .B1(n15410), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n12667), .ZN(n12668) );
  OAI211_X1 U16100 ( .C1(n12678), .C2(n12670), .A(n12669), .B(n12668), .ZN(
        n12671) );
  INV_X1 U16101 ( .A(n12671), .ZN(n12672) );
  AOI222_X1 U16102 ( .A1(n12673), .A2(n12672), .B1(n12673), .B2(n19651), .C1(
        n12672), .C2(n19651), .ZN(n12675) );
  NAND2_X1 U16103 ( .A1(n12670), .A2(n12678), .ZN(n12674) );
  NAND2_X1 U16104 ( .A1(n12675), .A2(n12674), .ZN(n12676) );
  NAND2_X1 U16105 ( .A1(n12676), .A2(n15610), .ZN(n12704) );
  OAI21_X1 U16106 ( .B1(n12699), .B2(n10141), .A(n15531), .ZN(n12701) );
  NAND2_X1 U16107 ( .A1(n12678), .A2(n12677), .ZN(n12698) );
  INV_X1 U16108 ( .A(n12679), .ZN(n12680) );
  AOI22_X1 U16109 ( .A1(n12683), .A2(n12682), .B1(n12681), .B2(n12680), .ZN(
        n12687) );
  NAND2_X1 U16110 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  AND2_X1 U16111 ( .A1(n12687), .A2(n12686), .ZN(n19673) );
  INV_X1 U16112 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n12688) );
  NAND2_X1 U16113 ( .A1(n12689), .A2(n12688), .ZN(n12695) );
  NAND2_X1 U16114 ( .A1(n19683), .A2(n12690), .ZN(n12692) );
  OAI22_X1 U16115 ( .A1(n12693), .A2(n12692), .B1(n10739), .B2(n12691), .ZN(
        n12694) );
  AOI21_X1 U16116 ( .B1(n12696), .B2(n12695), .A(n12694), .ZN(n12697) );
  OAI211_X1 U16117 ( .C1(n12699), .C2(n12698), .A(n19673), .B(n12697), .ZN(
        n12700) );
  AOI21_X1 U16118 ( .B1(n12702), .B2(n12701), .A(n12700), .ZN(n12703) );
  AND2_X1 U16119 ( .A1(n12704), .A2(n12703), .ZN(n16175) );
  NAND2_X1 U16120 ( .A1(n16175), .A2(n13184), .ZN(n12705) );
  NAND2_X1 U16121 ( .A1(n12705), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12709) );
  OR2_X1 U16122 ( .A1(n12706), .A2(n19493), .ZN(n19682) );
  AOI21_X1 U16123 ( .B1(n10718), .B2(n12707), .A(n19682), .ZN(n12708) );
  NOR2_X1 U16124 ( .A1(n19550), .A2(n12317), .ZN(n12711) );
  OAI21_X1 U16125 ( .B1(n12711), .B2(n19639), .A(n12710), .ZN(P2_U3593) );
  INV_X1 U16126 ( .A(n12712), .ZN(n12967) );
  INV_X1 U16127 ( .A(n12713), .ZN(n12714) );
  INV_X1 U16128 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12716) );
  INV_X1 U16129 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n12715) );
  OAI22_X1 U16130 ( .A1(n14677), .A2(n12716), .B1(n19927), .B2(n12715), .ZN(
        n12717) );
  AOI21_X1 U16131 ( .B1(n12967), .B2(n19916), .A(n12717), .ZN(n12722) );
  OR2_X1 U16132 ( .A1(n12719), .A2(n12718), .ZN(n19953) );
  NAND3_X1 U16133 ( .A1(n19953), .A2(n12720), .A3(n19917), .ZN(n12721) );
  OAI211_X1 U16134 ( .C1(n12974), .C2(n19967), .A(n12722), .B(n12721), .ZN(
        P1_U2997) );
  NAND2_X1 U16135 ( .A1(n12724), .A2(n12723), .ZN(n12726) );
  XNOR2_X1 U16136 ( .A(n12726), .B(n12725), .ZN(n12743) );
  MUX2_X1 U16137 ( .A(n12729), .B(n12728), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n12735) );
  XNOR2_X1 U16138 ( .A(n12731), .B(n12730), .ZN(n19640) );
  INV_X1 U16139 ( .A(n19640), .ZN(n18901) );
  NOR2_X1 U16140 ( .A1(n12737), .A2(n19016), .ZN(n12732) );
  AOI21_X1 U16141 ( .B1(n16150), .B2(n18901), .A(n12732), .ZN(n12733) );
  OAI21_X1 U16142 ( .B1(n12532), .B2(n16158), .A(n12733), .ZN(n12734) );
  AOI211_X1 U16143 ( .C1(n12741), .C2(n16154), .A(n12735), .B(n12734), .ZN(
        n12736) );
  OAI21_X1 U16144 ( .B1(n12743), .B2(n16152), .A(n12736), .ZN(P2_U3043) );
  OAI22_X1 U16145 ( .A1(n16121), .A2(n12760), .B1(n12737), .B2(n19016), .ZN(
        n12738) );
  AOI21_X1 U16146 ( .B1(n16107), .B2(n12758), .A(n12738), .ZN(n12739) );
  OAI21_X1 U16147 ( .B1(n12532), .B2(n16117), .A(n12739), .ZN(n12740) );
  AOI21_X1 U16148 ( .B1(n12741), .B2(n16114), .A(n12740), .ZN(n12742) );
  OAI21_X1 U16149 ( .B1(n12743), .B2(n18982), .A(n12742), .ZN(P2_U3011) );
  NAND2_X1 U16150 ( .A1(n12744), .A2(n12628), .ZN(n12747) );
  INV_X1 U16151 ( .A(n12745), .ZN(n12746) );
  AND2_X1 U16152 ( .A1(n12747), .A2(n12746), .ZN(n18739) );
  INV_X1 U16153 ( .A(n18739), .ZN(n12755) );
  AND2_X1 U16154 ( .A1(n12750), .A2(n12748), .ZN(n12752) );
  AND2_X1 U16155 ( .A1(n12751), .A2(n12748), .ZN(n12749) );
  OAI211_X1 U16156 ( .C1(n12752), .C2(n12751), .A(n14907), .B(n13006), .ZN(
        n12754) );
  NAND2_X1 U16157 ( .A1(n12420), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12753) );
  OAI211_X1 U16158 ( .C1(n12755), .C2(n12420), .A(n12754), .B(n12753), .ZN(
        P2_U2875) );
  NAND2_X1 U16159 ( .A1(n18814), .A2(n12756), .ZN(n12757) );
  XNOR2_X1 U16160 ( .A(n12758), .B(n12757), .ZN(n12766) );
  OAI22_X1 U16161 ( .A1(n12737), .A2(n18792), .B1(n12759), .B2(n18810), .ZN(
        n12762) );
  OAI22_X1 U16162 ( .A1(n12760), .A2(n18742), .B1(n18842), .B2(n19640), .ZN(
        n12761) );
  AOI211_X1 U16163 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n18856), .A(n12762), .B(
        n12761), .ZN(n12764) );
  NAND2_X1 U16164 ( .A1(n19636), .A2(n18857), .ZN(n12763) );
  OAI211_X1 U16165 ( .C1(n18822), .C2(n12532), .A(n12764), .B(n12763), .ZN(
        n12765) );
  AOI21_X1 U16166 ( .B1(n12766), .B2(n18818), .A(n12765), .ZN(n12767) );
  INV_X1 U16167 ( .A(n12767), .ZN(P2_U2852) );
  INV_X1 U16168 ( .A(DATAI_2_), .ZN(n12769) );
  NAND2_X1 U16169 ( .A1(n19965), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12768) );
  OAI21_X1 U16170 ( .B1(n19965), .B2(n12769), .A(n12768), .ZN(n19862) );
  INV_X1 U16171 ( .A(n19862), .ZN(n19991) );
  INV_X1 U16172 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19864) );
  OAI222_X1 U16173 ( .A1(n9576), .A2(n12974), .B1(n19991), .B2(n14601), .C1(
        n15730), .C2(n19864), .ZN(P1_U2902) );
  NOR2_X1 U16174 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20570), .ZN(n12818) );
  INV_X1 U16175 ( .A(n12770), .ZN(n19975) );
  AND3_X1 U16176 ( .A1(n12784), .A2(n12772), .A3(n12771), .ZN(n12773) );
  AND2_X1 U16177 ( .A1(n12484), .A2(n12773), .ZN(n12775) );
  AND2_X1 U16178 ( .A1(n12775), .A2(n12774), .ZN(n14062) );
  INV_X1 U16179 ( .A(n14062), .ZN(n14843) );
  XNOR2_X1 U16180 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12780) );
  NAND2_X1 U16181 ( .A1(n12776), .A2(n12785), .ZN(n12798) );
  INV_X1 U16182 ( .A(n14844), .ZN(n14839) );
  NAND2_X1 U16183 ( .A1(n14839), .A2(n9710), .ZN(n12796) );
  NAND2_X1 U16184 ( .A1(n14844), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12799) );
  NAND2_X1 U16185 ( .A1(n12796), .A2(n12799), .ZN(n12777) );
  NAND2_X1 U16186 ( .A1(n12798), .A2(n12777), .ZN(n12779) );
  INV_X1 U16187 ( .A(n12777), .ZN(n14850) );
  NAND3_X1 U16188 ( .A1(n14062), .A2(n12801), .A3(n14850), .ZN(n12778) );
  OAI211_X1 U16189 ( .C1(n15558), .C2(n12780), .A(n12779), .B(n12778), .ZN(
        n12781) );
  AOI21_X1 U16190 ( .B1(n19975), .B2(n14843), .A(n12781), .ZN(n14854) );
  INV_X1 U16191 ( .A(n14854), .ZN(n12795) );
  INV_X1 U16192 ( .A(n12782), .ZN(n12787) );
  NOR2_X1 U16193 ( .A1(n15605), .A2(n20585), .ZN(n12783) );
  AND2_X1 U16194 ( .A1(n12822), .A2(n12783), .ZN(n15582) );
  NAND3_X1 U16195 ( .A1(n12785), .A2(n15558), .A3(n12784), .ZN(n12786) );
  OAI21_X1 U16196 ( .B1(n12787), .B2(n15582), .A(n12786), .ZN(n12794) );
  OAI211_X1 U16197 ( .C1(n12927), .C2(n11974), .A(n12789), .B(n12788), .ZN(
        n12790) );
  INV_X1 U16198 ( .A(n12790), .ZN(n12791) );
  AND2_X1 U16199 ( .A1(n12792), .A2(n12791), .ZN(n12793) );
  MUX2_X1 U16200 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n12795), .S(
        n15561), .Z(n15567) );
  AOI22_X1 U16201 ( .A1(n12818), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15567), .B2(n20570), .ZN(n12812) );
  XNOR2_X1 U16202 ( .A(n12796), .B(n11518), .ZN(n12797) );
  NAND2_X1 U16203 ( .A1(n12798), .A2(n12797), .ZN(n12808) );
  NAND2_X1 U16204 ( .A1(n12799), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12800) );
  NAND2_X1 U16205 ( .A1(n11715), .A2(n12800), .ZN(n14856) );
  NAND3_X1 U16206 ( .A1(n14062), .A2(n12801), .A3(n14856), .ZN(n12807) );
  INV_X1 U16207 ( .A(n15558), .ZN(n14060) );
  INV_X1 U16208 ( .A(n12802), .ZN(n12805) );
  NAND2_X1 U16209 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12803) );
  NAND2_X1 U16210 ( .A1(n11518), .A2(n12803), .ZN(n12804) );
  NAND3_X1 U16211 ( .A1(n14060), .A2(n12805), .A3(n12804), .ZN(n12806) );
  NAND3_X1 U16212 ( .A1(n12808), .A2(n12807), .A3(n12806), .ZN(n12809) );
  AOI21_X1 U16213 ( .B1(n20255), .B2(n14843), .A(n12809), .ZN(n14859) );
  NOR2_X1 U16214 ( .A1(n15561), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12810) );
  AOI21_X1 U16215 ( .B1(n14859), .B2(n15561), .A(n12810), .ZN(n15555) );
  AOI22_X1 U16216 ( .A1(n12818), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20570), .B2(n15555), .ZN(n12811) );
  NOR2_X1 U16217 ( .A1(n12812), .A2(n12811), .ZN(n15570) );
  INV_X1 U16218 ( .A(n12813), .ZN(n14838) );
  NAND2_X1 U16219 ( .A1(n15570), .A2(n14838), .ZN(n12830) );
  INV_X1 U16220 ( .A(n20134), .ZN(n20384) );
  OR2_X1 U16221 ( .A1(n12814), .A2(n20384), .ZN(n12815) );
  XNOR2_X1 U16222 ( .A(n12815), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19760) );
  INV_X1 U16223 ( .A(n12484), .ZN(n12816) );
  NAND2_X1 U16224 ( .A1(n19760), .A2(n12816), .ZN(n15915) );
  NAND2_X1 U16225 ( .A1(n15915), .A2(n15561), .ZN(n12821) );
  INV_X1 U16226 ( .A(n15561), .ZN(n12817) );
  AOI21_X1 U16227 ( .B1(n12817), .B2(n15917), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n12820) );
  AND2_X1 U16228 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12818), .ZN(
        n12819) );
  AOI21_X1 U16229 ( .B1(n12821), .B2(n12820), .A(n12819), .ZN(n15579) );
  INV_X1 U16230 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19709) );
  AND3_X1 U16231 ( .A1(n12830), .A2(n15579), .A3(n19709), .ZN(n12823) );
  NAND2_X1 U16232 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12829), .ZN(n15926) );
  INV_X1 U16233 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20386) );
  NAND2_X1 U16234 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20386), .ZN(n12857) );
  INV_X1 U16235 ( .A(n12857), .ZN(n14836) );
  NOR2_X1 U16236 ( .A1(n12770), .A2(n14836), .ZN(n12827) );
  NAND2_X1 U16237 ( .A1(n20053), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20098) );
  NOR2_X1 U16238 ( .A1(n20098), .A2(n20509), .ZN(n12825) );
  AND2_X1 U16239 ( .A1(n20098), .A2(n20518), .ZN(n20514) );
  MUX2_X1 U16240 ( .A(n12825), .B(n20514), .S(n12824), .Z(n12826) );
  OAI21_X1 U16241 ( .B1(n12827), .B2(n12826), .A(n19963), .ZN(n12828) );
  OAI21_X1 U16242 ( .B1(n19963), .B2(n20256), .A(n12828), .ZN(P1_U3476) );
  NAND3_X1 U16243 ( .A1(n12830), .A2(n15579), .A3(n12829), .ZN(n15588) );
  INV_X1 U16244 ( .A(n15588), .ZN(n12832) );
  INV_X1 U16245 ( .A(n12253), .ZN(n14063) );
  OAI22_X1 U16246 ( .A1(n20052), .A2(n20509), .B1(n14063), .B2(n14836), .ZN(
        n12831) );
  OAI21_X1 U16247 ( .B1(n12832), .B2(n12831), .A(n19963), .ZN(n12833) );
  OAI21_X1 U16248 ( .B1(n19963), .B2(n20428), .A(n12833), .ZN(P1_U3478) );
  XNOR2_X1 U16249 ( .A(n12835), .B(n12834), .ZN(n18983) );
  OAI21_X1 U16250 ( .B1(n12837), .B2(n12844), .A(n12836), .ZN(n18981) );
  OR2_X1 U16251 ( .A1(n12839), .A2(n12838), .ZN(n12841) );
  NAND2_X1 U16252 ( .A1(n12841), .A2(n12840), .ZN(n18824) );
  INV_X1 U16253 ( .A(n12842), .ZN(n16161) );
  NOR2_X1 U16254 ( .A1(n10842), .A2(n19016), .ZN(n12843) );
  AOI221_X1 U16255 ( .B1(n16161), .B2(n12844), .C1(n16151), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n12843), .ZN(n12850) );
  INV_X1 U16256 ( .A(n12845), .ZN(n12846) );
  AOI21_X1 U16257 ( .B1(n12848), .B2(n12847), .A(n12846), .ZN(n18987) );
  NAND2_X1 U16258 ( .A1(n18987), .A2(n19004), .ZN(n12849) );
  OAI211_X1 U16259 ( .C1(n18995), .C2(n18824), .A(n12850), .B(n12849), .ZN(
        n12851) );
  AOI21_X1 U16260 ( .B1(n16154), .B2(n18981), .A(n12851), .ZN(n12852) );
  OAI21_X1 U16261 ( .B1(n16152), .B2(n18983), .A(n12852), .ZN(P2_U3042) );
  INV_X1 U16262 ( .A(n19963), .ZN(n12862) );
  INV_X1 U16263 ( .A(n12854), .ZN(n12853) );
  OAI22_X1 U16264 ( .A1(n20475), .A2(n20053), .B1(n20232), .B2(n20098), .ZN(
        n12856) );
  INV_X1 U16265 ( .A(n19969), .ZN(n12855) );
  NAND2_X1 U16266 ( .A1(n12856), .A2(n20356), .ZN(n12859) );
  AOI21_X1 U16267 ( .B1(n19969), .B2(n20055), .A(n20509), .ZN(n12858) );
  AOI22_X1 U16268 ( .A1(n12859), .A2(n12858), .B1(n12857), .B2(n20255), .ZN(
        n12861) );
  NAND2_X1 U16269 ( .A1(n12862), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12860) );
  OAI21_X1 U16270 ( .B1(n12862), .B2(n12861), .A(n12860), .ZN(P1_U3475) );
  AND2_X1 U16271 ( .A1(n12864), .A2(n12863), .ZN(n12865) );
  OR2_X1 U16272 ( .A1(n12627), .A2(n12865), .ZN(n15369) );
  NOR2_X1 U16273 ( .A1(n12420), .A2(n15369), .ZN(n12869) );
  AOI211_X1 U16274 ( .C1(n12867), .C2(n12866), .A(n14929), .B(n12750), .ZN(
        n12868) );
  AOI211_X1 U16275 ( .C1(n12420), .C2(P2_EBX_REG_10__SCAN_IN), .A(n12869), .B(
        n12868), .ZN(n12870) );
  INV_X1 U16276 ( .A(n12870), .ZN(P2_U2877) );
  NAND2_X1 U16277 ( .A1(n12872), .A2(n12871), .ZN(n12882) );
  NAND2_X1 U16278 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12874) );
  INV_X1 U16279 ( .A(n12874), .ZN(n12873) );
  INV_X1 U16280 ( .A(n12915), .ZN(n12946) );
  INV_X1 U16281 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12875) );
  NAND2_X1 U16282 ( .A1(n12875), .A2(n12874), .ZN(n12876) );
  NAND2_X1 U16283 ( .A1(n12946), .A2(n12876), .ZN(n19776) );
  AOI22_X1 U16284 ( .A1(n19776), .A2(n13946), .B1(n13953), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12878) );
  NAND2_X1 U16285 ( .A1(n13900), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12877) );
  OAI211_X1 U16286 ( .C1(n12944), .C2(n11518), .A(n12878), .B(n12877), .ZN(
        n12879) );
  INV_X1 U16287 ( .A(n12879), .ZN(n12880) );
  OR2_X1 U16288 ( .A1(n12882), .A2(n12881), .ZN(n12883) );
  AND2_X1 U16289 ( .A1(n13095), .A2(n12883), .ZN(n19786) );
  INV_X1 U16290 ( .A(n19786), .ZN(n12911) );
  INV_X1 U16291 ( .A(n12884), .ZN(n12887) );
  INV_X1 U16292 ( .A(n12999), .ZN(n12885) );
  AOI21_X1 U16293 ( .B1(n12887), .B2(n12886), .A(n12885), .ZN(n19935) );
  AOI22_X1 U16294 ( .A1(n19792), .A2(n19935), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14520), .ZN(n12888) );
  OAI21_X1 U16295 ( .B1(n12911), .B2(n14530), .A(n12888), .ZN(P1_U2869) );
  OR2_X1 U16296 ( .A1(n12889), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12890) );
  AND2_X1 U16297 ( .A1(n12891), .A2(n12890), .ZN(n19918) );
  INV_X1 U16298 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n12892) );
  OAI22_X1 U16299 ( .A1(n19955), .A2(n12893), .B1(n19927), .B2(n12892), .ZN(
        n12900) );
  NOR2_X1 U16300 ( .A1(n12895), .A2(n12894), .ZN(n12898) );
  INV_X1 U16301 ( .A(n12896), .ZN(n12897) );
  MUX2_X1 U16302 ( .A(n12898), .B(n12897), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n12899) );
  AOI211_X1 U16303 ( .C1(n19952), .C2(n19918), .A(n12900), .B(n12899), .ZN(
        n12901) );
  INV_X1 U16304 ( .A(n12901), .ZN(P1_U3030) );
  OAI21_X1 U16305 ( .B1(n12904), .B2(n12903), .A(n12902), .ZN(n19937) );
  INV_X1 U16306 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n12905) );
  NOR2_X1 U16307 ( .A1(n19927), .A2(n12905), .ZN(n19934) );
  AOI21_X1 U16308 ( .B1(n19914), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n19934), .ZN(n12906) );
  OAI21_X1 U16309 ( .B1(n19912), .B2(n19776), .A(n12906), .ZN(n12907) );
  AOI21_X1 U16310 ( .B1(n19786), .B2(n15781), .A(n12907), .ZN(n12908) );
  OAI21_X1 U16311 ( .B1(n19937), .B2(n19708), .A(n12908), .ZN(P1_U2996) );
  INV_X1 U16312 ( .A(DATAI_3_), .ZN(n12910) );
  NAND2_X1 U16313 ( .A1(n19965), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12909) );
  OAI21_X1 U16314 ( .B1(n19965), .B2(n12910), .A(n12909), .ZN(n19865) );
  INV_X1 U16315 ( .A(n19865), .ZN(n19996) );
  INV_X1 U16316 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20744) );
  OAI222_X1 U16317 ( .A1(n9576), .A2(n12911), .B1(n19996), .B2(n14601), .C1(
        n15730), .C2(n20744), .ZN(P1_U2901) );
  NAND2_X1 U16318 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20670), .ZN(n15587) );
  NOR2_X1 U16319 ( .A1(n15587), .A2(n20571), .ZN(n12914) );
  NAND2_X1 U16320 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20571), .ZN(n12912) );
  OAI21_X1 U16321 ( .B1(n12912), .B2(n13952), .A(n19927), .ZN(n12913) );
  NAND2_X1 U16322 ( .A1(n13855), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13858) );
  INV_X1 U16323 ( .A(n13858), .ZN(n12920) );
  NAND2_X1 U16324 ( .A1(n13929), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12921) );
  INV_X1 U16325 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14319) );
  XNOR2_X1 U16326 ( .A(n12921), .B(n14319), .ZN(n13957) );
  NOR2_X1 U16327 ( .A1(n13957), .A2(n20570), .ZN(n12922) );
  OR2_X1 U16328 ( .A1(n12934), .A2(n12923), .ZN(n12924) );
  OR2_X1 U16329 ( .A1(n12925), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12928) );
  NAND2_X1 U16330 ( .A1(n19747), .A2(n13915), .ZN(n14418) );
  NOR2_X1 U16331 ( .A1(n12934), .A2(n12927), .ZN(n19780) );
  INV_X1 U16332 ( .A(n19780), .ZN(n19762) );
  INV_X1 U16333 ( .A(n12928), .ZN(n12931) );
  NAND2_X1 U16334 ( .A1(n12929), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12932) );
  NAND2_X1 U16335 ( .A1(n12932), .A2(n19972), .ZN(n12930) );
  AND2_X1 U16336 ( .A1(n20666), .A2(n20055), .ZN(n12933) );
  AOI22_X1 U16337 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(n19774), .B1(n19773), .B2(
        n12935), .ZN(n12938) );
  AND2_X1 U16338 ( .A1(n13957), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12936) );
  OAI21_X1 U16339 ( .B1(n19779), .B2(n19778), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12937) );
  OAI211_X1 U16340 ( .C1(n19762), .C2(n14063), .A(n12938), .B(n12937), .ZN(
        n12939) );
  AOI21_X1 U16341 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n14418), .A(n12939), .ZN(
        n12940) );
  OAI21_X1 U16342 ( .B1(n12941), .B2(n19766), .A(n12940), .ZN(P1_U2840) );
  NAND2_X1 U16343 ( .A1(n20573), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12943) );
  NAND2_X1 U16344 ( .A1(n13900), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12942) );
  OAI211_X1 U16345 ( .C1(n12944), .C2(n15917), .A(n12943), .B(n12942), .ZN(
        n12949) );
  INV_X1 U16346 ( .A(n13100), .ZN(n12948) );
  INV_X1 U16347 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U16348 ( .A1(n12946), .A2(n12945), .ZN(n12947) );
  NAND2_X1 U16349 ( .A1(n12948), .A2(n12947), .ZN(n19911) );
  MUX2_X1 U16350 ( .A(n12949), .B(n19911), .S(n13946), .Z(n12950) );
  AOI21_X1 U16351 ( .B1(n12951), .B2(n13706), .A(n12950), .ZN(n13096) );
  XNOR2_X1 U16352 ( .A(n13097), .B(n13095), .ZN(n19907) );
  INV_X1 U16353 ( .A(n19907), .ZN(n13002) );
  INV_X1 U16354 ( .A(DATAI_4_), .ZN(n12953) );
  NAND2_X1 U16355 ( .A1(n19965), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12952) );
  OAI21_X1 U16356 ( .B1(n19965), .B2(n12953), .A(n12952), .ZN(n20002) );
  AOI22_X1 U16357 ( .A1(n15727), .A2(n20002), .B1(P1_EAX_REG_4__SCAN_IN), .B2(
        n14604), .ZN(n12954) );
  OAI21_X1 U16358 ( .B1(n13002), .B2(n9576), .A(n12954), .ZN(P1_U2900) );
  INV_X1 U16359 ( .A(n13915), .ZN(n19725) );
  AOI22_X1 U16360 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n19774), .B1(n19725), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n12960) );
  MUX2_X1 U16361 ( .A(n19778), .B(n19779), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n12957) );
  NAND2_X1 U16362 ( .A1(n15639), .A2(n12892), .ZN(n12966) );
  OAI21_X1 U16363 ( .B1(n19762), .B2(n12955), .A(n12966), .ZN(n12956) );
  AOI211_X1 U16364 ( .C1(n19773), .C2(n12958), .A(n12957), .B(n12956), .ZN(
        n12959) );
  OAI211_X1 U16365 ( .C1(n19766), .C2(n19921), .A(n12960), .B(n12959), .ZN(
        P1_U2839) );
  XNOR2_X1 U16366 ( .A(n13006), .B(n13007), .ZN(n12965) );
  OR2_X1 U16367 ( .A1(n12961), .A2(n12745), .ZN(n12962) );
  AND2_X1 U16368 ( .A1(n9677), .A2(n12962), .ZN(n18728) );
  INV_X1 U16369 ( .A(n18728), .ZN(n16062) );
  MUX2_X1 U16370 ( .A(n12963), .B(n16062), .S(n14918), .Z(n12964) );
  OAI21_X1 U16371 ( .B1(n12965), .B2(n14929), .A(n12964), .ZN(P2_U2874) );
  NAND2_X1 U16372 ( .A1(n12966), .A2(n13915), .ZN(n19775) );
  NAND2_X1 U16373 ( .A1(n19775), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U16374 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19779), .B1(
        n19778), .B2(n12967), .ZN(n12969) );
  NAND2_X1 U16375 ( .A1(n19774), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12968) );
  NAND3_X1 U16376 ( .A1(n12970), .A2(n12969), .A3(n12968), .ZN(n12972) );
  NAND2_X1 U16377 ( .A1(n15639), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19790) );
  OAI22_X1 U16378 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n19790), .B1(n19761), 
        .B2(n19954), .ZN(n12971) );
  AOI211_X1 U16379 ( .C1(n19780), .C2(n19975), .A(n12972), .B(n12971), .ZN(
        n12973) );
  OAI21_X1 U16380 ( .B1(n19766), .B2(n12974), .A(n12973), .ZN(P1_U2838) );
  INV_X1 U16381 ( .A(n12975), .ZN(n12976) );
  NAND2_X1 U16382 ( .A1(n12977), .A2(n12976), .ZN(n12978) );
  OAI21_X1 U16383 ( .B1(n12979), .B2(n12978), .A(n13961), .ZN(n18828) );
  INV_X1 U16384 ( .A(n19647), .ZN(n13086) );
  OR2_X1 U16385 ( .A1(n12981), .A2(n12980), .ZN(n12983) );
  NAND2_X1 U16386 ( .A1(n12983), .A2(n12982), .ZN(n19649) );
  XNOR2_X1 U16387 ( .A(n19647), .B(n19649), .ZN(n18910) );
  XNOR2_X1 U16388 ( .A(n19654), .B(n19658), .ZN(n18915) );
  INV_X1 U16389 ( .A(n12985), .ZN(n18924) );
  NAND2_X1 U16390 ( .A1(n19663), .A2(n18924), .ZN(n18923) );
  NAND2_X1 U16391 ( .A1(n18915), .A2(n18923), .ZN(n18914) );
  OAI21_X1 U16392 ( .B1(n19658), .B2(n18847), .A(n18914), .ZN(n18909) );
  NAND2_X1 U16393 ( .A1(n18910), .A2(n18909), .ZN(n18908) );
  OAI21_X1 U16394 ( .B1(n13086), .B2(n19649), .A(n18908), .ZN(n18903) );
  XNOR2_X1 U16395 ( .A(n19636), .B(n19640), .ZN(n18904) );
  NAND2_X1 U16396 ( .A1(n18903), .A2(n18904), .ZN(n18902) );
  OAI21_X1 U16397 ( .B1(n18901), .B2(n19636), .A(n18902), .ZN(n12986) );
  NAND2_X1 U16398 ( .A1(n12986), .A2(n18824), .ZN(n18898) );
  XOR2_X1 U16399 ( .A(n18828), .B(n18898), .Z(n12997) );
  NAND2_X1 U16400 ( .A1(n12988), .A2(n12987), .ZN(n12990) );
  INV_X1 U16401 ( .A(n18824), .ZN(n12992) );
  AOI22_X1 U16402 ( .A1(n18921), .A2(n12992), .B1(n18920), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n12996) );
  AND2_X1 U16403 ( .A1(n13985), .A2(n19050), .ZN(n12993) );
  AND2_X1 U16404 ( .A1(n19050), .A2(n19043), .ZN(n12994) );
  NAND2_X1 U16405 ( .A1(n15005), .A2(n13212), .ZN(n18874) );
  INV_X1 U16406 ( .A(n15004), .ZN(n13058) );
  NAND2_X1 U16407 ( .A1(n18874), .A2(n13058), .ZN(n12995) );
  OAI211_X1 U16408 ( .C1(n12997), .C2(n18868), .A(n12996), .B(n12995), .ZN(
        P2_U2915) );
  NAND2_X1 U16409 ( .A1(n12999), .A2(n12998), .ZN(n13000) );
  NAND2_X1 U16410 ( .A1(n13122), .A2(n13000), .ZN(n19928) );
  INV_X1 U16411 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13001) );
  OAI222_X1 U16412 ( .A1(n19928), .A2(n14528), .B1(n14530), .B2(n13002), .C1(
        n13001), .C2(n19797), .ZN(P1_U2868) );
  AND2_X1 U16413 ( .A1(n9677), .A2(n13004), .ZN(n13005) );
  OR2_X1 U16414 ( .A1(n13003), .A2(n13005), .ZN(n15313) );
  OAI211_X1 U16415 ( .C1(n9676), .C2(n13010), .A(n10036), .B(n14907), .ZN(
        n13012) );
  NAND2_X1 U16416 ( .A1(n12420), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13011) );
  OAI211_X1 U16417 ( .C1(n15313), .C2(n12420), .A(n13012), .B(n13011), .ZN(
        P2_U2873) );
  INV_X1 U16418 ( .A(n19087), .ZN(n19147) );
  OAI21_X1 U16419 ( .B1(n19216), .B2(n19220), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13020) );
  NAND2_X1 U16420 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n12670), .ZN(
        n19221) );
  INV_X1 U16421 ( .A(n19221), .ZN(n13013) );
  NAND2_X1 U16422 ( .A1(n13125), .A2(n13013), .ZN(n13019) );
  OAI21_X1 U16423 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n12317), .ZN(n16166) );
  INV_X1 U16424 ( .A(n16166), .ZN(n19684) );
  INV_X1 U16425 ( .A(n13014), .ZN(n13015) );
  NAND2_X1 U16426 ( .A1(n19684), .A2(n13015), .ZN(n13016) );
  NOR3_X2 U16427 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19489), .ZN(n19214) );
  AOI211_X1 U16428 ( .C1(n13023), .C2(n19639), .A(n19642), .B(n19214), .ZN(
        n13018) );
  INV_X1 U16429 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14098) );
  AOI22_X1 U16430 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19047), .ZN(n19398) );
  AOI22_X1 U16431 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19047), .ZN(n19505) );
  AOI22_X1 U16432 ( .A1(n19216), .A2(n19502), .B1(n19220), .B2(n19453), .ZN(
        n13027) );
  OAI21_X1 U16433 ( .B1(n13023), .B2(n19214), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13024) );
  OAI21_X1 U16434 ( .B1(n19221), .B2(n19305), .A(n13024), .ZN(n19215) );
  NAND2_X1 U16435 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19392), .ZN(n19033) );
  AND2_X1 U16436 ( .A1(n10217), .A2(n19049), .ZN(n19494) );
  AOI22_X1 U16437 ( .A1(n19215), .A2(n13025), .B1(n19494), .B2(n19214), .ZN(
        n13026) );
  OAI211_X1 U16438 ( .C1(n19219), .C2(n14098), .A(n13027), .B(n13026), .ZN(
        P2_U3096) );
  XNOR2_X1 U16439 ( .A(n13190), .B(n13189), .ZN(n13033) );
  INV_X1 U16440 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13031) );
  OR2_X1 U16441 ( .A1(n13003), .A2(n13029), .ZN(n13030) );
  NAND2_X1 U16442 ( .A1(n13028), .A2(n13030), .ZN(n18707) );
  MUX2_X1 U16443 ( .A(n13031), .B(n18707), .S(n14918), .Z(n13032) );
  OAI21_X1 U16444 ( .B1(n13033), .B2(n14929), .A(n13032), .ZN(P2_U2872) );
  INV_X1 U16445 ( .A(n19499), .ZN(n13035) );
  OAI21_X1 U16446 ( .B1(n13035), .B2(n19066), .A(n19642), .ZN(n13045) );
  INV_X1 U16447 ( .A(n13045), .ZN(n13039) );
  NAND2_X1 U16448 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19651), .ZN(
        n19334) );
  INV_X1 U16449 ( .A(n19334), .ZN(n19333) );
  NAND2_X1 U16450 ( .A1(n19333), .A2(n10817), .ZN(n13044) );
  INV_X1 U16451 ( .A(n13042), .ZN(n13036) );
  NAND2_X1 U16452 ( .A1(n13036), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13037) );
  NOR3_X2 U16453 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19666), .A3(
        n19334), .ZN(n19306) );
  AOI21_X1 U16454 ( .B1(n13037), .B2(n19639), .A(n19306), .ZN(n13038) );
  INV_X1 U16455 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13048) );
  NOR2_X2 U16456 ( .A1(n19395), .A2(n19066), .ZN(n19329) );
  INV_X1 U16457 ( .A(n19329), .ZN(n13056) );
  INV_X1 U16458 ( .A(n19494), .ZN(n19385) );
  INV_X1 U16459 ( .A(n19306), .ZN(n13055) );
  OAI22_X1 U16460 ( .A1(n19505), .A2(n13056), .B1(n19385), .B2(n13055), .ZN(
        n13041) );
  AOI21_X1 U16461 ( .B1(n19297), .B2(n19502), .A(n13041), .ZN(n13047) );
  OAI21_X1 U16462 ( .B1(n13042), .B2(n19306), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13043) );
  OAI21_X1 U16463 ( .B1(n13045), .B2(n13044), .A(n13043), .ZN(n19298) );
  NAND2_X1 U16464 ( .A1(n19298), .A2(n13025), .ZN(n13046) );
  OAI211_X1 U16465 ( .C1(n19302), .C2(n13048), .A(n13047), .B(n13046), .ZN(
        P2_U3120) );
  INV_X1 U16466 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16467 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19047), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19048), .ZN(n19404) );
  AOI22_X1 U16468 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19047), .ZN(n19510) );
  INV_X1 U16469 ( .A(n19506), .ZN(n19399) );
  OAI22_X1 U16470 ( .A1(n19510), .A2(n13056), .B1(n19399), .B2(n13055), .ZN(
        n13049) );
  AOI21_X1 U16471 ( .B1(n19297), .B2(n19507), .A(n13049), .ZN(n13052) );
  NAND2_X1 U16472 ( .A1(n19298), .A2(n13050), .ZN(n13051) );
  OAI211_X1 U16473 ( .C1(n19302), .C2(n13053), .A(n13052), .B(n13051), .ZN(
        P2_U3121) );
  INV_X1 U16474 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U16475 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19047), .ZN(n19422) );
  AOI22_X1 U16476 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19047), .ZN(n19526) );
  NAND2_X1 U16477 ( .A1(n13054), .A2(n19049), .ZN(n19417) );
  OAI22_X1 U16478 ( .A1(n19526), .A2(n13056), .B1(n13055), .B2(n19417), .ZN(
        n13057) );
  AOI21_X1 U16479 ( .B1(n19297), .B2(n19523), .A(n13057), .ZN(n13060) );
  NAND2_X1 U16480 ( .A1(n13058), .A2(n19392), .ZN(n19418) );
  NAND2_X1 U16481 ( .A1(n19298), .A2(n19522), .ZN(n13059) );
  OAI211_X1 U16482 ( .C1(n19302), .C2(n13061), .A(n13060), .B(n13059), .ZN(
        P2_U3124) );
  XNOR2_X1 U16483 ( .A(n13063), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13064) );
  XNOR2_X1 U16484 ( .A(n13062), .B(n13064), .ZN(n13145) );
  INV_X1 U16485 ( .A(n19945), .ZN(n13070) );
  NAND2_X1 U16486 ( .A1(n19924), .A2(n13065), .ZN(n15912) );
  INV_X1 U16487 ( .A(n13072), .ZN(n15870) );
  NOR2_X1 U16488 ( .A1(n15870), .A2(n19946), .ZN(n13068) );
  INV_X1 U16489 ( .A(n13066), .ZN(n13071) );
  OAI21_X1 U16490 ( .B1(n14823), .B2(n13071), .A(n13067), .ZN(n19923) );
  AOI211_X1 U16491 ( .C1(n19950), .C2(n13069), .A(n13068), .B(n19923), .ZN(
        n15907) );
  OAI21_X1 U16492 ( .B1(n13070), .B2(n15912), .A(n15907), .ZN(n15888) );
  AOI21_X1 U16493 ( .B1(n13071), .B2(n19945), .A(n14784), .ZN(n15869) );
  NOR2_X1 U16494 ( .A1(n15869), .A2(n13072), .ZN(n15892) );
  AOI22_X1 U16495 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15888), .B1(
        n15892), .B2(n15890), .ZN(n13075) );
  XOR2_X1 U16496 ( .A(n13073), .B(n9631), .Z(n13112) );
  INV_X1 U16497 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20600) );
  NOR2_X1 U16498 ( .A1(n19927), .A2(n20600), .ZN(n13139) );
  AOI21_X1 U16499 ( .B1(n13112), .B2(n19936), .A(n13139), .ZN(n13074) );
  OAI211_X1 U16500 ( .C1(n13145), .C2(n19925), .A(n13075), .B(n13074), .ZN(
        P1_U3025) );
  AOI22_X1 U16501 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18838), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n18856), .ZN(n13080) );
  AOI22_X1 U16502 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n18853), .B1(n13076), 
        .B2(n18852), .ZN(n13079) );
  NAND2_X1 U16503 ( .A1(n19005), .A2(n18854), .ZN(n13078) );
  NAND2_X1 U16504 ( .A1(n19649), .A2(n18855), .ZN(n13077) );
  NAND4_X1 U16505 ( .A1(n13080), .A2(n13079), .A3(n13078), .A4(n13077), .ZN(
        n13085) );
  INV_X1 U16506 ( .A(n13974), .ZN(n13083) );
  NOR2_X1 U16507 ( .A1(n18830), .A2(n13081), .ZN(n13180) );
  INV_X1 U16508 ( .A(n13180), .ZN(n13082) );
  AOI221_X1 U16509 ( .B1(n13083), .B2(n13180), .C1(n13974), .C2(n13082), .A(
        n19555), .ZN(n13084) );
  AOI211_X1 U16510 ( .C1(n13086), .C2(n18857), .A(n13085), .B(n13084), .ZN(
        n13087) );
  INV_X1 U16511 ( .A(n13087), .ZN(P2_U2853) );
  NAND2_X1 U16512 ( .A1(n13088), .A2(n13706), .ZN(n13094) );
  NAND2_X1 U16513 ( .A1(n13099), .A2(n13114), .ZN(n13090) );
  INV_X1 U16514 ( .A(n13221), .ZN(n13089) );
  NAND2_X1 U16515 ( .A1(n13090), .A2(n13089), .ZN(n13141) );
  NAND2_X1 U16516 ( .A1(n13141), .A2(n13797), .ZN(n13091) );
  OAI21_X1 U16517 ( .B1(n13114), .B2(n13670), .A(n13091), .ZN(n13092) );
  AOI21_X1 U16518 ( .B1(n13900), .B2(P1_EAX_REG_6__SCAN_IN), .A(n13092), .ZN(
        n13093) );
  NAND2_X1 U16519 ( .A1(n13094), .A2(n13093), .ZN(n13105) );
  INV_X1 U16520 ( .A(n13105), .ZN(n13108) );
  INV_X1 U16521 ( .A(n13098), .ZN(n13104) );
  INV_X1 U16522 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13102) );
  OAI21_X1 U16523 ( .B1(n13100), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13099), .ZN(n15791) );
  AOI22_X1 U16524 ( .A1(n15791), .A2(n13946), .B1(n13953), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13101) );
  OAI21_X1 U16525 ( .B1(n13793), .B2(n13102), .A(n13101), .ZN(n13103) );
  INV_X1 U16526 ( .A(n13106), .ZN(n13107) );
  AOI21_X1 U16527 ( .B1(n13108), .B2(n13107), .A(n13227), .ZN(n13143) );
  INV_X1 U16528 ( .A(n13143), .ZN(n13156) );
  AOI22_X1 U16529 ( .A1(n13112), .A2(n19792), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14520), .ZN(n13109) );
  OAI21_X1 U16530 ( .B1(n13156), .B2(n14530), .A(n13109), .ZN(P1_U2866) );
  NAND3_X1 U16531 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n13147) );
  NOR2_X1 U16532 ( .A1(n12892), .A2(n13147), .ZN(n13146) );
  NAND2_X1 U16533 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n13146), .ZN(n13111) );
  NOR2_X1 U16534 ( .A1(n20600), .A2(n13111), .ZN(n19749) );
  OAI21_X1 U16535 ( .B1(n19747), .B2(n19749), .A(n13915), .ZN(n19754) );
  OR2_X1 U16536 ( .A1(n19747), .A2(n19749), .ZN(n13110) );
  OAI22_X1 U16537 ( .A1(n13141), .A2(n19751), .B1(n13111), .B2(n13110), .ZN(
        n13116) );
  AOI22_X1 U16538 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n19774), .B1(n19773), .B2(
        n13112), .ZN(n13113) );
  OAI211_X1 U16539 ( .C1(n19728), .C2(n13114), .A(n13113), .B(n19927), .ZN(
        n13115) );
  AOI211_X1 U16540 ( .C1(P1_REIP_REG_6__SCAN_IN), .C2(n19754), .A(n13116), .B(
        n13115), .ZN(n13117) );
  OAI21_X1 U16541 ( .B1(n13156), .B2(n15657), .A(n13117), .ZN(P1_U2834) );
  AND2_X1 U16542 ( .A1(n13119), .A2(n13118), .ZN(n13120) );
  NOR2_X1 U16543 ( .A1(n13106), .A2(n13120), .ZN(n15788) );
  INV_X1 U16544 ( .A(n15788), .ZN(n13159) );
  INV_X1 U16545 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13124) );
  AND2_X1 U16546 ( .A1(n13122), .A2(n13121), .ZN(n13123) );
  OR2_X1 U16547 ( .A1(n13123), .A2(n9631), .ZN(n15905) );
  OAI222_X1 U16548 ( .A1(n13159), .A2(n14530), .B1(n13124), .B2(n19797), .C1(
        n14528), .C2(n15905), .ZN(P1_U2867) );
  NOR2_X2 U16549 ( .A1(n19395), .A2(n19303), .ZN(n19375) );
  OAI21_X1 U16550 ( .B1(n19380), .B2(n19375), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13130) );
  INV_X1 U16551 ( .A(n13125), .ZN(n13127) );
  NAND2_X1 U16552 ( .A1(n13127), .A2(n13126), .ZN(n19148) );
  OR2_X1 U16553 ( .A1(n12670), .A2(n19148), .ZN(n13129) );
  NAND3_X1 U16554 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n10817), .ZN(n19390) );
  NOR2_X1 U16555 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19390), .ZN(
        n19373) );
  AOI211_X1 U16556 ( .C1(n13132), .C2(n19639), .A(n19642), .B(n19373), .ZN(
        n13128) );
  INV_X1 U16557 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14105) );
  AOI22_X1 U16558 ( .A1(n19375), .A2(n19502), .B1(n19380), .B2(n19453), .ZN(
        n13136) );
  INV_X1 U16559 ( .A(n13131), .ZN(n13134) );
  OAI21_X1 U16560 ( .B1(n13132), .B2(n19373), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13133) );
  OAI21_X1 U16561 ( .B1(n13134), .B2(n19148), .A(n13133), .ZN(n19374) );
  AOI22_X1 U16562 ( .A1(n19374), .A2(n13025), .B1(n19494), .B2(n19373), .ZN(
        n13135) );
  OAI211_X1 U16563 ( .C1(n19379), .C2(n14105), .A(n13136), .B(n13135), .ZN(
        P2_U3144) );
  INV_X1 U16564 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14140) );
  AOI22_X1 U16565 ( .A1(n19375), .A2(n19507), .B1(n19380), .B2(n19461), .ZN(
        n13138) );
  AOI22_X1 U16566 ( .A1(n19374), .A2(n13050), .B1(n19373), .B2(n19506), .ZN(
        n13137) );
  OAI211_X1 U16567 ( .C1(n19379), .C2(n14140), .A(n13138), .B(n13137), .ZN(
        P2_U3145) );
  AOI21_X1 U16568 ( .B1(n19914), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13139), .ZN(n13140) );
  OAI21_X1 U16569 ( .B1(n19912), .B2(n13141), .A(n13140), .ZN(n13142) );
  AOI21_X1 U16570 ( .B1(n13143), .B2(n15781), .A(n13142), .ZN(n13144) );
  OAI21_X1 U16571 ( .B1(n13145), .B2(n19708), .A(n13144), .ZN(P1_U2993) );
  OAI21_X1 U16572 ( .B1(n19747), .B2(n13146), .A(n13915), .ZN(n19767) );
  NOR3_X1 U16573 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n13147), .A3(n19790), .ZN(
        n13149) );
  NOR2_X1 U16574 ( .A1(n15791), .A2(n19751), .ZN(n13148) );
  AOI211_X1 U16575 ( .C1(n19767), .C2(P1_REIP_REG_5__SCAN_IN), .A(n13149), .B(
        n13148), .ZN(n13153) );
  AOI22_X1 U16576 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(n19774), .ZN(n13150) );
  OAI211_X1 U16577 ( .C1(n19761), .C2(n15905), .A(n19927), .B(n13150), .ZN(
        n13151) );
  INV_X1 U16578 ( .A(n13151), .ZN(n13152) );
  OAI211_X1 U16579 ( .C1(n19766), .C2(n13159), .A(n13153), .B(n13152), .ZN(
        P1_U2835) );
  INV_X1 U16580 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19873) );
  INV_X1 U16581 ( .A(DATAI_6_), .ZN(n13155) );
  NAND2_X1 U16582 ( .A1(n19965), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13154) );
  OAI21_X1 U16583 ( .B1(n19965), .B2(n13155), .A(n13154), .ZN(n19871) );
  INV_X1 U16584 ( .A(n19871), .ZN(n20010) );
  OAI222_X1 U16585 ( .A1(n13156), .A2(n9576), .B1(n15730), .B2(n19873), .C1(
        n14601), .C2(n20010), .ZN(P1_U2898) );
  INV_X1 U16586 ( .A(DATAI_5_), .ZN(n13158) );
  NAND2_X1 U16587 ( .A1(n19965), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13157) );
  OAI21_X1 U16588 ( .B1(n19965), .B2(n13158), .A(n13157), .ZN(n19869) );
  INV_X1 U16589 ( .A(n19869), .ZN(n20006) );
  OAI222_X1 U16590 ( .A1(n9576), .A2(n13159), .B1(n20006), .B2(n14601), .C1(
        n15730), .C2(n13102), .ZN(P1_U2899) );
  OAI21_X1 U16591 ( .B1(n13161), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13160), .ZN(n13179) );
  XOR2_X1 U16592 ( .A(n13162), .B(n13164), .Z(n13177) );
  INV_X1 U16593 ( .A(n13268), .ZN(n16160) );
  AOI21_X1 U16594 ( .B1(n15263), .B2(n16160), .A(n16151), .ZN(n13267) );
  NAND3_X1 U16595 ( .A1(n13268), .A2(n16161), .A3(n13166), .ZN(n13266) );
  NAND2_X1 U16596 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n18980), .ZN(n13165) );
  OAI211_X1 U16597 ( .C1(n13267), .C2(n13166), .A(n13266), .B(n13165), .ZN(
        n13171) );
  OAI21_X1 U16598 ( .B1(n13169), .B2(n13168), .A(n13167), .ZN(n18804) );
  OAI22_X1 U16599 ( .A1(n13175), .A2(n16158), .B1(n18995), .B2(n18804), .ZN(
        n13170) );
  AOI211_X1 U16600 ( .C1(n13177), .C2(n18999), .A(n13171), .B(n13170), .ZN(
        n13172) );
  OAI21_X1 U16601 ( .B1(n18994), .B2(n13179), .A(n13172), .ZN(P2_U3040) );
  OAI22_X1 U16602 ( .A1(n10855), .A2(n19016), .B1(n18992), .B2(n18799), .ZN(
        n13173) );
  AOI21_X1 U16603 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18979), .A(
        n13173), .ZN(n13174) );
  OAI21_X1 U16604 ( .B1(n16117), .B2(n13175), .A(n13174), .ZN(n13176) );
  AOI21_X1 U16605 ( .B1(n13177), .B2(n16102), .A(n13176), .ZN(n13178) );
  OAI21_X1 U16606 ( .B1(n18984), .B2(n13179), .A(n13178), .ZN(P2_U3008) );
  OAI21_X1 U16607 ( .B1(n13183), .B2(n13181), .A(n13180), .ZN(n18850) );
  OAI21_X1 U16608 ( .B1(n18814), .B2(n13182), .A(n18850), .ZN(n15411) );
  INV_X1 U16609 ( .A(n13183), .ZN(n18858) );
  AOI22_X1 U16610 ( .A1(n18830), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18858), .B2(n18814), .ZN(n15404) );
  NOR2_X1 U16611 ( .A1(n15404), .A2(n13184), .ZN(n15409) );
  INV_X1 U16612 ( .A(n16167), .ZN(n15413) );
  INV_X1 U16613 ( .A(n19634), .ZN(n15526) );
  OAI22_X1 U16614 ( .A1(n19647), .A2(n15413), .B1(n13185), .B2(n15526), .ZN(
        n13186) );
  AOI21_X1 U16615 ( .B1(n15411), .B2(n15409), .A(n13186), .ZN(n13187) );
  MUX2_X1 U16616 ( .A(n13187), .B(n12581), .S(n15414), .Z(n13188) );
  INV_X1 U16617 ( .A(n13188), .ZN(P2_U3599) );
  AOI22_X1 U16618 ( .A1(n10344), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U16619 ( .A1(n10432), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U16620 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13192) );
  AOI22_X1 U16621 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13191) );
  NAND4_X1 U16622 ( .A1(n13194), .A2(n13193), .A3(n13192), .A4(n13191), .ZN(
        n13201) );
  AOI22_X1 U16623 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U16624 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U16625 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14122), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13197) );
  AOI22_X1 U16626 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13196) );
  NAND4_X1 U16627 ( .A1(n13199), .A2(n13198), .A3(n13197), .A4(n13196), .ZN(
        n13200) );
  NAND2_X1 U16628 ( .A1(n9580), .A2(n13465), .ZN(n13355) );
  OAI21_X1 U16629 ( .B1(n9580), .B2(n13465), .A(n13355), .ZN(n13219) );
  NAND2_X1 U16630 ( .A1(n13028), .A2(n13203), .ZN(n13204) );
  NAND2_X1 U16631 ( .A1(n13339), .A2(n13204), .ZN(n18695) );
  NOR2_X1 U16632 ( .A1(n18695), .A2(n12420), .ZN(n13205) );
  AOI21_X1 U16633 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n12420), .A(n13205), .ZN(
        n13206) );
  OAI21_X1 U16634 ( .B1(n13219), .B2(n14929), .A(n13206), .ZN(P2_U2871) );
  NOR2_X1 U16635 ( .A1(n13208), .A2(n9662), .ZN(n13209) );
  OR2_X1 U16636 ( .A1(n13207), .A2(n13209), .ZN(n18696) );
  INV_X1 U16637 ( .A(n18696), .ZN(n13217) );
  OAI22_X1 U16638 ( .A1(n15005), .A2(n18928), .B1(n18892), .B2(n13210), .ZN(
        n13216) );
  INV_X1 U16639 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n13214) );
  INV_X1 U16640 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n13213) );
  OAI22_X1 U16641 ( .A1(n15008), .A2(n13214), .B1(n15006), .B2(n13213), .ZN(
        n13215) );
  AOI211_X1 U16642 ( .C1(n18921), .C2(n13217), .A(n13216), .B(n13215), .ZN(
        n13218) );
  OAI21_X1 U16643 ( .B1(n13219), .B2(n18868), .A(n13218), .ZN(P2_U2903) );
  NAND2_X1 U16644 ( .A1(n13220), .A2(n13706), .ZN(n13226) );
  INV_X1 U16645 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13223) );
  OAI21_X1 U16646 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13221), .A(
        n13289), .ZN(n19752) );
  NAND2_X1 U16647 ( .A1(n19752), .A2(n13797), .ZN(n13222) );
  OAI21_X1 U16648 ( .B1(n13223), .B2(n13670), .A(n13222), .ZN(n13224) );
  AOI21_X1 U16649 ( .B1(n13900), .B2(P1_EAX_REG_7__SCAN_IN), .A(n13224), .ZN(
        n13225) );
  NAND2_X1 U16650 ( .A1(n13226), .A2(n13225), .ZN(n13228) );
  OR2_X1 U16651 ( .A1(n13227), .A2(n13228), .ZN(n13229) );
  AND2_X1 U16652 ( .A1(n13297), .A2(n13229), .ZN(n19756) );
  OR2_X1 U16653 ( .A1(n13232), .A2(n13231), .ZN(n13233) );
  NAND2_X1 U16654 ( .A1(n13230), .A2(n13233), .ZN(n19750) );
  OAI22_X1 U16655 ( .A1(n19750), .A2(n14528), .B1(n13234), .B2(n19797), .ZN(
        n13235) );
  AOI21_X1 U16656 ( .B1(n19756), .B2(n19793), .A(n13235), .ZN(n13236) );
  INV_X1 U16657 ( .A(n13236), .ZN(P1_U2865) );
  INV_X1 U16658 ( .A(n13355), .ZN(n13432) );
  AOI22_X1 U16659 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13240) );
  AOI22_X1 U16660 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10384), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U16661 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U16662 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13237) );
  NAND4_X1 U16663 ( .A1(n13240), .A2(n13239), .A3(n13238), .A4(n13237), .ZN(
        n13246) );
  AOI22_X1 U16664 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10437), .B1(
        n14120), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16665 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n14121), .ZN(n13243) );
  AOI22_X1 U16666 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14122), .ZN(n13242) );
  AOI22_X1 U16667 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13241) );
  NAND4_X1 U16668 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        n13245) );
  NOR2_X1 U16669 ( .A1(n13246), .A2(n13245), .ZN(n13354) );
  INV_X1 U16670 ( .A(n13354), .ZN(n13247) );
  OR2_X1 U16671 ( .A1(n13355), .A2(n13354), .ZN(n13356) );
  OAI21_X1 U16672 ( .B1(n13432), .B2(n13247), .A(n13356), .ZN(n13343) );
  NOR2_X1 U16673 ( .A1(n13207), .A2(n13248), .ZN(n13249) );
  NOR2_X1 U16674 ( .A1(n13385), .A2(n13249), .ZN(n18681) );
  OAI22_X1 U16675 ( .A1(n15005), .A2(n18919), .B1(n18892), .B2(n13250), .ZN(
        n13254) );
  INV_X1 U16676 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13252) );
  INV_X1 U16677 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n13251) );
  OAI22_X1 U16678 ( .A1(n15008), .A2(n13252), .B1(n15006), .B2(n13251), .ZN(
        n13253) );
  AOI211_X1 U16679 ( .C1(n18921), .C2(n18681), .A(n13254), .B(n13253), .ZN(
        n13255) );
  OAI21_X1 U16680 ( .B1(n13343), .B2(n18868), .A(n13255), .ZN(P2_U2902) );
  INV_X1 U16681 ( .A(n19756), .ZN(n13258) );
  INV_X1 U16682 ( .A(DATAI_7_), .ZN(n13257) );
  NAND2_X1 U16683 ( .A1(n19965), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13256) );
  OAI21_X1 U16684 ( .B1(n19965), .B2(n13257), .A(n13256), .ZN(n19874) );
  INV_X1 U16685 ( .A(n19874), .ZN(n20019) );
  INV_X1 U16686 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n19876) );
  OAI222_X1 U16687 ( .A1(n9576), .A2(n13258), .B1(n20019), .B2(n14601), .C1(
        n15730), .C2(n19876), .ZN(P1_U2897) );
  NAND2_X1 U16688 ( .A1(n13309), .A2(n13310), .ZN(n13260) );
  XNOR2_X1 U16689 ( .A(n13259), .B(n13260), .ZN(n16103) );
  INV_X1 U16690 ( .A(n16103), .ZN(n13278) );
  INV_X1 U16691 ( .A(n13261), .ZN(n13263) );
  NAND2_X1 U16692 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  XNOR2_X1 U16693 ( .A(n13265), .B(n13264), .ZN(n16100) );
  NAND2_X1 U16694 ( .A1(n16100), .A2(n16154), .ZN(n13277) );
  NAND2_X1 U16695 ( .A1(n13267), .A2(n13266), .ZN(n13320) );
  NAND3_X1 U16696 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13268), .A3(
        n16161), .ZN(n13316) );
  XNOR2_X1 U16697 ( .A(n13270), .B(n13269), .ZN(n18891) );
  INV_X1 U16698 ( .A(n18891), .ZN(n13272) );
  NOR2_X1 U16699 ( .A1(n10861), .A2(n19016), .ZN(n13271) );
  AOI21_X1 U16700 ( .B1(n16150), .B2(n13272), .A(n13271), .ZN(n13274) );
  INV_X1 U16701 ( .A(n18793), .ZN(n16101) );
  NAND2_X1 U16702 ( .A1(n16101), .A2(n19004), .ZN(n13273) );
  OAI211_X1 U16703 ( .C1(n13316), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n13274), .B(n13273), .ZN(n13275) );
  AOI21_X1 U16704 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n13320), .A(
        n13275), .ZN(n13276) );
  OAI211_X1 U16705 ( .C1(n13278), .C2(n16152), .A(n13277), .B(n13276), .ZN(
        P2_U3039) );
  AOI22_X1 U16706 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U16707 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16708 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U16709 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13279) );
  NAND4_X1 U16710 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n13288) );
  AOI22_X1 U16711 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13286) );
  AOI22_X1 U16712 ( .A1(n13861), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11574), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13285) );
  AOI22_X1 U16713 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13284) );
  AOI22_X1 U16714 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13283) );
  NAND4_X1 U16715 ( .A1(n13286), .A2(n13285), .A3(n13284), .A4(n13283), .ZN(
        n13287) );
  OAI21_X1 U16716 ( .B1(n13288), .B2(n13287), .A(n13706), .ZN(n13294) );
  XNOR2_X1 U16717 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n13289), .ZN(
        n19739) );
  INV_X1 U16718 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13290) );
  OAI22_X1 U16719 ( .A1(n19739), .A2(n13952), .B1(n13670), .B2(n13290), .ZN(
        n13291) );
  INV_X1 U16720 ( .A(n13291), .ZN(n13293) );
  NAND2_X1 U16721 ( .A1(n13900), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13292) );
  NAND2_X1 U16722 ( .A1(n13297), .A2(n13296), .ZN(n13298) );
  AND2_X1 U16723 ( .A1(n13379), .A2(n13298), .ZN(n19743) );
  INV_X1 U16724 ( .A(n19743), .ZN(n13306) );
  INV_X1 U16725 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13302) );
  INV_X1 U16726 ( .A(n13230), .ZN(n13301) );
  INV_X1 U16727 ( .A(n13299), .ZN(n13300) );
  OAI21_X1 U16728 ( .B1(n13301), .B2(n13300), .A(n9751), .ZN(n19741) );
  OAI222_X1 U16729 ( .A1(n13306), .A2(n14530), .B1(n19797), .B2(n13302), .C1(
        n19741), .C2(n14528), .ZN(P1_U2864) );
  INV_X1 U16730 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13305) );
  INV_X1 U16731 ( .A(DATAI_8_), .ZN(n20783) );
  NAND2_X1 U16732 ( .A1(n19966), .A2(n20783), .ZN(n13304) );
  INV_X1 U16733 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16256) );
  NAND2_X1 U16734 ( .A1(n19965), .A2(n16256), .ZN(n13303) );
  AND2_X1 U16735 ( .A1(n13304), .A2(n13303), .ZN(n19877) );
  INV_X1 U16736 ( .A(n19877), .ZN(n14564) );
  OAI222_X1 U16737 ( .A1(n13306), .A2(n9576), .B1(n13305), .B2(n15730), .C1(
        n14564), .C2(n14601), .ZN(P1_U2896) );
  XNOR2_X1 U16738 ( .A(n13308), .B(n13307), .ZN(n16096) );
  NAND2_X1 U16739 ( .A1(n13259), .A2(n13309), .ZN(n13311) );
  NAND2_X1 U16740 ( .A1(n13311), .A2(n13310), .ZN(n13315) );
  AND2_X1 U16741 ( .A1(n13313), .A2(n13312), .ZN(n13314) );
  XNOR2_X1 U16742 ( .A(n13315), .B(n13314), .ZN(n16095) );
  NOR2_X1 U16743 ( .A1(n10875), .A2(n19016), .ZN(n13319) );
  AOI221_X1 U16744 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(n11169), .C2(n13317), .A(
        n13316), .ZN(n13318) );
  AOI211_X1 U16745 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n13320), .A(
        n13319), .B(n13318), .ZN(n13327) );
  OR2_X1 U16746 ( .A1(n13322), .A2(n13321), .ZN(n13324) );
  NAND2_X1 U16747 ( .A1(n13324), .A2(n13323), .ZN(n18889) );
  INV_X1 U16748 ( .A(n18889), .ZN(n13325) );
  AOI22_X1 U16749 ( .A1(n19004), .A2(n18783), .B1(n16150), .B2(n13325), .ZN(
        n13326) );
  OAI211_X1 U16750 ( .C1(n16095), .C2(n16152), .A(n13327), .B(n13326), .ZN(
        n13328) );
  INV_X1 U16751 ( .A(n13328), .ZN(n13329) );
  OAI21_X1 U16752 ( .B1(n16096), .B2(n18994), .A(n13329), .ZN(P2_U3038) );
  XNOR2_X1 U16753 ( .A(n13331), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13332) );
  XNOR2_X1 U16754 ( .A(n13330), .B(n13332), .ZN(n15891) );
  INV_X1 U16755 ( .A(n19739), .ZN(n13334) );
  INV_X2 U16756 ( .A(n19927), .ZN(n19913) );
  AOI22_X1 U16757 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13333) );
  OAI21_X1 U16758 ( .B1(n19912), .B2(n13334), .A(n13333), .ZN(n13335) );
  AOI21_X1 U16759 ( .B1(n19743), .B2(n15781), .A(n13335), .ZN(n13336) );
  OAI21_X1 U16760 ( .B1(n15891), .B2(n19708), .A(n13336), .ZN(P1_U2991) );
  NAND2_X1 U16761 ( .A1(n13339), .A2(n13338), .ZN(n13340) );
  NAND2_X1 U16762 ( .A1(n13337), .A2(n13340), .ZN(n18688) );
  NOR2_X1 U16763 ( .A1(n18688), .A2(n12420), .ZN(n13341) );
  AOI21_X1 U16764 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n12420), .A(n13341), .ZN(
        n13342) );
  OAI21_X1 U16765 ( .B1(n13343), .B2(n14929), .A(n13342), .ZN(P2_U2870) );
  AOI22_X1 U16766 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10864), .B1(
        n10344), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13347) );
  AOI22_X1 U16767 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10432), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U16768 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13345) );
  AOI22_X1 U16769 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13344) );
  NAND4_X1 U16770 ( .A1(n13347), .A2(n13346), .A3(n13345), .A4(n13344), .ZN(
        n13353) );
  AOI22_X1 U16771 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10437), .B1(
        n14120), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13351) );
  AOI22_X1 U16772 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n14121), .ZN(n13350) );
  AOI22_X1 U16773 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n14122), .ZN(n13349) );
  AOI22_X1 U16774 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13348) );
  NAND4_X1 U16775 ( .A1(n13351), .A2(n13350), .A3(n13349), .A4(n13348), .ZN(
        n13352) );
  NOR2_X1 U16776 ( .A1(n13353), .A2(n13352), .ZN(n13357) );
  OR2_X1 U16777 ( .A1(n13357), .A2(n13354), .ZN(n13430) );
  NOR2_X1 U16778 ( .A1(n13355), .A2(n13430), .ZN(n13435) );
  AOI21_X1 U16779 ( .B1(n13357), .B2(n13356), .A(n13435), .ZN(n13358) );
  INV_X1 U16780 ( .A(n13358), .ZN(n13394) );
  NAND2_X1 U16781 ( .A1(n13337), .A2(n13359), .ZN(n13360) );
  AND2_X1 U16782 ( .A1(n9622), .A2(n13360), .ZN(n18673) );
  NOR2_X1 U16783 ( .A1(n14918), .A2(n18667), .ZN(n13361) );
  AOI21_X1 U16784 ( .B1(n18673), .B2(n14918), .A(n13361), .ZN(n13362) );
  OAI21_X1 U16785 ( .B1(n13394), .B2(n14929), .A(n13362), .ZN(P2_U2869) );
  XOR2_X1 U16786 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n13363), .Z(n19726) );
  AOI22_X1 U16787 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U16788 ( .A1(n13861), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11574), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U16789 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U16790 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13364) );
  NAND4_X1 U16791 ( .A1(n13367), .A2(n13366), .A3(n13365), .A4(n13364), .ZN(
        n13373) );
  AOI22_X1 U16792 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13371) );
  AOI22_X1 U16793 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13370) );
  AOI22_X1 U16794 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13369) );
  AOI22_X1 U16795 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13368) );
  NAND4_X1 U16796 ( .A1(n13371), .A2(n13370), .A3(n13369), .A4(n13368), .ZN(
        n13372) );
  NOR2_X1 U16797 ( .A1(n13373), .A2(n13372), .ZN(n13376) );
  NAND2_X1 U16798 ( .A1(n13900), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13375) );
  NAND2_X1 U16799 ( .A1(n13953), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13374) );
  OAI211_X1 U16800 ( .C1(n13607), .C2(n13376), .A(n13375), .B(n13374), .ZN(
        n13377) );
  AOI21_X1 U16801 ( .B1(n19726), .B2(n13946), .A(n13377), .ZN(n13378) );
  AND2_X1 U16802 ( .A1(n13379), .A2(n13378), .ZN(n13380) );
  OR2_X1 U16803 ( .A1(n13380), .A2(n13409), .ZN(n13450) );
  INV_X1 U16804 ( .A(DATAI_9_), .ZN(n13382) );
  NAND2_X1 U16805 ( .A1(n19965), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13381) );
  OAI21_X1 U16806 ( .B1(n19965), .B2(n13382), .A(n13381), .ZN(n19879) );
  AOI22_X1 U16807 ( .A1(n15727), .A2(n19879), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14604), .ZN(n13383) );
  OAI21_X1 U16808 ( .B1(n13450), .B2(n9576), .A(n13383), .ZN(P1_U2895) );
  OR2_X1 U16809 ( .A1(n13385), .A2(n13384), .ZN(n13386) );
  NAND2_X1 U16810 ( .A1(n13386), .A2(n13436), .ZN(n18676) );
  INV_X1 U16811 ( .A(n18676), .ZN(n13392) );
  OAI22_X1 U16812 ( .A1(n15005), .A2(n19029), .B1(n18892), .B2(n13387), .ZN(
        n13391) );
  INV_X1 U16813 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n13389) );
  INV_X1 U16814 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n13388) );
  OAI22_X1 U16815 ( .A1(n15008), .A2(n13389), .B1(n15006), .B2(n13388), .ZN(
        n13390) );
  AOI211_X1 U16816 ( .C1(n18921), .C2(n13392), .A(n13391), .B(n13390), .ZN(
        n13393) );
  OAI21_X1 U16817 ( .B1(n13394), .B2(n18868), .A(n13393), .ZN(P2_U2901) );
  AOI22_X1 U16818 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U16819 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13397) );
  AOI22_X1 U16820 ( .A1(n13861), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U16821 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13395) );
  NAND4_X1 U16822 ( .A1(n13398), .A2(n13397), .A3(n13396), .A4(n13395), .ZN(
        n13404) );
  AOI22_X1 U16823 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U16824 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13401) );
  AOI22_X1 U16825 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13400) );
  AOI22_X1 U16826 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13399) );
  NAND4_X1 U16827 ( .A1(n13402), .A2(n13401), .A3(n13400), .A4(n13399), .ZN(
        n13403) );
  NOR2_X1 U16828 ( .A1(n13404), .A2(n13403), .ZN(n13408) );
  XNOR2_X1 U16829 ( .A(n13405), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14713) );
  NAND2_X1 U16830 ( .A1(n14713), .A2(n13946), .ZN(n13407) );
  AOI22_X1 U16831 ( .A1(n13900), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13953), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13406) );
  OAI211_X1 U16832 ( .C1(n13408), .C2(n13607), .A(n13407), .B(n13406), .ZN(
        n13410) );
  OAI21_X1 U16833 ( .B1(n13409), .B2(n13410), .A(n13561), .ZN(n13475) );
  INV_X1 U16834 ( .A(DATAI_10_), .ZN(n13412) );
  NAND2_X1 U16835 ( .A1(n19965), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13411) );
  OAI21_X1 U16836 ( .B1(n19965), .B2(n13412), .A(n13411), .ZN(n19882) );
  AOI22_X1 U16837 ( .A1(n15727), .A2(n19882), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14604), .ZN(n13413) );
  OAI21_X1 U16838 ( .B1(n13475), .B2(n9576), .A(n13413), .ZN(P1_U2894) );
  AOI22_X1 U16839 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U16840 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10432), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U16841 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U16842 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13414) );
  NAND4_X1 U16843 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13429) );
  AOI22_X1 U16844 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n14121), .ZN(n13427) );
  OAI22_X1 U16845 ( .A1(n13419), .A2(n9623), .B1(n13418), .B2(n14185), .ZN(
        n13423) );
  INV_X1 U16846 ( .A(n14123), .ZN(n13421) );
  INV_X1 U16847 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14183) );
  INV_X1 U16848 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n20809) );
  INV_X1 U16849 ( .A(n14122), .ZN(n13420) );
  OAI22_X1 U16850 ( .A1(n13421), .A2(n14183), .B1(n20809), .B2(n13420), .ZN(
        n13422) );
  NOR2_X1 U16851 ( .A1(n13423), .A2(n13422), .ZN(n13426) );
  NAND2_X1 U16852 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13425) );
  NAND2_X1 U16853 ( .A1(n10437), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13424) );
  NAND4_X1 U16854 ( .A1(n13427), .A2(n13426), .A3(n13425), .A4(n13424), .ZN(
        n13428) );
  OR2_X1 U16855 ( .A1(n13429), .A2(n13428), .ZN(n13434) );
  INV_X1 U16856 ( .A(n13434), .ZN(n13431) );
  NOR2_X1 U16857 ( .A1(n13431), .A2(n13430), .ZN(n13464) );
  AND2_X1 U16858 ( .A1(n13432), .A2(n13464), .ZN(n13470) );
  INV_X1 U16859 ( .A(n13470), .ZN(n13433) );
  OAI21_X1 U16860 ( .B1(n13435), .B2(n13434), .A(n13433), .ZN(n14930) );
  XNOR2_X1 U16861 ( .A(n13437), .B(n13436), .ZN(n18665) );
  INV_X1 U16862 ( .A(n18665), .ZN(n13443) );
  OAI22_X1 U16863 ( .A1(n15005), .A2(n19034), .B1(n18892), .B2(n13438), .ZN(
        n13442) );
  INV_X1 U16864 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n13440) );
  INV_X1 U16865 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n13439) );
  OAI22_X1 U16866 ( .A1(n15008), .A2(n13440), .B1(n15006), .B2(n13439), .ZN(
        n13441) );
  AOI211_X1 U16867 ( .C1(n18921), .C2(n13443), .A(n13442), .B(n13441), .ZN(
        n13444) );
  OAI21_X1 U16868 ( .B1(n14930), .B2(n18868), .A(n13444), .ZN(P2_U2900) );
  INV_X1 U16869 ( .A(n13446), .ZN(n13448) );
  NOR2_X1 U16870 ( .A1(n13448), .A2(n13447), .ZN(n13449) );
  XNOR2_X1 U16871 ( .A(n13445), .B(n13449), .ZN(n15878) );
  AOI22_X1 U16872 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n13451) );
  OAI21_X1 U16873 ( .B1(n19912), .B2(n19726), .A(n13451), .ZN(n13452) );
  AOI21_X1 U16874 ( .B1(n19794), .B2(n15781), .A(n13452), .ZN(n13453) );
  OAI21_X1 U16875 ( .B1(n15878), .B2(n19708), .A(n13453), .ZN(P1_U2990) );
  AOI22_X1 U16876 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U16877 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10432), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U16878 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U16879 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13454) );
  NAND4_X1 U16880 ( .A1(n13457), .A2(n13456), .A3(n13455), .A4(n13454), .ZN(
        n13463) );
  AOI22_X1 U16881 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10437), .B1(
        n14120), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13461) );
  AOI22_X1 U16882 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n14121), .ZN(n13460) );
  AOI22_X1 U16883 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n14122), .ZN(n13459) );
  AOI22_X1 U16884 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13458) );
  NAND4_X1 U16885 ( .A1(n13461), .A2(n13460), .A3(n13459), .A4(n13458), .ZN(
        n13462) );
  OR2_X1 U16886 ( .A1(n13463), .A2(n13462), .ZN(n13469) );
  AND2_X1 U16887 ( .A1(n13469), .A2(n13464), .ZN(n13466) );
  AND2_X1 U16888 ( .A1(n13466), .A2(n13465), .ZN(n13467) );
  NAND2_X1 U16889 ( .A1(n13468), .A2(n13467), .ZN(n14068) );
  OAI21_X1 U16890 ( .B1(n13470), .B2(n13469), .A(n14068), .ZN(n15013) );
  INV_X1 U16891 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n13473) );
  OAI21_X1 U16892 ( .B1(n14925), .B2(n13472), .A(n13471), .ZN(n15081) );
  MUX2_X1 U16893 ( .A(n13473), .B(n15081), .S(n14918), .Z(n13474) );
  OAI21_X1 U16894 ( .B1(n15013), .B2(n14929), .A(n13474), .ZN(P2_U2867) );
  INV_X1 U16895 ( .A(n13475), .ZN(n14715) );
  AND2_X1 U16896 ( .A1(n15881), .A2(n13476), .ZN(n13477) );
  OR2_X1 U16897 ( .A1(n13477), .A2(n13510), .ZN(n15874) );
  OAI22_X1 U16898 ( .A1(n15874), .A2(n14528), .B1(n13478), .B2(n19797), .ZN(
        n13479) );
  AOI21_X1 U16899 ( .B1(n14715), .B2(n19793), .A(n13479), .ZN(n13480) );
  INV_X1 U16900 ( .A(n13480), .ZN(P1_U2862) );
  INV_X1 U16901 ( .A(n13482), .ZN(n13483) );
  NAND2_X1 U16902 ( .A1(n13481), .A2(n13483), .ZN(n14672) );
  NAND2_X1 U16903 ( .A1(n13484), .A2(n14672), .ZN(n14684) );
  NAND2_X1 U16904 ( .A1(n14684), .A2(n13485), .ZN(n13487) );
  AOI22_X1 U16905 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n14814), .B2(n14777), .ZN(n13486) );
  XNOR2_X1 U16906 ( .A(n13487), .B(n13486), .ZN(n15763) );
  XNOR2_X1 U16907 ( .A(n10083), .B(n14513), .ZN(n15714) );
  INV_X1 U16908 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20612) );
  NOR2_X1 U16909 ( .A1(n19927), .A2(n20612), .ZN(n13492) );
  AOI21_X1 U16910 ( .B1(n14784), .B2(n13488), .A(n19948), .ZN(n13489) );
  OAI21_X1 U16911 ( .B1(n14823), .B2(n13490), .A(n13489), .ZN(n15850) );
  MUX2_X1 U16912 ( .A(n14813), .B(n15850), .S(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n13491) );
  AOI211_X1 U16913 ( .C1(n19936), .C2(n15714), .A(n13492), .B(n13491), .ZN(
        n13493) );
  OAI21_X1 U16914 ( .B1(n15763), .B2(n19925), .A(n13493), .ZN(P1_U3017) );
  INV_X1 U16915 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13496) );
  OAI21_X1 U16916 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13494), .A(
        n13587), .ZN(n15776) );
  NAND2_X1 U16917 ( .A1(n15776), .A2(n13797), .ZN(n13495) );
  OAI21_X1 U16918 ( .B1(n13496), .B2(n13670), .A(n13495), .ZN(n13497) );
  AOI21_X1 U16919 ( .B1(n13900), .B2(P1_EAX_REG_11__SCAN_IN), .A(n13497), .ZN(
        n13498) );
  AOI21_X1 U16920 ( .B1(n13498), .B2(n13561), .A(n9625), .ZN(n14430) );
  AOI22_X1 U16921 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13502) );
  AOI22_X1 U16922 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11574), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13501) );
  AOI22_X1 U16923 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13500) );
  AOI22_X1 U16924 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13499) );
  NAND4_X1 U16925 ( .A1(n13502), .A2(n13501), .A3(n13500), .A4(n13499), .ZN(
        n13508) );
  AOI22_X1 U16926 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13506) );
  AOI22_X1 U16927 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13505) );
  AOI22_X1 U16928 ( .A1(n13879), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13504) );
  AOI22_X1 U16929 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13503) );
  NAND4_X1 U16930 ( .A1(n13506), .A2(n13505), .A3(n13504), .A4(n13503), .ZN(
        n13507) );
  OR2_X1 U16931 ( .A1(n13508), .A2(n13507), .ZN(n13509) );
  NAND2_X1 U16932 ( .A1(n13706), .A2(n13509), .ZN(n14429) );
  XNOR2_X1 U16933 ( .A(n14430), .B(n14429), .ZN(n15773) );
  INV_X1 U16934 ( .A(n15773), .ZN(n13518) );
  INV_X1 U16935 ( .A(n13510), .ZN(n13512) );
  INV_X1 U16936 ( .A(n14526), .ZN(n13511) );
  AOI21_X1 U16937 ( .B1(n13513), .B2(n13512), .A(n13511), .ZN(n15859) );
  AOI22_X1 U16938 ( .A1(n15859), .A2(n19792), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14520), .ZN(n13514) );
  OAI21_X1 U16939 ( .B1(n13518), .B2(n14530), .A(n13514), .ZN(P1_U2861) );
  INV_X1 U16940 ( .A(DATAI_11_), .ZN(n20693) );
  NAND2_X1 U16941 ( .A1(n19966), .A2(n20693), .ZN(n13516) );
  NAND2_X1 U16942 ( .A1(n19965), .A2(n12299), .ZN(n13515) );
  AND2_X1 U16943 ( .A1(n13516), .A2(n13515), .ZN(n19885) );
  AOI22_X1 U16944 ( .A1(n15727), .A2(n19885), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14604), .ZN(n13517) );
  OAI21_X1 U16945 ( .B1(n13518), .B2(n9576), .A(n13517), .ZN(P1_U2893) );
  NAND3_X1 U16946 ( .A1(n16864), .A2(n15523), .A3(n15525), .ZN(n17951) );
  NOR2_X1 U16947 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17951), .ZN(n13519) );
  NAND3_X1 U16948 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18542)
         );
  INV_X1 U16949 ( .A(n18247), .ZN(n18000) );
  OAI21_X1 U16950 ( .B1(n13519), .B2(n18542), .A(n18000), .ZN(n17957) );
  INV_X1 U16951 ( .A(n17957), .ZN(n13520) );
  NOR2_X1 U16952 ( .A1(n17584), .A2(n18605), .ZN(n15512) );
  AOI21_X1 U16953 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15512), .ZN(n15513) );
  NOR2_X1 U16954 ( .A1(n13520), .A2(n15513), .ZN(n13522) );
  NOR2_X1 U16955 ( .A1(n18543), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n17999) );
  OR2_X1 U16956 ( .A1(n17999), .A2(n13520), .ZN(n15511) );
  OR2_X1 U16957 ( .A1(n18298), .A2(n15511), .ZN(n13521) );
  MUX2_X1 U16958 ( .A(n13522), .B(n13521), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NAND2_X1 U16959 ( .A1(n13523), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13989) );
  OAI21_X1 U16960 ( .B1(n13523), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n13989), .ZN(n15932) );
  AOI21_X1 U16961 ( .B1(n18979), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n13524), .ZN(n13527) );
  NAND2_X1 U16962 ( .A1(n13525), .A2(n18988), .ZN(n13526) );
  OAI211_X1 U16963 ( .C1(n15932), .C2(n18992), .A(n13527), .B(n13526), .ZN(
        n13528) );
  AOI21_X1 U16964 ( .B1(n13529), .B2(n16114), .A(n13528), .ZN(n13530) );
  OAI21_X1 U16965 ( .B1(n13531), .B2(n18982), .A(n13530), .ZN(P2_U2986) );
  NAND2_X1 U16966 ( .A1(n13532), .A2(n13543), .ZN(n13547) );
  NAND2_X1 U16967 ( .A1(n13547), .A2(n18999), .ZN(n13546) );
  OR2_X1 U16968 ( .A1(n13533), .A2(n13534), .ZN(n13535) );
  NAND2_X1 U16969 ( .A1(n13536), .A2(n13535), .ZN(n15979) );
  XNOR2_X1 U16970 ( .A(n14957), .B(n13537), .ZN(n15973) );
  INV_X1 U16971 ( .A(n15973), .ZN(n14952) );
  NAND2_X1 U16972 ( .A1(n18980), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n13550) );
  OAI21_X1 U16973 ( .B1(n13538), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n13550), .ZN(n13539) );
  AOI21_X1 U16974 ( .B1(n16150), .B2(n14952), .A(n13539), .ZN(n13540) );
  OAI21_X1 U16975 ( .B1(n15979), .B2(n16158), .A(n13540), .ZN(n13541) );
  AOI21_X1 U16976 ( .B1(n13542), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n13541), .ZN(n13545) );
  NAND2_X1 U16977 ( .A1(n15028), .A2(n13543), .ZN(n13552) );
  NAND3_X1 U16978 ( .A1(n13553), .A2(n16154), .A3(n13552), .ZN(n13544) );
  OAI211_X1 U16979 ( .C1(n13557), .C2(n13546), .A(n13545), .B(n13544), .ZN(
        P2_U3019) );
  NAND2_X1 U16980 ( .A1(n13547), .A2(n16102), .ZN(n13556) );
  AOI21_X1 U16981 ( .B1(n15031), .B2(n13548), .A(n13523), .ZN(n15975) );
  NAND2_X1 U16982 ( .A1(n18979), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13549) );
  OAI211_X1 U16983 ( .C1(n15979), .C2(n16117), .A(n13550), .B(n13549), .ZN(
        n13551) );
  AOI21_X1 U16984 ( .B1(n15975), .B2(n16107), .A(n13551), .ZN(n13555) );
  NAND3_X1 U16985 ( .A1(n13553), .A2(n16114), .A3(n13552), .ZN(n13554) );
  OAI211_X1 U16986 ( .C1(n13557), .C2(n13556), .A(n13555), .B(n13554), .ZN(
        P2_U2987) );
  NOR2_X1 U16987 ( .A1(n13559), .A2(n13558), .ZN(n13560) );
  XNOR2_X1 U16988 ( .A(n13858), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13919) );
  INV_X1 U16989 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13898) );
  NAND2_X1 U16990 ( .A1(n19913), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14725) );
  OAI21_X1 U16991 ( .B1(n14677), .B2(n13898), .A(n14725), .ZN(n13906) );
  XNOR2_X1 U16992 ( .A(n13562), .B(n14437), .ZN(n14703) );
  AOI22_X1 U16993 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13566) );
  AOI22_X1 U16994 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9594), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13565) );
  AOI22_X1 U16995 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13564) );
  AOI22_X1 U16996 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13563) );
  NAND4_X1 U16997 ( .A1(n13566), .A2(n13565), .A3(n13564), .A4(n13563), .ZN(
        n13572) );
  AOI22_X1 U16998 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13570) );
  AOI22_X1 U16999 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13569) );
  AOI22_X1 U17000 ( .A1(n13887), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13568) );
  AOI22_X1 U17001 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13567) );
  NAND4_X1 U17002 ( .A1(n13570), .A2(n13569), .A3(n13568), .A4(n13567), .ZN(
        n13571) );
  NOR2_X1 U17003 ( .A1(n13572), .A2(n13571), .ZN(n13575) );
  NAND2_X1 U17004 ( .A1(n13953), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13574) );
  NAND2_X1 U17005 ( .A1(n13900), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13573) );
  OAI211_X1 U17006 ( .C1(n13607), .C2(n13575), .A(n13574), .B(n13573), .ZN(
        n13576) );
  AOI21_X1 U17007 ( .B1(n14703), .B2(n13797), .A(n13576), .ZN(n14431) );
  AOI22_X1 U17008 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13821), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13580) );
  AOI22_X1 U17009 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U17010 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13578) );
  AOI22_X1 U17011 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n9594), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13577) );
  NAND4_X1 U17012 ( .A1(n13580), .A2(n13579), .A3(n13578), .A4(n13577), .ZN(
        n13586) );
  AOI22_X1 U17013 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13878), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13584) );
  AOI22_X1 U17014 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13861), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13583) );
  AOI22_X1 U17015 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13582) );
  AOI22_X1 U17016 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11582), .B1(
        n13881), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13581) );
  NAND4_X1 U17017 ( .A1(n13584), .A2(n13583), .A3(n13582), .A4(n13581), .ZN(
        n13585) );
  OAI21_X1 U17018 ( .B1(n13586), .B2(n13585), .A(n13706), .ZN(n13591) );
  XNOR2_X1 U17019 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n13587), .ZN(
        n15765) );
  OAI22_X1 U17020 ( .A1(n15765), .A2(n13952), .B1(n13670), .B2(n15699), .ZN(
        n13588) );
  INV_X1 U17021 ( .A(n13588), .ZN(n13590) );
  NAND2_X1 U17022 ( .A1(n13900), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n13589) );
  NOR2_X1 U17023 ( .A1(n14431), .A2(n14523), .ZN(n13592) );
  XOR2_X1 U17024 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n13593), .Z(
        n15759) );
  INV_X1 U17025 ( .A(n15759), .ZN(n13609) );
  AOI22_X1 U17026 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13597) );
  AOI22_X1 U17027 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U17028 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13595) );
  AOI22_X1 U17029 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13594) );
  NAND4_X1 U17030 ( .A1(n13597), .A2(n13596), .A3(n13595), .A4(n13594), .ZN(
        n13603) );
  AOI22_X1 U17031 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13601) );
  AOI22_X1 U17032 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U17033 ( .A1(n13731), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13599) );
  AOI22_X1 U17034 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13598) );
  NAND4_X1 U17035 ( .A1(n13601), .A2(n13600), .A3(n13599), .A4(n13598), .ZN(
        n13602) );
  NOR2_X1 U17036 ( .A1(n13603), .A2(n13602), .ZN(n13606) );
  NAND2_X1 U17037 ( .A1(n13900), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13605) );
  NAND2_X1 U17038 ( .A1(n13953), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13604) );
  OAI211_X1 U17039 ( .C1(n13607), .C2(n13606), .A(n13605), .B(n13604), .ZN(
        n13608) );
  AOI21_X1 U17040 ( .B1(n13609), .B2(n13797), .A(n13608), .ZN(n14599) );
  OR2_X1 U17041 ( .A1(n13610), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13611) );
  NAND2_X1 U17042 ( .A1(n13611), .A2(n13742), .ZN(n15753) );
  INV_X1 U17043 ( .A(n14061), .ZN(n14840) );
  AOI22_X1 U17044 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13615) );
  AOI22_X1 U17045 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13821), .B1(
        n13880), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13614) );
  AOI22_X1 U17046 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n9594), .B1(
        n13889), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13613) );
  AOI22_X1 U17047 ( .A1(n13887), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13612) );
  NAND4_X1 U17048 ( .A1(n13615), .A2(n13614), .A3(n13613), .A4(n13612), .ZN(
        n13621) );
  AOI22_X1 U17049 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13886), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13619) );
  AOI22_X1 U17050 ( .A1(n13861), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U17051 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13879), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13617) );
  AOI22_X1 U17052 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11582), .B1(
        n13881), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13616) );
  NAND4_X1 U17053 ( .A1(n13619), .A2(n13618), .A3(n13617), .A4(n13616), .ZN(
        n13620) );
  NOR2_X1 U17054 ( .A1(n13621), .A2(n13620), .ZN(n13624) );
  OAI21_X1 U17055 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20055), .A(
        n20573), .ZN(n13623) );
  NAND2_X1 U17056 ( .A1(n13900), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n13622) );
  OAI211_X1 U17057 ( .C1(n13949), .C2(n13624), .A(n13623), .B(n13622), .ZN(
        n13625) );
  OAI21_X1 U17058 ( .B1(n15753), .B2(n13952), .A(n13625), .ZN(n13626) );
  INV_X1 U17059 ( .A(n13626), .ZN(n14478) );
  AOI22_X1 U17060 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13630) );
  AOI22_X1 U17061 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13731), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13629) );
  AOI22_X1 U17062 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13628) );
  AOI22_X1 U17063 ( .A1(n13887), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13627) );
  NAND4_X1 U17064 ( .A1(n13630), .A2(n13629), .A3(n13628), .A4(n13627), .ZN(
        n13636) );
  AOI22_X1 U17065 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13634) );
  AOI22_X1 U17066 ( .A1(n13861), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13633) );
  AOI22_X1 U17067 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13632) );
  AOI22_X1 U17068 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13631) );
  NAND4_X1 U17069 ( .A1(n13634), .A2(n13633), .A3(n13632), .A4(n13631), .ZN(
        n13635) );
  NOR2_X1 U17070 ( .A1(n13636), .A2(n13635), .ZN(n13640) );
  NAND2_X1 U17071 ( .A1(n20573), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13637) );
  NAND2_X1 U17072 ( .A1(n13952), .A2(n13637), .ZN(n13638) );
  AOI21_X1 U17073 ( .B1(n13900), .B2(P1_EAX_REG_19__SCAN_IN), .A(n13638), .ZN(
        n13639) );
  OAI21_X1 U17074 ( .B1(n13949), .B2(n13640), .A(n13639), .ZN(n13642) );
  XNOR2_X1 U17075 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n13644), .ZN(
        n15653) );
  NAND2_X1 U17076 ( .A1(n15653), .A2(n13797), .ZN(n13641) );
  AND2_X1 U17077 ( .A1(n13642), .A2(n13641), .ZN(n14483) );
  INV_X1 U17078 ( .A(n14483), .ZN(n13674) );
  OR2_X1 U17079 ( .A1(n13643), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13645) );
  NAND2_X1 U17080 ( .A1(n13645), .A2(n13644), .ZN(n15665) );
  AOI22_X1 U17081 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13649) );
  AOI22_X1 U17082 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13648) );
  AOI22_X1 U17083 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13647) );
  AOI22_X1 U17084 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13646) );
  NAND4_X1 U17085 ( .A1(n13649), .A2(n13648), .A3(n13647), .A4(n13646), .ZN(
        n13655) );
  AOI22_X1 U17086 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13653) );
  AOI22_X1 U17087 ( .A1(n13861), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13652) );
  AOI22_X1 U17088 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13651) );
  AOI22_X1 U17089 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13650) );
  NAND4_X1 U17090 ( .A1(n13653), .A2(n13652), .A3(n13651), .A4(n13650), .ZN(
        n13654) );
  NOR2_X1 U17091 ( .A1(n13655), .A2(n13654), .ZN(n13658) );
  OAI21_X1 U17092 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20055), .A(
        n20573), .ZN(n13657) );
  NAND2_X1 U17093 ( .A1(n13900), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n13656) );
  OAI211_X1 U17094 ( .C1(n13949), .C2(n13658), .A(n13657), .B(n13656), .ZN(
        n13659) );
  OAI21_X1 U17095 ( .B1(n15665), .B2(n13952), .A(n13659), .ZN(n14492) );
  AOI22_X1 U17096 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U17097 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13662) );
  AOI22_X1 U17098 ( .A1(n13879), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U17099 ( .A1(n13838), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13660) );
  NAND4_X1 U17100 ( .A1(n13663), .A2(n13662), .A3(n13661), .A4(n13660), .ZN(
        n13669) );
  AOI22_X1 U17101 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13667) );
  AOI22_X1 U17102 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13666) );
  AOI22_X1 U17103 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13889), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13665) );
  AOI22_X1 U17104 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13664) );
  NAND4_X1 U17105 ( .A1(n13667), .A2(n13666), .A3(n13665), .A4(n13664), .ZN(
        n13668) );
  OAI21_X1 U17106 ( .B1(n13669), .B2(n13668), .A(n13896), .ZN(n13673) );
  XNOR2_X1 U17107 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n13676), .ZN(
        n14679) );
  OAI22_X1 U17108 ( .A1(n14679), .A2(n13952), .B1(n13670), .B2(n14425), .ZN(
        n13671) );
  AOI21_X1 U17109 ( .B1(n13900), .B2(P1_EAX_REG_17__SCAN_IN), .A(n13671), .ZN(
        n13672) );
  OR2_X1 U17110 ( .A1(n14492), .A2(n14414), .ZN(n14482) );
  OR2_X1 U17111 ( .A1(n13675), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13677) );
  NAND2_X1 U17112 ( .A1(n13677), .A2(n13676), .ZN(n15758) );
  AOI22_X1 U17113 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13681) );
  AOI22_X1 U17114 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13680) );
  AOI22_X1 U17115 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13889), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13679) );
  AOI22_X1 U17116 ( .A1(n13879), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13678) );
  NAND4_X1 U17117 ( .A1(n13681), .A2(n13680), .A3(n13679), .A4(n13678), .ZN(
        n13688) );
  AOI22_X1 U17118 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13686) );
  AOI22_X1 U17119 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13685) );
  AOI22_X1 U17120 ( .A1(n13887), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13684) );
  AOI22_X1 U17121 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11582), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13683) );
  NAND4_X1 U17122 ( .A1(n13686), .A2(n13685), .A3(n13684), .A4(n13683), .ZN(
        n13687) );
  NOR2_X1 U17123 ( .A1(n13688), .A2(n13687), .ZN(n13691) );
  OAI21_X1 U17124 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20055), .A(
        n20573), .ZN(n13690) );
  NAND2_X1 U17125 ( .A1(n13900), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n13689) );
  OAI211_X1 U17126 ( .C1(n13949), .C2(n13691), .A(n13690), .B(n13689), .ZN(
        n13692) );
  OAI21_X1 U17127 ( .B1(n15758), .B2(n13952), .A(n13692), .ZN(n14501) );
  NOR2_X1 U17128 ( .A1(n13693), .A2(n14501), .ZN(n14476) );
  AND2_X1 U17129 ( .A1(n14478), .A2(n14476), .ZN(n13709) );
  XNOR2_X1 U17130 ( .A(n13694), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15682) );
  AOI22_X1 U17131 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U17132 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13889), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U17133 ( .A1(n13861), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U17134 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11582), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13695) );
  NAND4_X1 U17135 ( .A1(n13698), .A2(n13697), .A3(n13696), .A4(n13695), .ZN(
        n13704) );
  AOI22_X1 U17136 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U17137 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U17138 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U17139 ( .A1(n13838), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13699) );
  NAND4_X1 U17140 ( .A1(n13702), .A2(n13701), .A3(n13700), .A4(n13699), .ZN(
        n13703) );
  OR2_X1 U17141 ( .A1(n13704), .A2(n13703), .ZN(n13705) );
  AOI22_X1 U17142 ( .A1(n13706), .A2(n13705), .B1(n13953), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13708) );
  NAND2_X1 U17143 ( .A1(n12512), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13707) );
  OAI211_X1 U17144 ( .C1(n15682), .C2(n13952), .A(n13708), .B(n13707), .ZN(
        n14510) );
  AND2_X1 U17145 ( .A1(n13709), .A2(n14510), .ZN(n13710) );
  OR2_X1 U17146 ( .A1(n13711), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13712) );
  NAND2_X1 U17147 ( .A1(n13712), .A2(n13773), .ZN(n15743) );
  AOI22_X1 U17148 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13716) );
  AOI22_X1 U17149 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13889), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U17150 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U17151 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13713) );
  NAND4_X1 U17152 ( .A1(n13716), .A2(n13715), .A3(n13714), .A4(n13713), .ZN(
        n13722) );
  AOI22_X1 U17153 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13720) );
  AOI22_X1 U17154 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13719) );
  AOI22_X1 U17155 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13718) );
  AOI22_X1 U17156 ( .A1(n13838), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13717) );
  NAND4_X1 U17157 ( .A1(n13720), .A2(n13719), .A3(n13718), .A4(n13717), .ZN(
        n13721) );
  NOR2_X1 U17158 ( .A1(n13722), .A2(n13721), .ZN(n13725) );
  OAI21_X1 U17159 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20055), .A(
        n20573), .ZN(n13724) );
  NAND2_X1 U17160 ( .A1(n12512), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n13723) );
  OAI211_X1 U17161 ( .C1(n13949), .C2(n13725), .A(n13724), .B(n13723), .ZN(
        n13726) );
  OAI21_X1 U17162 ( .B1(n15743), .B2(n13952), .A(n13726), .ZN(n15631) );
  INV_X1 U17163 ( .A(n15631), .ZN(n13746) );
  AOI22_X1 U17164 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13730) );
  AOI22_X1 U17165 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13729) );
  AOI22_X1 U17166 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13728) );
  AOI22_X1 U17167 ( .A1(n13887), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13727) );
  NAND4_X1 U17168 ( .A1(n13730), .A2(n13729), .A3(n13728), .A4(n13727), .ZN(
        n13737) );
  AOI22_X1 U17169 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13735) );
  AOI22_X1 U17170 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13731), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13734) );
  AOI22_X1 U17171 ( .A1(n13861), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13733) );
  AOI22_X1 U17172 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11582), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13732) );
  NAND4_X1 U17173 ( .A1(n13735), .A2(n13734), .A3(n13733), .A4(n13732), .ZN(
        n13736) );
  NOR2_X1 U17174 ( .A1(n13737), .A2(n13736), .ZN(n13741) );
  NAND2_X1 U17175 ( .A1(n20573), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13738) );
  NAND2_X1 U17176 ( .A1(n13952), .A2(n13738), .ZN(n13739) );
  AOI21_X1 U17177 ( .B1(n13900), .B2(P1_EAX_REG_21__SCAN_IN), .A(n13739), .ZN(
        n13740) );
  OAI21_X1 U17178 ( .B1(n13949), .B2(n13741), .A(n13740), .ZN(n13744) );
  XNOR2_X1 U17179 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n13742), .ZN(
        n15744) );
  NAND2_X1 U17180 ( .A1(n13797), .A2(n15744), .ZN(n13743) );
  NAND2_X1 U17181 ( .A1(n13744), .A2(n13743), .ZN(n15632) );
  AOI22_X1 U17182 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13751) );
  AOI22_X1 U17183 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13750) );
  AOI22_X1 U17184 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13749) );
  AOI22_X1 U17185 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11582), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13748) );
  NAND4_X1 U17186 ( .A1(n13751), .A2(n13750), .A3(n13749), .A4(n13748), .ZN(
        n13757) );
  AOI22_X1 U17187 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13755) );
  AOI22_X1 U17188 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13754) );
  AOI22_X1 U17189 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13753) );
  AOI22_X1 U17190 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13752) );
  NAND4_X1 U17191 ( .A1(n13755), .A2(n13754), .A3(n13753), .A4(n13752), .ZN(
        n13756) );
  NOR2_X1 U17192 ( .A1(n13757), .A2(n13756), .ZN(n13779) );
  AOI22_X1 U17193 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U17194 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13760) );
  AOI22_X1 U17195 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13759) );
  AOI22_X1 U17196 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13758) );
  NAND4_X1 U17197 ( .A1(n13761), .A2(n13760), .A3(n13759), .A4(n13758), .ZN(
        n13767) );
  AOI22_X1 U17198 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13765) );
  AOI22_X1 U17199 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13764) );
  AOI22_X1 U17200 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U17201 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13762) );
  NAND4_X1 U17202 ( .A1(n13765), .A2(n13764), .A3(n13763), .A4(n13762), .ZN(
        n13766) );
  NOR2_X1 U17203 ( .A1(n13767), .A2(n13766), .ZN(n13780) );
  XOR2_X1 U17204 ( .A(n13779), .B(n13780), .Z(n13768) );
  NAND2_X1 U17205 ( .A1(n13768), .A2(n13896), .ZN(n13772) );
  NAND2_X1 U17206 ( .A1(n20573), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13769) );
  NAND2_X1 U17207 ( .A1(n13952), .A2(n13769), .ZN(n13770) );
  AOI21_X1 U17208 ( .B1(n13900), .B2(P1_EAX_REG_23__SCAN_IN), .A(n13770), .ZN(
        n13771) );
  NAND2_X1 U17209 ( .A1(n13772), .A2(n13771), .ZN(n13775) );
  XNOR2_X1 U17210 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n13773), .ZN(
        n14653) );
  NAND2_X1 U17211 ( .A1(n14653), .A2(n13797), .ZN(n13774) );
  NAND2_X1 U17212 ( .A1(n13775), .A2(n13774), .ZN(n14392) );
  OR2_X1 U17213 ( .A1(n13777), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13778) );
  NAND2_X1 U17214 ( .A1(n13778), .A2(n13815), .ZN(n15736) );
  INV_X1 U17215 ( .A(n15736), .ZN(n13798) );
  NOR2_X1 U17216 ( .A1(n13780), .A2(n13779), .ZN(n13801) );
  AOI22_X1 U17217 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13784) );
  AOI22_X1 U17218 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13783) );
  AOI22_X1 U17219 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13782) );
  AOI22_X1 U17220 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13781) );
  NAND4_X1 U17221 ( .A1(n13784), .A2(n13783), .A3(n13782), .A4(n13781), .ZN(
        n13790) );
  AOI22_X1 U17222 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U17223 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13787) );
  AOI22_X1 U17224 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13786) );
  AOI22_X1 U17225 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13785) );
  NAND4_X1 U17226 ( .A1(n13788), .A2(n13787), .A3(n13786), .A4(n13785), .ZN(
        n13789) );
  OR2_X1 U17227 ( .A1(n13790), .A2(n13789), .ZN(n13800) );
  INV_X1 U17228 ( .A(n13800), .ZN(n13791) );
  XNOR2_X1 U17229 ( .A(n13801), .B(n13791), .ZN(n13795) );
  INV_X1 U17230 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14563) );
  NAND2_X1 U17231 ( .A1(n20573), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13792) );
  OAI211_X1 U17232 ( .C1(n13793), .C2(n14563), .A(n13952), .B(n13792), .ZN(
        n13794) );
  AOI21_X1 U17233 ( .B1(n13795), .B2(n13896), .A(n13794), .ZN(n13796) );
  AOI21_X1 U17234 ( .B1(n13798), .B2(n13797), .A(n13796), .ZN(n14462) );
  NAND2_X1 U17235 ( .A1(n13801), .A2(n13800), .ZN(n13819) );
  AOI22_X1 U17236 ( .A1(n13937), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13805) );
  AOI22_X1 U17237 ( .A1(n13861), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13804) );
  AOI22_X1 U17238 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13803) );
  AOI22_X1 U17239 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13802) );
  NAND4_X1 U17240 ( .A1(n13805), .A2(n13804), .A3(n13803), .A4(n13802), .ZN(
        n13812) );
  AOI22_X1 U17241 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U17242 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13806), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13809) );
  AOI22_X1 U17243 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U17244 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13807) );
  NAND4_X1 U17245 ( .A1(n13810), .A2(n13809), .A3(n13808), .A4(n13807), .ZN(
        n13811) );
  NOR2_X1 U17246 ( .A1(n13812), .A2(n13811), .ZN(n13820) );
  XOR2_X1 U17247 ( .A(n13819), .B(n13820), .Z(n13813) );
  NAND2_X1 U17248 ( .A1(n13813), .A2(n13896), .ZN(n13817) );
  INV_X1 U17249 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14646) );
  AOI21_X1 U17250 ( .B1(n14646), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13814) );
  AOI21_X1 U17251 ( .B1(n13900), .B2(P1_EAX_REG_25__SCAN_IN), .A(n13814), .ZN(
        n13816) );
  XNOR2_X1 U17252 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n13815), .ZN(
        n14650) );
  AOI22_X1 U17253 ( .A1(n13817), .A2(n13816), .B1(n13946), .B2(n14650), .ZN(
        n14378) );
  OAI21_X1 U17254 ( .B1(n13818), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n13852), .ZN(n14637) );
  NOR2_X1 U17255 ( .A1(n13820), .A2(n13819), .ZN(n13837) );
  AOI22_X1 U17256 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13825) );
  AOI22_X1 U17257 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13824) );
  AOI22_X1 U17258 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13823) );
  AOI22_X1 U17259 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13822) );
  NAND4_X1 U17260 ( .A1(n13825), .A2(n13824), .A3(n13823), .A4(n13822), .ZN(
        n13831) );
  AOI22_X1 U17261 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13829) );
  AOI22_X1 U17262 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13828) );
  AOI22_X1 U17263 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13827) );
  AOI22_X1 U17264 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13826) );
  NAND4_X1 U17265 ( .A1(n13829), .A2(n13828), .A3(n13827), .A4(n13826), .ZN(
        n13830) );
  OR2_X1 U17266 ( .A1(n13831), .A2(n13830), .ZN(n13836) );
  XNOR2_X1 U17267 ( .A(n13837), .B(n13836), .ZN(n13834) );
  AOI21_X1 U17268 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20573), .A(
        n13946), .ZN(n13833) );
  NAND2_X1 U17269 ( .A1(n12512), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n13832) );
  OAI211_X1 U17270 ( .C1(n13834), .C2(n13949), .A(n13833), .B(n13832), .ZN(
        n13835) );
  OAI21_X1 U17271 ( .B1(n13952), .B2(n14637), .A(n13835), .ZN(n14364) );
  NAND2_X1 U17272 ( .A1(n13837), .A2(n13836), .ZN(n13859) );
  AOI22_X1 U17273 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13842) );
  AOI22_X1 U17274 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U17275 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13881), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13840) );
  AOI22_X1 U17276 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13839) );
  NAND4_X1 U17277 ( .A1(n13842), .A2(n13841), .A3(n13840), .A4(n13839), .ZN(
        n13849) );
  AOI22_X1 U17278 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13847) );
  AOI22_X1 U17279 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13821), .B1(
        n13843), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17280 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13806), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U17281 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n13889), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13844) );
  NAND4_X1 U17282 ( .A1(n13847), .A2(n13846), .A3(n13845), .A4(n13844), .ZN(
        n13848) );
  NOR2_X1 U17283 ( .A1(n13849), .A2(n13848), .ZN(n13860) );
  XOR2_X1 U17284 ( .A(n13859), .B(n13860), .Z(n13850) );
  NAND2_X1 U17285 ( .A1(n13850), .A2(n13896), .ZN(n13854) );
  NOR2_X1 U17286 ( .A1(n20813), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13851) );
  AOI211_X1 U17287 ( .C1(n13900), .C2(P1_EAX_REG_27__SCAN_IN), .A(n13946), .B(
        n13851), .ZN(n13853) );
  AOI21_X1 U17288 ( .B1(n20813), .B2(n13852), .A(n13855), .ZN(n14629) );
  AOI22_X1 U17289 ( .A1(n13854), .A2(n13853), .B1(n13946), .B2(n14629), .ZN(
        n14356) );
  NAND2_X1 U17290 ( .A1(n14355), .A2(n14356), .ZN(n14345) );
  INV_X1 U17291 ( .A(n13855), .ZN(n13856) );
  INV_X1 U17292 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14348) );
  NAND2_X1 U17293 ( .A1(n13856), .A2(n14348), .ZN(n13857) );
  NAND2_X1 U17294 ( .A1(n13858), .A2(n13857), .ZN(n14621) );
  NOR2_X1 U17295 ( .A1(n13860), .A2(n13859), .ZN(n13877) );
  AOI22_X1 U17296 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13865) );
  AOI22_X1 U17297 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13864) );
  AOI22_X1 U17298 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13863) );
  AOI22_X1 U17299 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13862) );
  NAND4_X1 U17300 ( .A1(n13865), .A2(n13864), .A3(n13863), .A4(n13862), .ZN(
        n13871) );
  AOI22_X1 U17301 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13869) );
  AOI22_X1 U17302 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13868) );
  AOI22_X1 U17303 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13867) );
  AOI22_X1 U17304 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13866) );
  NAND4_X1 U17305 ( .A1(n13869), .A2(n13868), .A3(n13867), .A4(n13866), .ZN(
        n13870) );
  OR2_X1 U17306 ( .A1(n13871), .A2(n13870), .ZN(n13876) );
  XNOR2_X1 U17307 ( .A(n13877), .B(n13876), .ZN(n13874) );
  AOI21_X1 U17308 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20573), .A(
        n13946), .ZN(n13873) );
  NAND2_X1 U17309 ( .A1(n13900), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n13872) );
  OAI211_X1 U17310 ( .C1(n13874), .C2(n13949), .A(n13873), .B(n13872), .ZN(
        n13875) );
  OAI21_X1 U17311 ( .B1(n13952), .B2(n14621), .A(n13875), .ZN(n14347) );
  NAND2_X1 U17312 ( .A1(n13877), .A2(n13876), .ZN(n13930) );
  AOI22_X1 U17313 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U17314 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13879), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U17315 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11716), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13883) );
  AOI22_X1 U17316 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13882) );
  NAND4_X1 U17317 ( .A1(n13885), .A2(n13884), .A3(n13883), .A4(n13882), .ZN(
        n13895) );
  AOI22_X1 U17318 ( .A1(n13886), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U17319 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11612), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13892) );
  AOI22_X1 U17320 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13887), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13891) );
  AOI22_X1 U17321 ( .A1(n13889), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13890) );
  NAND4_X1 U17322 ( .A1(n13893), .A2(n13892), .A3(n13891), .A4(n13890), .ZN(
        n13894) );
  NOR2_X1 U17323 ( .A1(n13895), .A2(n13894), .ZN(n13931) );
  XOR2_X1 U17324 ( .A(n13930), .B(n13931), .Z(n13897) );
  NAND2_X1 U17325 ( .A1(n13897), .A2(n13896), .ZN(n13902) );
  AOI21_X1 U17326 ( .B1(n13898), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13899) );
  AOI21_X1 U17327 ( .B1(n13900), .B2(P1_EAX_REG_29__SCAN_IN), .A(n13899), .ZN(
        n13901) );
  AOI22_X1 U17328 ( .A1(n13902), .A2(n13901), .B1(n13946), .B2(n13919), .ZN(
        n13903) );
  NOR2_X1 U17329 ( .A1(n13908), .A2(n19967), .ZN(n13905) );
  OAI21_X1 U17330 ( .B1(n14730), .B2(n19708), .A(n13907), .ZN(P1_U2970) );
  NAND2_X1 U17331 ( .A1(n13909), .A2(n19965), .ZN(n15726) );
  INV_X1 U17332 ( .A(DATAI_29_), .ZN(n13912) );
  INV_X1 U17333 ( .A(n15721), .ZN(n14586) );
  INV_X1 U17334 ( .A(DATAI_13_), .ZN(n20754) );
  NAND2_X1 U17335 ( .A1(n19965), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13910) );
  OAI21_X1 U17336 ( .B1(n19965), .B2(n20754), .A(n13910), .ZN(n19890) );
  AOI22_X1 U17337 ( .A1(n14586), .A2(n19890), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n14604), .ZN(n13911) );
  OAI21_X1 U17338 ( .B1(n14589), .B2(n13912), .A(n13911), .ZN(n13913) );
  AOI21_X1 U17339 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14593), .A(n13913), .ZN(
        n13914) );
  OAI21_X1 U17340 ( .B1(n13908), .B2(n9576), .A(n13914), .ZN(P1_U2875) );
  INV_X1 U17341 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20625) );
  INV_X1 U17342 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20627) );
  INV_X1 U17343 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20623) );
  INV_X1 U17344 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20603) );
  NAND2_X1 U17345 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19749), .ZN(n19736) );
  NOR2_X1 U17346 ( .A1(n20603), .A2(n19736), .ZN(n19724) );
  NAND3_X1 U17347 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n19724), .ZN(n15697) );
  NAND2_X1 U17348 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14402) );
  NOR2_X1 U17349 ( .A1(n15697), .A2(n14402), .ZN(n14434) );
  INV_X1 U17350 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20621) );
  NAND2_X1 U17351 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14420) );
  NAND3_X1 U17352 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14417) );
  NAND2_X1 U17353 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15652) );
  NOR4_X1 U17354 ( .A1(n20621), .A2(n14420), .A3(n14417), .A4(n15652), .ZN(
        n14403) );
  NAND2_X1 U17355 ( .A1(n14434), .A2(n14403), .ZN(n14404) );
  NOR2_X1 U17356 ( .A1(n20623), .A2(n14404), .ZN(n15638) );
  NAND2_X1 U17357 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15638), .ZN(n14397) );
  OR2_X1 U17358 ( .A1(n20627), .A2(n14397), .ZN(n15621) );
  NOR2_X1 U17359 ( .A1(n20625), .A2(n15621), .ZN(n14385) );
  NAND3_X1 U17360 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .A3(n14385), .ZN(n13917) );
  NAND2_X1 U17361 ( .A1(n15639), .A2(n13917), .ZN(n14374) );
  NAND2_X1 U17362 ( .A1(n14374), .A2(n13915), .ZN(n14370) );
  AND2_X1 U17363 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n13918) );
  NOR2_X1 U17364 ( .A1(n19747), .A2(n13918), .ZN(n13916) );
  NOR2_X1 U17365 ( .A1(n14370), .A2(n13916), .ZN(n14350) );
  INV_X1 U17366 ( .A(n14350), .ZN(n13926) );
  NOR2_X1 U17367 ( .A1(n19747), .A2(n13917), .ZN(n14359) );
  NAND2_X1 U17368 ( .A1(n14359), .A2(n13918), .ZN(n14334) );
  AOI22_X1 U17369 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19779), .B1(
        n19778), .B2(n13919), .ZN(n13921) );
  NAND2_X1 U17370 ( .A1(n19774), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n13920) );
  OAI211_X1 U17371 ( .C1(n14334), .C2(P1_REIP_REG_29__SCAN_IN), .A(n13921), 
        .B(n13920), .ZN(n13925) );
  OAI21_X1 U17372 ( .B1(n14344), .B2(n13923), .A(n13922), .ZN(n14726) );
  NOR2_X1 U17373 ( .A1(n14726), .A2(n19761), .ZN(n13924) );
  AOI211_X1 U17374 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n13926), .A(n13925), 
        .B(n13924), .ZN(n13927) );
  OAI21_X1 U17375 ( .B1(n13908), .B2(n15657), .A(n13927), .ZN(P1_U2811) );
  OAI222_X1 U17376 ( .A1(n14530), .A2(n13908), .B1(n13928), .B2(n19797), .C1(
        n14726), .C2(n14528), .ZN(P1_U2843) );
  XNOR2_X1 U17377 ( .A(n13929), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14609) );
  NOR2_X1 U17378 ( .A1(n13931), .A2(n13930), .ZN(n13945) );
  AOI22_X1 U17379 ( .A1(n13878), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13886), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U17380 ( .A1(n13843), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13861), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13935) );
  AOI22_X1 U17381 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13889), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13934) );
  AOI22_X1 U17382 ( .A1(n13881), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13932), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13933) );
  NAND4_X1 U17383 ( .A1(n13936), .A2(n13935), .A3(n13934), .A4(n13933), .ZN(
        n13943) );
  AOI22_X1 U17384 ( .A1(n13821), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13937), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13941) );
  AOI22_X1 U17385 ( .A1(n13880), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11581), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13940) );
  AOI22_X1 U17386 ( .A1(n13887), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13838), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17387 ( .A1(n9594), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13888), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13938) );
  NAND4_X1 U17388 ( .A1(n13941), .A2(n13940), .A3(n13939), .A4(n13938), .ZN(
        n13942) );
  NOR2_X1 U17389 ( .A1(n13943), .A2(n13942), .ZN(n13944) );
  XOR2_X1 U17390 ( .A(n13945), .B(n13944), .Z(n13950) );
  AOI21_X1 U17391 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20573), .A(
        n13946), .ZN(n13948) );
  NAND2_X1 U17392 ( .A1(n12512), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13947) );
  OAI211_X1 U17393 ( .C1(n13950), .C2(n13949), .A(n13948), .B(n13947), .ZN(
        n13951) );
  OAI21_X1 U17394 ( .B1(n13952), .B2(n14609), .A(n13951), .ZN(n14328) );
  AOI22_X1 U17395 ( .A1(n12512), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13953), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13954) );
  AOI21_X1 U17396 ( .B1(n19914), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13955), .ZN(n13956) );
  OAI21_X1 U17397 ( .B1(n19912), .B2(n13957), .A(n13956), .ZN(n13958) );
  AOI21_X1 U17398 ( .B1(n14533), .B2(n15781), .A(n13958), .ZN(n13959) );
  OAI21_X1 U17399 ( .B1(n13960), .B2(n19708), .A(n13959), .ZN(P1_U2968) );
  XOR2_X1 U17400 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13961), .Z(n13966)
         );
  NAND2_X1 U17401 ( .A1(n12845), .A2(n13962), .ZN(n13963) );
  NAND2_X1 U17402 ( .A1(n13964), .A2(n13963), .ZN(n18821) );
  MUX2_X1 U17403 ( .A(n18821), .B(n11050), .S(n12420), .Z(n13965) );
  OAI21_X1 U17404 ( .B1(n13966), .B2(n14929), .A(n13965), .ZN(P2_U2882) );
  NOR2_X1 U17405 ( .A1(n14918), .A2(n18825), .ZN(n13967) );
  AOI21_X1 U17406 ( .B1(n18987), .B2(n14918), .A(n13967), .ZN(n13968) );
  OAI21_X1 U17407 ( .B1(n18828), .B2(n14929), .A(n13968), .ZN(P2_U2883) );
  OAI21_X1 U17408 ( .B1(n13971), .B2(n13970), .A(n13969), .ZN(n13972) );
  INV_X1 U17409 ( .A(n13972), .ZN(n18998) );
  AOI22_X1 U17410 ( .A1(n18979), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n18980), .B2(P2_REIP_REG_2__SCAN_IN), .ZN(n13973) );
  OAI21_X1 U17411 ( .B1(n18992), .B2(n13974), .A(n13973), .ZN(n13979) );
  OAI21_X1 U17412 ( .B1(n13977), .B2(n13976), .A(n13975), .ZN(n18993) );
  NOR2_X1 U17413 ( .A1(n18993), .A2(n18984), .ZN(n13978) );
  AOI211_X1 U17414 ( .C1(n18998), .C2(n16102), .A(n13979), .B(n13978), .ZN(
        n13980) );
  OAI21_X1 U17415 ( .B1(n10318), .B2(n16117), .A(n13980), .ZN(P2_U3012) );
  NAND2_X1 U17416 ( .A1(n13985), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14008) );
  XOR2_X1 U17417 ( .A(n14008), .B(n14009), .Z(n15949) );
  INV_X1 U17418 ( .A(n15949), .ZN(n13986) );
  INV_X1 U17419 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15147) );
  NAND3_X1 U17420 ( .A1(n15949), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10858), .ZN(n15014) );
  NAND2_X1 U17421 ( .A1(n14006), .A2(n15014), .ZN(n13987) );
  INV_X1 U17422 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13999) );
  AOI21_X1 U17423 ( .B1(n13999), .B2(n13989), .A(n13988), .ZN(n15954) );
  INV_X1 U17424 ( .A(n15954), .ZN(n14003) );
  INV_X1 U17425 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n13992) );
  NAND2_X1 U17426 ( .A1(n14022), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n13991) );
  NAND2_X1 U17427 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13990) );
  OAI211_X1 U17428 ( .C1(n13993), .C2(n13992), .A(n13991), .B(n13990), .ZN(
        n13994) );
  AOI21_X1 U17429 ( .B1(n13995), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13994), .ZN(n13996) );
  NAND2_X1 U17430 ( .A1(n18980), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15151) );
  INV_X1 U17431 ( .A(n14000), .ZN(n14001) );
  INV_X1 U17432 ( .A(n14004), .ZN(n14005) );
  OAI21_X1 U17433 ( .B1(n9565), .B2(n18982), .A(n14005), .ZN(P2_U2985) );
  NAND2_X1 U17434 ( .A1(n14009), .A2(n14008), .ZN(n14013) );
  INV_X1 U17435 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n14010) );
  NOR2_X1 U17436 ( .A1(n10468), .A2(n14010), .ZN(n14011) );
  XNOR2_X1 U17437 ( .A(n14013), .B(n14011), .ZN(n15943) );
  INV_X1 U17438 ( .A(n15943), .ZN(n14012) );
  INV_X1 U17439 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14044) );
  NOR2_X1 U17440 ( .A1(n14013), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14014) );
  MUX2_X1 U17441 ( .A(n14015), .B(n14014), .S(n13985), .Z(n15928) );
  NAND2_X1 U17442 ( .A1(n15928), .A2(n10858), .ZN(n14016) );
  XNOR2_X1 U17443 ( .A(n14016), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14017) );
  XNOR2_X1 U17444 ( .A(n14018), .B(n14017), .ZN(n14058) );
  NAND2_X1 U17445 ( .A1(n15021), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14019) );
  XNOR2_X1 U17446 ( .A(n14019), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14056) );
  AOI22_X1 U17447 ( .A1(n10247), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n14021) );
  NAND2_X1 U17448 ( .A1(n14022), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14020) );
  OAI211_X1 U17449 ( .C1(n14026), .C2(n14044), .A(n14021), .B(n14020), .ZN(
        n14314) );
  NAND2_X1 U17450 ( .A1(n14313), .A2(n14314), .ZN(n14028) );
  AOI22_X1 U17451 ( .A1(n10247), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14024) );
  NAND2_X1 U17452 ( .A1(n14022), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14023) );
  OAI211_X1 U17453 ( .C1(n14026), .C2(n14025), .A(n14024), .B(n14023), .ZN(
        n14027) );
  XNOR2_X1 U17454 ( .A(n14028), .B(n14027), .ZN(n15931) );
  INV_X1 U17455 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14029) );
  NOR2_X1 U17456 ( .A1(n19016), .A2(n14029), .ZN(n14047) );
  AOI21_X1 U17457 ( .B1(n18979), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14047), .ZN(n14030) );
  OAI21_X1 U17458 ( .B1(n14031), .B2(n18992), .A(n14030), .ZN(n14032) );
  INV_X1 U17459 ( .A(n14032), .ZN(n14033) );
  AOI21_X1 U17460 ( .B1(n14056), .B2(n16114), .A(n14035), .ZN(n14036) );
  INV_X1 U17461 ( .A(n15931), .ZN(n14054) );
  INV_X1 U17462 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n14037) );
  OR2_X1 U17463 ( .A1(n10827), .A2(n14037), .ZN(n14039) );
  AOI22_X1 U17464 ( .A1(n10987), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14038) );
  NAND2_X1 U17465 ( .A1(n14039), .A2(n14038), .ZN(n14933) );
  AOI222_X1 U17466 ( .A1(n10835), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14040), .C1(n10987), .C2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14307) );
  AOI222_X1 U17467 ( .A1(n10835), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n14040), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n10987), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n14041) );
  XNOR2_X1 U17468 ( .A(n14042), .B(n14041), .ZN(n15930) );
  INV_X1 U17469 ( .A(n14043), .ZN(n15148) );
  NAND3_X1 U17470 ( .A1(n15149), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15148), .ZN(n15135) );
  NOR3_X1 U17471 ( .A1(n15135), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14044), .ZN(n14051) );
  AOI21_X1 U17472 ( .B1(n14045), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15365), .ZN(n15134) );
  NOR2_X1 U17473 ( .A1(n15400), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14046) );
  OAI21_X1 U17474 ( .B1(n15134), .B2(n14046), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14049) );
  INV_X1 U17475 ( .A(n14047), .ZN(n14048) );
  NAND2_X1 U17476 ( .A1(n14049), .A2(n14048), .ZN(n14050) );
  OAI21_X1 U17477 ( .B1(n14054), .B2(n16158), .A(n14053), .ZN(n14055) );
  AOI21_X1 U17478 ( .B1(n14056), .B2(n16154), .A(n14055), .ZN(n14057) );
  INV_X1 U17479 ( .A(n15926), .ZN(n14059) );
  AOI22_X1 U17480 ( .A1(n15561), .A2(n19701), .B1(n14059), .B2(
        P1_FLUSH_REG_SCAN_IN), .ZN(n15914) );
  OAI21_X1 U17481 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20386), .A(n15914), 
        .ZN(n15918) );
  INV_X1 U17482 ( .A(n15918), .ZN(n14066) );
  AOI21_X1 U17483 ( .B1(n14060), .B2(n19700), .A(n14066), .ZN(n14067) );
  OAI22_X1 U17484 ( .A1(n14063), .A2(n14062), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14061), .ZN(n15556) );
  OAI22_X1 U17485 ( .A1(n20570), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14857), .ZN(n14064) );
  AOI21_X1 U17486 ( .B1(n15556), .B2(n19700), .A(n14064), .ZN(n14065) );
  OAI22_X1 U17487 ( .A1(n14067), .A2(n15559), .B1(n14066), .B2(n14065), .ZN(
        P1_U3474) );
  INV_X1 U17488 ( .A(n14068), .ZN(n14090) );
  AOI22_X1 U17489 ( .A1(n10344), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14072) );
  AOI22_X1 U17490 ( .A1(n10432), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14071) );
  AOI22_X1 U17491 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14070) );
  AOI22_X1 U17492 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14069) );
  NAND4_X1 U17493 ( .A1(n14072), .A2(n14071), .A3(n14070), .A4(n14069), .ZN(
        n14078) );
  AOI22_X1 U17494 ( .A1(n14120), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14076) );
  AOI22_X1 U17495 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14121), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14075) );
  AOI22_X1 U17496 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14122), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14074) );
  AOI22_X1 U17497 ( .A1(n13195), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14073) );
  NAND4_X1 U17498 ( .A1(n14076), .A2(n14075), .A3(n14074), .A4(n14073), .ZN(
        n14077) );
  NOR2_X1 U17499 ( .A1(n14078), .A2(n14077), .ZN(n14920) );
  AOI22_X1 U17500 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10864), .B1(
        n10344), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17501 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10432), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U17502 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14080) );
  AOI22_X1 U17503 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14079) );
  NAND4_X1 U17504 ( .A1(n14082), .A2(n14081), .A3(n14080), .A4(n14079), .ZN(
        n14088) );
  AOI22_X1 U17505 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10437), .B1(
        n14120), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U17506 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n14121), .ZN(n14085) );
  AOI22_X1 U17507 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n14122), .ZN(n14084) );
  AOI22_X1 U17508 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14083) );
  NAND4_X1 U17509 ( .A1(n14086), .A2(n14085), .A3(n14084), .A4(n14083), .ZN(
        n14087) );
  NOR2_X1 U17510 ( .A1(n14088), .A2(n14087), .ZN(n14910) );
  NOR2_X1 U17511 ( .A1(n14920), .A2(n14910), .ZN(n14089) );
  NAND2_X1 U17512 ( .A1(n14090), .A2(n14089), .ZN(n14131) );
  AOI22_X1 U17513 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14279), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14103) );
  AOI22_X1 U17514 ( .A1(n14297), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U17515 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14101) );
  INV_X1 U17516 ( .A(n9588), .ZN(n14292) );
  INV_X1 U17517 ( .A(n14093), .ZN(n14095) );
  NAND2_X1 U17518 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14094) );
  NAND2_X1 U17519 ( .A1(n14095), .A2(n14094), .ZN(n14286) );
  INV_X1 U17520 ( .A(n14282), .ZN(n14288) );
  INV_X1 U17521 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14096) );
  OR2_X1 U17522 ( .A1(n14288), .A2(n14096), .ZN(n14097) );
  OAI211_X1 U17523 ( .C1(n14292), .C2(n14098), .A(n14286), .B(n14097), .ZN(
        n14099) );
  INV_X1 U17524 ( .A(n14099), .ZN(n14100) );
  NAND4_X1 U17525 ( .A1(n14103), .A2(n14102), .A3(n14101), .A4(n14100), .ZN(
        n14113) );
  AOI22_X1 U17526 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14279), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U17527 ( .A1(n14297), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14110) );
  INV_X1 U17528 ( .A(n14104), .ZN(n14290) );
  AOI22_X1 U17529 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14109) );
  INV_X1 U17530 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19460) );
  INV_X1 U17531 ( .A(n14286), .ZN(n14264) );
  OR2_X1 U17532 ( .A1(n14288), .A2(n14105), .ZN(n14106) );
  OAI211_X1 U17533 ( .C1(n14292), .C2(n19460), .A(n14264), .B(n14106), .ZN(
        n14107) );
  INV_X1 U17534 ( .A(n14107), .ZN(n14108) );
  NAND4_X1 U17535 ( .A1(n14111), .A2(n14110), .A3(n14109), .A4(n14108), .ZN(
        n14112) );
  AND2_X1 U17536 ( .A1(n14113), .A2(n14112), .ZN(n14150) );
  NAND2_X1 U17537 ( .A1(n9573), .A2(n14150), .ZN(n14130) );
  AOI22_X1 U17538 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10432), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14119) );
  AOI22_X1 U17539 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10344), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U17540 ( .A1(n14114), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U17541 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14115), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14116) );
  NAND4_X1 U17542 ( .A1(n14119), .A2(n14118), .A3(n14117), .A4(n14116), .ZN(
        n14129) );
  AOI22_X1 U17543 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10437), .B1(
        n14120), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14127) );
  AOI22_X1 U17544 ( .A1(n10349), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n14121), .ZN(n14126) );
  AOI22_X1 U17545 ( .A1(n14123), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14122), .ZN(n14125) );
  AOI22_X1 U17546 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13195), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14124) );
  NAND4_X1 U17547 ( .A1(n14127), .A2(n14126), .A3(n14125), .A4(n14124), .ZN(
        n14128) );
  XNOR2_X1 U17548 ( .A(n14130), .B(n14151), .ZN(n14156) );
  XNOR2_X1 U17549 ( .A(n14131), .B(n14156), .ZN(n14903) );
  INV_X1 U17550 ( .A(n14150), .ZN(n14154) );
  NOR2_X1 U17551 ( .A1(n9573), .A2(n14154), .ZN(n14904) );
  INV_X1 U17552 ( .A(n14131), .ZN(n14132) );
  AOI22_X1 U17553 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14139) );
  AOI22_X1 U17554 ( .A1(n14279), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14138) );
  AOI22_X1 U17555 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14137) );
  OR2_X1 U17556 ( .A1(n14288), .A2(n14133), .ZN(n14134) );
  OAI211_X1 U17557 ( .C1(n14292), .C2(n10309), .A(n14286), .B(n14134), .ZN(
        n14135) );
  INV_X1 U17558 ( .A(n14135), .ZN(n14136) );
  NAND4_X1 U17559 ( .A1(n14139), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        n14149) );
  AOI22_X1 U17560 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U17561 ( .A1(n14279), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U17562 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14145) );
  INV_X1 U17563 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14142) );
  OR2_X1 U17564 ( .A1(n14288), .A2(n14140), .ZN(n14141) );
  OAI211_X1 U17565 ( .C1(n14292), .C2(n14142), .A(n14264), .B(n14141), .ZN(
        n14143) );
  INV_X1 U17566 ( .A(n14143), .ZN(n14144) );
  NAND4_X1 U17567 ( .A1(n14147), .A2(n14146), .A3(n14145), .A4(n14144), .ZN(
        n14148) );
  NAND2_X1 U17568 ( .A1(n14149), .A2(n14148), .ZN(n14157) );
  NAND2_X1 U17569 ( .A1(n14151), .A2(n14150), .ZN(n14158) );
  XOR2_X1 U17570 ( .A(n14157), .B(n14158), .Z(n14152) );
  NAND2_X1 U17571 ( .A1(n14152), .A2(n14201), .ZN(n14892) );
  INV_X1 U17572 ( .A(n14157), .ZN(n14153) );
  NAND2_X1 U17573 ( .A1(n19683), .A2(n14153), .ZN(n14894) );
  NOR2_X1 U17574 ( .A1(n14894), .A2(n14154), .ZN(n14155) );
  NOR2_X1 U17575 ( .A1(n14158), .A2(n14157), .ZN(n14176) );
  AOI22_X1 U17576 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14166) );
  AOI22_X1 U17577 ( .A1(n14279), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14165) );
  AOI22_X1 U17578 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14164) );
  INV_X1 U17579 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14161) );
  INV_X1 U17580 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14159) );
  OR2_X1 U17581 ( .A1(n14288), .A2(n14159), .ZN(n14160) );
  OAI211_X1 U17582 ( .C1(n14292), .C2(n14161), .A(n14286), .B(n14160), .ZN(
        n14162) );
  INV_X1 U17583 ( .A(n14162), .ZN(n14163) );
  NAND4_X1 U17584 ( .A1(n14166), .A2(n14165), .A3(n14164), .A4(n14163), .ZN(
        n14175) );
  AOI22_X1 U17585 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14279), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14173) );
  INV_X1 U17586 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n19265) );
  AOI22_X1 U17587 ( .A1(n14297), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14172) );
  AOI22_X1 U17588 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14171) );
  INV_X1 U17589 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14168) );
  INV_X1 U17590 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n19364) );
  OR2_X1 U17591 ( .A1(n14288), .A2(n19364), .ZN(n14167) );
  OAI211_X1 U17592 ( .C1(n14292), .C2(n14168), .A(n14264), .B(n14167), .ZN(
        n14169) );
  INV_X1 U17593 ( .A(n14169), .ZN(n14170) );
  NAND4_X1 U17594 ( .A1(n14173), .A2(n14172), .A3(n14171), .A4(n14170), .ZN(
        n14174) );
  AND2_X1 U17595 ( .A1(n14175), .A2(n14174), .ZN(n14178) );
  NAND2_X1 U17596 ( .A1(n14176), .A2(n14178), .ZN(n14226) );
  OAI211_X1 U17597 ( .C1(n14176), .C2(n14178), .A(n14201), .B(n14226), .ZN(
        n14180) );
  INV_X1 U17598 ( .A(n14180), .ZN(n14177) );
  INV_X1 U17599 ( .A(n14178), .ZN(n14179) );
  NOR2_X1 U17600 ( .A1(n9573), .A2(n14179), .ZN(n14886) );
  AOI22_X1 U17601 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U17602 ( .A1(n14279), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14189) );
  AOI22_X1 U17603 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14188) );
  OR2_X1 U17604 ( .A1(n14288), .A2(n14183), .ZN(n14184) );
  OAI211_X1 U17605 ( .C1(n14292), .C2(n14185), .A(n14286), .B(n14184), .ZN(
        n14186) );
  INV_X1 U17606 ( .A(n14186), .ZN(n14187) );
  NAND4_X1 U17607 ( .A1(n14190), .A2(n14189), .A3(n14188), .A4(n14187), .ZN(
        n14200) );
  AOI22_X1 U17608 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14198) );
  AOI22_X1 U17609 ( .A1(n14279), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14197) );
  AOI22_X1 U17610 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14196) );
  INV_X1 U17611 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14193) );
  OR2_X1 U17612 ( .A1(n14288), .A2(n14191), .ZN(n14192) );
  OAI211_X1 U17613 ( .C1(n14292), .C2(n14193), .A(n14264), .B(n14192), .ZN(
        n14194) );
  INV_X1 U17614 ( .A(n14194), .ZN(n14195) );
  NAND4_X1 U17615 ( .A1(n14198), .A2(n14197), .A3(n14196), .A4(n14195), .ZN(
        n14199) );
  AND2_X1 U17616 ( .A1(n14200), .A2(n14199), .ZN(n14203) );
  XNOR2_X1 U17617 ( .A(n14226), .B(n14203), .ZN(n14202) );
  NAND2_X1 U17618 ( .A1(n14202), .A2(n14201), .ZN(n14205) );
  INV_X1 U17619 ( .A(n14203), .ZN(n14225) );
  NOR2_X1 U17620 ( .A1(n9573), .A2(n14225), .ZN(n14878) );
  INV_X1 U17621 ( .A(n14204), .ZN(n14206) );
  NAND2_X1 U17622 ( .A1(n14877), .A2(n10080), .ZN(n14230) );
  AOI22_X1 U17623 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14213) );
  AOI22_X1 U17624 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14295), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14212) );
  AOI22_X1 U17625 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14211) );
  INV_X1 U17626 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14208) );
  NAND2_X1 U17627 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14207) );
  OAI211_X1 U17628 ( .C1(n14288), .C2(n14208), .A(n14207), .B(n14264), .ZN(
        n14209) );
  INV_X1 U17629 ( .A(n14209), .ZN(n14210) );
  NAND4_X1 U17630 ( .A1(n14213), .A2(n14212), .A3(n14211), .A4(n14210), .ZN(
        n14224) );
  AOI22_X1 U17631 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14222) );
  AOI22_X1 U17632 ( .A1(n14279), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14221) );
  AOI22_X1 U17633 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14220) );
  INV_X1 U17634 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14217) );
  INV_X1 U17635 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14215) );
  OR2_X1 U17636 ( .A1(n14288), .A2(n14215), .ZN(n14216) );
  OAI211_X1 U17637 ( .C1(n14292), .C2(n14217), .A(n14286), .B(n14216), .ZN(
        n14218) );
  INV_X1 U17638 ( .A(n14218), .ZN(n14219) );
  NAND4_X1 U17639 ( .A1(n14222), .A2(n14221), .A3(n14220), .A4(n14219), .ZN(
        n14223) );
  NAND2_X1 U17640 ( .A1(n14224), .A2(n14223), .ZN(n14232) );
  OR2_X1 U17641 ( .A1(n14226), .A2(n14225), .ZN(n14228) );
  NOR2_X1 U17642 ( .A1(n14228), .A2(n14232), .ZN(n14254) );
  AOI211_X1 U17643 ( .C1(n14232), .C2(n14228), .A(n14227), .B(n14254), .ZN(
        n14229) );
  NAND2_X1 U17644 ( .A1(n14230), .A2(n14229), .ZN(n14234) );
  INV_X1 U17645 ( .A(n14232), .ZN(n14233) );
  NAND2_X1 U17646 ( .A1(n19683), .A2(n14233), .ZN(n14872) );
  INV_X1 U17647 ( .A(n14234), .ZN(n14253) );
  AOI22_X1 U17648 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14242) );
  AOI22_X1 U17649 ( .A1(n14279), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U17650 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14240) );
  OR2_X1 U17651 ( .A1(n14288), .A2(n14235), .ZN(n14236) );
  OAI211_X1 U17652 ( .C1(n14292), .C2(n14237), .A(n14286), .B(n14236), .ZN(
        n14238) );
  INV_X1 U17653 ( .A(n14238), .ZN(n14239) );
  NAND4_X1 U17654 ( .A1(n14242), .A2(n14241), .A3(n14240), .A4(n14239), .ZN(
        n14252) );
  AOI22_X1 U17655 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14250) );
  AOI22_X1 U17656 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14249) );
  AOI22_X1 U17657 ( .A1(n14295), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14248) );
  OR2_X1 U17658 ( .A1(n14288), .A2(n14243), .ZN(n14244) );
  OAI211_X1 U17659 ( .C1(n14292), .C2(n14245), .A(n14264), .B(n14244), .ZN(
        n14246) );
  INV_X1 U17660 ( .A(n14246), .ZN(n14247) );
  NAND4_X1 U17661 ( .A1(n14250), .A2(n14249), .A3(n14248), .A4(n14247), .ZN(
        n14251) );
  AND2_X1 U17662 ( .A1(n14252), .A2(n14251), .ZN(n14867) );
  INV_X1 U17663 ( .A(n14254), .ZN(n14866) );
  NAND2_X1 U17664 ( .A1(n9573), .A2(n14867), .ZN(n14255) );
  NOR2_X1 U17665 ( .A1(n14866), .A2(n14255), .ZN(n14275) );
  AOI22_X1 U17666 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14279), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14262) );
  AOI22_X1 U17667 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14295), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14261) );
  AOI22_X1 U17668 ( .A1(n14297), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14260) );
  OR2_X1 U17669 ( .A1(n14288), .A2(n14256), .ZN(n14257) );
  OAI211_X1 U17670 ( .C1(n10528), .C2(n14290), .A(n14257), .B(n14286), .ZN(
        n14258) );
  INV_X1 U17671 ( .A(n14258), .ZN(n14259) );
  NAND4_X1 U17672 ( .A1(n14262), .A2(n14261), .A3(n14260), .A4(n14259), .ZN(
        n14273) );
  INV_X1 U17673 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n19296) );
  AOI22_X1 U17674 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14279), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14271) );
  AOI22_X1 U17675 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14295), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14270) );
  INV_X1 U17676 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n19277) );
  AOI22_X1 U17677 ( .A1(n14297), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14269) );
  NAND2_X1 U17678 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14265) );
  OAI211_X1 U17679 ( .C1(n14288), .C2(n14266), .A(n14265), .B(n14264), .ZN(
        n14267) );
  INV_X1 U17680 ( .A(n14267), .ZN(n14268) );
  NAND4_X1 U17681 ( .A1(n14271), .A2(n14270), .A3(n14269), .A4(n14268), .ZN(
        n14272) );
  AND2_X1 U17682 ( .A1(n14273), .A2(n14272), .ZN(n14274) );
  NAND2_X1 U17683 ( .A1(n14275), .A2(n14274), .ZN(n14276) );
  OAI21_X1 U17684 ( .B1(n14275), .B2(n14274), .A(n14276), .ZN(n14863) );
  INV_X1 U17685 ( .A(n14276), .ZN(n14277) );
  NOR2_X1 U17686 ( .A1(n14861), .A2(n14277), .ZN(n14305) );
  AOI22_X1 U17687 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14297), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14281) );
  AOI22_X1 U17688 ( .A1(n14279), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14278), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14280) );
  NAND2_X1 U17689 ( .A1(n14281), .A2(n14280), .ZN(n14303) );
  INV_X1 U17690 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14285) );
  AOI22_X1 U17691 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14263), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14284) );
  AOI21_X1 U17692 ( .B1(n14282), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n14286), .ZN(n14283) );
  OAI211_X1 U17693 ( .C1(n12645), .C2(n14285), .A(n14284), .B(n14283), .ZN(
        n14302) );
  INV_X1 U17694 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14287) );
  OAI21_X1 U17695 ( .B1(n14288), .B2(n14287), .A(n14286), .ZN(n14294) );
  INV_X1 U17696 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14291) );
  INV_X1 U17697 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14289) );
  OAI22_X1 U17698 ( .A1(n14292), .A2(n14291), .B1(n14290), .B2(n14289), .ZN(
        n14293) );
  AOI211_X1 U17699 ( .C1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n14295), .A(
        n14294), .B(n14293), .ZN(n14300) );
  AOI22_X1 U17700 ( .A1(n14092), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9579), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14299) );
  AOI22_X1 U17701 ( .A1(n14297), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14296), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14298) );
  NAND3_X1 U17702 ( .A1(n14300), .A2(n14299), .A3(n14298), .ZN(n14301) );
  OAI21_X1 U17703 ( .B1(n14303), .B2(n14302), .A(n14301), .ZN(n14304) );
  XNOR2_X1 U17704 ( .A(n14305), .B(n14304), .ZN(n14318) );
  MUX2_X1 U17705 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n12166), .Z(n18972) );
  INV_X1 U17706 ( .A(n18972), .ZN(n14309) );
  INV_X1 U17707 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14308) );
  OAI22_X1 U17708 ( .A1(n15005), .A2(n14309), .B1(n18892), .B2(n14308), .ZN(
        n14310) );
  AOI21_X1 U17709 ( .B1(n15945), .B2(n18921), .A(n14310), .ZN(n14312) );
  AOI22_X1 U17710 ( .A1(n18864), .A2(BUF2_REG_30__SCAN_IN), .B1(n18865), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14311) );
  OAI211_X1 U17711 ( .C1(n14318), .C2(n18868), .A(n14312), .B(n14311), .ZN(
        P2_U2889) );
  XOR2_X1 U17712 ( .A(n14314), .B(n14313), .Z(n14315) );
  NAND2_X1 U17713 ( .A1(n14315), .A2(n14918), .ZN(n14317) );
  NAND2_X1 U17714 ( .A1(n12420), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14316) );
  OAI211_X1 U17715 ( .C1(n14318), .C2(n14929), .A(n14317), .B(n14316), .ZN(
        P2_U2857) );
  NAND2_X1 U17716 ( .A1(n14533), .A2(n19755), .ZN(n14325) );
  INV_X1 U17717 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20638) );
  INV_X1 U17718 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20807) );
  NOR2_X1 U17719 ( .A1(n20638), .A2(n20807), .ZN(n14320) );
  OAI21_X1 U17720 ( .B1(n14320), .B2(n19747), .A(n14350), .ZN(n14335) );
  INV_X1 U17721 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14452) );
  OAI22_X1 U17722 ( .A1(n19728), .A2(n14319), .B1(n15629), .B2(n14452), .ZN(
        n14323) );
  INV_X1 U17723 ( .A(n14320), .ZN(n14321) );
  NOR3_X1 U17724 ( .A1(n14334), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14321), 
        .ZN(n14322) );
  AOI211_X1 U17725 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14335), .A(n14323), 
        .B(n14322), .ZN(n14324) );
  OAI211_X1 U17726 ( .C1(n14453), .C2(n19761), .A(n14325), .B(n14324), .ZN(
        P1_U2809) );
  AOI21_X1 U17727 ( .B1(n14328), .B2(n14327), .A(n14326), .ZN(n14611) );
  INV_X1 U17728 ( .A(n14611), .ZN(n14542) );
  INV_X1 U17729 ( .A(n14329), .ZN(n14330) );
  AOI22_X1 U17730 ( .A1(n13922), .A2(n14331), .B1(n14344), .B2(n14330), .ZN(
        n14333) );
  INV_X1 U17731 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14455) );
  NOR2_X1 U17732 ( .A1(n14334), .A2(n20638), .ZN(n14336) );
  OAI21_X1 U17733 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14336), .A(n14335), 
        .ZN(n14339) );
  INV_X1 U17734 ( .A(n14609), .ZN(n14337) );
  AOI22_X1 U17735 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19779), .B1(
        n19778), .B2(n14337), .ZN(n14338) );
  OAI211_X1 U17736 ( .C1(n15629), .C2(n14455), .A(n14339), .B(n14338), .ZN(
        n14340) );
  AOI21_X1 U17737 ( .B1(n14721), .B2(n19773), .A(n14340), .ZN(n14341) );
  OAI21_X1 U17738 ( .B1(n14542), .B2(n15657), .A(n14341), .ZN(P1_U2810) );
  NOR2_X1 U17739 ( .A1(n14357), .A2(n14342), .ZN(n14343) );
  OR2_X1 U17740 ( .A1(n14344), .A2(n14343), .ZN(n14737) );
  AOI21_X1 U17741 ( .B1(n14347), .B2(n14345), .A(n14346), .ZN(n14623) );
  NAND2_X1 U17742 ( .A1(n14623), .A2(n19755), .ZN(n14354) );
  OAI22_X1 U17743 ( .A1(n14348), .A2(n19728), .B1(n19751), .B2(n14621), .ZN(
        n14352) );
  AOI21_X1 U17744 ( .B1(n14359), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14349) );
  NOR2_X1 U17745 ( .A1(n14350), .A2(n14349), .ZN(n14351) );
  AOI211_X1 U17746 ( .C1(n19774), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14352), .B(
        n14351), .ZN(n14353) );
  OAI211_X1 U17747 ( .C1(n19761), .C2(n14737), .A(n14354), .B(n14353), .ZN(
        P1_U2812) );
  OAI21_X1 U17748 ( .B1(n14355), .B2(n14356), .A(n14345), .ZN(n14632) );
  AOI21_X1 U17749 ( .B1(n14358), .B2(n14365), .A(n14357), .ZN(n14749) );
  INV_X1 U17750 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20634) );
  AOI22_X1 U17751 ( .A1(n14629), .A2(n19778), .B1(n14359), .B2(n20634), .ZN(
        n14361) );
  AOI22_X1 U17752 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(n19774), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(n14370), .ZN(n14360) );
  OAI211_X1 U17753 ( .C1(n20813), .C2(n19728), .A(n14361), .B(n14360), .ZN(
        n14362) );
  AOI21_X1 U17754 ( .B1(n14749), .B2(n19773), .A(n14362), .ZN(n14363) );
  OAI21_X1 U17755 ( .B1(n14632), .B2(n15657), .A(n14363), .ZN(P1_U2813) );
  AOI21_X1 U17756 ( .B1(n14364), .B2(n14377), .A(n14355), .ZN(n14639) );
  INV_X1 U17757 ( .A(n14639), .ZN(n14558) );
  INV_X1 U17758 ( .A(n14365), .ZN(n14366) );
  AOI21_X1 U17759 ( .B1(n14367), .B2(n14383), .A(n14366), .ZN(n14760) );
  NAND2_X1 U17760 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14385), .ZN(n14373) );
  INV_X1 U17761 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14368) );
  OAI22_X1 U17762 ( .A1(n14368), .A2(n19728), .B1(n19751), .B2(n14637), .ZN(
        n14369) );
  AOI21_X1 U17763 ( .B1(n19774), .B2(P1_EBX_REG_26__SCAN_IN), .A(n14369), .ZN(
        n14372) );
  NAND2_X1 U17764 ( .A1(n14370), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14371) );
  OAI211_X1 U17765 ( .C1(n14374), .C2(n14373), .A(n14372), .B(n14371), .ZN(
        n14375) );
  AOI21_X1 U17766 ( .B1(n14760), .B2(n19773), .A(n14375), .ZN(n14376) );
  OAI21_X1 U17767 ( .B1(n14558), .B2(n15657), .A(n14376), .ZN(P1_U2814) );
  OAI21_X1 U17768 ( .B1(n9649), .B2(n14378), .A(n14377), .ZN(n14647) );
  INV_X1 U17769 ( .A(n14647), .ZN(n14379) );
  NAND2_X1 U17770 ( .A1(n14379), .A2(n19755), .ZN(n14390) );
  INV_X1 U17771 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14459) );
  OAI22_X1 U17772 ( .A1(n14646), .A2(n19728), .B1(n14459), .B2(n15629), .ZN(
        n14380) );
  AOI21_X1 U17773 ( .B1(n19778), .B2(n14650), .A(n14380), .ZN(n14389) );
  NAND2_X1 U17774 ( .A1(n14467), .A2(n14381), .ZN(n14382) );
  AND2_X1 U17775 ( .A1(n14383), .A2(n14382), .ZN(n15796) );
  AOI21_X1 U17776 ( .B1(n15639), .B2(n15621), .A(n19725), .ZN(n15620) );
  OAI21_X1 U17777 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n19747), .A(n15620), 
        .ZN(n14384) );
  AOI22_X1 U17778 ( .A1(n15796), .A2(n19773), .B1(P1_REIP_REG_25__SCAN_IN), 
        .B2(n14384), .ZN(n14388) );
  INV_X1 U17779 ( .A(n14385), .ZN(n14386) );
  OR3_X1 U17780 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n19747), .A3(n14386), .ZN(
        n14387) );
  NAND4_X1 U17781 ( .A1(n14390), .A2(n14389), .A3(n14388), .A4(n14387), .ZN(
        P1_U2815) );
  AOI21_X1 U17782 ( .B1(n14392), .B2(n15633), .A(n9624), .ZN(n14657) );
  INV_X1 U17783 ( .A(n14657), .ZN(n14572) );
  INV_X1 U17784 ( .A(n15636), .ZN(n14406) );
  AOI21_X1 U17785 ( .B1(n14406), .B2(n15635), .A(n14393), .ZN(n14394) );
  OR2_X1 U17786 ( .A1(n14394), .A2(n14465), .ZN(n14471) );
  INV_X1 U17787 ( .A(n14471), .ZN(n15804) );
  AOI22_X1 U17788 ( .A1(n14653), .A2(n19778), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n19774), .ZN(n14395) );
  OAI21_X1 U17789 ( .B1(n14396), .B2(n19728), .A(n14395), .ZN(n14399) );
  AOI221_X1 U17790 ( .B1(n19747), .B2(n20627), .C1(n14397), .C2(n20627), .A(
        n15620), .ZN(n14398) );
  AOI211_X1 U17791 ( .C1(n19773), .C2(n15804), .A(n14399), .B(n14398), .ZN(
        n14400) );
  OAI21_X1 U17792 ( .B1(n14572), .B2(n15657), .A(n14400), .ZN(P1_U2817) );
  XOR2_X1 U17793 ( .A(n15632), .B(n14401), .Z(n15745) );
  INV_X1 U17794 ( .A(n14418), .ZN(n14443) );
  NAND2_X1 U17795 ( .A1(n14418), .A2(n14419), .ZN(n15703) );
  OAI21_X1 U17796 ( .B1(n14403), .B2(n14443), .A(n15703), .ZN(n15648) );
  NOR3_X1 U17797 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n19747), .A3(n14404), 
        .ZN(n15637) );
  INV_X1 U17798 ( .A(n15744), .ZN(n14410) );
  AOI21_X1 U17799 ( .B1(n14407), .B2(n14405), .A(n14406), .ZN(n14788) );
  NAND2_X1 U17800 ( .A1(n14788), .A2(n19773), .ZN(n14409) );
  AOI22_X1 U17801 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(n19774), .ZN(n14408) );
  OAI211_X1 U17802 ( .C1(n14410), .C2(n19751), .A(n14409), .B(n14408), .ZN(
        n14411) );
  AOI211_X1 U17803 ( .C1(n15648), .C2(P1_REIP_REG_21__SCAN_IN), .A(n15637), 
        .B(n14411), .ZN(n14412) );
  OAI21_X1 U17804 ( .B1(n14577), .B2(n15657), .A(n14412), .ZN(P1_U2819) );
  NAND2_X1 U17805 ( .A1(n14413), .A2(n14510), .ZN(n14512) );
  INV_X1 U17806 ( .A(n14503), .ZN(n14416) );
  INV_X1 U17807 ( .A(n14414), .ZN(n14415) );
  NAND2_X1 U17808 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15672) );
  NAND4_X1 U17809 ( .A1(n15639), .A2(n14434), .A3(P1_REIP_REG_14__SCAN_IN), 
        .A4(P1_REIP_REG_13__SCAN_IN), .ZN(n15689) );
  NOR2_X1 U17810 ( .A1(n15672), .A2(n15689), .ZN(n15646) );
  INV_X1 U17811 ( .A(n14417), .ZN(n14421) );
  OAI21_X1 U17812 ( .B1(n14420), .B2(n14419), .A(n14418), .ZN(n15691) );
  OAI21_X1 U17813 ( .B1(n14421), .B2(n14443), .A(n15691), .ZN(n15663) );
  OAI21_X1 U17814 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15646), .A(n15663), 
        .ZN(n14428) );
  NAND2_X1 U17815 ( .A1(n14506), .A2(n14422), .ZN(n14423) );
  AND2_X1 U17816 ( .A1(n14494), .A2(n14423), .ZN(n15836) );
  AOI22_X1 U17817 ( .A1(n14679), .A2(n19778), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n19774), .ZN(n14424) );
  OAI211_X1 U17818 ( .C1(n19728), .C2(n14425), .A(n14424), .B(n19927), .ZN(
        n14426) );
  AOI21_X1 U17819 ( .B1(n15836), .B2(n19773), .A(n14426), .ZN(n14427) );
  OAI211_X1 U17820 ( .C1(n14682), .C2(n15657), .A(n14428), .B(n14427), .ZN(
        P1_U2823) );
  AOI21_X1 U17821 ( .B1(n14430), .B2(n9856), .A(n9625), .ZN(n14524) );
  NOR2_X1 U17822 ( .A1(n14524), .A2(n14523), .ZN(n14522) );
  INV_X1 U17823 ( .A(n14431), .ZN(n14433) );
  OAI21_X1 U17824 ( .B1(n14522), .B2(n14433), .A(n14432), .ZN(n14707) );
  INV_X1 U17825 ( .A(n15703), .ZN(n14440) );
  NAND2_X1 U17826 ( .A1(n15639), .A2(n14434), .ZN(n15690) );
  OAI22_X1 U17827 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15690), .B1(n14703), 
        .B2(n19751), .ZN(n14439) );
  AOI21_X1 U17828 ( .B1(n14435), .B2(n9671), .A(n10083), .ZN(n15852) );
  AOI22_X1 U17829 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n19774), .B1(n19773), 
        .B2(n15852), .ZN(n14436) );
  OAI211_X1 U17830 ( .C1(n19728), .C2(n14437), .A(n14436), .B(n19927), .ZN(
        n14438) );
  AOI211_X1 U17831 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n14440), .A(n14439), 
        .B(n14438), .ZN(n14441) );
  OAI21_X1 U17832 ( .B1(n14707), .B2(n15657), .A(n14441), .ZN(P1_U2827) );
  NAND2_X1 U17833 ( .A1(n14715), .A2(n19755), .ZN(n14451) );
  NOR2_X1 U17834 ( .A1(n19725), .A2(n15697), .ZN(n14442) );
  NOR2_X1 U17835 ( .A1(n14443), .A2(n14442), .ZN(n15707) );
  NAND2_X1 U17836 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n15707), .ZN(n14450) );
  INV_X1 U17837 ( .A(n14713), .ZN(n14445) );
  INV_X1 U17838 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20605) );
  NAND2_X1 U17839 ( .A1(n15639), .A2(n19724), .ZN(n19733) );
  NOR3_X1 U17840 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20605), .A3(n19733), 
        .ZN(n14444) );
  AOI21_X1 U17841 ( .B1(n19778), .B2(n14445), .A(n14444), .ZN(n14449) );
  AOI22_X1 U17842 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_10__SCAN_IN), .B2(n19774), .ZN(n14446) );
  OAI211_X1 U17843 ( .C1(n15874), .C2(n19761), .A(n14446), .B(n19927), .ZN(
        n14447) );
  INV_X1 U17844 ( .A(n14447), .ZN(n14448) );
  NAND4_X1 U17845 ( .A1(n14451), .A2(n14450), .A3(n14449), .A4(n14448), .ZN(
        P1_U2830) );
  OAI22_X1 U17846 ( .A1(n14453), .A2(n14528), .B1(n19797), .B2(n14452), .ZN(
        P1_U2841) );
  OAI222_X1 U17847 ( .A1(n14530), .A2(n14542), .B1(n14455), .B2(n19797), .C1(
        n14454), .C2(n14528), .ZN(P1_U2842) );
  INV_X1 U17848 ( .A(n14623), .ZN(n14549) );
  INV_X1 U17849 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14456) );
  OAI222_X1 U17850 ( .A1(n14530), .A2(n14549), .B1(n14456), .B2(n19797), .C1(
        n14737), .C2(n14528), .ZN(P1_U2844) );
  AOI22_X1 U17851 ( .A1(n14749), .A2(n19792), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14520), .ZN(n14457) );
  OAI21_X1 U17852 ( .B1(n14632), .B2(n14530), .A(n14457), .ZN(P1_U2845) );
  AOI22_X1 U17853 ( .A1(n14760), .A2(n19792), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14520), .ZN(n14458) );
  OAI21_X1 U17854 ( .B1(n14558), .B2(n14530), .A(n14458), .ZN(P1_U2846) );
  NOR2_X1 U17855 ( .A1(n19797), .A2(n14459), .ZN(n14460) );
  AOI21_X1 U17856 ( .B1(n15796), .B2(n19792), .A(n14460), .ZN(n14461) );
  OAI21_X1 U17857 ( .B1(n14647), .B2(n14530), .A(n14461), .ZN(P1_U2847) );
  NOR2_X1 U17858 ( .A1(n9624), .A2(n14462), .ZN(n14463) );
  OR2_X1 U17859 ( .A1(n9649), .A2(n14463), .ZN(n15731) );
  OR2_X1 U17860 ( .A1(n14465), .A2(n14464), .ZN(n14466) );
  NAND2_X1 U17861 ( .A1(n14467), .A2(n14466), .ZN(n15628) );
  OAI22_X1 U17862 ( .A1(n15628), .A2(n14528), .B1(n14468), .B2(n19797), .ZN(
        n14469) );
  INV_X1 U17863 ( .A(n14469), .ZN(n14470) );
  OAI21_X1 U17864 ( .B1(n15731), .B2(n14530), .A(n14470), .ZN(P1_U2848) );
  INV_X1 U17865 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14472) );
  OAI222_X1 U17866 ( .A1(n14530), .A2(n14572), .B1(n14472), .B2(n19797), .C1(
        n14471), .C2(n14528), .ZN(P1_U2849) );
  AOI22_X1 U17867 ( .A1(n14788), .A2(n19792), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14520), .ZN(n14473) );
  OAI21_X1 U17868 ( .B1(n14577), .B2(n14530), .A(n14473), .ZN(P1_U2851) );
  OR2_X1 U17869 ( .A1(n14488), .A2(n14474), .ZN(n14475) );
  NAND2_X1 U17870 ( .A1(n14405), .A2(n14475), .ZN(n15651) );
  INV_X1 U17871 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14481) );
  AND2_X1 U17872 ( .A1(n14413), .A2(n14510), .ZN(n14477) );
  AND2_X1 U17873 ( .A1(n14477), .A2(n14476), .ZN(n14485) );
  OR2_X1 U17874 ( .A1(n14485), .A2(n14478), .ZN(n14479) );
  INV_X1 U17875 ( .A(n15749), .ZN(n14480) );
  OAI222_X1 U17876 ( .A1(n14528), .A2(n15651), .B1(n14481), .B2(n19797), .C1(
        n14480), .C2(n14530), .ZN(P1_U2852) );
  NOR2_X1 U17877 ( .A1(n14503), .A2(n14482), .ZN(n14490) );
  NOR2_X1 U17878 ( .A1(n14490), .A2(n14483), .ZN(n14484) );
  INV_X1 U17879 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14489) );
  NOR2_X1 U17880 ( .A1(n14495), .A2(n14486), .ZN(n14487) );
  OR2_X1 U17881 ( .A1(n14488), .A2(n14487), .ZN(n15821) );
  OAI222_X1 U17882 ( .A1(n14530), .A2(n15658), .B1(n14489), .B2(n19797), .C1(
        n15821), .C2(n14528), .ZN(P1_U2853) );
  AOI21_X1 U17883 ( .B1(n14492), .B2(n14491), .A(n14490), .ZN(n15668) );
  AND2_X1 U17884 ( .A1(n14494), .A2(n14493), .ZN(n14496) );
  OR2_X1 U17885 ( .A1(n14496), .A2(n14495), .ZN(n15829) );
  OAI22_X1 U17886 ( .A1(n15829), .A2(n14528), .B1(n14497), .B2(n19797), .ZN(
        n14498) );
  AOI21_X1 U17887 ( .B1(n15668), .B2(n19793), .A(n14498), .ZN(n14499) );
  INV_X1 U17888 ( .A(n14499), .ZN(P1_U2854) );
  AOI22_X1 U17889 ( .A1(n15836), .A2(n19792), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14520), .ZN(n14500) );
  OAI21_X1 U17890 ( .B1(n14682), .B2(n14530), .A(n14500), .ZN(P1_U2855) );
  NAND2_X1 U17891 ( .A1(n14512), .A2(n14501), .ZN(n14502) );
  OR2_X1 U17892 ( .A1(n14518), .A2(n14504), .ZN(n14505) );
  NAND2_X1 U17893 ( .A1(n14506), .A2(n14505), .ZN(n15676) );
  OAI22_X1 U17894 ( .A1(n15676), .A2(n14528), .B1(n14507), .B2(n19797), .ZN(
        n14508) );
  AOI21_X1 U17895 ( .B1(n15754), .B2(n19793), .A(n14508), .ZN(n14509) );
  INV_X1 U17896 ( .A(n14509), .ZN(P1_U2856) );
  OR2_X1 U17897 ( .A1(n14413), .A2(n14510), .ZN(n14511) );
  NAND2_X1 U17898 ( .A1(n14512), .A2(n14511), .ZN(n15683) );
  INV_X1 U17899 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14519) );
  INV_X1 U17900 ( .A(n14513), .ZN(n14516) );
  INV_X1 U17901 ( .A(n14514), .ZN(n14515) );
  AOI21_X1 U17902 ( .B1(n10083), .B2(n14516), .A(n14515), .ZN(n14517) );
  OR2_X1 U17903 ( .A1(n14518), .A2(n14517), .ZN(n15681) );
  OAI222_X1 U17904 ( .A1(n15683), .A2(n14530), .B1(n14519), .B2(n19797), .C1(
        n14528), .C2(n15681), .ZN(P1_U2857) );
  AOI22_X1 U17905 ( .A1(n15852), .A2(n19792), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14520), .ZN(n14521) );
  OAI21_X1 U17906 ( .B1(n14707), .B2(n14530), .A(n14521), .ZN(P1_U2859) );
  AOI21_X1 U17907 ( .B1(n14524), .B2(n14523), .A(n14522), .ZN(n15764) );
  INV_X1 U17908 ( .A(n15764), .ZN(n14531) );
  INV_X1 U17909 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14529) );
  NAND2_X1 U17910 ( .A1(n14526), .A2(n14525), .ZN(n14527) );
  NAND2_X1 U17911 ( .A1(n9671), .A2(n14527), .ZN(n15698) );
  OAI222_X1 U17912 ( .A1(n14531), .A2(n14530), .B1(n14529), .B2(n19797), .C1(
        n14528), .C2(n15698), .ZN(P1_U2860) );
  INV_X1 U17913 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16226) );
  AOI22_X1 U17914 ( .A1(n15723), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14604), .ZN(n14534) );
  OAI211_X1 U17915 ( .C1(n15726), .C2(n16226), .A(n14535), .B(n14534), .ZN(
        P1_U2873) );
  INV_X1 U17916 ( .A(DATAI_14_), .ZN(n14537) );
  NAND2_X1 U17917 ( .A1(n19965), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14536) );
  OAI21_X1 U17918 ( .B1(n19965), .B2(n14537), .A(n14536), .ZN(n19893) );
  INV_X1 U17919 ( .A(n19893), .ZN(n14602) );
  INV_X1 U17920 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14538) );
  OAI22_X1 U17921 ( .A1(n15721), .A2(n14602), .B1(n15730), .B2(n14538), .ZN(
        n14539) );
  AOI21_X1 U17922 ( .B1(n15723), .B2(DATAI_30_), .A(n14539), .ZN(n14541) );
  NAND2_X1 U17923 ( .A1(n14593), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14540) );
  OAI211_X1 U17924 ( .C1(n14542), .C2(n9576), .A(n14541), .B(n14540), .ZN(
        P1_U2874) );
  INV_X1 U17925 ( .A(DATAI_28_), .ZN(n14546) );
  INV_X1 U17926 ( .A(DATAI_12_), .ZN(n14544) );
  NAND2_X1 U17927 ( .A1(n19965), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14543) );
  OAI21_X1 U17928 ( .B1(n19965), .B2(n14544), .A(n14543), .ZN(n19888) );
  AOI22_X1 U17929 ( .A1(n14586), .A2(n19888), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n14604), .ZN(n14545) );
  OAI21_X1 U17930 ( .B1(n14589), .B2(n14546), .A(n14545), .ZN(n14547) );
  AOI21_X1 U17931 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14593), .A(n14547), .ZN(
        n14548) );
  OAI21_X1 U17932 ( .B1(n14549), .B2(n9576), .A(n14548), .ZN(P1_U2876) );
  INV_X1 U17933 ( .A(DATAI_27_), .ZN(n14551) );
  AOI22_X1 U17934 ( .A1(n14586), .A2(n19885), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n14604), .ZN(n14550) );
  OAI21_X1 U17935 ( .B1(n14589), .B2(n14551), .A(n14550), .ZN(n14552) );
  AOI21_X1 U17936 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14593), .A(n14552), .ZN(
        n14553) );
  OAI21_X1 U17937 ( .B1(n14632), .B2(n9576), .A(n14553), .ZN(P1_U2877) );
  INV_X1 U17938 ( .A(DATAI_26_), .ZN(n14555) );
  AOI22_X1 U17939 ( .A1(n14586), .A2(n19882), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n14604), .ZN(n14554) );
  OAI21_X1 U17940 ( .B1(n14589), .B2(n14555), .A(n14554), .ZN(n14556) );
  AOI21_X1 U17941 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14593), .A(n14556), .ZN(
        n14557) );
  OAI21_X1 U17942 ( .B1(n14558), .B2(n9576), .A(n14557), .ZN(P1_U2878) );
  INV_X1 U17943 ( .A(DATAI_25_), .ZN(n14560) );
  AOI22_X1 U17944 ( .A1(n14586), .A2(n19879), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n14604), .ZN(n14559) );
  OAI21_X1 U17945 ( .B1(n14589), .B2(n14560), .A(n14559), .ZN(n14561) );
  AOI21_X1 U17946 ( .B1(n14593), .B2(BUF1_REG_25__SCAN_IN), .A(n14561), .ZN(
        n14562) );
  OAI21_X1 U17947 ( .B1(n14647), .B2(n9576), .A(n14562), .ZN(P1_U2879) );
  OAI22_X1 U17948 ( .A1(n15721), .A2(n14564), .B1(n15730), .B2(n14563), .ZN(
        n14565) );
  AOI21_X1 U17949 ( .B1(n15723), .B2(DATAI_24_), .A(n14565), .ZN(n14567) );
  NAND2_X1 U17950 ( .A1(n14593), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14566) );
  OAI211_X1 U17951 ( .C1(n15731), .C2(n9576), .A(n14567), .B(n14566), .ZN(
        P1_U2880) );
  INV_X1 U17952 ( .A(DATAI_23_), .ZN(n14569) );
  AOI22_X1 U17953 ( .A1(n14586), .A2(n19874), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n14604), .ZN(n14568) );
  OAI21_X1 U17954 ( .B1(n14589), .B2(n14569), .A(n14568), .ZN(n14570) );
  AOI21_X1 U17955 ( .B1(n14593), .B2(BUF1_REG_23__SCAN_IN), .A(n14570), .ZN(
        n14571) );
  OAI21_X1 U17956 ( .B1(n14572), .B2(n9576), .A(n14571), .ZN(P1_U2881) );
  INV_X1 U17957 ( .A(DATAI_21_), .ZN(n14574) );
  AOI22_X1 U17958 ( .A1(n14586), .A2(n19869), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n14604), .ZN(n14573) );
  OAI21_X1 U17959 ( .B1(n14589), .B2(n14574), .A(n14573), .ZN(n14575) );
  AOI21_X1 U17960 ( .B1(n14593), .B2(BUF1_REG_21__SCAN_IN), .A(n14575), .ZN(
        n14576) );
  OAI21_X1 U17961 ( .B1(n14577), .B2(n9576), .A(n14576), .ZN(P1_U2883) );
  INV_X1 U17962 ( .A(DATAI_19_), .ZN(n14579) );
  AOI22_X1 U17963 ( .A1(n14586), .A2(n19865), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n14604), .ZN(n14578) );
  OAI21_X1 U17964 ( .B1(n14589), .B2(n14579), .A(n14578), .ZN(n14580) );
  AOI21_X1 U17965 ( .B1(n14593), .B2(BUF1_REG_19__SCAN_IN), .A(n14580), .ZN(
        n14581) );
  OAI21_X1 U17966 ( .B1(n15658), .B2(n9576), .A(n14581), .ZN(P1_U2885) );
  INV_X1 U17967 ( .A(n15668), .ZN(n14585) );
  OAI22_X1 U17968 ( .A1(n15721), .A2(n19991), .B1(n15730), .B2(n19833), .ZN(
        n14582) );
  AOI21_X1 U17969 ( .B1(n15723), .B2(DATAI_18_), .A(n14582), .ZN(n14584) );
  NAND2_X1 U17970 ( .A1(n14593), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14583) );
  OAI211_X1 U17971 ( .C1(n14585), .C2(n9576), .A(n14584), .B(n14583), .ZN(
        P1_U2886) );
  INV_X1 U17972 ( .A(DATAI_17_), .ZN(n14588) );
  AOI22_X1 U17973 ( .A1(n14586), .A2(n19859), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n14604), .ZN(n14587) );
  OAI21_X1 U17974 ( .B1(n14589), .B2(n14588), .A(n14587), .ZN(n14590) );
  AOI21_X1 U17975 ( .B1(n14593), .B2(BUF1_REG_17__SCAN_IN), .A(n14590), .ZN(
        n14591) );
  OAI21_X1 U17976 ( .B1(n14682), .B2(n9576), .A(n14591), .ZN(P1_U2887) );
  INV_X1 U17977 ( .A(n15754), .ZN(n14596) );
  OAI22_X1 U17978 ( .A1(n15721), .A2(n19978), .B1(n15730), .B2(n20815), .ZN(
        n14592) );
  AOI21_X1 U17979 ( .B1(n15723), .B2(DATAI_16_), .A(n14592), .ZN(n14595) );
  NAND2_X1 U17980 ( .A1(n14593), .A2(BUF1_REG_16__SCAN_IN), .ZN(n14594) );
  OAI211_X1 U17981 ( .C1(n14596), .C2(n9576), .A(n14595), .B(n14594), .ZN(
        P1_U2888) );
  INV_X1 U17982 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19804) );
  INV_X1 U17983 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14597) );
  NOR2_X1 U17984 ( .A1(n19966), .A2(n14597), .ZN(n14598) );
  AOI21_X1 U17985 ( .B1(DATAI_15_), .B2(n19966), .A(n14598), .ZN(n19902) );
  OAI222_X1 U17986 ( .A1(n15683), .A2(n9576), .B1(n15730), .B2(n19804), .C1(
        n14601), .C2(n19902), .ZN(P1_U2889) );
  AOI21_X1 U17987 ( .B1(n14599), .B2(n14432), .A(n14413), .ZN(n15760) );
  INV_X1 U17988 ( .A(n15760), .ZN(n14603) );
  INV_X1 U17989 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14600) );
  OAI222_X1 U17990 ( .A1(n14603), .A2(n9576), .B1(n14602), .B2(n14601), .C1(
        n14600), .C2(n15730), .ZN(P1_U2890) );
  AOI22_X1 U17991 ( .A1(n15727), .A2(n19890), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14604), .ZN(n14605) );
  OAI21_X1 U17992 ( .B1(n14707), .B2(n9576), .A(n14605), .ZN(P1_U2891) );
  AOI21_X1 U17993 ( .B1(n14607), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14606), .ZN(n14722) );
  NOR2_X1 U17994 ( .A1(n19927), .A2(n20807), .ZN(n14720) );
  AOI21_X1 U17995 ( .B1(n19914), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14720), .ZN(n14608) );
  OAI21_X1 U17996 ( .B1(n19912), .B2(n14609), .A(n14608), .ZN(n14610) );
  AOI21_X1 U17997 ( .B1(n14611), .B2(n15781), .A(n14610), .ZN(n14612) );
  OAI21_X1 U17998 ( .B1(n14722), .B2(n19708), .A(n14612), .ZN(P1_U2969) );
  NAND2_X1 U17999 ( .A1(n14777), .A2(n14614), .ZN(n14633) );
  NAND2_X1 U18000 ( .A1(n14613), .A2(n14633), .ZN(n14618) );
  OAI21_X1 U18001 ( .B1(n14615), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14618), .ZN(n14617) );
  MUX2_X1 U18002 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14750), .S(
        n14764), .Z(n14616) );
  OAI211_X1 U18003 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14618), .A(
        n14617), .B(n14616), .ZN(n14619) );
  XNOR2_X1 U18004 ( .A(n14619), .B(n14731), .ZN(n14738) );
  INV_X1 U18005 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20636) );
  NOR2_X1 U18006 ( .A1(n19927), .A2(n20636), .ZN(n14732) );
  AOI21_X1 U18007 ( .B1(n19914), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14732), .ZN(n14620) );
  OAI21_X1 U18008 ( .B1(n19912), .B2(n14621), .A(n14620), .ZN(n14622) );
  AOI21_X1 U18009 ( .B1(n14623), .B2(n15781), .A(n14622), .ZN(n14624) );
  OAI21_X1 U18010 ( .B1(n19708), .B2(n14738), .A(n14624), .ZN(P1_U2971) );
  XNOR2_X1 U18011 ( .A(n14627), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14744) );
  NAND2_X1 U18012 ( .A1(n14744), .A2(n19917), .ZN(n14631) );
  NOR2_X1 U18013 ( .A1(n19927), .A2(n20634), .ZN(n14748) );
  NOR2_X1 U18014 ( .A1(n14677), .A2(n20813), .ZN(n14628) );
  AOI211_X1 U18015 ( .C1(n19916), .C2(n14629), .A(n14748), .B(n14628), .ZN(
        n14630) );
  OAI211_X1 U18016 ( .C1(n14764), .C2(n14613), .A(n14634), .B(n14633), .ZN(
        n14635) );
  XOR2_X1 U18017 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14635), .Z(
        n14762) );
  NAND2_X1 U18018 ( .A1(n19913), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14755) );
  NAND2_X1 U18019 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14636) );
  OAI211_X1 U18020 ( .C1(n19912), .C2(n14637), .A(n14755), .B(n14636), .ZN(
        n14638) );
  AOI21_X1 U18021 ( .B1(n14639), .B2(n15781), .A(n14638), .ZN(n14640) );
  OAI21_X1 U18022 ( .B1(n19708), .B2(n14762), .A(n14640), .ZN(P1_U2973) );
  NOR3_X1 U18023 ( .A1(n14613), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14643) );
  NAND2_X1 U18024 ( .A1(n14641), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14766) );
  NOR2_X1 U18025 ( .A1(n14766), .A2(n15793), .ZN(n14642) );
  MUX2_X1 U18026 ( .A(n14643), .B(n14642), .S(n14777), .Z(n14644) );
  XNOR2_X1 U18027 ( .A(n14644), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15795) );
  INV_X1 U18028 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14645) );
  OAI22_X1 U18029 ( .A1(n14677), .A2(n14646), .B1(n19927), .B2(n14645), .ZN(
        n14649) );
  NOR2_X1 U18030 ( .A1(n14647), .A2(n19967), .ZN(n14648) );
  AOI211_X1 U18031 ( .C1(n19916), .C2(n14650), .A(n14649), .B(n14648), .ZN(
        n14651) );
  OAI21_X1 U18032 ( .B1(n19708), .B2(n15795), .A(n14651), .ZN(P1_U2974) );
  XNOR2_X1 U18033 ( .A(n15769), .B(n15808), .ZN(n14652) );
  XNOR2_X1 U18034 ( .A(n14613), .B(n14652), .ZN(n15803) );
  INV_X1 U18035 ( .A(n14653), .ZN(n14655) );
  AOI22_X1 U18036 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14654) );
  OAI21_X1 U18037 ( .B1(n19912), .B2(n14655), .A(n14654), .ZN(n14656) );
  AOI21_X1 U18038 ( .B1(n14657), .B2(n15781), .A(n14656), .ZN(n14658) );
  OAI21_X1 U18039 ( .B1(n15803), .B2(n19708), .A(n14658), .ZN(P1_U2976) );
  AOI21_X1 U18040 ( .B1(n14764), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n14778), .ZN(n14776) );
  INV_X1 U18041 ( .A(n14776), .ZN(n14795) );
  NAND2_X1 U18042 ( .A1(n14764), .A2(n14798), .ZN(n14794) );
  OAI21_X1 U18043 ( .B1(n14764), .B2(n14798), .A(n14794), .ZN(n14659) );
  XNOR2_X1 U18044 ( .A(n14795), .B(n14659), .ZN(n15820) );
  INV_X1 U18045 ( .A(n15658), .ZN(n14663) );
  INV_X1 U18046 ( .A(n15653), .ZN(n14661) );
  AOI22_X1 U18047 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14660) );
  OAI21_X1 U18048 ( .B1(n19912), .B2(n14661), .A(n14660), .ZN(n14662) );
  AOI21_X1 U18049 ( .B1(n14663), .B2(n15781), .A(n14662), .ZN(n14664) );
  OAI21_X1 U18050 ( .B1(n15820), .B2(n19708), .A(n14664), .ZN(P1_U2980) );
  INV_X1 U18051 ( .A(n14778), .ZN(n14665) );
  OAI21_X1 U18052 ( .B1(n14667), .B2(n14666), .A(n14665), .ZN(n15830) );
  AOI22_X1 U18053 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14668) );
  OAI21_X1 U18054 ( .B1(n19912), .B2(n15665), .A(n14668), .ZN(n14669) );
  AOI21_X1 U18055 ( .B1(n15668), .B2(n15781), .A(n14669), .ZN(n14670) );
  OAI21_X1 U18056 ( .B1(n19708), .B2(n15830), .A(n14670), .ZN(P1_U2981) );
  NAND2_X1 U18057 ( .A1(n14764), .A2(n14815), .ZN(n14674) );
  OAI21_X1 U18058 ( .B1(n14809), .B2(n14672), .A(n14671), .ZN(n14673) );
  MUX2_X1 U18059 ( .A(n14764), .B(n14674), .S(n14673), .Z(n14675) );
  XNOR2_X1 U18060 ( .A(n14675), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15837) );
  NAND2_X1 U18061 ( .A1(n15837), .A2(n19917), .ZN(n14681) );
  INV_X1 U18062 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14676) );
  OAI22_X1 U18063 ( .A1(n14677), .A2(n14425), .B1(n19927), .B2(n14676), .ZN(
        n14678) );
  AOI21_X1 U18064 ( .B1(n19916), .B2(n14679), .A(n14678), .ZN(n14680) );
  OAI211_X1 U18065 ( .C1(n19967), .C2(n14682), .A(n14681), .B(n14680), .ZN(
        P1_U2982) );
  NOR2_X1 U18066 ( .A1(n14684), .A2(n14683), .ZN(n14810) );
  INV_X1 U18067 ( .A(n14685), .ZN(n14686) );
  NOR2_X1 U18068 ( .A1(n14810), .A2(n14686), .ZN(n14688) );
  AOI21_X1 U18069 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14764), .A(
        n14807), .ZN(n14687) );
  XNOR2_X1 U18070 ( .A(n14688), .B(n14687), .ZN(n15845) );
  INV_X1 U18071 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n14689) );
  NOR2_X1 U18072 ( .A1(n19927), .A2(n14689), .ZN(n15842) );
  AOI21_X1 U18073 ( .B1(n19914), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15842), .ZN(n14691) );
  NAND2_X1 U18074 ( .A1(n19916), .A2(n15682), .ZN(n14690) );
  OAI211_X1 U18075 ( .C1(n15683), .C2(n19967), .A(n14691), .B(n14690), .ZN(
        n14692) );
  AOI21_X1 U18076 ( .B1(n15845), .B2(n19917), .A(n14692), .ZN(n14693) );
  INV_X1 U18077 ( .A(n14693), .ZN(P1_U2984) );
  OAI21_X1 U18078 ( .B1(n13481), .B2(n14695), .A(n14694), .ZN(n14821) );
  INV_X1 U18079 ( .A(n14699), .ZN(n14696) );
  NAND2_X1 U18080 ( .A1(n14697), .A2(n14696), .ZN(n14822) );
  NOR2_X1 U18081 ( .A1(n14821), .A2(n14822), .ZN(n14698) );
  NOR2_X1 U18082 ( .A1(n14699), .A2(n14698), .ZN(n14701) );
  XNOR2_X1 U18083 ( .A(n14701), .B(n14700), .ZN(n15854) );
  NAND2_X1 U18084 ( .A1(n15854), .A2(n19917), .ZN(n14706) );
  INV_X1 U18085 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14702) );
  NOR2_X1 U18086 ( .A1(n19927), .A2(n14702), .ZN(n15851) );
  NOR2_X1 U18087 ( .A1(n19912), .A2(n14703), .ZN(n14704) );
  AOI211_X1 U18088 ( .C1(n19914), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15851), .B(n14704), .ZN(n14705) );
  OAI211_X1 U18089 ( .C1(n19967), .C2(n14707), .A(n14706), .B(n14705), .ZN(
        P1_U2986) );
  AND2_X1 U18090 ( .A1(n9582), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14710) );
  XNOR2_X1 U18091 ( .A(n13481), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14709) );
  MUX2_X1 U18092 ( .A(n14710), .B(n14709), .S(n14777), .Z(n14711) );
  NOR3_X1 U18093 ( .A1(n9582), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14777), .ZN(n15770) );
  NOR2_X1 U18094 ( .A1(n14711), .A2(n15770), .ZN(n15868) );
  AOI22_X1 U18095 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14712) );
  OAI21_X1 U18096 ( .B1(n19912), .B2(n14713), .A(n14712), .ZN(n14714) );
  AOI21_X1 U18097 ( .B1(n14715), .B2(n15781), .A(n14714), .ZN(n14716) );
  OAI21_X1 U18098 ( .B1(n15868), .B2(n19708), .A(n14716), .ZN(P1_U2989) );
  NAND3_X1 U18099 ( .A1(n14745), .A2(n11921), .A3(n14723), .ZN(n14724) );
  OAI211_X1 U18100 ( .C1(n14726), .C2(n19955), .A(n14725), .B(n14724), .ZN(
        n14727) );
  AOI21_X1 U18101 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14728), .A(
        n14727), .ZN(n14729) );
  NOR2_X1 U18102 ( .A1(n14756), .A2(n14731), .ZN(n14742) );
  INV_X1 U18103 ( .A(n14751), .ZN(n14741) );
  INV_X1 U18104 ( .A(n14732), .ZN(n14736) );
  NAND3_X1 U18105 ( .A1(n14745), .A2(n14734), .A3(n14733), .ZN(n14735) );
  OAI211_X1 U18106 ( .C1(n14737), .C2(n19955), .A(n14736), .B(n14735), .ZN(
        n14740) );
  NOR2_X1 U18107 ( .A1(n14738), .A2(n19925), .ZN(n14739) );
  INV_X1 U18108 ( .A(n14743), .ZN(P1_U3003) );
  INV_X1 U18109 ( .A(n14744), .ZN(n14754) );
  INV_X1 U18110 ( .A(n14745), .ZN(n14746) );
  NOR2_X1 U18111 ( .A1(n14746), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14747) );
  AOI211_X1 U18112 ( .C1(n14749), .C2(n19936), .A(n14748), .B(n14747), .ZN(
        n14753) );
  OR3_X1 U18113 ( .A1(n14751), .A2(n14756), .A3(n14750), .ZN(n14752) );
  INV_X1 U18114 ( .A(n14755), .ZN(n14759) );
  INV_X1 U18115 ( .A(n15792), .ZN(n15802) );
  AOI21_X1 U18116 ( .B1(n15802), .B2(n9715), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14757) );
  NOR2_X1 U18117 ( .A1(n14757), .A2(n14756), .ZN(n14758) );
  AOI211_X1 U18118 ( .C1(n14760), .C2(n19936), .A(n14759), .B(n14758), .ZN(
        n14761) );
  OAI21_X1 U18119 ( .B1(n14762), .B2(n19925), .A(n14761), .ZN(P1_U3005) );
  INV_X1 U18120 ( .A(n14613), .ZN(n14763) );
  NAND2_X1 U18121 ( .A1(n14763), .A2(n14766), .ZN(n14765) );
  MUX2_X1 U18122 ( .A(n14766), .B(n14765), .S(n14764), .Z(n14767) );
  XNOR2_X1 U18123 ( .A(n14767), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15733) );
  INV_X1 U18124 ( .A(n15733), .ZN(n14775) );
  NOR2_X1 U18125 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n14768), .ZN(
        n14770) );
  OAI21_X1 U18126 ( .B1(n14770), .B2(n14769), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14774) );
  NOR3_X1 U18127 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15808), .A3(
        n15792), .ZN(n14772) );
  NOR2_X1 U18128 ( .A1(n15628), .A2(n19955), .ZN(n14771) );
  AOI211_X1 U18129 ( .C1(n19913), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14772), 
        .B(n14771), .ZN(n14773) );
  OAI211_X1 U18130 ( .C1(n14775), .C2(n19925), .A(n14774), .B(n14773), .ZN(
        P1_U3007) );
  NAND2_X1 U18131 ( .A1(n14776), .A2(n14796), .ZN(n14779) );
  NAND2_X1 U18132 ( .A1(n14778), .A2(n14777), .ZN(n14793) );
  AOI22_X1 U18133 ( .A1(n14779), .A2(n14793), .B1(n14787), .B2(n14794), .ZN(
        n14780) );
  XNOR2_X1 U18134 ( .A(n14780), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15748) );
  INV_X1 U18135 ( .A(n14781), .ZN(n14786) );
  NOR2_X1 U18136 ( .A1(n19947), .A2(n14785), .ZN(n14782) );
  AOI22_X1 U18137 ( .A1(n14784), .A2(n14783), .B1(n10093), .B2(n14782), .ZN(
        n14802) );
  OAI21_X1 U18138 ( .B1(n14785), .B2(n14801), .A(n14802), .ZN(n15853) );
  NAND2_X1 U18139 ( .A1(n14786), .A2(n15853), .ZN(n15826) );
  NOR2_X1 U18140 ( .A1(n14787), .A2(n15826), .ZN(n15814) );
  AOI22_X1 U18141 ( .A1(n14788), .A2(n19936), .B1(n19913), .B2(
        P1_REIP_REG_21__SCAN_IN), .ZN(n14789) );
  OAI21_X1 U18142 ( .B1(n20808), .B2(n14790), .A(n14789), .ZN(n14791) );
  AOI21_X1 U18143 ( .B1(n15814), .B2(n20808), .A(n14791), .ZN(n14792) );
  OAI21_X1 U18144 ( .B1(n15748), .B2(n19925), .A(n14792), .ZN(P1_U3010) );
  OAI22_X1 U18145 ( .A1(n14795), .A2(n14794), .B1(n14798), .B2(n14793), .ZN(
        n14797) );
  XNOR2_X1 U18146 ( .A(n14797), .B(n14796), .ZN(n15750) );
  INV_X1 U18147 ( .A(n15750), .ZN(n14806) );
  NOR2_X1 U18148 ( .A1(n15651), .A2(n19955), .ZN(n14800) );
  NOR3_X1 U18149 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14798), .A3(
        n15826), .ZN(n14799) );
  AOI211_X1 U18150 ( .C1(n19913), .C2(P1_REIP_REG_20__SCAN_IN), .A(n14800), 
        .B(n14799), .ZN(n14805) );
  AOI21_X1 U18151 ( .B1(n14802), .B2(n14801), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14803) );
  OAI21_X1 U18152 ( .B1(n15819), .B2(n14803), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14804) );
  OAI211_X1 U18153 ( .C1(n14806), .C2(n19925), .A(n14805), .B(n14804), .ZN(
        P1_U3011) );
  INV_X1 U18154 ( .A(n14807), .ZN(n14808) );
  OAI21_X1 U18155 ( .B1(n14810), .B2(n14809), .A(n14808), .ZN(n14811) );
  XOR2_X1 U18156 ( .A(n14812), .B(n14811), .Z(n15755) );
  INV_X1 U18157 ( .A(n14813), .ZN(n15828) );
  NOR2_X1 U18158 ( .A1(n15828), .A2(n14814), .ZN(n15844) );
  OAI21_X1 U18159 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15844), .ZN(n14816) );
  AOI21_X1 U18160 ( .B1(n14814), .B2(n15889), .A(n15850), .ZN(n15849) );
  OAI22_X1 U18161 ( .A1(n15835), .A2(n14816), .B1(n15849), .B2(n14815), .ZN(
        n14819) );
  INV_X1 U18162 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14817) );
  OAI22_X1 U18163 ( .A1(n15676), .A2(n19955), .B1(n19927), .B2(n14817), .ZN(
        n14818) );
  AOI211_X1 U18164 ( .C1(n15755), .C2(n19952), .A(n14819), .B(n14818), .ZN(
        n14820) );
  INV_X1 U18165 ( .A(n14820), .ZN(P1_U3015) );
  NAND2_X1 U18166 ( .A1(n14826), .A2(n15892), .ZN(n14834) );
  XOR2_X1 U18167 ( .A(n14822), .B(n14821), .Z(n15768) );
  OR2_X1 U18168 ( .A1(n15768), .A2(n19925), .ZN(n14833) );
  INV_X1 U18169 ( .A(n15860), .ZN(n14825) );
  AOI21_X1 U18170 ( .B1(n14825), .B2(n14824), .A(n14823), .ZN(n14828) );
  AOI21_X1 U18171 ( .B1(n15870), .B2(n14826), .A(n19946), .ZN(n14827) );
  NOR3_X1 U18172 ( .A1(n14828), .A2(n19948), .A3(n14827), .ZN(n15865) );
  OAI21_X1 U18173 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n13070), .A(
        n15865), .ZN(n14831) );
  INV_X1 U18174 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n14829) );
  OAI22_X1 U18175 ( .A1(n15698), .A2(n19955), .B1(n19927), .B2(n14829), .ZN(
        n14830) );
  AOI21_X1 U18176 ( .B1(n14831), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14830), .ZN(n14832) );
  OAI211_X1 U18177 ( .C1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n14834), .A(
        n14833), .B(n14832), .ZN(P1_U3019) );
  OAI21_X1 U18178 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20053), .A(n20514), 
        .ZN(n14835) );
  OAI21_X1 U18179 ( .B1(n14836), .B2(n12955), .A(n14835), .ZN(n14837) );
  MUX2_X1 U18180 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14837), .S(
        n19963), .Z(P1_U3477) );
  INV_X1 U18181 ( .A(n12955), .ZN(n20471) );
  NAND3_X1 U18182 ( .A1(n14840), .A2(n14839), .A3(n14838), .ZN(n14841) );
  OAI21_X1 U18183 ( .B1(n15558), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n14841), .ZN(n14842) );
  AOI21_X1 U18184 ( .B1(n20471), .B2(n14843), .A(n14842), .ZN(n15560) );
  INV_X1 U18185 ( .A(n19700), .ZN(n15913) );
  AOI22_X1 U18186 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19951), .B2(n12023), .ZN(
        n14852) );
  INV_X1 U18187 ( .A(n14852), .ZN(n14846) );
  NOR2_X1 U18188 ( .A1(n20570), .A2(n19947), .ZN(n14851) );
  NOR3_X1 U18189 ( .A1(n12813), .A2(n14844), .A3(n14857), .ZN(n14845) );
  AOI21_X1 U18190 ( .B1(n14846), .B2(n14851), .A(n14845), .ZN(n14847) );
  OAI21_X1 U18191 ( .B1(n15560), .B2(n15913), .A(n14847), .ZN(n14848) );
  MUX2_X1 U18192 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14848), .S(
        n15918), .Z(P1_U3473) );
  INV_X1 U18193 ( .A(n14857), .ZN(n14849) );
  AOI22_X1 U18194 ( .A1(n14852), .A2(n14851), .B1(n14850), .B2(n14849), .ZN(
        n14853) );
  OAI21_X1 U18195 ( .B1(n14854), .B2(n15913), .A(n14853), .ZN(n14855) );
  MUX2_X1 U18196 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14855), .S(
        n15918), .Z(P1_U3472) );
  INV_X1 U18197 ( .A(n14856), .ZN(n14858) );
  OAI22_X1 U18198 ( .A1(n14859), .A2(n15913), .B1(n14858), .B2(n14857), .ZN(
        n14860) );
  MUX2_X1 U18199 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14860), .S(
        n15918), .Z(P1_U3469) );
  MUX2_X1 U18200 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n15931), .S(n14918), .Z(
        P2_U2856) );
  INV_X1 U18201 ( .A(n14861), .ZN(n14932) );
  NAND2_X1 U18202 ( .A1(n14862), .A2(n14863), .ZN(n14931) );
  NAND3_X1 U18203 ( .A1(n14932), .A2(n14907), .A3(n14931), .ZN(n14865) );
  NAND2_X1 U18204 ( .A1(n12420), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14864) );
  OAI211_X1 U18205 ( .C1(n12420), .C2(n15146), .A(n14865), .B(n14864), .ZN(
        P2_U2858) );
  NAND2_X1 U18206 ( .A1(n14234), .A2(n14866), .ZN(n14868) );
  XNOR2_X1 U18207 ( .A(n14868), .B(n14867), .ZN(n14945) );
  NAND2_X1 U18208 ( .A1(n12420), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14870) );
  NAND2_X1 U18209 ( .A1(n13525), .A2(n14918), .ZN(n14869) );
  OAI211_X1 U18210 ( .C1(n14945), .C2(n14929), .A(n14870), .B(n14869), .ZN(
        P2_U2859) );
  AOI21_X1 U18211 ( .B1(n14873), .B2(n14872), .A(n14871), .ZN(n14946) );
  NAND2_X1 U18212 ( .A1(n14946), .A2(n14907), .ZN(n14875) );
  NAND2_X1 U18213 ( .A1(n12420), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14874) );
  OAI211_X1 U18214 ( .C1(n12420), .C2(n15979), .A(n14875), .B(n14874), .ZN(
        P2_U2860) );
  OAI21_X1 U18215 ( .B1(n14876), .B2(n14878), .A(n14877), .ZN(n14963) );
  NOR2_X1 U18216 ( .A1(n14879), .A2(n14880), .ZN(n14881) );
  OR2_X1 U18217 ( .A1(n13533), .A2(n14881), .ZN(n15980) );
  NOR2_X1 U18218 ( .A1(n15980), .A2(n12420), .ZN(n14882) );
  AOI21_X1 U18219 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n12420), .A(n14882), .ZN(
        n14883) );
  OAI21_X1 U18220 ( .B1(n14963), .B2(n14929), .A(n14883), .ZN(P2_U2861) );
  OAI21_X1 U18221 ( .B1(n14884), .B2(n14886), .A(n14885), .ZN(n14974) );
  AND2_X1 U18222 ( .A1(n14897), .A2(n14887), .ZN(n14888) );
  OR2_X1 U18223 ( .A1(n14888), .A2(n14879), .ZN(n15999) );
  MUX2_X1 U18224 ( .A(n15999), .B(n14889), .S(n12420), .Z(n14890) );
  OAI21_X1 U18225 ( .B1(n14974), .B2(n14929), .A(n14890), .ZN(P2_U2862) );
  AOI21_X1 U18226 ( .B1(n14891), .B2(n14892), .A(n9605), .ZN(n14893) );
  XOR2_X1 U18227 ( .A(n14894), .B(n14893), .Z(n14982) );
  NAND2_X1 U18228 ( .A1(n14901), .A2(n14895), .ZN(n14896) );
  AND2_X1 U18229 ( .A1(n14897), .A2(n14896), .ZN(n16009) );
  NOR2_X1 U18230 ( .A1(n14918), .A2(n14898), .ZN(n14899) );
  AOI21_X1 U18231 ( .B1(n14918), .B2(n16009), .A(n14899), .ZN(n14900) );
  OAI21_X1 U18232 ( .B1(n14982), .B2(n14929), .A(n14900), .ZN(P2_U2863) );
  OAI21_X1 U18233 ( .B1(n14902), .B2(n14913), .A(n14901), .ZN(n16039) );
  NOR2_X1 U18234 ( .A1(n14903), .A2(n14904), .ZN(n14906) );
  NOR2_X1 U18235 ( .A1(n14906), .A2(n14905), .ZN(n16025) );
  NAND2_X1 U18236 ( .A1(n16025), .A2(n14907), .ZN(n14909) );
  NAND2_X1 U18237 ( .A1(n12420), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14908) );
  OAI211_X1 U18238 ( .C1(n16039), .C2(n12420), .A(n14909), .B(n14908), .ZN(
        P2_U2864) );
  OR2_X1 U18239 ( .A1(n14068), .A2(n14920), .ZN(n14921) );
  INV_X1 U18240 ( .A(n14921), .ZN(n14912) );
  INV_X1 U18241 ( .A(n14910), .ZN(n14911) );
  OAI21_X1 U18242 ( .B1(n14912), .B2(n14911), .A(n14131), .ZN(n14992) );
  AOI21_X1 U18243 ( .B1(n14915), .B2(n14914), .A(n14913), .ZN(n16048) );
  INV_X1 U18244 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n14916) );
  NOR2_X1 U18245 ( .A1(n14918), .A2(n14916), .ZN(n14917) );
  AOI21_X1 U18246 ( .B1(n16048), .B2(n14918), .A(n14917), .ZN(n14919) );
  OAI21_X1 U18247 ( .B1(n14992), .B2(n14929), .A(n14919), .ZN(P2_U2865) );
  INV_X1 U18248 ( .A(n14920), .ZN(n14922) );
  OAI21_X1 U18249 ( .B1(n14090), .B2(n14922), .A(n14921), .ZN(n14999) );
  MUX2_X1 U18250 ( .A(n15213), .B(n11112), .S(n12420), .Z(n14923) );
  OAI21_X1 U18251 ( .B1(n14999), .B2(n14929), .A(n14923), .ZN(P2_U2866) );
  AND2_X1 U18252 ( .A1(n9622), .A2(n14924), .ZN(n14926) );
  OR2_X1 U18253 ( .A1(n14926), .A2(n14925), .ZN(n15235) );
  NOR2_X1 U18254 ( .A1(n15235), .A2(n12420), .ZN(n14927) );
  AOI21_X1 U18255 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n12420), .A(n14927), .ZN(
        n14928) );
  OAI21_X1 U18256 ( .B1(n14930), .B2(n14929), .A(n14928), .ZN(P2_U2868) );
  NAND3_X1 U18257 ( .A1(n14932), .A2(n18922), .A3(n14931), .ZN(n14939) );
  INV_X1 U18258 ( .A(n15005), .ZN(n16024) );
  AOI22_X1 U18259 ( .A1(n16024), .A2(n18875), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n18920), .ZN(n14938) );
  AOI22_X1 U18260 ( .A1(n18864), .A2(BUF2_REG_29__SCAN_IN), .B1(n18865), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14937) );
  INV_X1 U18261 ( .A(n15152), .ZN(n15950) );
  NAND2_X1 U18262 ( .A1(n15950), .A2(n18921), .ZN(n14936) );
  NAND4_X1 U18263 ( .A1(n14939), .A2(n14938), .A3(n14937), .A4(n14936), .ZN(
        P2_U2890) );
  INV_X1 U18264 ( .A(n15969), .ZN(n14942) );
  OAI22_X1 U18265 ( .A1(n15005), .A2(n18878), .B1(n18892), .B2(n14940), .ZN(
        n14941) );
  AOI21_X1 U18266 ( .B1(n18921), .B2(n14942), .A(n14941), .ZN(n14944) );
  AOI22_X1 U18267 ( .A1(n18864), .A2(BUF2_REG_28__SCAN_IN), .B1(n18865), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14943) );
  OAI211_X1 U18268 ( .C1(n14945), .C2(n18868), .A(n14944), .B(n14943), .ZN(
        P2_U2891) );
  INV_X1 U18269 ( .A(n14946), .ZN(n14954) );
  OAI22_X1 U18270 ( .A1(n15005), .A2(n18882), .B1(n18892), .B2(n14947), .ZN(
        n14951) );
  INV_X1 U18271 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n14949) );
  INV_X1 U18272 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n14948) );
  OAI22_X1 U18273 ( .A1(n15008), .A2(n14949), .B1(n15006), .B2(n14948), .ZN(
        n14950) );
  AOI211_X1 U18274 ( .C1(n18921), .C2(n14952), .A(n14951), .B(n14950), .ZN(
        n14953) );
  OAI21_X1 U18275 ( .B1(n14954), .B2(n18868), .A(n14953), .ZN(P2_U2892) );
  OR2_X1 U18276 ( .A1(n14965), .A2(n14955), .ZN(n14956) );
  NAND2_X1 U18277 ( .A1(n14957), .A2(n14956), .ZN(n15986) );
  INV_X1 U18278 ( .A(n15986), .ZN(n15164) );
  OAI22_X1 U18279 ( .A1(n15005), .A2(n18883), .B1(n18892), .B2(n14958), .ZN(
        n14961) );
  INV_X1 U18280 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n14959) );
  INV_X1 U18281 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16233) );
  OAI22_X1 U18282 ( .A1(n15008), .A2(n14959), .B1(n15006), .B2(n16233), .ZN(
        n14960) );
  AOI211_X1 U18283 ( .C1(n18921), .C2(n15164), .A(n14961), .B(n14960), .ZN(
        n14962) );
  OAI21_X1 U18284 ( .B1(n14963), .B2(n18868), .A(n14962), .ZN(P2_U2893) );
  AND2_X1 U18285 ( .A1(n14977), .A2(n14964), .ZN(n14966) );
  OR2_X1 U18286 ( .A1(n14966), .A2(n14965), .ZN(n15993) );
  INV_X1 U18287 ( .A(n15993), .ZN(n14972) );
  OAI22_X1 U18288 ( .A1(n15005), .A2(n18887), .B1(n18892), .B2(n14967), .ZN(
        n14971) );
  INV_X1 U18289 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n14969) );
  INV_X1 U18290 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14968) );
  OAI22_X1 U18291 ( .A1(n15008), .A2(n14969), .B1(n15006), .B2(n14968), .ZN(
        n14970) );
  AOI211_X1 U18292 ( .C1(n18921), .C2(n14972), .A(n14971), .B(n14970), .ZN(
        n14973) );
  OAI21_X1 U18293 ( .B1(n14974), .B2(n18868), .A(n14973), .ZN(P2_U2894) );
  NAND2_X1 U18294 ( .A1(n16013), .A2(n14975), .ZN(n14976) );
  NAND2_X1 U18295 ( .A1(n14977), .A2(n14976), .ZN(n16006) );
  INV_X1 U18296 ( .A(n16006), .ZN(n15187) );
  OAI22_X1 U18297 ( .A1(n15005), .A2(n18888), .B1(n18892), .B2(n14978), .ZN(
        n14979) );
  AOI21_X1 U18298 ( .B1(n18921), .B2(n15187), .A(n14979), .ZN(n14981) );
  AOI22_X1 U18299 ( .A1(n18864), .A2(BUF2_REG_24__SCAN_IN), .B1(n18865), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14980) );
  OAI211_X1 U18300 ( .C1(n14982), .C2(n18868), .A(n14981), .B(n14980), .ZN(
        P2_U2895) );
  OR2_X1 U18301 ( .A1(n12233), .A2(n14983), .ZN(n14985) );
  INV_X1 U18302 ( .A(n16011), .ZN(n14984) );
  NAND2_X1 U18303 ( .A1(n14985), .A2(n14984), .ZN(n15553) );
  INV_X1 U18304 ( .A(n15553), .ZN(n15204) );
  OAI22_X1 U18305 ( .A1(n15005), .A2(n19044), .B1(n18892), .B2(n14986), .ZN(
        n14990) );
  INV_X1 U18306 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n14988) );
  INV_X1 U18307 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14987) );
  OAI22_X1 U18308 ( .A1(n15008), .A2(n14988), .B1(n15006), .B2(n14987), .ZN(
        n14989) );
  AOI211_X1 U18309 ( .C1(n18921), .C2(n15204), .A(n14990), .B(n14989), .ZN(
        n14991) );
  OAI21_X1 U18310 ( .B1(n14992), .B2(n18868), .A(n14991), .ZN(P2_U2897) );
  OAI22_X1 U18311 ( .A1(n15005), .A2(n19040), .B1(n18892), .B2(n14993), .ZN(
        n14997) );
  INV_X1 U18312 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14995) );
  INV_X1 U18313 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14994) );
  OAI22_X1 U18314 ( .A1(n15008), .A2(n14995), .B1(n15006), .B2(n14994), .ZN(
        n14996) );
  AOI211_X1 U18315 ( .C1(n18921), .C2(n15210), .A(n14997), .B(n14996), .ZN(
        n14998) );
  OAI21_X1 U18316 ( .B1(n14999), .B2(n18868), .A(n14998), .ZN(P2_U2898) );
  NOR2_X1 U18317 ( .A1(n15001), .A2(n15000), .ZN(n15002) );
  OR2_X1 U18318 ( .A1(n12234), .A2(n15002), .ZN(n18650) );
  INV_X1 U18319 ( .A(n18650), .ZN(n15011) );
  OAI22_X1 U18320 ( .A1(n15005), .A2(n15004), .B1(n18892), .B2(n15003), .ZN(
        n15010) );
  INV_X1 U18321 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n15007) );
  OAI22_X1 U18322 ( .A1(n15008), .A2(n15007), .B1(n15006), .B2(n16242), .ZN(
        n15009) );
  AOI211_X1 U18323 ( .C1(n18921), .C2(n15011), .A(n15010), .B(n15009), .ZN(
        n15012) );
  OAI21_X1 U18324 ( .B1(n15013), .B2(n18868), .A(n15012), .ZN(P2_U2899) );
  NAND2_X1 U18325 ( .A1(n15015), .A2(n15014), .ZN(n15020) );
  INV_X1 U18326 ( .A(n15016), .ZN(n15017) );
  NOR2_X1 U18327 ( .A1(n15018), .A2(n15017), .ZN(n15019) );
  XNOR2_X1 U18328 ( .A(n15020), .B(n15019), .ZN(n15145) );
  XOR2_X1 U18329 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15021), .Z(
        n15143) );
  XNOR2_X1 U18330 ( .A(n13988), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15940) );
  INV_X1 U18331 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n15022) );
  NOR2_X1 U18332 ( .A1(n19016), .A2(n15022), .ZN(n15136) );
  AOI21_X1 U18333 ( .B1(n18979), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15136), .ZN(n15024) );
  NAND2_X1 U18334 ( .A1(n14315), .A2(n18988), .ZN(n15023) );
  OAI211_X1 U18335 ( .C1(n15940), .C2(n18992), .A(n15024), .B(n15023), .ZN(
        n15025) );
  AOI21_X1 U18336 ( .B1(n15143), .B2(n16114), .A(n15025), .ZN(n15026) );
  OAI21_X1 U18337 ( .B1(n15145), .B2(n18982), .A(n15026), .ZN(P2_U2984) );
  OR2_X1 U18338 ( .A1(n15175), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15027) );
  NAND2_X1 U18339 ( .A1(n15028), .A2(n15027), .ZN(n15167) );
  NOR2_X1 U18340 ( .A1(n15173), .A2(n15169), .ZN(n15030) );
  XNOR2_X1 U18341 ( .A(n15030), .B(n15029), .ZN(n15156) );
  NAND2_X1 U18342 ( .A1(n15156), .A2(n16102), .ZN(n15035) );
  OAI21_X1 U18343 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n9678), .A(
        n15031), .ZN(n15933) );
  OAI22_X1 U18344 ( .A1(n19611), .A2(n19016), .B1(n18992), .B2(n15933), .ZN(
        n15033) );
  OAI22_X1 U18345 ( .A1(n15980), .A2(n16117), .B1(n9904), .B2(n16121), .ZN(
        n15032) );
  NOR2_X1 U18346 ( .A1(n15033), .A2(n15032), .ZN(n15034) );
  OAI211_X1 U18347 ( .C1(n18984), .C2(n15167), .A(n15035), .B(n15034), .ZN(
        P2_U2988) );
  XNOR2_X1 U18348 ( .A(n15037), .B(n15192), .ZN(n15038) );
  XNOR2_X1 U18349 ( .A(n15036), .B(n15038), .ZN(n15185) );
  NOR2_X1 U18350 ( .A1(n16041), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15040) );
  OR2_X1 U18351 ( .A1(n15039), .A2(n15040), .ZN(n15196) );
  AOI22_X1 U18352 ( .A1(n16009), .A2(n18988), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18979), .ZN(n15045) );
  OAI21_X1 U18353 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n15041), .A(
        n15042), .ZN(n15934) );
  OAI22_X1 U18354 ( .A1(n19607), .A2(n19016), .B1(n18992), .B2(n15934), .ZN(
        n15043) );
  INV_X1 U18355 ( .A(n15043), .ZN(n15044) );
  OAI211_X1 U18356 ( .C1(n15196), .C2(n18984), .A(n15045), .B(n15044), .ZN(
        n15046) );
  AOI21_X1 U18357 ( .B1(n15185), .B2(n16102), .A(n15046), .ZN(n15047) );
  INV_X1 U18358 ( .A(n15047), .ZN(P2_U2990) );
  INV_X1 U18359 ( .A(n15048), .ZN(n15343) );
  INV_X1 U18360 ( .A(n15322), .ZN(n15049) );
  NOR2_X1 U18361 ( .A1(n15344), .A2(n15049), .ZN(n15050) );
  OAI211_X1 U18362 ( .C1(n15052), .C2(n15343), .A(n15051), .B(n15050), .ZN(
        n15053) );
  NAND2_X1 U18363 ( .A1(n15053), .A2(n15323), .ZN(n15307) );
  INV_X1 U18364 ( .A(n15305), .ZN(n15054) );
  OAI21_X1 U18365 ( .B1(n15307), .B2(n15054), .A(n15304), .ZN(n15290) );
  INV_X1 U18366 ( .A(n15288), .ZN(n15055) );
  OAI21_X1 U18367 ( .B1(n15290), .B2(n15055), .A(n15287), .ZN(n15130) );
  INV_X1 U18368 ( .A(n15129), .ZN(n15057) );
  OAI21_X1 U18369 ( .B1(n15130), .B2(n15057), .A(n15056), .ZN(n15115) );
  NAND2_X1 U18370 ( .A1(n15059), .A2(n15058), .ZN(n15116) );
  NOR2_X1 U18371 ( .A1(n15115), .A2(n15116), .ZN(n15114) );
  INV_X1 U18372 ( .A(n15059), .ZN(n15060) );
  NOR2_X1 U18373 ( .A1(n15114), .A2(n15060), .ZN(n15106) );
  INV_X1 U18374 ( .A(n15103), .ZN(n15061) );
  NOR2_X1 U18375 ( .A1(n15106), .A2(n15061), .ZN(n15092) );
  NAND2_X1 U18376 ( .A1(n15092), .A2(n15090), .ZN(n15076) );
  INV_X1 U18377 ( .A(n15078), .ZN(n15062) );
  AOI21_X1 U18378 ( .B1(n15076), .B2(n15063), .A(n15062), .ZN(n15067) );
  NAND2_X1 U18379 ( .A1(n15065), .A2(n15064), .ZN(n15066) );
  XNOR2_X1 U18380 ( .A(n15067), .B(n15066), .ZN(n15221) );
  INV_X1 U18381 ( .A(n15198), .ZN(n16040) );
  AOI21_X1 U18382 ( .B1(n15068), .B2(n15085), .A(n16040), .ZN(n15218) );
  NAND2_X1 U18383 ( .A1(n18980), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15212) );
  OAI21_X1 U18384 ( .B1(n16121), .B2(n15069), .A(n15212), .ZN(n15070) );
  AOI21_X1 U18385 ( .B1(n16107), .B2(n15071), .A(n15070), .ZN(n15072) );
  OAI21_X1 U18386 ( .B1(n15213), .B2(n16117), .A(n15072), .ZN(n15073) );
  AOI21_X1 U18387 ( .B1(n15218), .B2(n16114), .A(n15073), .ZN(n15074) );
  OAI21_X1 U18388 ( .B1(n15221), .B2(n18982), .A(n15074), .ZN(P2_U2993) );
  NAND2_X1 U18389 ( .A1(n15076), .A2(n15075), .ZN(n15080) );
  NAND2_X1 U18390 ( .A1(n15078), .A2(n15077), .ZN(n15079) );
  XNOR2_X1 U18391 ( .A(n15080), .B(n15079), .ZN(n15233) );
  INV_X1 U18392 ( .A(n15081), .ZN(n18653) );
  NOR2_X1 U18393 ( .A1(n19016), .A2(n19601), .ZN(n15226) );
  AOI21_X1 U18394 ( .B1(n18979), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15226), .ZN(n15082) );
  OAI21_X1 U18395 ( .B1(n18992), .B2(n15083), .A(n15082), .ZN(n15087) );
  INV_X1 U18396 ( .A(n15269), .ZN(n16140) );
  NOR2_X2 U18397 ( .A1(n15339), .A2(n15332), .ZN(n15340) );
  OAI21_X1 U18398 ( .B1(n15095), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15085), .ZN(n15229) );
  NOR2_X1 U18399 ( .A1(n15229), .A2(n18984), .ZN(n15086) );
  AOI211_X1 U18400 ( .C1(n18988), .C2(n18653), .A(n15087), .B(n15086), .ZN(
        n15088) );
  NAND2_X1 U18401 ( .A1(n15090), .A2(n15089), .ZN(n15094) );
  INV_X1 U18402 ( .A(n15104), .ZN(n15091) );
  NOR2_X1 U18403 ( .A1(n15092), .A2(n15091), .ZN(n15093) );
  XOR2_X1 U18404 ( .A(n15094), .B(n15093), .Z(n15244) );
  AOI21_X1 U18405 ( .B1(n15096), .B2(n15108), .A(n15095), .ZN(n15242) );
  OAI22_X1 U18406 ( .A1(n16121), .A2(n15098), .B1(n19016), .B2(n15097), .ZN(
        n15099) );
  AOI21_X1 U18407 ( .B1(n18657), .B2(n16107), .A(n15099), .ZN(n15100) );
  OAI21_X1 U18408 ( .B1(n15235), .B2(n16117), .A(n15100), .ZN(n15101) );
  AOI21_X1 U18409 ( .B1(n15242), .B2(n16114), .A(n15101), .ZN(n15102) );
  OAI21_X1 U18410 ( .B1(n15244), .B2(n18982), .A(n15102), .ZN(P2_U2995) );
  NAND2_X1 U18411 ( .A1(n15104), .A2(n15103), .ZN(n15105) );
  XNOR2_X1 U18412 ( .A(n15106), .B(n15105), .ZN(n15245) );
  NAND2_X1 U18413 ( .A1(n15122), .A2(n15247), .ZN(n15107) );
  NAND2_X1 U18414 ( .A1(n15108), .A2(n15107), .ZN(n15257) );
  AOI22_X1 U18415 ( .A1(n18673), .A2(n18988), .B1(n18979), .B2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15111) );
  OAI22_X1 U18416 ( .A1(n19598), .A2(n19016), .B1(n18992), .B2(n18671), .ZN(
        n15109) );
  INV_X1 U18417 ( .A(n15109), .ZN(n15110) );
  OAI211_X1 U18418 ( .C1(n15257), .C2(n18984), .A(n15111), .B(n15110), .ZN(
        n15112) );
  AOI21_X1 U18419 ( .B1(n15245), .B2(n16102), .A(n15112), .ZN(n15113) );
  INV_X1 U18420 ( .A(n15113), .ZN(P2_U2996) );
  AOI21_X1 U18421 ( .B1(n15116), .B2(n15115), .A(n15114), .ZN(n15264) );
  INV_X1 U18422 ( .A(n18688), .ZN(n15121) );
  OAI22_X1 U18423 ( .A1(n16121), .A2(n15117), .B1(n10984), .B2(n19016), .ZN(
        n15120) );
  INV_X1 U18424 ( .A(n15118), .ZN(n18684) );
  NOR2_X1 U18425 ( .A1(n18684), .A2(n18992), .ZN(n15119) );
  AOI211_X1 U18426 ( .C1(n15121), .C2(n18988), .A(n15120), .B(n15119), .ZN(
        n15125) );
  NAND2_X1 U18427 ( .A1(n15268), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15259) );
  INV_X1 U18428 ( .A(n15259), .ZN(n15123) );
  OAI211_X1 U18429 ( .C1(n15123), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16114), .B(n15122), .ZN(n15124) );
  OAI211_X1 U18430 ( .C1(n15264), .C2(n18982), .A(n15125), .B(n15124), .ZN(
        P2_U2997) );
  XNOR2_X1 U18431 ( .A(n15268), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15133) );
  INV_X1 U18432 ( .A(n18695), .ZN(n15128) );
  INV_X1 U18433 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18701) );
  NAND2_X1 U18434 ( .A1(n18980), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15279) );
  OAI21_X1 U18435 ( .B1(n16121), .B2(n18701), .A(n15279), .ZN(n15127) );
  NOR2_X1 U18436 ( .A1(n18694), .A2(n18992), .ZN(n15126) );
  AOI211_X1 U18437 ( .C1(n15128), .C2(n18988), .A(n15127), .B(n15126), .ZN(
        n15132) );
  XNOR2_X1 U18438 ( .A(n15130), .B(n15129), .ZN(n15282) );
  NAND2_X1 U18439 ( .A1(n15282), .A2(n16102), .ZN(n15131) );
  OAI211_X1 U18440 ( .C1(n15133), .C2(n18984), .A(n15132), .B(n15131), .ZN(
        P2_U2998) );
  INV_X1 U18441 ( .A(n14315), .ZN(n15141) );
  NAND2_X1 U18442 ( .A1(n15134), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15140) );
  NOR2_X1 U18443 ( .A1(n15135), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15137) );
  OAI211_X1 U18444 ( .C1(n15141), .C2(n16158), .A(n15140), .B(n15139), .ZN(
        n15142) );
  AOI21_X1 U18445 ( .B1(n15143), .B2(n16154), .A(n15142), .ZN(n15144) );
  OAI21_X1 U18446 ( .B1(n15145), .B2(n16152), .A(n15144), .ZN(P2_U3016) );
  INV_X1 U18447 ( .A(n15146), .ZN(n15951) );
  NAND3_X1 U18448 ( .A1(n15149), .A2(n15148), .A3(n15147), .ZN(n15150) );
  OAI211_X1 U18449 ( .C1(n18995), .C2(n15152), .A(n15151), .B(n15150), .ZN(
        n15153) );
  NAND2_X1 U18450 ( .A1(n15156), .A2(n18999), .ZN(n15166) );
  INV_X1 U18451 ( .A(n15186), .ZN(n15157) );
  AOI21_X1 U18452 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15157), .A(
        n15365), .ZN(n15179) );
  AOI211_X1 U18453 ( .C1(n15159), .C2(n9814), .A(n15158), .B(n15176), .ZN(
        n15161) );
  NOR2_X1 U18454 ( .A1(n19016), .A2(n19611), .ZN(n15160) );
  AOI211_X1 U18455 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n15179), .A(
        n15161), .B(n15160), .ZN(n15162) );
  OAI21_X1 U18456 ( .B1(n15980), .B2(n16158), .A(n15162), .ZN(n15163) );
  AOI21_X1 U18457 ( .B1(n16150), .B2(n15164), .A(n15163), .ZN(n15165) );
  OAI211_X1 U18458 ( .C1(n15167), .C2(n18994), .A(n15166), .B(n15165), .ZN(
        P2_U3020) );
  INV_X1 U18459 ( .A(n15169), .ZN(n15172) );
  OR2_X1 U18460 ( .A1(n15169), .A2(n15168), .ZN(n15170) );
  AOI22_X1 U18461 ( .A1(n15173), .A2(n15172), .B1(n15171), .B2(n15170), .ZN(
        n16032) );
  INV_X1 U18462 ( .A(n16032), .ZN(n15184) );
  NOR2_X1 U18463 ( .A1(n15039), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15174) );
  NOR2_X1 U18464 ( .A1(n15175), .A2(n15174), .ZN(n16031) );
  NOR2_X1 U18465 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15176), .ZN(
        n15178) );
  INV_X1 U18466 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19609) );
  NOR2_X1 U18467 ( .A1(n19609), .A2(n19016), .ZN(n15177) );
  AOI211_X1 U18468 ( .C1(n15179), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15178), .B(n15177), .ZN(n15181) );
  INV_X1 U18469 ( .A(n15999), .ZN(n16030) );
  NAND2_X1 U18470 ( .A1(n19004), .A2(n16030), .ZN(n15180) );
  OAI211_X1 U18471 ( .C1(n18995), .C2(n15993), .A(n15181), .B(n15180), .ZN(
        n15182) );
  AOI21_X1 U18472 ( .B1(n16031), .B2(n16154), .A(n15182), .ZN(n15183) );
  OAI21_X1 U18473 ( .B1(n15184), .B2(n16152), .A(n15183), .ZN(P2_U3021) );
  NAND2_X1 U18474 ( .A1(n15185), .A2(n18999), .ZN(n15195) );
  INV_X1 U18475 ( .A(n16009), .ZN(n15190) );
  NAND2_X1 U18476 ( .A1(n15186), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15189) );
  AOI22_X1 U18477 ( .A1(n16150), .A2(n15187), .B1(n18980), .B2(
        P2_REIP_REG_24__SCAN_IN), .ZN(n15188) );
  OAI211_X1 U18478 ( .C1(n15190), .C2(n16158), .A(n15189), .B(n15188), .ZN(
        n15191) );
  AOI21_X1 U18479 ( .B1(n15193), .B2(n15192), .A(n15191), .ZN(n15194) );
  OAI211_X1 U18480 ( .C1(n15196), .C2(n18994), .A(n15195), .B(n15194), .ZN(
        P2_U3022) );
  XNOR2_X1 U18481 ( .A(n15198), .B(n15197), .ZN(n16045) );
  NAND2_X1 U18482 ( .A1(n15200), .A2(n15199), .ZN(n15202) );
  XOR2_X1 U18483 ( .A(n15202), .B(n15201), .Z(n16046) );
  NOR2_X1 U18484 ( .A1(n19604), .A2(n19016), .ZN(n15203) );
  AOI221_X1 U18485 ( .B1(n16124), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), 
        .C1(n16129), .C2(n15197), .A(n15203), .ZN(n15206) );
  AOI22_X1 U18486 ( .A1(n16048), .A2(n19004), .B1(n16150), .B2(n15204), .ZN(
        n15205) );
  OAI211_X1 U18487 ( .C1(n16046), .C2(n16152), .A(n15206), .B(n15205), .ZN(
        n15207) );
  INV_X1 U18488 ( .A(n15207), .ZN(n15208) );
  OAI21_X1 U18489 ( .B1(n18994), .B2(n16045), .A(n15208), .ZN(P2_U3024) );
  OAI21_X1 U18490 ( .B1(n15209), .B2(n15400), .A(n15366), .ZN(n15217) );
  NAND2_X1 U18491 ( .A1(n16150), .A2(n15210), .ZN(n15211) );
  OAI211_X1 U18492 ( .C1(n15213), .C2(n16158), .A(n15212), .B(n15211), .ZN(
        n15216) );
  NOR3_X1 U18493 ( .A1(n15385), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15214), .ZN(n15215) );
  AOI211_X1 U18494 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15217), .A(
        n15216), .B(n15215), .ZN(n15220) );
  NAND2_X1 U18495 ( .A1(n15218), .A2(n16154), .ZN(n15219) );
  OAI211_X1 U18496 ( .C1(n15221), .C2(n16152), .A(n15220), .B(n15219), .ZN(
        P2_U3025) );
  AND2_X1 U18497 ( .A1(n15366), .A2(n15222), .ZN(n15246) );
  NOR2_X1 U18498 ( .A1(n15223), .A2(n15385), .ZN(n15224) );
  NAND2_X1 U18499 ( .A1(n15224), .A2(n15247), .ZN(n15248) );
  OAI21_X1 U18500 ( .B1(n15365), .B2(n15246), .A(n15248), .ZN(n15234) );
  NAND2_X1 U18501 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15224), .ZN(
        n15240) );
  XNOR2_X1 U18502 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15228) );
  NOR2_X1 U18503 ( .A1(n18995), .A2(n18650), .ZN(n15225) );
  AOI211_X1 U18504 ( .C1(n18653), .C2(n19004), .A(n15226), .B(n15225), .ZN(
        n15227) );
  OAI21_X1 U18505 ( .B1(n15240), .B2(n15228), .A(n15227), .ZN(n15231) );
  NOR2_X1 U18506 ( .A1(n15229), .A2(n18994), .ZN(n15230) );
  AOI211_X1 U18507 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15234), .A(
        n15231), .B(n15230), .ZN(n15232) );
  OAI21_X1 U18508 ( .B1(n15233), .B2(n16152), .A(n15232), .ZN(P2_U3026) );
  NAND2_X1 U18509 ( .A1(n15234), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15239) );
  INV_X1 U18510 ( .A(n15235), .ZN(n18663) );
  NOR2_X1 U18511 ( .A1(n18995), .A2(n18665), .ZN(n15237) );
  NOR2_X1 U18512 ( .A1(n15097), .A2(n19016), .ZN(n15236) );
  AOI211_X1 U18513 ( .C1(n18663), .C2(n19004), .A(n15237), .B(n15236), .ZN(
        n15238) );
  OAI211_X1 U18514 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15240), .A(
        n15239), .B(n15238), .ZN(n15241) );
  AOI21_X1 U18515 ( .B1(n15242), .B2(n16154), .A(n15241), .ZN(n15243) );
  OAI21_X1 U18516 ( .B1(n15244), .B2(n16152), .A(n15243), .ZN(P2_U3027) );
  NAND2_X1 U18517 ( .A1(n15245), .A2(n18999), .ZN(n15256) );
  INV_X1 U18518 ( .A(n15246), .ZN(n15254) );
  NOR2_X1 U18519 ( .A1(n15365), .A2(n15247), .ZN(n15253) );
  NAND2_X1 U18520 ( .A1(n18673), .A2(n19004), .ZN(n15251) );
  INV_X1 U18521 ( .A(n15248), .ZN(n15249) );
  AOI21_X1 U18522 ( .B1(n18980), .B2(P2_REIP_REG_18__SCAN_IN), .A(n15249), 
        .ZN(n15250) );
  OAI211_X1 U18523 ( .C1(n18995), .C2(n18676), .A(n15251), .B(n15250), .ZN(
        n15252) );
  AOI21_X1 U18524 ( .B1(n15254), .B2(n15253), .A(n15252), .ZN(n15255) );
  OAI211_X1 U18525 ( .C1(n15257), .C2(n18994), .A(n15256), .B(n15255), .ZN(
        P2_U3028) );
  INV_X1 U18526 ( .A(n15258), .ZN(n19000) );
  OAI21_X1 U18527 ( .B1(n16154), .B2(n19000), .A(n15259), .ZN(n15262) );
  INV_X1 U18528 ( .A(n15260), .ZN(n15261) );
  INV_X1 U18529 ( .A(n15366), .ZN(n15388) );
  AOI21_X1 U18530 ( .B1(n15261), .B2(n15263), .A(n15388), .ZN(n15299) );
  OAI211_X1 U18531 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n19006), .A(
        n15262), .B(n15299), .ZN(n15278) );
  AOI21_X1 U18532 ( .B1(n20764), .B2(n15263), .A(n15278), .ZN(n15276) );
  INV_X1 U18533 ( .A(n15264), .ZN(n15267) );
  AOI22_X1 U18534 ( .A1(n16150), .A2(n18681), .B1(n18980), .B2(
        P2_REIP_REG_17__SCAN_IN), .ZN(n15265) );
  OAI21_X1 U18535 ( .B1(n18688), .B2(n16158), .A(n15265), .ZN(n15266) );
  AOI21_X1 U18536 ( .B1(n15267), .B2(n18999), .A(n15266), .ZN(n15274) );
  INV_X1 U18537 ( .A(n15268), .ZN(n15286) );
  OR2_X1 U18538 ( .A1(n15286), .A2(n18994), .ZN(n15272) );
  NOR2_X1 U18539 ( .A1(n15380), .A2(n15385), .ZN(n16141) );
  NAND2_X1 U18540 ( .A1(n15269), .A2(n16141), .ZN(n15330) );
  NOR2_X1 U18541 ( .A1(n15270), .A2(n15330), .ZN(n15291) );
  NAND2_X1 U18542 ( .A1(n15291), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15271) );
  NAND2_X1 U18543 ( .A1(n15272), .A2(n15271), .ZN(n15277) );
  NAND3_X1 U18544 ( .A1(n15277), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15275), .ZN(n15273) );
  OAI211_X1 U18545 ( .C1(n15276), .C2(n15275), .A(n15274), .B(n15273), .ZN(
        P2_U3029) );
  INV_X1 U18546 ( .A(n15277), .ZN(n15285) );
  NAND2_X1 U18547 ( .A1(n15278), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15284) );
  NOR2_X1 U18548 ( .A1(n18695), .A2(n16158), .ZN(n15281) );
  OAI21_X1 U18549 ( .B1(n18995), .B2(n18696), .A(n15279), .ZN(n15280) );
  AOI211_X1 U18550 ( .C1(n15282), .C2(n18999), .A(n15281), .B(n15280), .ZN(
        n15283) );
  OAI211_X1 U18551 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15285), .A(
        n15284), .B(n15283), .ZN(P2_U3030) );
  NAND2_X1 U18552 ( .A1(n15288), .A2(n15287), .ZN(n15289) );
  XNOR2_X1 U18553 ( .A(n15290), .B(n15289), .ZN(n16054) );
  NAND2_X1 U18554 ( .A1(n15291), .A2(n15298), .ZN(n15297) );
  INV_X1 U18555 ( .A(n18707), .ZN(n16053) );
  NOR2_X1 U18556 ( .A1(n11091), .A2(n19016), .ZN(n15295) );
  XNOR2_X1 U18557 ( .A(n15293), .B(n15292), .ZN(n18871) );
  NOR2_X1 U18558 ( .A1(n18995), .A2(n18871), .ZN(n15294) );
  AOI211_X1 U18559 ( .C1(n16053), .C2(n19004), .A(n15295), .B(n15294), .ZN(
        n15296) );
  OAI211_X1 U18560 ( .C1(n15299), .C2(n15298), .A(n15297), .B(n15296), .ZN(
        n15300) );
  AOI21_X1 U18561 ( .B1(n16054), .B2(n18999), .A(n15300), .ZN(n15301) );
  OAI21_X1 U18562 ( .B1(n16052), .B2(n18994), .A(n15301), .ZN(P2_U3031) );
  INV_X1 U18563 ( .A(n15302), .ZN(n15303) );
  OAI21_X1 U18564 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15327), .A(
        n15303), .ZN(n16058) );
  NAND2_X1 U18565 ( .A1(n15305), .A2(n15304), .ZN(n15306) );
  XNOR2_X1 U18566 ( .A(n15307), .B(n15306), .ZN(n16057) );
  NOR3_X1 U18567 ( .A1(n15332), .A2(n15333), .A3(n15330), .ZN(n15312) );
  NOR2_X1 U18568 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15330), .ZN(
        n15347) );
  NOR2_X1 U18569 ( .A1(n15380), .A2(n16140), .ZN(n15308) );
  OAI21_X1 U18570 ( .B1(n15308), .B2(n15400), .A(n15366), .ZN(n15348) );
  NOR2_X1 U18571 ( .A1(n15347), .A2(n15348), .ZN(n15334) );
  OAI21_X1 U18572 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15330), .A(
        n15334), .ZN(n15310) );
  NOR2_X1 U18573 ( .A1(n10962), .A2(n19016), .ZN(n15309) );
  AOI221_X1 U18574 ( .B1(n15312), .B2(n15311), .C1(n15310), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n15309), .ZN(n15319) );
  INV_X1 U18575 ( .A(n15313), .ZN(n18719) );
  OR2_X1 U18576 ( .A1(n15315), .A2(n15314), .ZN(n15316) );
  NAND2_X1 U18577 ( .A1(n15316), .A2(n15292), .ZN(n18873) );
  INV_X1 U18578 ( .A(n18873), .ZN(n15317) );
  AOI22_X1 U18579 ( .A1(n19004), .A2(n18719), .B1(n16150), .B2(n15317), .ZN(
        n15318) );
  OAI211_X1 U18580 ( .C1(n16057), .C2(n16152), .A(n15319), .B(n15318), .ZN(
        n15320) );
  INV_X1 U18581 ( .A(n15320), .ZN(n15321) );
  OAI21_X1 U18582 ( .B1(n16058), .B2(n18994), .A(n15321), .ZN(P2_U3032) );
  NAND2_X1 U18583 ( .A1(n15323), .A2(n15322), .ZN(n15324) );
  XNOR2_X1 U18584 ( .A(n15325), .B(n15324), .ZN(n16063) );
  NOR2_X1 U18585 ( .A1(n15340), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15326) );
  NAND2_X1 U18586 ( .A1(n9626), .A2(n16154), .ZN(n15338) );
  AOI21_X1 U18587 ( .B1(n15328), .B2(n15351), .A(n15314), .ZN(n18876) );
  INV_X1 U18588 ( .A(n18876), .ZN(n15329) );
  OAI22_X1 U18589 ( .A1(n18995), .A2(n15329), .B1(n10936), .B2(n19016), .ZN(
        n15336) );
  OR2_X1 U18590 ( .A1(n15330), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15331) );
  OAI22_X1 U18591 ( .A1(n15334), .A2(n15333), .B1(n15332), .B2(n15331), .ZN(
        n15335) );
  AOI211_X1 U18592 ( .C1(n18728), .C2(n19004), .A(n15336), .B(n15335), .ZN(
        n15337) );
  OAI211_X1 U18593 ( .C1(n16063), .C2(n16152), .A(n15338), .B(n15337), .ZN(
        P2_U3033) );
  INV_X1 U18594 ( .A(n15339), .ZN(n16078) );
  INV_X1 U18595 ( .A(n15340), .ZN(n15341) );
  OAI21_X1 U18596 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16078), .A(
        n15341), .ZN(n16069) );
  NOR2_X1 U18597 ( .A1(n15344), .A2(n15343), .ZN(n15345) );
  XNOR2_X1 U18598 ( .A(n15342), .B(n15345), .ZN(n16068) );
  NOR2_X1 U18599 ( .A1(n10932), .A2(n19016), .ZN(n15346) );
  AOI211_X1 U18600 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15348), .A(
        n15347), .B(n15346), .ZN(n15355) );
  OR2_X1 U18601 ( .A1(n15350), .A2(n15349), .ZN(n15352) );
  NAND2_X1 U18602 ( .A1(n15352), .A2(n15351), .ZN(n18879) );
  INV_X1 U18603 ( .A(n18879), .ZN(n15353) );
  AOI22_X1 U18604 ( .A1(n19004), .A2(n18739), .B1(n16150), .B2(n15353), .ZN(
        n15354) );
  OAI211_X1 U18605 ( .C1(n16068), .C2(n16152), .A(n15355), .B(n15354), .ZN(
        n15356) );
  INV_X1 U18606 ( .A(n15356), .ZN(n15357) );
  OAI21_X1 U18607 ( .B1(n16069), .B2(n18994), .A(n15357), .ZN(P2_U3034) );
  INV_X1 U18608 ( .A(n15358), .ZN(n15379) );
  NAND2_X1 U18609 ( .A1(n15379), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16079) );
  OAI21_X1 U18610 ( .B1(n15379), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16079), .ZN(n16083) );
  OR2_X1 U18611 ( .A1(n15359), .A2(n15391), .ZN(n15364) );
  INV_X1 U18612 ( .A(n15360), .ZN(n15361) );
  AND2_X1 U18613 ( .A1(n15362), .A2(n15361), .ZN(n15363) );
  XNOR2_X1 U18614 ( .A(n15364), .B(n15363), .ZN(n16082) );
  AOI21_X1 U18615 ( .B1(n15366), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15365), .ZN(n16136) );
  NOR2_X1 U18616 ( .A1(n10905), .A2(n19016), .ZN(n15367) );
  AOI221_X1 U18617 ( .B1(n16136), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n16141), .C2(n15368), .A(n15367), .ZN(n15375) );
  OR2_X1 U18618 ( .A1(n15371), .A2(n15370), .ZN(n15372) );
  NAND2_X1 U18619 ( .A1(n15372), .A2(n16134), .ZN(n18884) );
  INV_X1 U18620 ( .A(n18884), .ZN(n15373) );
  AOI22_X1 U18621 ( .A1(n19004), .A2(n18764), .B1(n16150), .B2(n15373), .ZN(
        n15374) );
  OAI211_X1 U18622 ( .C1(n16082), .C2(n16152), .A(n15375), .B(n15374), .ZN(
        n15376) );
  INV_X1 U18623 ( .A(n15376), .ZN(n15377) );
  OAI21_X1 U18624 ( .B1(n16083), .B2(n18994), .A(n15377), .ZN(P2_U3036) );
  INV_X1 U18625 ( .A(n15378), .ZN(n15381) );
  AOI21_X1 U18626 ( .B1(n15381), .B2(n15380), .A(n15379), .ZN(n16091) );
  INV_X1 U18627 ( .A(n16091), .ZN(n15395) );
  AOI21_X1 U18628 ( .B1(n15382), .B2(n13323), .A(n15370), .ZN(n18885) );
  NAND2_X1 U18629 ( .A1(n16150), .A2(n18885), .ZN(n15384) );
  NAND2_X1 U18630 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18980), .ZN(n15383) );
  OAI211_X1 U18631 ( .C1(n18776), .C2(n16158), .A(n15384), .B(n15383), .ZN(
        n15387) );
  NOR2_X1 U18632 ( .A1(n15385), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15386) );
  AOI211_X1 U18633 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15388), .A(
        n15387), .B(n15386), .ZN(n15394) );
  INV_X1 U18634 ( .A(n15391), .ZN(n15389) );
  NAND2_X1 U18635 ( .A1(n15359), .A2(n15389), .ZN(n16088) );
  OAI21_X1 U18636 ( .B1(n15392), .B2(n15391), .A(n15390), .ZN(n16087) );
  NAND3_X1 U18637 ( .A1(n16088), .A2(n18999), .A3(n16087), .ZN(n15393) );
  OAI211_X1 U18638 ( .C1(n15395), .C2(n18994), .A(n15394), .B(n15393), .ZN(
        P2_U3037) );
  NOR2_X1 U18639 ( .A1(n16152), .A2(n15396), .ZN(n15397) );
  AOI211_X1 U18640 ( .C1(n19004), .C2(n12340), .A(n15398), .B(n15397), .ZN(
        n15403) );
  AOI22_X1 U18641 ( .A1(n16154), .A2(n15399), .B1(n16150), .B2(n18924), .ZN(
        n15402) );
  MUX2_X1 U18642 ( .A(n15400), .B(n19001), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n15401) );
  NAND3_X1 U18643 ( .A1(n15403), .A2(n15402), .A3(n15401), .ZN(P2_U3046) );
  NAND2_X1 U18644 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15404), .ZN(n15407) );
  NAND2_X1 U18645 ( .A1(n15405), .A2(n19634), .ZN(n15406) );
  OAI211_X1 U18646 ( .C1(n12414), .C2(n15413), .A(n15407), .B(n15406), .ZN(
        n15408) );
  MUX2_X1 U18647 ( .A(n15408), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15414), .Z(P2_U3601) );
  INV_X1 U18648 ( .A(n15409), .ZN(n15412) );
  OAI222_X1 U18649 ( .A1(n15413), .A2(n19654), .B1(n15412), .B2(n15411), .C1(
        n15526), .C2(n15410), .ZN(n15415) );
  INV_X1 U18650 ( .A(n15414), .ZN(n15532) );
  MUX2_X1 U18651 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15415), .S(
        n15532), .Z(P2_U3600) );
  INV_X1 U18652 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16727) );
  INV_X1 U18653 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16724) );
  INV_X1 U18654 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16678) );
  INV_X1 U18655 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16771) );
  NOR3_X1 U18656 ( .A1(n15416), .A2(n17991), .A3(n17976), .ZN(n15418) );
  INV_X1 U18657 ( .A(n18591), .ZN(n15520) );
  NAND3_X1 U18658 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .ZN(n16907) );
  NOR3_X1 U18659 ( .A1(n16906), .A2(n16595), .A3(n16907), .ZN(n16856) );
  NAND4_X1 U18660 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(P3_EBX_REG_2__SCAN_IN), .ZN(n16973) );
  NOR2_X1 U18661 ( .A1(n16616), .A2(n16973), .ZN(n15420) );
  NAND4_X1 U18662 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .A3(n16856), .A4(n15420), .ZN(n16874) );
  NAND3_X1 U18663 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n16858) );
  NOR3_X1 U18664 ( .A1(n16857), .A2(n16874), .A3(n16858), .ZN(n16839) );
  NAND2_X1 U18665 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16839), .ZN(n16824) );
  NOR2_X1 U18666 ( .A1(n16825), .A2(n16824), .ZN(n16811) );
  NAND2_X1 U18667 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16811), .ZN(n16810) );
  NAND2_X1 U18668 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16797), .ZN(n16796) );
  NOR2_X1 U18669 ( .A1(n17991), .A2(n16796), .ZN(n16783) );
  NAND2_X1 U18670 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16783), .ZN(n16772) );
  NAND2_X1 U18671 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16744), .ZN(n16738) );
  NAND2_X1 U18672 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16743), .ZN(n16728) );
  NOR3_X1 U18673 ( .A1(n16727), .A2(n16724), .A3(n16728), .ZN(n16716) );
  NAND2_X1 U18674 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16716), .ZN(n15496) );
  AND2_X1 U18675 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16715) );
  NAND2_X1 U18676 ( .A1(n17144), .A2(n16995), .ZN(n16990) );
  INV_X1 U18677 ( .A(n16716), .ZN(n16721) );
  NAND2_X1 U18678 ( .A1(n16984), .A2(n16721), .ZN(n16726) );
  OAI21_X1 U18679 ( .B1(n16715), .B2(n16990), .A(n16726), .ZN(n16713) );
  AOI22_X1 U18680 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15424) );
  AOI22_X1 U18681 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15423) );
  AOI22_X1 U18682 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U18683 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15421) );
  NAND4_X1 U18684 ( .A1(n15424), .A2(n15423), .A3(n15422), .A4(n15421), .ZN(
        n15430) );
  AOI22_X1 U18685 ( .A1(n11393), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15428) );
  AOI22_X1 U18686 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15427) );
  AOI22_X1 U18687 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15426) );
  AOI22_X1 U18688 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15425) );
  NAND4_X1 U18689 ( .A1(n15428), .A2(n15427), .A3(n15426), .A4(n15425), .ZN(
        n15429) );
  NOR2_X1 U18690 ( .A1(n15430), .A2(n15429), .ZN(n15494) );
  AOI22_X1 U18691 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15434) );
  AOI22_X1 U18692 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15433) );
  AOI22_X1 U18693 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15432) );
  AOI22_X1 U18694 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15431) );
  NAND4_X1 U18695 ( .A1(n15434), .A2(n15433), .A3(n15432), .A4(n15431), .ZN(
        n15440) );
  AOI22_X1 U18696 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15438) );
  AOI22_X1 U18697 ( .A1(n16862), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15437) );
  AOI22_X1 U18698 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15436) );
  AOI22_X1 U18699 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15435) );
  NAND4_X1 U18700 ( .A1(n15438), .A2(n15437), .A3(n15436), .A4(n15435), .ZN(
        n15439) );
  NOR2_X1 U18701 ( .A1(n15440), .A2(n15439), .ZN(n16723) );
  AOI22_X1 U18702 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n16899), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n16953), .ZN(n15444) );
  AOI22_X1 U18703 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n16881), .ZN(n15443) );
  AOI22_X1 U18704 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9574), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n15502), .ZN(n15442) );
  AOI22_X1 U18705 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n16945), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n16926), .ZN(n15441) );
  NAND4_X1 U18706 ( .A1(n15444), .A2(n15443), .A3(n15442), .A4(n15441), .ZN(
        n15450) );
  AOI22_X1 U18707 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U18708 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11393), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n16927), .ZN(n15447) );
  AOI22_X1 U18709 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15446) );
  AOI22_X1 U18710 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n9575), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15445) );
  NAND4_X1 U18711 ( .A1(n15448), .A2(n15447), .A3(n15446), .A4(n15445), .ZN(
        n15449) );
  NOR2_X1 U18712 ( .A1(n15450), .A2(n15449), .ZN(n16734) );
  AOI22_X1 U18713 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15461) );
  AOI22_X1 U18714 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15460) );
  AOI22_X1 U18715 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15451) );
  OAI21_X1 U18716 ( .B1(n16746), .B2(n15452), .A(n15451), .ZN(n15458) );
  AOI22_X1 U18717 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15456) );
  AOI22_X1 U18718 ( .A1(n16862), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15455) );
  AOI22_X1 U18719 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15454) );
  AOI22_X1 U18720 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15453) );
  NAND4_X1 U18721 ( .A1(n15456), .A2(n15455), .A3(n15454), .A4(n15453), .ZN(
        n15457) );
  AOI211_X1 U18722 ( .C1(n16954), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n15458), .B(n15457), .ZN(n15459) );
  NAND3_X1 U18723 ( .A1(n15461), .A2(n15460), .A3(n15459), .ZN(n16740) );
  AOI22_X1 U18724 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U18725 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U18726 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15462) );
  OAI21_X1 U18727 ( .B1(n16864), .B2(n16966), .A(n15462), .ZN(n15468) );
  AOI22_X1 U18728 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U18729 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15465) );
  AOI22_X1 U18730 ( .A1(n11393), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15464) );
  AOI22_X1 U18731 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15463) );
  NAND4_X1 U18732 ( .A1(n15466), .A2(n15465), .A3(n15464), .A4(n15463), .ZN(
        n15467) );
  AOI211_X1 U18733 ( .C1(n16934), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n15468), .B(n15467), .ZN(n15469) );
  NAND3_X1 U18734 ( .A1(n15471), .A2(n15470), .A3(n15469), .ZN(n16741) );
  NAND2_X1 U18735 ( .A1(n16740), .A2(n16741), .ZN(n16739) );
  NOR2_X1 U18736 ( .A1(n16734), .A2(n16739), .ZN(n16733) );
  AOI22_X1 U18737 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15481) );
  AOI22_X1 U18738 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15480) );
  AOI22_X1 U18739 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15472) );
  OAI21_X1 U18740 ( .B1(n16746), .B2(n16985), .A(n15472), .ZN(n15478) );
  AOI22_X1 U18741 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U18742 ( .A1(n16862), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15475) );
  AOI22_X1 U18743 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15474) );
  AOI22_X1 U18744 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15473) );
  NAND4_X1 U18745 ( .A1(n15476), .A2(n15475), .A3(n15474), .A4(n15473), .ZN(
        n15477) );
  AOI211_X1 U18746 ( .C1(n16934), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n15478), .B(n15477), .ZN(n15479) );
  NAND3_X1 U18747 ( .A1(n15481), .A2(n15480), .A3(n15479), .ZN(n16730) );
  NAND2_X1 U18748 ( .A1(n16733), .A2(n16730), .ZN(n16729) );
  NOR2_X1 U18749 ( .A1(n16723), .A2(n16729), .ZN(n16722) );
  AOI22_X1 U18750 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15493) );
  AOI22_X1 U18751 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15492) );
  INV_X1 U18752 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U18753 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15482) );
  OAI21_X1 U18754 ( .B1(n15484), .B2(n15483), .A(n15482), .ZN(n15490) );
  AOI22_X1 U18755 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15488) );
  AOI22_X1 U18756 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15487) );
  AOI22_X1 U18757 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15486) );
  AOI22_X1 U18758 ( .A1(n15502), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15485) );
  NAND4_X1 U18759 ( .A1(n15488), .A2(n15487), .A3(n15486), .A4(n15485), .ZN(
        n15489) );
  AOI211_X1 U18760 ( .C1(n16953), .C2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n15490), .B(n15489), .ZN(n15491) );
  NAND3_X1 U18761 ( .A1(n15493), .A2(n15492), .A3(n15491), .ZN(n16719) );
  NAND2_X1 U18762 ( .A1(n16722), .A2(n16719), .ZN(n16718) );
  NOR2_X1 U18763 ( .A1(n15494), .A2(n16718), .ZN(n16712) );
  AOI21_X1 U18764 ( .B1(n15494), .B2(n16718), .A(n16712), .ZN(n17012) );
  AOI22_X1 U18765 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16713), .B1(n17012), 
        .B2(n16993), .ZN(n15495) );
  OAI21_X1 U18766 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15496), .A(n15495), .ZN(
        P3_U2675) );
  AOI22_X1 U18767 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U18768 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15499) );
  AOI22_X1 U18769 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15498) );
  AOI22_X1 U18770 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15497) );
  NAND4_X1 U18771 ( .A1(n15500), .A2(n15499), .A3(n15498), .A4(n15497), .ZN(
        n15508) );
  AOI22_X1 U18772 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15506) );
  AOI22_X1 U18773 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15505) );
  AOI22_X1 U18774 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U18775 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15503) );
  NAND4_X1 U18776 ( .A1(n15506), .A2(n15505), .A3(n15504), .A4(n15503), .ZN(
        n15507) );
  NOR2_X1 U18777 ( .A1(n15508), .A2(n15507), .ZN(n17089) );
  INV_X1 U18778 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16875) );
  NOR3_X1 U18779 ( .A1(n16875), .A2(n16874), .A3(n16990), .ZN(n15509) );
  NOR2_X1 U18780 ( .A1(n16993), .A2(n15509), .ZN(n16892) );
  AOI22_X1 U18781 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16892), .B1(n15509), 
        .B2(n16876), .ZN(n15510) );
  OAI21_X1 U18782 ( .B1(n17089), .B2(n16984), .A(n15510), .ZN(P3_U2690) );
  NAND2_X1 U18783 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18109) );
  AOI221_X1 U18784 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18109), .C1(n15512), 
        .C2(n18109), .A(n15511), .ZN(n17956) );
  INV_X1 U18785 ( .A(n15513), .ZN(n15514) );
  INV_X1 U18786 ( .A(n18298), .ZN(n18245) );
  NAND2_X1 U18787 ( .A1(n18405), .A2(n18245), .ZN(n18133) );
  OAI211_X1 U18788 ( .C1(n18298), .C2(n15514), .A(n17957), .B(n18133), .ZN(
        n17954) );
  AOI22_X1 U18789 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17956), .B1(
        n17954), .B2(n20820), .ZN(P3_U2865) );
  INV_X1 U18790 ( .A(n15515), .ZN(n15518) );
  INV_X1 U18791 ( .A(n18468), .ZN(n18597) );
  OAI211_X1 U18792 ( .C1(n17152), .C2(n15611), .A(n18430), .B(n18608), .ZN(
        n15517) );
  OAI211_X1 U18793 ( .C1(n15520), .C2(n15519), .A(n15518), .B(n15517), .ZN(
        n18422) );
  INV_X1 U18794 ( .A(n18422), .ZN(n18433) );
  NAND2_X1 U18795 ( .A1(n18603), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17959) );
  INV_X1 U18796 ( .A(n18542), .ZN(n18455) );
  NAND2_X1 U18797 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18455), .ZN(n15521) );
  INV_X1 U18798 ( .A(n18556), .ZN(n18571) );
  AOI21_X1 U18799 ( .B1(n15523), .B2(n15525), .A(n15522), .ZN(n18432) );
  NAND3_X1 U18800 ( .A1(n18573), .A2(n18571), .A3(n18432), .ZN(n15524) );
  OAI21_X1 U18801 ( .B1(n18573), .B2(n15525), .A(n15524), .ZN(P3_U3284) );
  NOR4_X1 U18802 ( .A1(n15528), .A2(n15527), .A3(n9573), .A4(n15526), .ZN(
        n15529) );
  NAND2_X1 U18803 ( .A1(n15532), .A2(n15529), .ZN(n15530) );
  OAI21_X1 U18804 ( .B1(n15532), .B2(n15531), .A(n15530), .ZN(P2_U3595) );
  INV_X1 U18805 ( .A(n17865), .ZN(n15536) );
  OAI21_X1 U18806 ( .B1(n15536), .B2(n16211), .A(n15533), .ZN(n15534) );
  AOI21_X1 U18807 ( .B1(n16189), .B2(n17945), .A(n15534), .ZN(n15599) );
  INV_X1 U18808 ( .A(n15535), .ZN(n16188) );
  OAI22_X1 U18809 ( .A1(n16188), .A2(n15536), .B1(n16190), .B2(n17939), .ZN(
        n15600) );
  INV_X1 U18810 ( .A(n17836), .ZN(n17756) );
  AOI21_X1 U18811 ( .B1(n17756), .B2(n17638), .A(n15537), .ZN(n16214) );
  OAI22_X1 U18812 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17929), .B1(
        n16214), .B2(n9563), .ZN(n15538) );
  NOR3_X1 U18813 ( .A1(n17936), .A2(n15600), .A3(n15538), .ZN(n15542) );
  NOR2_X1 U18814 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17528), .ZN(
        n16205) );
  INV_X1 U18815 ( .A(n16205), .ZN(n15539) );
  OAI221_X1 U18816 ( .B1(n16207), .B2(n9570), .C1(n16207), .C2(n16215), .A(
        n15539), .ZN(n15540) );
  XNOR2_X1 U18817 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n15540), .ZN(
        n16194) );
  AOI22_X1 U18818 ( .A1(n9578), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n17850), 
        .B2(n16194), .ZN(n15541) );
  OAI221_X1 U18819 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15599), 
        .C1(n16191), .C2(n15542), .A(n15541), .ZN(P3_U2833) );
  OAI21_X1 U18820 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n15544), .A(
        n15543), .ZN(n16051) );
  INV_X1 U18821 ( .A(n16051), .ZN(n15546) );
  AOI211_X1 U18822 ( .C1(n15546), .C2(n9914), .A(n15935), .B(n19555), .ZN(
        n15551) );
  AOI22_X1 U18823 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18853), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n18856), .ZN(n15548) );
  NAND2_X1 U18824 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18859), .ZN(
        n15547) );
  OAI211_X1 U18825 ( .C1(n18810), .C2(n15549), .A(n15548), .B(n15547), .ZN(
        n15550) );
  AOI211_X1 U18826 ( .C1(n18854), .C2(n16048), .A(n15551), .B(n15550), .ZN(
        n15552) );
  OAI21_X1 U18827 ( .B1(n15553), .B2(n18842), .A(n15552), .ZN(P2_U2833) );
  NOR2_X1 U18828 ( .A1(n15554), .A2(n15587), .ZN(n15595) );
  INV_X1 U18829 ( .A(n15555), .ZN(n15569) );
  INV_X1 U18830 ( .A(n15556), .ZN(n15557) );
  OAI211_X1 U18831 ( .C1(n15559), .C2(n15558), .A(n15557), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15563) );
  INV_X1 U18832 ( .A(n15560), .ZN(n15562) );
  OAI211_X1 U18833 ( .C1(n15563), .C2(n20507), .A(n15562), .B(n15561), .ZN(
        n15565) );
  NAND2_X1 U18834 ( .A1(n15563), .A2(n20507), .ZN(n15564) );
  NAND2_X1 U18835 ( .A1(n15565), .A2(n15564), .ZN(n15566) );
  AOI222_X1 U18836 ( .A1(n15567), .A2(n20256), .B1(n15567), .B2(n15566), .C1(
        n20256), .C2(n15566), .ZN(n15568) );
  AOI222_X1 U18837 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15569), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15568), .C1(n15569), 
        .C2(n15568), .ZN(n15571) );
  AOI21_X1 U18838 ( .B1(n15571), .B2(n19964), .A(n15570), .ZN(n15581) );
  NOR2_X1 U18839 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15575) );
  INV_X1 U18840 ( .A(n15572), .ZN(n15573) );
  OAI211_X1 U18841 ( .C1(n15576), .C2(n15575), .A(n15574), .B(n15573), .ZN(
        n15577) );
  INV_X1 U18842 ( .A(n15577), .ZN(n15578) );
  AND2_X1 U18843 ( .A1(n15579), .A2(n15578), .ZN(n15580) );
  AND3_X1 U18844 ( .A1(n20055), .A2(n19823), .A3(n15582), .ZN(n15583) );
  AOI221_X1 U18845 ( .B1(n15585), .B2(n15584), .C1(n20666), .C2(n15584), .A(
        n15583), .ZN(n15921) );
  OAI221_X1 U18846 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15586), 
        .A(n15921), .ZN(n15927) );
  NAND2_X1 U18847 ( .A1(n15927), .A2(n20571), .ZN(n15594) );
  INV_X1 U18848 ( .A(n15586), .ZN(n15590) );
  OAI211_X1 U18849 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20666), .A(n15588), 
        .B(n15587), .ZN(n15589) );
  AOI21_X1 U18850 ( .B1(n15591), .B2(n15590), .A(n15589), .ZN(n15592) );
  AND2_X1 U18851 ( .A1(n15927), .A2(n15592), .ZN(n15593) );
  OAI22_X1 U18852 ( .A1(n15595), .A2(n15594), .B1(n15593), .B2(n20571), .ZN(
        P1_U3161) );
  NAND2_X1 U18853 ( .A1(n15597), .A2(n15596), .ZN(n15598) );
  XNOR2_X1 U18854 ( .A(n15598), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16187) );
  NOR2_X1 U18855 ( .A1(n15601), .A2(n15600), .ZN(n15602) );
  MUX2_X1 U18856 ( .A(n10084), .B(n15602), .S(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n15603) );
  NAND2_X1 U18857 ( .A1(n9578), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16179) );
  OAI211_X1 U18858 ( .C1(n16187), .C2(n17870), .A(n15603), .B(n16179), .ZN(
        P3_U2832) );
  INV_X1 U18859 ( .A(HOLD), .ZN(n20581) );
  NAND2_X1 U18860 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20576) );
  OAI21_X1 U18861 ( .B1(n20581), .B2(n19698), .A(n20576), .ZN(n15604) );
  OAI21_X1 U18862 ( .B1(n20581), .B2(n20592), .A(n15604), .ZN(n15606) );
  NOR2_X1 U18863 ( .A1(n19698), .A2(n20666), .ZN(n20584) );
  INV_X1 U18864 ( .A(n20584), .ZN(n20575) );
  NAND3_X1 U18865 ( .A1(n15606), .A2(n15605), .A3(n20575), .ZN(P1_U3195) );
  INV_X1 U18866 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16302) );
  NOR2_X1 U18867 ( .A1(n19801), .A2(n16302), .ZN(P1_U2905) );
  NOR2_X1 U18868 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15607) );
  NOR3_X1 U18869 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12317), .A3(n19685), 
        .ZN(n19553) );
  NOR4_X1 U18870 ( .A1(n15608), .A2(n15607), .A3(n19553), .A4(n15609), .ZN(
        P2_U3178) );
  AOI221_X1 U18871 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15609), .C1(n19670), .C2(
        n15609), .A(n19392), .ZN(n19667) );
  INV_X1 U18872 ( .A(n19667), .ZN(n19664) );
  NOR2_X1 U18873 ( .A1(n15610), .A2(n19664), .ZN(P2_U3047) );
  NAND3_X1 U18874 ( .A1(n15611), .A2(n18430), .A3(n18608), .ZN(n15613) );
  AOI221_X4 U18875 ( .B1(n15614), .B2(n15613), .C1(n15612), .C2(n15613), .A(
        n18450), .ZN(n17000) );
  INV_X1 U18876 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20802) );
  AOI22_X1 U18877 ( .A1(n17147), .A2(BUF2_REG_0__SCAN_IN), .B1(n17146), .B2(
        n15617), .ZN(n15618) );
  OAI221_X1 U18878 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17142), .C1(n20802), 
        .C2(n17000), .A(n15618), .ZN(P3_U2735) );
  AOI22_X1 U18879 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_24__SCAN_IN), .B2(n19774), .ZN(n15619) );
  OAI21_X1 U18880 ( .B1(n15620), .B2(n20625), .A(n15619), .ZN(n15624) );
  NAND2_X1 U18881 ( .A1(n15639), .A2(n20625), .ZN(n15622) );
  OAI22_X1 U18882 ( .A1(n15736), .A2(n19751), .B1(n15622), .B2(n15621), .ZN(
        n15623) );
  NOR2_X1 U18883 ( .A1(n15624), .A2(n15623), .ZN(n15625) );
  OAI21_X1 U18884 ( .B1(n15731), .B2(n15657), .A(n15625), .ZN(n15626) );
  INV_X1 U18885 ( .A(n15626), .ZN(n15627) );
  OAI21_X1 U18886 ( .B1(n19761), .B2(n15628), .A(n15627), .ZN(P1_U2816) );
  OAI22_X1 U18887 ( .A1(n15743), .A2(n19751), .B1(n15713), .B2(n15629), .ZN(
        n15630) );
  AOI21_X1 U18888 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19779), .A(
        n15630), .ZN(n15643) );
  OAI21_X1 U18889 ( .B1(n14401), .B2(n15632), .A(n15631), .ZN(n15634) );
  AND2_X1 U18890 ( .A1(n15634), .A2(n15633), .ZN(n15740) );
  XNOR2_X1 U18891 ( .A(n15636), .B(n15635), .ZN(n15812) );
  AOI22_X1 U18892 ( .A1(n15740), .A2(n19755), .B1(n19773), .B2(n15812), .ZN(
        n15642) );
  OAI21_X1 U18893 ( .B1(n15637), .B2(n15648), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15641) );
  INV_X1 U18894 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20823) );
  NAND3_X1 U18895 ( .A1(n15639), .A2(n15638), .A3(n20823), .ZN(n15640) );
  NAND4_X1 U18896 ( .A1(n15643), .A2(n15642), .A3(n15641), .A4(n15640), .ZN(
        P1_U2818) );
  INV_X1 U18897 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15644) );
  OAI22_X1 U18898 ( .A1(n15644), .A2(n19728), .B1(n15753), .B2(n19751), .ZN(
        n15645) );
  AOI21_X1 U18899 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n19774), .A(n15645), .ZN(
        n15650) );
  NAND2_X1 U18900 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n15646), .ZN(n15671) );
  OAI21_X1 U18901 ( .B1(n15652), .B2(n15671), .A(n20621), .ZN(n15647) );
  AOI22_X1 U18902 ( .A1(n15749), .A2(n19755), .B1(n15648), .B2(n15647), .ZN(
        n15649) );
  OAI211_X1 U18903 ( .C1(n19761), .C2(n15651), .A(n15650), .B(n15649), .ZN(
        P1_U2820) );
  OAI21_X1 U18904 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15652), .ZN(n15662) );
  AOI22_X1 U18905 ( .A1(n15653), .A2(n19778), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n19774), .ZN(n15654) );
  OAI211_X1 U18906 ( .C1(n19728), .C2(n15655), .A(n15654), .B(n19927), .ZN(
        n15656) );
  AOI21_X1 U18907 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n15663), .A(n15656), 
        .ZN(n15661) );
  OAI22_X1 U18908 ( .A1(n15658), .A2(n15657), .B1(n19761), .B2(n15821), .ZN(
        n15659) );
  INV_X1 U18909 ( .A(n15659), .ZN(n15660) );
  OAI211_X1 U18910 ( .C1(n15671), .C2(n15662), .A(n15661), .B(n15660), .ZN(
        P1_U2821) );
  AOI22_X1 U18911 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(n19774), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n15663), .ZN(n15664) );
  OAI21_X1 U18912 ( .B1(n15665), .B2(n19751), .A(n15664), .ZN(n15666) );
  AOI211_X1 U18913 ( .C1(n19779), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19913), .B(n15666), .ZN(n15670) );
  INV_X1 U18914 ( .A(n15829), .ZN(n15667) );
  AOI22_X1 U18915 ( .A1(n15668), .A2(n19755), .B1(n19773), .B2(n15667), .ZN(
        n15669) );
  OAI211_X1 U18916 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15671), .A(n15670), 
        .B(n15669), .ZN(P1_U2822) );
  OAI21_X1 U18917 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15672), .ZN(n15680) );
  NOR2_X1 U18918 ( .A1(n15691), .A2(n14817), .ZN(n15678) );
  AOI22_X1 U18919 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_16__SCAN_IN), .B2(n19774), .ZN(n15675) );
  INV_X1 U18920 ( .A(n15758), .ZN(n15673) );
  AOI21_X1 U18921 ( .B1(n19778), .B2(n15673), .A(n19913), .ZN(n15674) );
  OAI211_X1 U18922 ( .C1(n19761), .C2(n15676), .A(n15675), .B(n15674), .ZN(
        n15677) );
  AOI211_X1 U18923 ( .C1(n15754), .C2(n19755), .A(n15678), .B(n15677), .ZN(
        n15679) );
  OAI21_X1 U18924 ( .B1(n15689), .B2(n15680), .A(n15679), .ZN(P1_U2824) );
  INV_X1 U18925 ( .A(n15681), .ZN(n15843) );
  AOI22_X1 U18926 ( .A1(n15682), .A2(n19778), .B1(n19773), .B2(n15843), .ZN(
        n15688) );
  INV_X1 U18927 ( .A(n15683), .ZN(n15686) );
  AOI22_X1 U18928 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_15__SCAN_IN), .B2(n19774), .ZN(n15684) );
  OAI211_X1 U18929 ( .C1(n15691), .C2(n14689), .A(n15684), .B(n19927), .ZN(
        n15685) );
  AOI21_X1 U18930 ( .B1(n15686), .B2(n19755), .A(n15685), .ZN(n15687) );
  OAI211_X1 U18931 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15689), .A(n15688), 
        .B(n15687), .ZN(P1_U2825) );
  AOI22_X1 U18932 ( .A1(n15759), .A2(n19778), .B1(n19773), .B2(n15714), .ZN(
        n15696) );
  AOI22_X1 U18933 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(n19774), .ZN(n15695) );
  OAI21_X1 U18934 ( .B1(n14702), .B2(n15690), .A(n20612), .ZN(n15693) );
  INV_X1 U18935 ( .A(n15691), .ZN(n15692) );
  AOI22_X1 U18936 ( .A1(n15760), .A2(n19755), .B1(n15693), .B2(n15692), .ZN(
        n15694) );
  NAND4_X1 U18937 ( .A1(n15696), .A2(n15695), .A3(n15694), .A4(n19927), .ZN(
        P1_U2826) );
  NOR2_X1 U18938 ( .A1(n19747), .A2(n15697), .ZN(n15705) );
  AOI21_X1 U18939 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15705), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15704) );
  OAI22_X1 U18940 ( .A1(n15699), .A2(n19728), .B1(n19761), .B2(n15698), .ZN(
        n15700) );
  AOI211_X1 U18941 ( .C1(n19774), .C2(P1_EBX_REG_12__SCAN_IN), .A(n19913), .B(
        n15700), .ZN(n15702) );
  AOI22_X1 U18942 ( .A1(n15765), .A2(n19778), .B1(n19755), .B2(n15764), .ZN(
        n15701) );
  OAI211_X1 U18943 ( .C1(n15704), .C2(n15703), .A(n15702), .B(n15701), .ZN(
        P1_U2828) );
  INV_X1 U18944 ( .A(n15776), .ZN(n15706) );
  INV_X1 U18945 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20609) );
  AOI22_X1 U18946 ( .A1(n15706), .A2(n19778), .B1(n15705), .B2(n20609), .ZN(
        n15711) );
  AOI22_X1 U18947 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_11__SCAN_IN), .B2(n19774), .ZN(n15710) );
  AOI21_X1 U18948 ( .B1(n15859), .B2(n19773), .A(n19913), .ZN(n15709) );
  AOI22_X1 U18949 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15707), .B1(n19755), 
        .B2(n15773), .ZN(n15708) );
  NAND4_X1 U18950 ( .A1(n15711), .A2(n15710), .A3(n15709), .A4(n15708), .ZN(
        P1_U2829) );
  AOI22_X1 U18951 ( .A1(n15740), .A2(n19793), .B1(n19792), .B2(n15812), .ZN(
        n15712) );
  OAI21_X1 U18952 ( .B1(n19797), .B2(n15713), .A(n15712), .ZN(P1_U2850) );
  AOI22_X1 U18953 ( .A1(n15760), .A2(n19793), .B1(n19792), .B2(n15714), .ZN(
        n15715) );
  OAI21_X1 U18954 ( .B1(n19797), .B2(n15716), .A(n15715), .ZN(P1_U2858) );
  OAI22_X1 U18955 ( .A1(n15721), .A2(n20010), .B1(n15730), .B2(n19841), .ZN(
        n15717) );
  INV_X1 U18956 ( .A(n15717), .ZN(n15719) );
  AOI22_X1 U18957 ( .A1(n15740), .A2(n15728), .B1(n15723), .B2(DATAI_22_), 
        .ZN(n15718) );
  OAI211_X1 U18958 ( .C1(n15726), .C2(n14987), .A(n15719), .B(n15718), .ZN(
        P1_U2882) );
  INV_X1 U18959 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16242) );
  INV_X1 U18960 ( .A(n20002), .ZN(n15720) );
  OAI22_X1 U18961 ( .A1(n15721), .A2(n15720), .B1(n15730), .B2(n19837), .ZN(
        n15722) );
  INV_X1 U18962 ( .A(n15722), .ZN(n15725) );
  AOI22_X1 U18963 ( .A1(n15749), .A2(n15728), .B1(n15723), .B2(DATAI_20_), 
        .ZN(n15724) );
  OAI211_X1 U18964 ( .C1(n15726), .C2(n16242), .A(n15725), .B(n15724), .ZN(
        P1_U2884) );
  INV_X1 U18965 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20786) );
  AOI22_X1 U18966 ( .A1(n15764), .A2(n15728), .B1(n19888), .B2(n15727), .ZN(
        n15729) );
  OAI21_X1 U18967 ( .B1(n15730), .B2(n20786), .A(n15729), .ZN(P1_U2892) );
  AOI22_X1 U18968 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n15735) );
  INV_X1 U18969 ( .A(n15731), .ZN(n15732) );
  AOI22_X1 U18970 ( .A1(n15733), .A2(n19917), .B1(n15781), .B2(n15732), .ZN(
        n15734) );
  OAI211_X1 U18971 ( .C1(n19912), .C2(n15736), .A(n15735), .B(n15734), .ZN(
        P1_U2975) );
  AOI22_X1 U18972 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15742) );
  NAND2_X1 U18973 ( .A1(n15738), .A2(n15737), .ZN(n15739) );
  XNOR2_X1 U18974 ( .A(n15739), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15811) );
  AOI22_X1 U18975 ( .A1(n19917), .A2(n15811), .B1(n15740), .B2(n15781), .ZN(
        n15741) );
  OAI211_X1 U18976 ( .C1(n19912), .C2(n15743), .A(n15742), .B(n15741), .ZN(
        P1_U2977) );
  AOI22_X1 U18977 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15747) );
  AOI22_X1 U18978 ( .A1(n15745), .A2(n15781), .B1(n19916), .B2(n15744), .ZN(
        n15746) );
  OAI211_X1 U18979 ( .C1(n19708), .C2(n15748), .A(n15747), .B(n15746), .ZN(
        P1_U2978) );
  AOI22_X1 U18980 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15752) );
  AOI22_X1 U18981 ( .A1(n15750), .A2(n19917), .B1(n15781), .B2(n15749), .ZN(
        n15751) );
  OAI211_X1 U18982 ( .C1(n19912), .C2(n15753), .A(n15752), .B(n15751), .ZN(
        P1_U2979) );
  AOI22_X1 U18983 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15757) );
  AOI22_X1 U18984 ( .A1(n15755), .A2(n19917), .B1(n15781), .B2(n15754), .ZN(
        n15756) );
  OAI211_X1 U18985 ( .C1(n19912), .C2(n15758), .A(n15757), .B(n15756), .ZN(
        P1_U2983) );
  AOI22_X1 U18986 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U18987 ( .A1(n15760), .A2(n15781), .B1(n15759), .B2(n19916), .ZN(
        n15761) );
  OAI211_X1 U18988 ( .C1(n15763), .C2(n19708), .A(n15762), .B(n15761), .ZN(
        P1_U2985) );
  AOI22_X1 U18989 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15767) );
  AOI22_X1 U18990 ( .A1(n19916), .A2(n15765), .B1(n15781), .B2(n15764), .ZN(
        n15766) );
  OAI211_X1 U18991 ( .C1(n15768), .C2(n19708), .A(n15767), .B(n15766), .ZN(
        P1_U2987) );
  AOI22_X1 U18992 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15775) );
  NOR3_X1 U18993 ( .A1(n13481), .A2(n15769), .A3(n12057), .ZN(n15771) );
  NOR2_X1 U18994 ( .A1(n15771), .A2(n15770), .ZN(n15772) );
  XNOR2_X1 U18995 ( .A(n15772), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15862) );
  AOI22_X1 U18996 ( .A1(n19917), .A2(n15862), .B1(n15781), .B2(n15773), .ZN(
        n15774) );
  OAI211_X1 U18997 ( .C1(n19912), .C2(n15776), .A(n15775), .B(n15774), .ZN(
        P1_U2988) );
  AOI22_X1 U18998 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15783) );
  NAND2_X1 U18999 ( .A1(n15779), .A2(n15778), .ZN(n15780) );
  XNOR2_X1 U19000 ( .A(n15777), .B(n15780), .ZN(n15898) );
  AOI22_X1 U19001 ( .A1(n15898), .A2(n19917), .B1(n15781), .B2(n19756), .ZN(
        n15782) );
  OAI211_X1 U19002 ( .C1(n19912), .C2(n19752), .A(n15783), .B(n15782), .ZN(
        P1_U2992) );
  AOI22_X1 U19003 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15790) );
  OR2_X1 U19004 ( .A1(n15785), .A2(n15784), .ZN(n15786) );
  AND2_X1 U19005 ( .A1(n15787), .A2(n15786), .ZN(n15908) );
  AOI22_X1 U19006 ( .A1(n15908), .A2(n19917), .B1(n15781), .B2(n15788), .ZN(
        n15789) );
  OAI211_X1 U19007 ( .C1(n19912), .C2(n15791), .A(n15790), .B(n15789), .ZN(
        P1_U2994) );
  INV_X1 U19008 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15800) );
  NOR4_X1 U19009 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15793), .A3(
        n15808), .A4(n15792), .ZN(n15794) );
  AOI21_X1 U19010 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n19913), .A(n15794), 
        .ZN(n15799) );
  INV_X1 U19011 ( .A(n15795), .ZN(n15797) );
  AOI22_X1 U19012 ( .A1(n15797), .A2(n19952), .B1(n19936), .B2(n15796), .ZN(
        n15798) );
  OAI211_X1 U19013 ( .C1(n15801), .C2(n15800), .A(n15799), .B(n15798), .ZN(
        P1_U3006) );
  AOI22_X1 U19014 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n19913), .B1(n15802), 
        .B2(n15808), .ZN(n15807) );
  INV_X1 U19015 ( .A(n15803), .ZN(n15805) );
  AOI22_X1 U19016 ( .A1(n15805), .A2(n19952), .B1(n19936), .B2(n15804), .ZN(
        n15806) );
  OAI211_X1 U19017 ( .C1(n15809), .C2(n15808), .A(n15807), .B(n15806), .ZN(
        P1_U3008) );
  AOI22_X1 U19018 ( .A1(n15811), .A2(n19952), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15810), .ZN(n15818) );
  NAND2_X1 U19019 ( .A1(n19913), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15817) );
  NAND2_X1 U19020 ( .A1(n15812), .A2(n19936), .ZN(n15816) );
  OAI211_X1 U19021 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15814), .B(n15813), .ZN(
        n15815) );
  NAND4_X1 U19022 ( .A1(n15818), .A2(n15817), .A3(n15816), .A4(n15815), .ZN(
        P1_U3009) );
  AOI22_X1 U19023 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15819), .B1(
        n19913), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15825) );
  INV_X1 U19024 ( .A(n15820), .ZN(n15823) );
  INV_X1 U19025 ( .A(n15821), .ZN(n15822) );
  AOI22_X1 U19026 ( .A1(n15823), .A2(n19952), .B1(n19936), .B2(n15822), .ZN(
        n15824) );
  OAI211_X1 U19027 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15826), .A(
        n15825), .B(n15824), .ZN(P1_U3012) );
  AOI21_X1 U19028 ( .B1(n15889), .B2(n15827), .A(n15850), .ZN(n15841) );
  NOR3_X1 U19029 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15828), .A3(
        n15827), .ZN(n15832) );
  OAI22_X1 U19030 ( .A1(n15830), .A2(n19925), .B1(n19955), .B2(n15829), .ZN(
        n15831) );
  AOI211_X1 U19031 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n19913), .A(n15832), 
        .B(n15831), .ZN(n15833) );
  OAI21_X1 U19032 ( .B1(n15841), .B2(n15834), .A(n15833), .ZN(P1_U3013) );
  AOI21_X1 U19033 ( .B1(n15835), .B2(n15844), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15840) );
  AOI22_X1 U19034 ( .A1(n15837), .A2(n19952), .B1(n19936), .B2(n15836), .ZN(
        n15839) );
  NAND2_X1 U19035 ( .A1(n19913), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15838) );
  OAI211_X1 U19036 ( .C1(n15841), .C2(n15840), .A(n15839), .B(n15838), .ZN(
        P1_U3014) );
  AOI21_X1 U19037 ( .B1(n15843), .B2(n19936), .A(n15842), .ZN(n15847) );
  AOI22_X1 U19038 ( .A1(n15845), .A2(n19952), .B1(n15844), .B2(n15848), .ZN(
        n15846) );
  OAI211_X1 U19039 ( .C1(n15849), .C2(n15848), .A(n15847), .B(n15846), .ZN(
        P1_U3016) );
  INV_X1 U19040 ( .A(n15850), .ZN(n15858) );
  AOI21_X1 U19041 ( .B1(n15852), .B2(n19936), .A(n15851), .ZN(n15856) );
  AOI22_X1 U19042 ( .A1(n15854), .A2(n19952), .B1(n15857), .B2(n15853), .ZN(
        n15855) );
  OAI211_X1 U19043 ( .C1(n15858), .C2(n15857), .A(n15856), .B(n15855), .ZN(
        P1_U3018) );
  AOI22_X1 U19044 ( .A1(n15859), .A2(n19936), .B1(n19913), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15864) );
  NOR2_X1 U19045 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15860), .ZN(
        n15861) );
  AOI22_X1 U19046 ( .A1(n15862), .A2(n19952), .B1(n15861), .B2(n15892), .ZN(
        n15863) );
  OAI211_X1 U19047 ( .C1(n15865), .C2(n11912), .A(n15864), .B(n15863), .ZN(
        P1_U3020) );
  NAND2_X1 U19048 ( .A1(n15870), .A2(n15871), .ZN(n15867) );
  OAI21_X1 U19049 ( .B1(n19923), .B2(n15867), .A(n15866), .ZN(n15887) );
  INV_X1 U19050 ( .A(n15868), .ZN(n15876) );
  INV_X1 U19051 ( .A(n15869), .ZN(n15903) );
  NAND3_X1 U19052 ( .A1(n15871), .A2(n15870), .A3(n15903), .ZN(n15883) );
  AOI221_X1 U19053 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n12057), .C2(n11905), .A(
        n15883), .ZN(n15872) );
  AOI21_X1 U19054 ( .B1(n19913), .B2(P1_REIP_REG_10__SCAN_IN), .A(n15872), 
        .ZN(n15873) );
  OAI21_X1 U19055 ( .B1(n15874), .B2(n19955), .A(n15873), .ZN(n15875) );
  AOI21_X1 U19056 ( .B1(n15876), .B2(n19952), .A(n15875), .ZN(n15877) );
  OAI21_X1 U19057 ( .B1(n12057), .B2(n15887), .A(n15877), .ZN(P1_U3021) );
  INV_X1 U19058 ( .A(n15878), .ZN(n15885) );
  NAND2_X1 U19059 ( .A1(n9751), .A2(n15879), .ZN(n15880) );
  AND2_X1 U19060 ( .A1(n15881), .A2(n15880), .ZN(n19791) );
  AOI22_X1 U19061 ( .A1(n19791), .A2(n19936), .B1(n19913), .B2(
        P1_REIP_REG_9__SCAN_IN), .ZN(n15882) );
  OAI21_X1 U19062 ( .B1(n15883), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15882), .ZN(n15884) );
  AOI21_X1 U19063 ( .B1(n15885), .B2(n19952), .A(n15884), .ZN(n15886) );
  OAI21_X1 U19064 ( .B1(n11905), .B2(n15887), .A(n15886), .ZN(P1_U3022) );
  AOI21_X1 U19065 ( .B1(n15890), .B2(n15889), .A(n15888), .ZN(n15900) );
  INV_X1 U19066 ( .A(n15891), .ZN(n15895) );
  NAND2_X1 U19067 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15892), .ZN(
        n15902) );
  AOI221_X1 U19068 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n11902), .C2(n15901), .A(
        n15902), .ZN(n15894) );
  OAI22_X1 U19069 ( .A1(n19741), .A2(n19955), .B1(n20603), .B2(n19927), .ZN(
        n15893) );
  AOI211_X1 U19070 ( .C1(n15895), .C2(n19952), .A(n15894), .B(n15893), .ZN(
        n15896) );
  OAI21_X1 U19071 ( .B1(n15900), .B2(n11902), .A(n15896), .ZN(P1_U3023) );
  INV_X1 U19072 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20757) );
  OAI22_X1 U19073 ( .A1(n19750), .A2(n19955), .B1(n20757), .B2(n19927), .ZN(
        n15897) );
  AOI21_X1 U19074 ( .B1(n15898), .B2(n19952), .A(n15897), .ZN(n15899) );
  OAI221_X1 U19075 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15902), .C1(
        n15901), .C2(n15900), .A(n15899), .ZN(P1_U3024) );
  NAND2_X1 U19076 ( .A1(n19922), .A2(n15903), .ZN(n19938) );
  INV_X1 U19077 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n15904) );
  OAI22_X1 U19078 ( .A1(n19955), .A2(n15905), .B1(n19927), .B2(n15904), .ZN(
        n15906) );
  INV_X1 U19079 ( .A(n15906), .ZN(n15911) );
  INV_X1 U19080 ( .A(n15907), .ZN(n15909) );
  AOI22_X1 U19081 ( .A1(n15909), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n15908), .B2(n19952), .ZN(n15910) );
  OAI211_X1 U19082 ( .C1(n15912), .C2(n19938), .A(n15911), .B(n15910), .ZN(
        P1_U3026) );
  OR3_X1 U19083 ( .A1(n15915), .A2(n15914), .A3(n15913), .ZN(n15916) );
  OAI21_X1 U19084 ( .B1(n15918), .B2(n15917), .A(n15916), .ZN(P1_U3468) );
  NAND2_X1 U19085 ( .A1(n20386), .A2(n20666), .ZN(n15925) );
  NAND4_X1 U19086 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20573), .A4(n20666), .ZN(n15919) );
  AND2_X1 U19087 ( .A1(n15920), .A2(n15919), .ZN(n20572) );
  AOI21_X1 U19088 ( .B1(n20572), .B2(n15922), .A(n15921), .ZN(n15924) );
  AOI21_X1 U19089 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n15927), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15923) );
  AOI211_X1 U19090 ( .C1(n20670), .C2(n15925), .A(n15924), .B(n15923), .ZN(
        P1_U3162) );
  OAI221_X1 U19091 ( .B1(n20386), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20386), 
        .C2(n15927), .A(n15926), .ZN(P1_U3466) );
  AOI22_X1 U19092 ( .A1(n15928), .A2(n18852), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n18853), .ZN(n15939) );
  AOI22_X1 U19093 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18859), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n15929), .ZN(n15938) );
  AOI22_X1 U19094 ( .A1(n18855), .A2(n15930), .B1(n18854), .B2(n15931), .ZN(
        n15937) );
  INV_X1 U19095 ( .A(n15932), .ZN(n15962) );
  INV_X1 U19096 ( .A(n15933), .ZN(n15983) );
  AOI21_X1 U19097 ( .B1(n16035), .B2(n15042), .A(n9678), .ZN(n16029) );
  INV_X1 U19098 ( .A(n15934), .ZN(n16002) );
  AOI21_X1 U19099 ( .B1(n20721), .B2(n15543), .A(n15041), .ZN(n16036) );
  NOR2_X1 U19100 ( .A1(n18830), .A2(n15935), .ZN(n16016) );
  NOR2_X1 U19101 ( .A1(n16036), .A2(n16016), .ZN(n16015) );
  NOR2_X1 U19102 ( .A1(n16002), .A2(n16001), .ZN(n16000) );
  NOR2_X1 U19103 ( .A1(n18830), .A2(n16000), .ZN(n15995) );
  NOR2_X1 U19104 ( .A1(n16029), .A2(n15995), .ZN(n15994) );
  NOR2_X1 U19105 ( .A1(n15962), .A2(n15961), .ZN(n15960) );
  NAND4_X1 U19106 ( .A1(n18818), .A2(n15952), .A3(n15940), .A4(n18814), .ZN(
        n15936) );
  NAND4_X1 U19107 ( .A1(n15939), .A2(n15938), .A3(n15937), .A4(n15936), .ZN(
        P2_U2824) );
  XNOR2_X1 U19108 ( .A(n15941), .B(n15940), .ZN(n15948) );
  AOI22_X1 U19109 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18856), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18853), .ZN(n15942) );
  OAI21_X1 U19110 ( .B1(n15943), .B2(n18810), .A(n15942), .ZN(n15944) );
  AOI21_X1 U19111 ( .B1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18859), .A(
        n15944), .ZN(n15947) );
  AOI22_X1 U19112 ( .A1(n14315), .A2(n18854), .B1(n15945), .B2(n18855), .ZN(
        n15946) );
  OAI211_X1 U19113 ( .C1(n19555), .C2(n15948), .A(n15947), .B(n15946), .ZN(
        P2_U2825) );
  AOI22_X1 U19114 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n18856), .B1(n15949), 
        .B2(n18852), .ZN(n15959) );
  AOI22_X1 U19115 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n18853), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18859), .ZN(n15958) );
  AOI22_X1 U19116 ( .A1(n15951), .A2(n18854), .B1(n15950), .B2(n18855), .ZN(
        n15957) );
  AOI21_X1 U19117 ( .B1(n15954), .B2(n15953), .A(n15952), .ZN(n15955) );
  NAND2_X1 U19118 ( .A1(n18818), .A2(n15955), .ZN(n15956) );
  NAND4_X1 U19119 ( .A1(n15959), .A2(n15958), .A3(n15957), .A4(n15956), .ZN(
        P2_U2826) );
  AOI211_X1 U19120 ( .C1(n15962), .C2(n15961), .A(n15960), .B(n19555), .ZN(
        n15967) );
  AOI22_X1 U19121 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n18853), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n18856), .ZN(n15964) );
  NAND2_X1 U19122 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18859), .ZN(
        n15963) );
  OAI211_X1 U19123 ( .C1(n18810), .C2(n15965), .A(n15964), .B(n15963), .ZN(
        n15966) );
  AOI211_X1 U19124 ( .C1(n18854), .C2(n13525), .A(n15967), .B(n15966), .ZN(
        n15968) );
  OAI21_X1 U19125 ( .B1(n15969), .B2(n18842), .A(n15968), .ZN(P2_U2827) );
  AOI22_X1 U19126 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n18853), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n18856), .ZN(n15972) );
  AOI22_X1 U19127 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18838), .B1(
        n15970), .B2(n18852), .ZN(n15971) );
  OAI211_X1 U19128 ( .C1(n15973), .C2(n18842), .A(n15972), .B(n15971), .ZN(
        n15977) );
  AOI211_X1 U19129 ( .C1(n15975), .C2(n9906), .A(n15974), .B(n19555), .ZN(
        n15976) );
  NOR2_X1 U19130 ( .A1(n15977), .A2(n15976), .ZN(n15978) );
  OAI21_X1 U19131 ( .B1(n15979), .B2(n18822), .A(n15978), .ZN(P2_U2828) );
  INV_X1 U19132 ( .A(n15980), .ZN(n15989) );
  AOI211_X1 U19133 ( .C1(n15983), .C2(n15982), .A(n15981), .B(n19555), .ZN(
        n15988) );
  AOI22_X1 U19134 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n18853), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n18856), .ZN(n15985) );
  OAI211_X1 U19135 ( .C1(n15986), .C2(n18842), .A(n15985), .B(n15984), .ZN(
        n15987) );
  AOI211_X1 U19136 ( .C1(n18854), .C2(n15989), .A(n15988), .B(n15987), .ZN(
        n15990) );
  INV_X1 U19137 ( .A(n15990), .ZN(P2_U2829) );
  AOI22_X1 U19138 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n18853), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n18856), .ZN(n15992) );
  AOI22_X1 U19139 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18838), .B1(
        n9638), .B2(n18852), .ZN(n15991) );
  OAI211_X1 U19140 ( .C1(n15993), .C2(n18842), .A(n15992), .B(n15991), .ZN(
        n15997) );
  AOI211_X1 U19141 ( .C1(n16029), .C2(n15995), .A(n15994), .B(n19555), .ZN(
        n15996) );
  NOR2_X1 U19142 ( .A1(n15997), .A2(n15996), .ZN(n15998) );
  OAI21_X1 U19143 ( .B1(n15999), .B2(n18822), .A(n15998), .ZN(P2_U2830) );
  AOI211_X1 U19144 ( .C1(n16002), .C2(n16001), .A(n16000), .B(n19555), .ZN(
        n16008) );
  AOI22_X1 U19145 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n18853), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n18856), .ZN(n16005) );
  AOI22_X1 U19146 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18838), .B1(
        n16003), .B2(n18852), .ZN(n16004) );
  OAI211_X1 U19147 ( .C1(n16006), .C2(n18842), .A(n16005), .B(n16004), .ZN(
        n16007) );
  AOI211_X1 U19148 ( .C1(n18854), .C2(n16009), .A(n16008), .B(n16007), .ZN(
        n16010) );
  INV_X1 U19149 ( .A(n16010), .ZN(P2_U2831) );
  OR2_X1 U19150 ( .A1(n16012), .A2(n16011), .ZN(n16014) );
  AND2_X1 U19151 ( .A1(n16014), .A2(n16013), .ZN(n16123) );
  AOI211_X1 U19152 ( .C1(n16036), .C2(n16016), .A(n16015), .B(n19555), .ZN(
        n16021) );
  AOI22_X1 U19153 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n18853), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n18856), .ZN(n16018) );
  NAND2_X1 U19154 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18859), .ZN(
        n16017) );
  OAI211_X1 U19155 ( .C1(n18810), .C2(n16019), .A(n16018), .B(n16017), .ZN(
        n16020) );
  AOI211_X1 U19156 ( .C1(n18855), .C2(n16123), .A(n16021), .B(n16020), .ZN(
        n16022) );
  OAI21_X1 U19157 ( .B1(n16039), .B2(n18822), .A(n16022), .ZN(P2_U2832) );
  AOI22_X1 U19158 ( .A1(n16024), .A2(n16023), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n18920), .ZN(n16028) );
  AOI22_X1 U19159 ( .A1(n18864), .A2(BUF2_REG_23__SCAN_IN), .B1(n18865), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16027) );
  AOI22_X1 U19160 ( .A1(n16025), .A2(n18922), .B1(n18921), .B2(n16123), .ZN(
        n16026) );
  NAND3_X1 U19161 ( .A1(n16028), .A2(n16027), .A3(n16026), .ZN(P2_U2896) );
  AOI22_X1 U19162 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n18980), .B1(n16107), 
        .B2(n16029), .ZN(n16034) );
  AOI222_X1 U19163 ( .A1(n16032), .A2(n16102), .B1(n16114), .B2(n16031), .C1(
        n18988), .C2(n16030), .ZN(n16033) );
  OAI211_X1 U19164 ( .C1(n16035), .C2(n16121), .A(n16034), .B(n16033), .ZN(
        P2_U2989) );
  AOI22_X1 U19165 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n18980), .B1(n16107), 
        .B2(n16036), .ZN(n16044) );
  XOR2_X1 U19166 ( .A(n16037), .B(n16038), .Z(n16127) );
  INV_X1 U19167 ( .A(n16039), .ZN(n16126) );
  AOI21_X1 U19168 ( .B1(n16040), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16042) );
  NOR2_X1 U19169 ( .A1(n16042), .A2(n16041), .ZN(n16125) );
  AOI222_X1 U19170 ( .A1(n16127), .A2(n16102), .B1(n18988), .B2(n16126), .C1(
        n16114), .C2(n16125), .ZN(n16043) );
  OAI211_X1 U19171 ( .C1(n20721), .C2(n16121), .A(n16044), .B(n16043), .ZN(
        P2_U2991) );
  AOI22_X1 U19172 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18979), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18980), .ZN(n16050) );
  OAI22_X1 U19173 ( .A1(n16046), .A2(n18982), .B1(n18984), .B2(n16045), .ZN(
        n16047) );
  AOI21_X1 U19174 ( .B1(n18988), .B2(n16048), .A(n16047), .ZN(n16049) );
  OAI211_X1 U19175 ( .C1(n18992), .C2(n16051), .A(n16050), .B(n16049), .ZN(
        P2_U2992) );
  AOI22_X1 U19176 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n18980), .B1(n16107), 
        .B2(n18703), .ZN(n16055) );
  AOI22_X1 U19177 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n18980), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18979), .ZN(n16061) );
  OAI22_X1 U19178 ( .A1(n16058), .A2(n18984), .B1(n18982), .B2(n16057), .ZN(
        n16059) );
  AOI21_X1 U19179 ( .B1(n18988), .B2(n18719), .A(n16059), .ZN(n16060) );
  OAI211_X1 U19180 ( .C1(n18992), .C2(n18716), .A(n16061), .B(n16060), .ZN(
        P2_U3000) );
  AOI22_X1 U19181 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n18980), .B1(n16107), 
        .B2(n18724), .ZN(n16066) );
  OAI22_X1 U19182 ( .A1(n16063), .A2(n18982), .B1(n16117), .B2(n16062), .ZN(
        n16064) );
  AOI21_X1 U19183 ( .B1(n9626), .B2(n16114), .A(n16064), .ZN(n16065) );
  OAI211_X1 U19184 ( .C1(n16067), .C2(n16121), .A(n16066), .B(n16065), .ZN(
        P2_U3001) );
  AOI22_X1 U19185 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18979), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18980), .ZN(n16072) );
  OAI22_X1 U19186 ( .A1(n16069), .A2(n18984), .B1(n16068), .B2(n18982), .ZN(
        n16070) );
  AOI21_X1 U19187 ( .B1(n18988), .B2(n18739), .A(n16070), .ZN(n16071) );
  OAI211_X1 U19188 ( .C1(n18992), .C2(n18738), .A(n16072), .B(n16071), .ZN(
        P2_U3002) );
  AOI22_X1 U19189 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18980), .B1(n16107), 
        .B2(n18753), .ZN(n16081) );
  NAND2_X1 U19190 ( .A1(n16074), .A2(n16073), .ZN(n16077) );
  NAND2_X1 U19191 ( .A1(n10088), .A2(n16075), .ZN(n16076) );
  XNOR2_X1 U19192 ( .A(n16077), .B(n16076), .ZN(n16139) );
  INV_X1 U19193 ( .A(n18756), .ZN(n16138) );
  AOI21_X1 U19194 ( .B1(n11075), .B2(n16079), .A(n16078), .ZN(n16137) );
  AOI222_X1 U19195 ( .A1(n16139), .A2(n16102), .B1(n18988), .B2(n16138), .C1(
        n16114), .C2(n16137), .ZN(n16080) );
  OAI211_X1 U19196 ( .C1(n18743), .C2(n16121), .A(n16081), .B(n16080), .ZN(
        P2_U3003) );
  AOI22_X1 U19197 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n18980), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18979), .ZN(n16086) );
  OAI22_X1 U19198 ( .A1(n16083), .A2(n18984), .B1(n16082), .B2(n18982), .ZN(
        n16084) );
  AOI21_X1 U19199 ( .B1(n18988), .B2(n18764), .A(n16084), .ZN(n16085) );
  OAI211_X1 U19200 ( .C1(n18992), .C2(n18761), .A(n16086), .B(n16085), .ZN(
        P2_U3004) );
  AOI22_X1 U19201 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18980), .B1(n16107), 
        .B2(n18772), .ZN(n16093) );
  NAND3_X1 U19202 ( .A1(n16088), .A2(n16102), .A3(n16087), .ZN(n16089) );
  OAI21_X1 U19203 ( .B1(n16117), .B2(n18776), .A(n16089), .ZN(n16090) );
  AOI21_X1 U19204 ( .B1(n16091), .B2(n16114), .A(n16090), .ZN(n16092) );
  OAI211_X1 U19205 ( .C1(n16094), .C2(n16121), .A(n16093), .B(n16092), .ZN(
        P2_U3005) );
  AOI22_X1 U19206 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18979), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18980), .ZN(n16099) );
  OAI22_X1 U19207 ( .A1(n16096), .A2(n18984), .B1(n16095), .B2(n18982), .ZN(
        n16097) );
  AOI21_X1 U19208 ( .B1(n18988), .B2(n18783), .A(n16097), .ZN(n16098) );
  OAI211_X1 U19209 ( .C1(n18992), .C2(n18781), .A(n16099), .B(n16098), .ZN(
        P2_U3006) );
  AOI22_X1 U19210 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n18980), .B1(n16107), 
        .B2(n18788), .ZN(n16105) );
  AOI222_X1 U19211 ( .A1(n16103), .A2(n16102), .B1(n18988), .B2(n16101), .C1(
        n16100), .C2(n16114), .ZN(n16104) );
  OAI211_X1 U19212 ( .C1(n16106), .C2(n16121), .A(n16105), .B(n16104), .ZN(
        P2_U3007) );
  AOI22_X1 U19213 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18980), .B1(n16107), 
        .B2(n18816), .ZN(n16120) );
  XNOR2_X1 U19214 ( .A(n16108), .B(n16109), .ZN(n16153) );
  OR2_X1 U19215 ( .A1(n16153), .A2(n18982), .ZN(n16116) );
  NOR2_X1 U19216 ( .A1(n16111), .A2(n16110), .ZN(n16113) );
  XNOR2_X1 U19217 ( .A(n16113), .B(n16112), .ZN(n16155) );
  NAND2_X1 U19218 ( .A1(n16155), .A2(n16114), .ZN(n16115) );
  OAI211_X1 U19219 ( .C1(n16117), .C2(n18821), .A(n16116), .B(n16115), .ZN(
        n16118) );
  INV_X1 U19220 ( .A(n16118), .ZN(n16119) );
  OAI211_X1 U19221 ( .C1(n16122), .C2(n16121), .A(n16120), .B(n16119), .ZN(
        P2_U3009) );
  AOI22_X1 U19222 ( .A1(n16124), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n16150), .B2(n16123), .ZN(n16133) );
  AOI222_X1 U19223 ( .A1(n16127), .A2(n18999), .B1(n19004), .B2(n16126), .C1(
        n16154), .C2(n16125), .ZN(n16132) );
  NAND2_X1 U19224 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n18980), .ZN(n16131) );
  OAI211_X1 U19225 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n16129), .B(n16128), .ZN(
        n16130) );
  NAND4_X1 U19226 ( .A1(n16133), .A2(n16132), .A3(n16131), .A4(n16130), .ZN(
        P2_U3023) );
  AOI21_X1 U19227 ( .B1(n16135), .B2(n16134), .A(n15349), .ZN(n18880) );
  AOI22_X1 U19228 ( .A1(n16136), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16150), .B2(n18880), .ZN(n16145) );
  AOI222_X1 U19229 ( .A1(n16139), .A2(n18999), .B1(n19004), .B2(n16138), .C1(
        n16154), .C2(n16137), .ZN(n16144) );
  NAND2_X1 U19230 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18980), .ZN(n16143) );
  OAI211_X1 U19231 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16141), .B(n16140), .ZN(
        n16142) );
  NAND4_X1 U19232 ( .A1(n16145), .A2(n16144), .A3(n16143), .A4(n16142), .ZN(
        P2_U3035) );
  INV_X1 U19233 ( .A(n16146), .ZN(n16149) );
  INV_X1 U19234 ( .A(n16147), .ZN(n16148) );
  AOI21_X1 U19235 ( .B1(n16149), .B2(n12840), .A(n16148), .ZN(n18896) );
  AOI22_X1 U19236 ( .A1(n16151), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n16150), .B2(n18896), .ZN(n16165) );
  OR2_X1 U19237 ( .A1(n16153), .A2(n16152), .ZN(n16157) );
  NAND2_X1 U19238 ( .A1(n16155), .A2(n16154), .ZN(n16156) );
  OAI211_X1 U19239 ( .C1(n18821), .C2(n16158), .A(n16157), .B(n16156), .ZN(
        n16159) );
  INV_X1 U19240 ( .A(n16159), .ZN(n16164) );
  NAND2_X1 U19241 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18980), .ZN(n16163) );
  OAI211_X1 U19242 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n16161), .B(n16160), .ZN(n16162) );
  NAND4_X1 U19243 ( .A1(n16165), .A2(n16164), .A3(n16163), .A4(n16162), .ZN(
        P2_U3041) );
  AND2_X1 U19244 ( .A1(n19550), .A2(n19680), .ZN(n19554) );
  INV_X1 U19245 ( .A(n19554), .ZN(n16170) );
  OAI21_X1 U19246 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16167), .A(n16166), 
        .ZN(n16169) );
  AOI211_X1 U19247 ( .C1(n16170), .C2(n16169), .A(n16168), .B(n19553), .ZN(
        n16173) );
  AND3_X1 U19248 ( .A1(n16171), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19660) );
  OAI21_X1 U19249 ( .B1(n19550), .B2(n19660), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16172) );
  OAI211_X1 U19250 ( .C1(n16175), .C2(n16174), .A(n16173), .B(n16172), .ZN(
        P2_U3176) );
  INV_X1 U19251 ( .A(n17524), .ZN(n17482) );
  OAI22_X1 U19252 ( .A1(n16190), .A2(n17628), .B1(n16188), .B2(n17482), .ZN(
        n16182) );
  AOI21_X1 U19253 ( .B1(n9987), .B2(n16177), .A(n16176), .ZN(n16181) );
  OAI21_X1 U19254 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n9682), .A(
        n16178), .ZN(n16353) );
  OAI21_X1 U19255 ( .B1(n17460), .B2(n16353), .A(n16179), .ZN(n16180) );
  AOI211_X1 U19256 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n16182), .A(
        n16181), .B(n16180), .ZN(n16186) );
  INV_X1 U19257 ( .A(n17821), .ZN(n17481) );
  INV_X1 U19258 ( .A(n17466), .ZN(n17824) );
  AOI22_X1 U19259 ( .A1(n17481), .A2(n17612), .B1(n17524), .B2(n17824), .ZN(
        n17520) );
  NOR3_X1 U19260 ( .A1(n17630), .A2(n17652), .A3(n17424), .ZN(n17280) );
  NAND3_X1 U19261 ( .A1(n16184), .A2(n17280), .A3(n16183), .ZN(n16185) );
  OAI211_X1 U19262 ( .C1(n16187), .C2(n17529), .A(n16186), .B(n16185), .ZN(
        P3_U2800) );
  AOI211_X1 U19263 ( .C1(n16191), .C2(n16211), .A(n16188), .B(n17482), .ZN(
        n16193) );
  INV_X1 U19264 ( .A(n16189), .ZN(n16212) );
  AOI211_X1 U19265 ( .C1(n16212), .C2(n16191), .A(n16190), .B(n17628), .ZN(
        n16192) );
  AOI211_X1 U19266 ( .C1(n16194), .C2(n17516), .A(n16193), .B(n16192), .ZN(
        n16202) );
  NAND2_X1 U19267 ( .A1(n9578), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16201) );
  AOI21_X1 U19268 ( .B1(n16371), .B2(n16195), .A(n9682), .ZN(n16367) );
  OAI21_X1 U19269 ( .B1(n16196), .B2(n17473), .A(n16367), .ZN(n16200) );
  OAI221_X1 U19270 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18273), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16198), .A(n16197), .ZN(
        n16199) );
  NAND4_X1 U19271 ( .A1(n16202), .A2(n16201), .A3(n16200), .A4(n16199), .ZN(
        P3_U2801) );
  OAI22_X1 U19272 ( .A1(n17821), .A2(n9776), .B1(n17466), .B2(n17823), .ZN(
        n17732) );
  AOI21_X1 U19273 ( .B1(n17733), .B2(n17732), .A(n17651), .ZN(n17681) );
  NOR2_X1 U19274 ( .A1(n17681), .A2(n9563), .ZN(n17720) );
  AND2_X1 U19275 ( .A1(n16215), .A2(n16203), .ZN(n17262) );
  AOI22_X1 U19276 ( .A1(n9578), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17720), 
        .B2(n17262), .ZN(n16222) );
  NAND3_X1 U19277 ( .A1(n16204), .A2(n17932), .A3(n16205), .ZN(n16221) );
  AOI21_X1 U19278 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17528), .A(
        n16205), .ZN(n17266) );
  NAND3_X1 U19279 ( .A1(n9570), .A2(n17850), .A3(n17266), .ZN(n16220) );
  NOR2_X1 U19280 ( .A1(n16204), .A2(n17266), .ZN(n17265) );
  INV_X1 U19281 ( .A(n16207), .ZN(n16209) );
  NAND2_X1 U19282 ( .A1(n16209), .A2(n16208), .ZN(n16210) );
  NOR2_X1 U19283 ( .A1(n17265), .A2(n16210), .ZN(n16218) );
  INV_X1 U19284 ( .A(n17823), .ZN(n17768) );
  AOI22_X1 U19285 ( .A1(n18439), .A2(n16212), .B1(n17768), .B2(n16211), .ZN(
        n16213) );
  NAND3_X1 U19286 ( .A1(n16214), .A2(n16213), .A3(n17900), .ZN(n16217) );
  NAND4_X1 U19287 ( .A1(n16222), .A2(n16221), .A3(n16220), .A4(n16219), .ZN(
        P3_U2834) );
  INV_X1 U19288 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n20699) );
  NOR4_X1 U19289 ( .A1(P3_BE_N_REG_0__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .A4(n20699), .ZN(n16224) );
  NOR4_X1 U19290 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16223) );
  NAND3_X1 U19291 ( .A1(n16224), .A2(n16223), .A3(U215), .ZN(U213) );
  INV_X1 U19292 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n18929) );
  OAI222_X1 U19293 ( .A1(U212), .A2(n18929), .B1(n16259), .B2(n16226), .C1(
        U214), .C2(n16302), .ZN(U216) );
  INV_X1 U19294 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n18932) );
  INV_X1 U19295 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16227) );
  INV_X1 U19296 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n20782) );
  OAI222_X1 U19297 ( .A1(U212), .A2(n18932), .B1(n16259), .B2(n16227), .C1(
        U214), .C2(n20782), .ZN(U217) );
  INV_X1 U19298 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16229) );
  AOI22_X1 U19299 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16257), .ZN(n16228) );
  OAI21_X1 U19300 ( .B1(n16229), .B2(n16259), .A(n16228), .ZN(U218) );
  AOI222_X1 U19301 ( .A1(n16257), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(n16268), 
        .B2(BUF1_REG_28__SCAN_IN), .C1(n16266), .C2(P1_DATAO_REG_28__SCAN_IN), 
        .ZN(n16230) );
  INV_X1 U19302 ( .A(n16230), .ZN(U219) );
  AOI22_X1 U19303 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16257), .ZN(n16231) );
  OAI21_X1 U19304 ( .B1(n14948), .B2(n16259), .A(n16231), .ZN(U220) );
  AOI22_X1 U19305 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16257), .ZN(n16232) );
  OAI21_X1 U19306 ( .B1(n16233), .B2(n16259), .A(n16232), .ZN(U221) );
  AOI22_X1 U19307 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16257), .ZN(n16234) );
  OAI21_X1 U19308 ( .B1(n14968), .B2(n16259), .A(n16234), .ZN(U222) );
  INV_X1 U19309 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16236) );
  AOI22_X1 U19310 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16257), .ZN(n16235) );
  OAI21_X1 U19311 ( .B1(n16236), .B2(n16259), .A(n16235), .ZN(U223) );
  INV_X1 U19312 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16238) );
  AOI22_X1 U19313 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16257), .ZN(n16237) );
  OAI21_X1 U19314 ( .B1(n16238), .B2(n16259), .A(n16237), .ZN(U224) );
  AOI22_X1 U19315 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16257), .ZN(n16239) );
  OAI21_X1 U19316 ( .B1(n14987), .B2(n16259), .A(n16239), .ZN(U225) );
  AOI222_X1 U19317 ( .A1(n16257), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(n16268), 
        .B2(BUF1_REG_21__SCAN_IN), .C1(n16266), .C2(P1_DATAO_REG_21__SCAN_IN), 
        .ZN(n16240) );
  INV_X1 U19318 ( .A(n16240), .ZN(U226) );
  AOI22_X1 U19319 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16257), .ZN(n16241) );
  OAI21_X1 U19320 ( .B1(n16242), .B2(n16259), .A(n16241), .ZN(U227) );
  AOI22_X1 U19321 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16257), .ZN(n16243) );
  OAI21_X1 U19322 ( .B1(n13439), .B2(n16259), .A(n16243), .ZN(U228) );
  AOI22_X1 U19323 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16257), .ZN(n16244) );
  OAI21_X1 U19324 ( .B1(n13388), .B2(n16259), .A(n16244), .ZN(U229) );
  AOI22_X1 U19325 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16257), .ZN(n16245) );
  OAI21_X1 U19326 ( .B1(n13251), .B2(n16259), .A(n16245), .ZN(U230) );
  AOI22_X1 U19327 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16257), .ZN(n16246) );
  OAI21_X1 U19328 ( .B1(n13213), .B2(n16259), .A(n16246), .ZN(U231) );
  AOI22_X1 U19329 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16257), .ZN(n16247) );
  OAI21_X1 U19330 ( .B1(n14597), .B2(n16259), .A(n16247), .ZN(U232) );
  INV_X1 U19331 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16249) );
  AOI22_X1 U19332 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16257), .ZN(n16248) );
  OAI21_X1 U19333 ( .B1(n16249), .B2(n16259), .A(n16248), .ZN(U233) );
  INV_X1 U19334 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16251) );
  AOI22_X1 U19335 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16257), .ZN(n16250) );
  OAI21_X1 U19336 ( .B1(n16251), .B2(n16259), .A(n16250), .ZN(U234) );
  AOI22_X1 U19337 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16257), .ZN(n16252) );
  OAI21_X1 U19338 ( .B1(n12359), .B2(n16259), .A(n16252), .ZN(U235) );
  INV_X1 U19339 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16281) );
  INV_X1 U19340 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n20702) );
  OAI222_X1 U19341 ( .A1(U212), .A2(n16281), .B1(n16259), .B2(n12299), .C1(
        U214), .C2(n20702), .ZN(U236) );
  INV_X1 U19342 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n20685) );
  AOI22_X1 U19343 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n16268), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16257), .ZN(n16253) );
  OAI21_X1 U19344 ( .B1(n20685), .B2(U214), .A(n16253), .ZN(U237) );
  INV_X1 U19345 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16279) );
  AOI22_X1 U19346 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16268), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16266), .ZN(n16254) );
  OAI21_X1 U19347 ( .B1(n16279), .B2(U212), .A(n16254), .ZN(U238) );
  AOI22_X1 U19348 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16257), .ZN(n16255) );
  OAI21_X1 U19349 ( .B1(n16256), .B2(n16259), .A(n16255), .ZN(U239) );
  AOI22_X1 U19350 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16266), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16257), .ZN(n16258) );
  OAI21_X1 U19351 ( .B1(n16260), .B2(n16259), .A(n16258), .ZN(U240) );
  INV_X1 U19352 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16276) );
  AOI22_X1 U19353 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16268), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16266), .ZN(n16261) );
  OAI21_X1 U19354 ( .B1(n16276), .B2(U212), .A(n16261), .ZN(U241) );
  INV_X1 U19355 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16275) );
  AOI22_X1 U19356 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16268), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16266), .ZN(n16262) );
  OAI21_X1 U19357 ( .B1(n16275), .B2(U212), .A(n16262), .ZN(U242) );
  INV_X1 U19358 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16274) );
  AOI22_X1 U19359 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n16268), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16266), .ZN(n16263) );
  OAI21_X1 U19360 ( .B1(n16274), .B2(U212), .A(n16263), .ZN(U243) );
  INV_X1 U19361 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16273) );
  AOI22_X1 U19362 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16268), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16266), .ZN(n16264) );
  OAI21_X1 U19363 ( .B1(n16273), .B2(U212), .A(n16264), .ZN(U244) );
  INV_X1 U19364 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16272) );
  AOI22_X1 U19365 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16268), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16266), .ZN(n16265) );
  OAI21_X1 U19366 ( .B1(n16272), .B2(U212), .A(n16265), .ZN(U245) );
  INV_X1 U19367 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16271) );
  AOI22_X1 U19368 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16268), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16266), .ZN(n16267) );
  OAI21_X1 U19369 ( .B1(n16271), .B2(U212), .A(n16267), .ZN(U246) );
  INV_X1 U19370 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16270) );
  AOI22_X1 U19371 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16268), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16266), .ZN(n16269) );
  OAI21_X1 U19372 ( .B1(n16270), .B2(U212), .A(n16269), .ZN(U247) );
  INV_X1 U19373 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n17961) );
  AOI22_X1 U19374 ( .A1(n16298), .A2(n16270), .B1(n17961), .B2(U215), .ZN(U251) );
  INV_X1 U19375 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n17966) );
  AOI22_X1 U19376 ( .A1(n16298), .A2(n16271), .B1(n17966), .B2(U215), .ZN(U252) );
  INV_X1 U19377 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n20714) );
  AOI22_X1 U19378 ( .A1(n16298), .A2(n16272), .B1(n20714), .B2(U215), .ZN(U253) );
  INV_X1 U19379 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n17972) );
  AOI22_X1 U19380 ( .A1(n16298), .A2(n16273), .B1(n17972), .B2(U215), .ZN(U254) );
  INV_X1 U19381 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n17978) );
  AOI22_X1 U19382 ( .A1(n16300), .A2(n16274), .B1(n17978), .B2(U215), .ZN(U255) );
  INV_X1 U19383 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n17982) );
  AOI22_X1 U19384 ( .A1(n16298), .A2(n16275), .B1(n17982), .B2(U215), .ZN(U256) );
  INV_X1 U19385 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n17987) );
  AOI22_X1 U19386 ( .A1(n16298), .A2(n16276), .B1(n17987), .B2(U215), .ZN(U257) );
  INV_X1 U19387 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16277) );
  AOI22_X1 U19388 ( .A1(n16300), .A2(n16277), .B1(n17992), .B2(U215), .ZN(U258) );
  INV_X1 U19389 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16278) );
  INV_X1 U19390 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U19391 ( .A1(n16298), .A2(n16278), .B1(n17115), .B2(U215), .ZN(U259) );
  INV_X1 U19392 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U19393 ( .A1(n16300), .A2(n16279), .B1(n17110), .B2(U215), .ZN(U260) );
  OAI22_X1 U19394 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16300), .ZN(n16280) );
  INV_X1 U19395 ( .A(n16280), .ZN(U261) );
  INV_X1 U19396 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U19397 ( .A1(n16298), .A2(n16281), .B1(n17101), .B2(U215), .ZN(U262) );
  INV_X1 U19398 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16282) );
  INV_X1 U19399 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U19400 ( .A1(n16300), .A2(n16282), .B1(n17097), .B2(U215), .ZN(U263) );
  INV_X1 U19401 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16283) );
  INV_X1 U19402 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U19403 ( .A1(n16298), .A2(n16283), .B1(n17092), .B2(U215), .ZN(U264) );
  OAI22_X1 U19404 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16298), .ZN(n16284) );
  INV_X1 U19405 ( .A(n16284), .ZN(U265) );
  OAI22_X1 U19406 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16298), .ZN(n16285) );
  INV_X1 U19407 ( .A(n16285), .ZN(U266) );
  OAI22_X1 U19408 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16298), .ZN(n16286) );
  INV_X1 U19409 ( .A(n16286), .ZN(U267) );
  OAI22_X1 U19410 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16298), .ZN(n16287) );
  INV_X1 U19411 ( .A(n16287), .ZN(U268) );
  OAI22_X1 U19412 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16298), .ZN(n16288) );
  INV_X1 U19413 ( .A(n16288), .ZN(U269) );
  OAI22_X1 U19414 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16298), .ZN(n16289) );
  INV_X1 U19415 ( .A(n16289), .ZN(U270) );
  OAI22_X1 U19416 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16298), .ZN(n16290) );
  INV_X1 U19417 ( .A(n16290), .ZN(U271) );
  OAI22_X1 U19418 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16298), .ZN(n16291) );
  INV_X1 U19419 ( .A(n16291), .ZN(U272) );
  OAI22_X1 U19420 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16300), .ZN(n16292) );
  INV_X1 U19421 ( .A(n16292), .ZN(U273) );
  OAI22_X1 U19422 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16298), .ZN(n16293) );
  INV_X1 U19423 ( .A(n16293), .ZN(U274) );
  INV_X1 U19424 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16294) );
  INV_X1 U19425 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n17963) );
  AOI22_X1 U19426 ( .A1(n16300), .A2(n16294), .B1(n17963), .B2(U215), .ZN(U275) );
  OAI22_X1 U19427 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16298), .ZN(n16295) );
  INV_X1 U19428 ( .A(n16295), .ZN(U276) );
  INV_X1 U19429 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16296) );
  AOI22_X1 U19430 ( .A1(n16298), .A2(n16296), .B1(n14959), .B2(U215), .ZN(U277) );
  OAI22_X1 U19431 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16298), .ZN(n16297) );
  INV_X1 U19432 ( .A(n16297), .ZN(U278) );
  INV_X1 U19433 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n20748) );
  INV_X1 U19434 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17977) );
  AOI22_X1 U19435 ( .A1(n16298), .A2(n20748), .B1(n17977), .B2(U215), .ZN(U279) );
  OAI22_X1 U19436 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16300), .ZN(n16299) );
  INV_X1 U19437 ( .A(n16299), .ZN(U280) );
  INV_X1 U19438 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n17986) );
  AOI22_X1 U19439 ( .A1(n16300), .A2(n18932), .B1(n17986), .B2(U215), .ZN(U281) );
  INV_X1 U19440 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17994) );
  AOI22_X1 U19441 ( .A1(n16300), .A2(n18929), .B1(n17994), .B2(U215), .ZN(U282) );
  INV_X1 U19442 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16301) );
  AOI222_X1 U19443 ( .A1(n16302), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n18929), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16301), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16303) );
  INV_X2 U19444 ( .A(n16305), .ZN(n16304) );
  INV_X1 U19445 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18496) );
  INV_X1 U19446 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19588) );
  AOI22_X1 U19447 ( .A1(n16304), .A2(n18496), .B1(n19588), .B2(n16305), .ZN(
        U347) );
  INV_X1 U19448 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18494) );
  INV_X1 U19449 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19587) );
  AOI22_X1 U19450 ( .A1(n16303), .A2(n18494), .B1(n19587), .B2(n16305), .ZN(
        U348) );
  INV_X1 U19451 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18492) );
  INV_X1 U19452 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19586) );
  AOI22_X1 U19453 ( .A1(n16304), .A2(n18492), .B1(n19586), .B2(n16305), .ZN(
        U349) );
  INV_X1 U19454 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18490) );
  INV_X1 U19455 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19585) );
  AOI22_X1 U19456 ( .A1(n16304), .A2(n18490), .B1(n19585), .B2(n16305), .ZN(
        U350) );
  INV_X1 U19457 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18488) );
  INV_X1 U19458 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19584) );
  AOI22_X1 U19459 ( .A1(n16304), .A2(n18488), .B1(n19584), .B2(n16305), .ZN(
        U351) );
  INV_X1 U19460 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18486) );
  INV_X1 U19461 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19583) );
  AOI22_X1 U19462 ( .A1(n16304), .A2(n18486), .B1(n19583), .B2(n16305), .ZN(
        U352) );
  INV_X1 U19463 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18484) );
  INV_X1 U19464 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19582) );
  AOI22_X1 U19465 ( .A1(n16304), .A2(n18484), .B1(n19582), .B2(n16305), .ZN(
        U353) );
  INV_X1 U19466 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18481) );
  AOI22_X1 U19467 ( .A1(n16304), .A2(n18481), .B1(n19581), .B2(n16305), .ZN(
        U354) );
  INV_X1 U19468 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18535) );
  INV_X1 U19469 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19621) );
  AOI22_X1 U19470 ( .A1(n16304), .A2(n18535), .B1(n19621), .B2(n16305), .ZN(
        U355) );
  INV_X1 U19471 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20722) );
  INV_X1 U19472 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19618) );
  AOI22_X1 U19473 ( .A1(n16304), .A2(n20722), .B1(n19618), .B2(n16305), .ZN(
        U356) );
  INV_X1 U19474 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18529) );
  INV_X1 U19475 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19617) );
  AOI22_X1 U19476 ( .A1(n16304), .A2(n18529), .B1(n19617), .B2(n16305), .ZN(
        U357) );
  INV_X1 U19477 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18527) );
  INV_X1 U19478 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19614) );
  AOI22_X1 U19479 ( .A1(n16304), .A2(n18527), .B1(n19614), .B2(n16305), .ZN(
        U358) );
  INV_X1 U19480 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18525) );
  INV_X1 U19481 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19612) );
  AOI22_X1 U19482 ( .A1(n16304), .A2(n18525), .B1(n19612), .B2(n16305), .ZN(
        U359) );
  INV_X1 U19483 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18523) );
  INV_X1 U19484 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19610) );
  AOI22_X1 U19485 ( .A1(n16304), .A2(n18523), .B1(n19610), .B2(n16305), .ZN(
        U360) );
  INV_X1 U19486 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18521) );
  INV_X1 U19487 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19608) );
  AOI22_X1 U19488 ( .A1(n16304), .A2(n18521), .B1(n19608), .B2(n16305), .ZN(
        U361) );
  INV_X1 U19489 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18519) );
  INV_X1 U19490 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19606) );
  AOI22_X1 U19491 ( .A1(n16304), .A2(n18519), .B1(n19606), .B2(n16305), .ZN(
        U362) );
  INV_X1 U19492 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18517) );
  INV_X1 U19493 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19605) );
  AOI22_X1 U19494 ( .A1(n16304), .A2(n18517), .B1(n19605), .B2(n16305), .ZN(
        U363) );
  INV_X1 U19495 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18515) );
  INV_X1 U19496 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19603) );
  AOI22_X1 U19497 ( .A1(n16304), .A2(n18515), .B1(n19603), .B2(n16305), .ZN(
        U364) );
  INV_X1 U19498 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18480) );
  INV_X1 U19499 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19580) );
  AOI22_X1 U19500 ( .A1(n16304), .A2(n18480), .B1(n19580), .B2(n16305), .ZN(
        U365) );
  INV_X1 U19501 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18513) );
  INV_X1 U19502 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20761) );
  AOI22_X1 U19503 ( .A1(n16304), .A2(n18513), .B1(n20761), .B2(n16305), .ZN(
        U366) );
  INV_X1 U19504 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18511) );
  INV_X1 U19505 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19600) );
  AOI22_X1 U19506 ( .A1(n16304), .A2(n18511), .B1(n19600), .B2(n16305), .ZN(
        U367) );
  INV_X1 U19507 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18509) );
  INV_X1 U19508 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19599) );
  AOI22_X1 U19509 ( .A1(n16304), .A2(n18509), .B1(n19599), .B2(n16305), .ZN(
        U368) );
  INV_X1 U19510 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18506) );
  INV_X1 U19511 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19597) );
  AOI22_X1 U19512 ( .A1(n16304), .A2(n18506), .B1(n19597), .B2(n16305), .ZN(
        U369) );
  INV_X1 U19513 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18505) );
  INV_X1 U19514 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19596) );
  AOI22_X1 U19515 ( .A1(n16304), .A2(n18505), .B1(n19596), .B2(n16305), .ZN(
        U370) );
  INV_X1 U19516 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18503) );
  INV_X1 U19517 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19594) );
  AOI22_X1 U19518 ( .A1(n16303), .A2(n18503), .B1(n19594), .B2(n16305), .ZN(
        U371) );
  INV_X1 U19519 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18500) );
  INV_X1 U19520 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19593) );
  AOI22_X1 U19521 ( .A1(n16304), .A2(n18500), .B1(n19593), .B2(n16305), .ZN(
        U372) );
  INV_X1 U19522 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18499) );
  INV_X1 U19523 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19592) );
  AOI22_X1 U19524 ( .A1(n16304), .A2(n18499), .B1(n19592), .B2(n16305), .ZN(
        U373) );
  INV_X1 U19525 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20700) );
  INV_X1 U19526 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19591) );
  AOI22_X1 U19527 ( .A1(n16304), .A2(n20700), .B1(n19591), .B2(n16305), .ZN(
        U374) );
  INV_X1 U19528 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18498) );
  INV_X1 U19529 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19590) );
  AOI22_X1 U19530 ( .A1(n16303), .A2(n18498), .B1(n19590), .B2(n16305), .ZN(
        U375) );
  INV_X1 U19531 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20727) );
  INV_X1 U19532 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19579) );
  AOI22_X1 U19533 ( .A1(n16303), .A2(n20727), .B1(n19579), .B2(n16305), .ZN(
        U376) );
  INV_X1 U19534 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16306) );
  NAND2_X1 U19535 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18478), .ZN(n18470) );
  OR2_X1 U19536 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n18462) );
  OAI21_X1 U19537 ( .B1(n18475), .B2(n18470), .A(n18462), .ZN(n18541) );
  OAI21_X1 U19538 ( .B1(n18475), .B2(n16306), .A(n18459), .ZN(P3_U2633) );
  INV_X1 U19539 ( .A(n18617), .ZN(n16308) );
  OAI21_X1 U19540 ( .B1(n16313), .B2(n17151), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16307) );
  OAI21_X1 U19541 ( .B1(n16308), .B2(n18603), .A(n16307), .ZN(P3_U2634) );
  AOI21_X1 U19542 ( .B1(n18475), .B2(n18478), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16309) );
  AOI22_X1 U19543 ( .A1(n18532), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16309), 
        .B2(n18612), .ZN(P3_U2635) );
  NOR2_X1 U19544 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18460) );
  OAI21_X1 U19545 ( .B1(n18460), .B2(BS16), .A(n18541), .ZN(n18539) );
  OAI21_X1 U19546 ( .B1(n18541), .B2(n20687), .A(n18539), .ZN(P3_U2636) );
  INV_X1 U19547 ( .A(n16310), .ZN(n16311) );
  NOR3_X1 U19548 ( .A1(n16313), .A2(n16312), .A3(n16311), .ZN(n18428) );
  NOR2_X1 U19549 ( .A1(n18428), .A2(n18450), .ZN(n18595) );
  INV_X1 U19550 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17952) );
  OAI21_X1 U19551 ( .B1(n18595), .B2(n17952), .A(n16314), .ZN(P3_U2637) );
  INV_X1 U19552 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18587) );
  INV_X1 U19553 ( .A(P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20780) );
  INV_X1 U19554 ( .A(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20678) );
  NAND2_X1 U19555 ( .A1(n20780), .A2(n20678), .ZN(n20822) );
  OR4_X1 U19556 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16315) );
  AOI211_X1 U19557 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(n20822), .B(n16315), .ZN(n16323) );
  NOR4_X1 U19558 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16322) );
  NOR4_X1 U19559 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16321) );
  NOR4_X1 U19560 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16319) );
  NOR4_X1 U19561 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16318) );
  NOR4_X1 U19562 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16317) );
  NOR4_X1 U19563 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16316) );
  AND4_X1 U19564 ( .A1(n16319), .A2(n16318), .A3(n16317), .A4(n16316), .ZN(
        n16320) );
  NAND4_X1 U19565 ( .A1(n16323), .A2(n16322), .A3(n16321), .A4(n16320), .ZN(
        n18586) );
  INV_X1 U19566 ( .A(n18586), .ZN(n18584) );
  INV_X1 U19567 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n20741) );
  NAND2_X1 U19568 ( .A1(n18584), .A2(n20741), .ZN(n18583) );
  NOR3_X1 U19569 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A3(n18583), .ZN(n16325) );
  AOI21_X1 U19570 ( .B1(P3_BYTEENABLE_REG_1__SCAN_IN), .B2(n18586), .A(n16325), 
        .ZN(n16324) );
  OAI21_X1 U19571 ( .B1(n18587), .B2(n18586), .A(n16324), .ZN(P3_U2638) );
  NAND2_X1 U19572 ( .A1(n18584), .A2(n18587), .ZN(n18577) );
  AOI21_X1 U19573 ( .B1(P3_BYTEENABLE_REG_3__SCAN_IN), .B2(n18586), .A(n16325), 
        .ZN(n16326) );
  OAI21_X1 U19574 ( .B1(P3_DATAWIDTH_REG_1__SCAN_IN), .B2(n18577), .A(n16326), 
        .ZN(P3_U2639) );
  NAND2_X1 U19575 ( .A1(n16445), .A2(n16771), .ZN(n16444) );
  NAND2_X1 U19576 ( .A1(n16435), .A2(n16678), .ZN(n16424) );
  NAND2_X1 U19577 ( .A1(n16414), .A2(n16724), .ZN(n16404) );
  NOR2_X1 U19578 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16404), .ZN(n16391) );
  INV_X1 U19579 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16387) );
  NAND2_X1 U19580 ( .A1(n16391), .A2(n16387), .ZN(n16386) );
  NOR2_X1 U19581 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16386), .ZN(n16373) );
  INV_X1 U19582 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16714) );
  NAND2_X1 U19583 ( .A1(n16373), .A2(n16714), .ZN(n16352) );
  NOR2_X1 U19584 ( .A1(n16663), .A2(n16352), .ZN(n16359) );
  INV_X1 U19585 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16330) );
  INV_X1 U19586 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18536) );
  INV_X1 U19587 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18524) );
  INV_X1 U19588 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18520) );
  INV_X1 U19589 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18516) );
  INV_X1 U19590 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18514) );
  NOR3_X1 U19591 ( .A1(n18516), .A2(n18514), .A3(n16432), .ZN(n16421) );
  NAND3_X1 U19592 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16327), .A3(n16421), 
        .ZN(n16401) );
  NOR2_X1 U19593 ( .A1(n18520), .A2(n16401), .ZN(n16405) );
  NAND2_X1 U19594 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16405), .ZN(n16400) );
  NOR2_X1 U19595 ( .A1(n18524), .A2(n16400), .ZN(n16332) );
  NAND2_X1 U19596 ( .A1(n16590), .A2(n16332), .ZN(n16383) );
  NAND2_X1 U19597 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16372) );
  NOR2_X1 U19598 ( .A1(n16383), .A2(n16372), .ZN(n16362) );
  NAND2_X1 U19599 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16362), .ZN(n16331) );
  NOR3_X1 U19600 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18536), .A3(n16331), 
        .ZN(n16329) );
  INV_X1 U19601 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16682) );
  OAI22_X1 U19602 ( .A1(n9983), .A2(n16658), .B1(n16682), .B2(n16638), .ZN(
        n16328) );
  AOI211_X1 U19603 ( .C1(n16359), .C2(n16330), .A(n16329), .B(n16328), .ZN(
        n16351) );
  NOR2_X1 U19604 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16331), .ZN(n16357) );
  INV_X1 U19605 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18531) );
  OR2_X1 U19606 ( .A1(n16664), .A2(n16332), .ZN(n16399) );
  NAND2_X1 U19607 ( .A1(n16674), .A2(n16399), .ZN(n16396) );
  AOI221_X1 U19608 ( .B1(n18531), .B2(n16590), .C1(n16372), .C2(n16590), .A(
        n16396), .ZN(n16355) );
  INV_X1 U19609 ( .A(n16355), .ZN(n16369) );
  OAI21_X1 U19610 ( .B1(n16357), .B2(n16369), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16350) );
  INV_X1 U19611 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16335) );
  NOR2_X1 U19612 ( .A1(n16333), .A2(n17618), .ZN(n16338) );
  NAND2_X1 U19613 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16338), .ZN(
        n16336) );
  AOI21_X1 U19614 ( .B1(n16335), .B2(n16336), .A(n16334), .ZN(n17259) );
  OAI21_X1 U19615 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16338), .A(
        n16336), .ZN(n17275) );
  INV_X1 U19616 ( .A(n17275), .ZN(n16382) );
  INV_X1 U19617 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16340) );
  NOR2_X1 U19618 ( .A1(n16337), .A2(n17618), .ZN(n16345) );
  INV_X1 U19619 ( .A(n16345), .ZN(n16343) );
  NOR2_X1 U19620 ( .A1(n17304), .A2(n16343), .ZN(n17257) );
  INV_X1 U19621 ( .A(n17257), .ZN(n16339) );
  AOI21_X1 U19622 ( .B1(n16340), .B2(n16339), .A(n16338), .ZN(n17290) );
  INV_X1 U19623 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16342) );
  NAND2_X1 U19624 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16345), .ZN(
        n16341) );
  AOI21_X1 U19625 ( .B1(n16342), .B2(n16341), .A(n17257), .ZN(n17297) );
  INV_X1 U19626 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17313) );
  OAI22_X1 U19627 ( .A1(n17313), .A2(n16343), .B1(n16345), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17310) );
  INV_X1 U19628 ( .A(n17310), .ZN(n16413) );
  INV_X1 U19629 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17325) );
  INV_X1 U19630 ( .A(n16347), .ZN(n16344) );
  NOR2_X1 U19631 ( .A1(n17346), .A2(n16344), .ZN(n17322) );
  INV_X1 U19632 ( .A(n17322), .ZN(n17295) );
  AOI21_X1 U19633 ( .B1(n17325), .B2(n17295), .A(n16345), .ZN(n17323) );
  INV_X1 U19634 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16437) );
  NAND2_X1 U19635 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16347), .ZN(
        n16346) );
  AOI21_X1 U19636 ( .B1(n16437), .B2(n16346), .A(n17322), .ZN(n17344) );
  XOR2_X1 U19637 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16347), .Z(
        n17353) );
  NOR2_X1 U19638 ( .A1(n17344), .A2(n16434), .ZN(n16433) );
  NOR2_X1 U19639 ( .A1(n16433), .A2(n10012), .ZN(n16423) );
  NOR2_X1 U19640 ( .A1(n17323), .A2(n16423), .ZN(n16422) );
  NOR2_X1 U19641 ( .A1(n16422), .A2(n10012), .ZN(n16412) );
  NOR2_X1 U19642 ( .A1(n17290), .A2(n16393), .ZN(n16392) );
  NOR2_X1 U19643 ( .A1(n9635), .A2(n10012), .ZN(n16366) );
  NAND4_X1 U19644 ( .A1(n10001), .A2(n18452), .A3(n16365), .A4(n16353), .ZN(
        n16349) );
  NAND3_X1 U19645 ( .A1(n16351), .A2(n16350), .A3(n16349), .ZN(P3_U2640) );
  NAND2_X1 U19646 ( .A1(n16672), .A2(n16352), .ZN(n16363) );
  NOR2_X1 U19647 ( .A1(n16365), .A2(n10012), .ZN(n16354) );
  XNOR2_X1 U19648 ( .A(n16354), .B(n16353), .ZN(n16358) );
  OAI22_X1 U19649 ( .A1(n16355), .A2(n18536), .B1(n9987), .B2(n16658), .ZN(
        n16356) );
  OAI21_X1 U19650 ( .B1(n16673), .B2(n16359), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16360) );
  OAI211_X1 U19651 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16363), .A(n16361), .B(
        n16360), .ZN(P3_U2641) );
  AOI22_X1 U19652 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16673), .B1(n16362), 
        .B2(n18531), .ZN(n16370) );
  INV_X1 U19653 ( .A(n16373), .ZN(n16364) );
  AOI21_X1 U19654 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16364), .A(n16363), .ZN(
        n16368) );
  OAI21_X1 U19655 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(P3_REIP_REG_27__SCAN_IN), 
        .A(n16372), .ZN(n16379) );
  AOI22_X1 U19656 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16603), .B1(
        n16673), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16378) );
  AOI211_X1 U19657 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16386), .A(n16373), .B(
        n16663), .ZN(n16376) );
  AOI211_X1 U19658 ( .C1(n17259), .C2(n16374), .A(n9635), .B(n16659), .ZN(
        n16375) );
  AOI211_X1 U19659 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16396), .A(n16376), 
        .B(n16375), .ZN(n16377) );
  OAI211_X1 U19660 ( .C1(n16383), .C2(n16379), .A(n16378), .B(n16377), .ZN(
        P3_U2643) );
  INV_X1 U19661 ( .A(n16396), .ZN(n16390) );
  INV_X1 U19662 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18526) );
  AOI211_X1 U19663 ( .C1(n16382), .C2(n16381), .A(n16380), .B(n16659), .ZN(
        n16385) );
  OAI22_X1 U19664 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16383), .B1(n16387), 
        .B2(n16638), .ZN(n16384) );
  AOI211_X1 U19665 ( .C1(n16603), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16385), .B(n16384), .ZN(n16389) );
  OAI211_X1 U19666 ( .C1(n16391), .C2(n16387), .A(n16672), .B(n16386), .ZN(
        n16388) );
  OAI211_X1 U19667 ( .C1(n16390), .C2(n18526), .A(n16389), .B(n16388), .ZN(
        P3_U2644) );
  AOI22_X1 U19668 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16603), .B1(
        n16673), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16398) );
  AOI211_X1 U19669 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16404), .A(n16391), .B(
        n16663), .ZN(n16395) );
  AOI211_X1 U19670 ( .C1(n17290), .C2(n16393), .A(n16392), .B(n16659), .ZN(
        n16394) );
  AOI211_X1 U19671 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16396), .A(n16395), 
        .B(n16394), .ZN(n16397) );
  OAI211_X1 U19672 ( .C1(n16400), .C2(n16399), .A(n16398), .B(n16397), .ZN(
        P3_U2645) );
  AOI22_X1 U19673 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16603), .B1(
        n16673), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16409) );
  NOR2_X1 U19674 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16664), .ZN(n16418) );
  INV_X1 U19675 ( .A(n16401), .ZN(n16417) );
  OAI21_X1 U19676 ( .B1(n16417), .B2(n16664), .A(n16674), .ZN(n16410) );
  AOI211_X1 U19677 ( .C1(n17297), .C2(n16402), .A(n9996), .B(n16659), .ZN(
        n16403) );
  AOI221_X1 U19678 ( .B1(n16418), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16410), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n16403), .ZN(n16408) );
  OAI211_X1 U19679 ( .C1(n16414), .C2(n16724), .A(n16672), .B(n16404), .ZN(
        n16407) );
  INV_X1 U19680 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18522) );
  NAND3_X1 U19681 ( .A1(n16590), .A2(n16405), .A3(n18522), .ZN(n16406) );
  NAND4_X1 U19682 ( .A1(n16409), .A2(n16408), .A3(n16407), .A4(n16406), .ZN(
        P3_U2646) );
  INV_X1 U19683 ( .A(n16410), .ZN(n16429) );
  AOI22_X1 U19684 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16603), .B1(
        n16673), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16420) );
  AOI211_X1 U19685 ( .C1(n16413), .C2(n16412), .A(n16411), .B(n16659), .ZN(
        n16416) );
  AOI211_X1 U19686 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16424), .A(n16414), .B(
        n16663), .ZN(n16415) );
  AOI211_X1 U19687 ( .C1(n16418), .C2(n16417), .A(n16416), .B(n16415), .ZN(
        n16419) );
  OAI211_X1 U19688 ( .C1(n16429), .C2(n18520), .A(n16420), .B(n16419), .ZN(
        P3_U2647) );
  NAND2_X1 U19689 ( .A1(n16421), .A2(n16473), .ZN(n16430) );
  INV_X1 U19690 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18518) );
  AOI211_X1 U19691 ( .C1(n17323), .C2(n16423), .A(n16422), .B(n16659), .ZN(
        n16427) );
  OAI211_X1 U19692 ( .C1(n16435), .C2(n16678), .A(n16672), .B(n16424), .ZN(
        n16425) );
  OAI21_X1 U19693 ( .B1(n16678), .B2(n16638), .A(n16425), .ZN(n16426) );
  AOI211_X1 U19694 ( .C1(n16603), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16427), .B(n16426), .ZN(n16428) );
  OAI221_X1 U19695 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n16430), .C1(n18518), 
        .C2(n16429), .A(n16428), .ZN(P3_U2648) );
  NOR2_X1 U19696 ( .A1(n16432), .A2(n16500), .ZN(n16431) );
  NAND2_X1 U19697 ( .A1(n16431), .A2(n18514), .ZN(n16449) );
  NOR4_X1 U19698 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n18514), .A3(n16432), 
        .A4(n16500), .ZN(n16441) );
  AOI211_X1 U19699 ( .C1(n17344), .C2(n16434), .A(n16433), .B(n16659), .ZN(
        n16440) );
  AOI211_X1 U19700 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16444), .A(n16435), .B(
        n16663), .ZN(n16439) );
  INV_X1 U19701 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16436) );
  OAI22_X1 U19702 ( .A1(n16437), .A2(n16658), .B1(n16638), .B2(n16436), .ZN(
        n16438) );
  NOR4_X1 U19703 ( .A1(n16441), .A2(n16440), .A3(n16439), .A4(n16438), .ZN(
        n16442) );
  OAI221_X1 U19704 ( .B1(n18516), .B2(n16451), .C1(n18516), .C2(n16449), .A(
        n16442), .ZN(P3_U2649) );
  AOI211_X1 U19705 ( .C1(n17353), .C2(n16443), .A(n10010), .B(n16659), .ZN(
        n16448) );
  OAI211_X1 U19706 ( .C1(n16445), .C2(n16771), .A(n16672), .B(n16444), .ZN(
        n16446) );
  OAI21_X1 U19707 ( .B1(n16771), .B2(n16638), .A(n16446), .ZN(n16447) );
  AOI211_X1 U19708 ( .C1(n16603), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16448), .B(n16447), .ZN(n16450) );
  OAI211_X1 U19709 ( .C1(n16451), .C2(n18514), .A(n16450), .B(n16449), .ZN(
        P3_U2650) );
  OAI21_X1 U19710 ( .B1(n16452), .B2(n16508), .A(n16671), .ZN(n16481) );
  AOI211_X1 U19711 ( .C1(n17376), .C2(n16454), .A(n16453), .B(n16659), .ZN(
        n16459) );
  OAI211_X1 U19712 ( .C1(n16466), .C2(n16457), .A(n16672), .B(n16455), .ZN(
        n16456) );
  OAI211_X1 U19713 ( .C1(n16638), .C2(n16457), .A(n17852), .B(n16456), .ZN(
        n16458) );
  AOI211_X1 U19714 ( .C1(n16603), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16459), .B(n16458), .ZN(n16463) );
  OAI211_X1 U19715 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16461), .B(n16460), .ZN(n16462) );
  OAI211_X1 U19716 ( .C1(n16481), .C2(n18510), .A(n16463), .B(n16462), .ZN(
        P3_U2652) );
  AOI211_X1 U19717 ( .C1(n17389), .C2(n16465), .A(n16464), .B(n16659), .ZN(
        n16470) );
  AOI211_X1 U19718 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16476), .A(n16466), .B(
        n16663), .ZN(n16469) );
  INV_X1 U19719 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17393) );
  INV_X1 U19720 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16467) );
  OAI22_X1 U19721 ( .A1(n17393), .A2(n16658), .B1(n16638), .B2(n16467), .ZN(
        n16468) );
  NOR4_X1 U19722 ( .A1(n9578), .A2(n16470), .A3(n16469), .A4(n16468), .ZN(
        n16471) );
  OAI221_X1 U19723 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16472), .C1(n18508), 
        .C2(n16481), .A(n16471), .ZN(P3_U2653) );
  NAND2_X1 U19724 ( .A1(n16485), .A2(n16473), .ZN(n16482) );
  INV_X1 U19725 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18507) );
  AOI211_X1 U19726 ( .C1(n17404), .C2(n16475), .A(n16474), .B(n16659), .ZN(
        n16479) );
  OAI211_X1 U19727 ( .C1(n16486), .C2(n16825), .A(n16672), .B(n16476), .ZN(
        n16477) );
  OAI211_X1 U19728 ( .C1(n16638), .C2(n16825), .A(n17852), .B(n16477), .ZN(
        n16478) );
  AOI211_X1 U19729 ( .C1(n16603), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16479), .B(n16478), .ZN(n16480) );
  OAI221_X1 U19730 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n16482), .C1(n18507), 
        .C2(n16481), .A(n16480), .ZN(P3_U2654) );
  NAND2_X1 U19731 ( .A1(n16671), .A2(n16508), .ZN(n16503) );
  AOI211_X1 U19732 ( .C1(n17417), .C2(n10085), .A(n16483), .B(n16659), .ZN(
        n16484) );
  AOI211_X1 U19733 ( .C1(n16673), .C2(P3_EBX_REG_16__SCAN_IN), .A(n9578), .B(
        n16484), .ZN(n16490) );
  AOI211_X1 U19734 ( .C1(n18504), .C2(n18502), .A(n16485), .B(n16500), .ZN(
        n16488) );
  AOI211_X1 U19735 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16494), .A(n16486), .B(
        n16663), .ZN(n16487) );
  AOI211_X1 U19736 ( .C1(n16603), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16488), .B(n16487), .ZN(n16489) );
  OAI211_X1 U19737 ( .C1(n18504), .C2(n16503), .A(n16490), .B(n16489), .ZN(
        P3_U2655) );
  NOR2_X1 U19738 ( .A1(n16638), .A2(n16857), .ZN(n16498) );
  OAI21_X1 U19739 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17416), .A(
        n16491), .ZN(n17425) );
  INV_X1 U19740 ( .A(n16492), .ZN(n17457) );
  NOR2_X1 U19741 ( .A1(n17618), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16647) );
  INV_X1 U19742 ( .A(n16647), .ZN(n16552) );
  OAI21_X1 U19743 ( .B1(n17457), .B2(n16552), .A(n10001), .ZN(n16529) );
  OAI21_X1 U19744 ( .B1(n17413), .B2(n10012), .A(n16529), .ZN(n16493) );
  XOR2_X1 U19745 ( .A(n17425), .B(n16493), .Z(n16496) );
  OAI211_X1 U19746 ( .C1(n16505), .C2(n16857), .A(n16672), .B(n16494), .ZN(
        n16495) );
  OAI211_X1 U19747 ( .C1(n16659), .C2(n16496), .A(n17852), .B(n16495), .ZN(
        n16497) );
  AOI211_X1 U19748 ( .C1(n16603), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16498), .B(n16497), .ZN(n16499) );
  OAI221_X1 U19749 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16500), .C1(n18502), 
        .C2(n16503), .A(n16499), .ZN(P3_U2656) );
  INV_X1 U19750 ( .A(n17443), .ZN(n17463) );
  INV_X1 U19751 ( .A(n17535), .ZN(n17521) );
  NOR2_X1 U19752 ( .A1(n17521), .A2(n17618), .ZN(n16564) );
  NAND2_X1 U19753 ( .A1(n16501), .A2(n16564), .ZN(n16550) );
  INV_X1 U19754 ( .A(n16550), .ZN(n16538) );
  NAND2_X1 U19755 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16538), .ZN(
        n16537) );
  INV_X1 U19756 ( .A(n16537), .ZN(n17459) );
  NAND2_X1 U19757 ( .A1(n17463), .A2(n17459), .ZN(n16513) );
  AOI21_X1 U19758 ( .B1(n17442), .B2(n16513), .A(n17416), .ZN(n17445) );
  OAI21_X1 U19759 ( .B1(n17463), .B2(n10012), .A(n16529), .ZN(n16520) );
  XNOR2_X1 U19760 ( .A(n17445), .B(n16520), .ZN(n16511) );
  AOI21_X1 U19761 ( .B1(n16515), .B2(P3_EBX_REG_14__SCAN_IN), .A(n16663), .ZN(
        n16502) );
  AOI21_X1 U19762 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16673), .A(n16502), .ZN(
        n16504) );
  INV_X1 U19763 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18501) );
  OAI22_X1 U19764 ( .A1(n16505), .A2(n16504), .B1(n16503), .B2(n18501), .ZN(
        n16506) );
  AOI211_X1 U19765 ( .C1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n16603), .A(
        n9578), .B(n16506), .ZN(n16510) );
  NOR2_X1 U19766 ( .A1(n16664), .A2(n16507), .ZN(n16517) );
  NAND3_X1 U19767 ( .A1(n16517), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n16508), 
        .ZN(n16509) );
  OAI211_X1 U19768 ( .C1(n16659), .C2(n16511), .A(n16510), .B(n16509), .ZN(
        P3_U2657) );
  AOI22_X1 U19769 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16603), .B1(
        n16673), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16524) );
  INV_X1 U19770 ( .A(n16525), .ZN(n16512) );
  AOI21_X1 U19771 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n16512), .A(n16663), .ZN(
        n16516) );
  INV_X1 U19772 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16528) );
  NOR2_X1 U19773 ( .A1(n16528), .A2(n16537), .ZN(n16527) );
  OAI21_X1 U19774 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16527), .A(
        n16513), .ZN(n17461) );
  NAND2_X1 U19775 ( .A1(n10001), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16660) );
  NAND2_X1 U19776 ( .A1(n18452), .A2(n16660), .ZN(n16661) );
  AOI211_X1 U19777 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n10001), .A(
        n17461), .B(n16661), .ZN(n16514) );
  AOI211_X1 U19778 ( .C1(n16516), .C2(n16515), .A(n9578), .B(n16514), .ZN(
        n16523) );
  INV_X1 U19779 ( .A(n16517), .ZN(n16519) );
  OAI21_X1 U19780 ( .B1(n16532), .B2(n16664), .A(n16674), .ZN(n16545) );
  NOR2_X1 U19781 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16664), .ZN(n16531) );
  NOR2_X1 U19782 ( .A1(n16545), .A2(n16531), .ZN(n16518) );
  MUX2_X1 U19783 ( .A(n16519), .B(n16518), .S(P3_REIP_REG_13__SCAN_IN), .Z(
        n16522) );
  NAND3_X1 U19784 ( .A1(n18452), .A2(n17461), .A3(n16520), .ZN(n16521) );
  NAND4_X1 U19785 ( .A1(n16524), .A2(n16523), .A3(n16522), .A4(n16521), .ZN(
        P3_U2658) );
  AOI211_X1 U19786 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16546), .A(n16525), .B(
        n16663), .ZN(n16526) );
  AOI21_X1 U19787 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16673), .A(n16526), .ZN(
        n16535) );
  AOI21_X1 U19788 ( .B1(n16528), .B2(n16537), .A(n16527), .ZN(n17472) );
  XNOR2_X1 U19789 ( .A(n17472), .B(n16529), .ZN(n16530) );
  AOI22_X1 U19790 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16603), .B1(
        n18452), .B2(n16530), .ZN(n16534) );
  AOI22_X1 U19791 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16545), .B1(n16532), 
        .B2(n16531), .ZN(n16533) );
  NAND4_X1 U19792 ( .A1(n16535), .A2(n16534), .A3(n16533), .A4(n17852), .ZN(
        P3_U2659) );
  OAI21_X1 U19793 ( .B1(n16664), .B2(n16536), .A(n18497), .ZN(n16544) );
  OAI21_X1 U19794 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16538), .A(
        n16537), .ZN(n17484) );
  OAI21_X1 U19795 ( .B1(n16539), .B2(n16552), .A(n10001), .ZN(n16541) );
  AOI21_X1 U19796 ( .B1(n17484), .B2(n16541), .A(n16659), .ZN(n16540) );
  OAI21_X1 U19797 ( .B1(n17484), .B2(n16541), .A(n16540), .ZN(n16542) );
  OAI211_X1 U19798 ( .C1(n17483), .C2(n16658), .A(n17852), .B(n16542), .ZN(
        n16543) );
  AOI21_X1 U19799 ( .B1(n16545), .B2(n16544), .A(n16543), .ZN(n16548) );
  OAI211_X1 U19800 ( .C1(n16553), .C2(n16906), .A(n16672), .B(n16546), .ZN(
        n16547) );
  OAI211_X1 U19801 ( .C1(n16906), .C2(n16638), .A(n16548), .B(n16547), .ZN(
        P3_U2660) );
  INV_X1 U19802 ( .A(n16564), .ZN(n16600) );
  NOR2_X1 U19803 ( .A1(n16549), .A2(n16600), .ZN(n16565) );
  OAI21_X1 U19804 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16565), .A(
        n16550), .ZN(n17499) );
  INV_X1 U19805 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17508) );
  NOR2_X1 U19806 ( .A1(n17521), .A2(n16552), .ZN(n16585) );
  NAND2_X1 U19807 ( .A1(n16551), .A2(n16585), .ZN(n16563) );
  OAI21_X1 U19808 ( .B1(n17508), .B2(n16563), .A(n10001), .ZN(n16567) );
  XNOR2_X1 U19809 ( .A(n17499), .B(n16567), .ZN(n16562) );
  AOI211_X1 U19810 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16572), .A(n16553), .B(
        n16663), .ZN(n16560) );
  NOR3_X1 U19811 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16664), .A3(n16554), .ZN(
        n16571) );
  INV_X1 U19812 ( .A(n16674), .ZN(n16588) );
  AOI21_X1 U19813 ( .B1(n16554), .B2(n16590), .A(n16588), .ZN(n16580) );
  INV_X1 U19814 ( .A(n16580), .ZN(n16555) );
  OAI21_X1 U19815 ( .B1(n16571), .B2(n16555), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16558) );
  INV_X1 U19816 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18495) );
  NAND3_X1 U19817 ( .A1(n16590), .A2(n16556), .A3(n18495), .ZN(n16557) );
  OAI211_X1 U19818 ( .C1(n16658), .C2(n17497), .A(n16558), .B(n16557), .ZN(
        n16559) );
  AOI211_X1 U19819 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16673), .A(n16560), .B(
        n16559), .ZN(n16561) );
  OAI211_X1 U19820 ( .C1(n16659), .C2(n16562), .A(n16561), .B(n17852), .ZN(
        P3_U2661) );
  AND2_X1 U19821 ( .A1(n10001), .A2(n16563), .ZN(n16568) );
  NAND2_X1 U19822 ( .A1(n16551), .A2(n16564), .ZN(n16575) );
  AOI21_X1 U19823 ( .B1(n17508), .B2(n16575), .A(n16565), .ZN(n17512) );
  INV_X1 U19824 ( .A(n17512), .ZN(n16566) );
  AOI221_X1 U19825 ( .B1(n16568), .B2(n17512), .C1(n16567), .C2(n16566), .A(
        n16659), .ZN(n16570) );
  OAI22_X1 U19826 ( .A1(n16580), .A2(n18493), .B1(n16638), .B2(n16923), .ZN(
        n16569) );
  NOR4_X1 U19827 ( .A1(n9578), .A2(n16571), .A3(n16570), .A4(n16569), .ZN(
        n16574) );
  OAI211_X1 U19828 ( .C1(n16577), .C2(n16923), .A(n16672), .B(n16572), .ZN(
        n16573) );
  OAI211_X1 U19829 ( .C1(n16658), .C2(n17508), .A(n16574), .B(n16573), .ZN(
        P3_U2662) );
  AOI21_X1 U19830 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16585), .A(
        n10012), .ZN(n16576) );
  NOR3_X1 U19831 ( .A1(n17521), .A2(n17546), .A3(n17618), .ZN(n16586) );
  OAI21_X1 U19832 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16586), .A(
        n16575), .ZN(n17530) );
  XOR2_X1 U19833 ( .A(n16576), .B(n17530), .Z(n16584) );
  AOI211_X1 U19834 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16594), .A(n16577), .B(
        n16663), .ZN(n16582) );
  AOI21_X1 U19835 ( .B1(n16590), .B2(n16578), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n16579) );
  OAI22_X1 U19836 ( .A1(n16580), .A2(n16579), .B1(n17534), .B2(n16658), .ZN(
        n16581) );
  AOI211_X1 U19837 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16673), .A(n16582), .B(
        n16581), .ZN(n16583) );
  OAI211_X1 U19838 ( .C1(n16659), .C2(n16584), .A(n16583), .B(n17852), .ZN(
        P3_U2663) );
  NOR2_X1 U19839 ( .A1(n16585), .A2(n10012), .ZN(n16601) );
  AOI21_X1 U19840 ( .B1(n17546), .B2(n16600), .A(n16586), .ZN(n17543) );
  XNOR2_X1 U19841 ( .A(n16601), .B(n17543), .ZN(n16587) );
  OAI21_X1 U19842 ( .B1(n16587), .B2(n16659), .A(n17852), .ZN(n16593) );
  NOR3_X1 U19843 ( .A1(n16664), .A2(n18482), .A3(n16644), .ZN(n16628) );
  NAND3_X1 U19844 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n16628), .ZN(n16609) );
  XNOR2_X1 U19845 ( .A(n18489), .B(n18487), .ZN(n16591) );
  AOI21_X1 U19846 ( .B1(n16590), .B2(n16589), .A(n16588), .ZN(n16612) );
  OAI22_X1 U19847 ( .A1(n16609), .A2(n16591), .B1(n18489), .B2(n16612), .ZN(
        n16592) );
  AOI211_X1 U19848 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16673), .A(n16593), .B(
        n16592), .ZN(n16597) );
  OAI211_X1 U19849 ( .C1(n16598), .C2(n16595), .A(n16672), .B(n16594), .ZN(
        n16596) );
  OAI211_X1 U19850 ( .C1(n16658), .C2(n17546), .A(n16597), .B(n16596), .ZN(
        P3_U2664) );
  AOI211_X1 U19851 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16615), .A(n16598), .B(
        n16663), .ZN(n16607) );
  NOR2_X1 U19852 ( .A1(n16599), .A2(n17618), .ZN(n16610) );
  OAI21_X1 U19853 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16610), .A(
        n16600), .ZN(n17556) );
  NAND3_X1 U19854 ( .A1(n17556), .A2(n16601), .A3(n18452), .ZN(n16605) );
  AOI211_X1 U19855 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n10001), .A(
        n17556), .B(n16661), .ZN(n16602) );
  AOI211_X1 U19856 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16603), .A(
        n9578), .B(n16602), .ZN(n16604) );
  NAND2_X1 U19857 ( .A1(n16605), .A2(n16604), .ZN(n16606) );
  AOI211_X1 U19858 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16673), .A(n16607), .B(
        n16606), .ZN(n16608) );
  OAI221_X1 U19859 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16609), .C1(n18487), 
        .C2(n16612), .A(n16608), .ZN(P3_U2665) );
  INV_X1 U19860 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16619) );
  AOI21_X1 U19861 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16628), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n16613) );
  NAND2_X1 U19862 ( .A1(n17560), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16620) );
  AOI21_X1 U19863 ( .B1(n16619), .B2(n16620), .A(n16610), .ZN(n17568) );
  OAI21_X1 U19864 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16620), .A(
        n10001), .ZN(n16621) );
  XOR2_X1 U19865 ( .A(n17568), .B(n16621), .Z(n16611) );
  OAI22_X1 U19866 ( .A1(n16613), .A2(n16612), .B1(n16659), .B2(n16611), .ZN(
        n16614) );
  AOI211_X1 U19867 ( .C1(n16673), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9578), .B(
        n16614), .ZN(n16618) );
  OAI211_X1 U19868 ( .C1(n16624), .C2(n16616), .A(n16672), .B(n16615), .ZN(
        n16617) );
  OAI211_X1 U19869 ( .C1(n16658), .C2(n16619), .A(n16618), .B(n16617), .ZN(
        P3_U2666) );
  NOR2_X1 U19870 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17583), .ZN(
        n17577) );
  NOR2_X1 U19871 ( .A1(n17583), .A2(n17618), .ZN(n16633) );
  OAI21_X1 U19872 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16633), .A(
        n16620), .ZN(n17586) );
  INV_X1 U19873 ( .A(n17586), .ZN(n16622) );
  OAI221_X1 U19874 ( .B1(n16622), .B2(n16621), .C1(n17586), .C2(n10001), .A(
        n17852), .ZN(n16623) );
  AOI21_X1 U19875 ( .B1(n17577), .B2(n16647), .A(n16623), .ZN(n16631) );
  NOR2_X1 U19876 ( .A1(n17960), .A2(n18616), .ZN(n16670) );
  AOI211_X1 U19877 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16635), .A(n16624), .B(
        n16663), .ZN(n16625) );
  AOI221_X1 U19878 ( .B1(n16926), .B2(n16670), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n16670), .A(n16625), .ZN(
        n16630) );
  OAI21_X1 U19879 ( .B1(n16626), .B2(n16664), .A(n16674), .ZN(n16641) );
  INV_X1 U19880 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18483) );
  INV_X1 U19881 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16855) );
  OAI22_X1 U19882 ( .A1(n17585), .A2(n16658), .B1(n16638), .B2(n16855), .ZN(
        n16627) );
  AOI221_X1 U19883 ( .B1(n16641), .B2(P3_REIP_REG_4__SCAN_IN), .C1(n16628), 
        .C2(n18483), .A(n16627), .ZN(n16629) );
  OAI211_X1 U19884 ( .C1(n16632), .C2(n16631), .A(n16630), .B(n16629), .ZN(
        P3_U2667) );
  INV_X1 U19885 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16643) );
  NOR2_X1 U19886 ( .A1(n16664), .A2(n16644), .ZN(n16640) );
  NAND2_X1 U19887 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16646) );
  AOI21_X1 U19888 ( .B1(n16643), .B2(n16646), .A(n16633), .ZN(n17596) );
  OAI21_X1 U19889 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16646), .A(
        n10001), .ZN(n16649) );
  XNOR2_X1 U19890 ( .A(n17596), .B(n16649), .ZN(n16634) );
  AOI21_X1 U19891 ( .B1(n18551), .B2(n18420), .A(n16926), .ZN(n18547) );
  AOI22_X1 U19892 ( .A1(n18452), .A2(n16634), .B1(n18547), .B2(n16670), .ZN(
        n16637) );
  OAI211_X1 U19893 ( .C1(n16650), .C2(n20694), .A(n16672), .B(n16635), .ZN(
        n16636) );
  OAI211_X1 U19894 ( .C1(n20694), .C2(n16638), .A(n16637), .B(n16636), .ZN(
        n16639) );
  AOI221_X1 U19895 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n16641), .C1(n16640), 
        .C2(n16641), .A(n16639), .ZN(n16642) );
  OAI21_X1 U19896 ( .B1(n16643), .B2(n16658), .A(n16642), .ZN(P3_U2668) );
  INV_X1 U19897 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17610) );
  INV_X1 U19898 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18479) );
  AOI21_X1 U19899 ( .B1(n18587), .B2(n18479), .A(n16664), .ZN(n16645) );
  AOI22_X1 U19900 ( .A1(n16673), .A2(P3_EBX_REG_2__SCAN_IN), .B1(n16645), .B2(
        n16644), .ZN(n16656) );
  OAI21_X1 U19901 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16646), .ZN(n17606) );
  NOR2_X1 U19902 ( .A1(n16647), .A2(n17606), .ZN(n16648) );
  OAI22_X1 U19903 ( .A1(n16649), .A2(n16648), .B1(n10001), .B2(n17606), .ZN(
        n16654) );
  INV_X1 U19904 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n20703) );
  INV_X1 U19905 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n16989) );
  NAND2_X1 U19906 ( .A1(n20703), .A2(n16989), .ZN(n16662) );
  AOI211_X1 U19907 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16662), .A(n16650), .B(
        n16663), .ZN(n16653) );
  NAND2_X1 U19908 ( .A1(n18560), .A2(n18392), .ZN(n18416) );
  NAND2_X1 U19909 ( .A1(n18420), .A2(n18416), .ZN(n18554) );
  INV_X1 U19910 ( .A(n16670), .ZN(n16651) );
  OAI22_X1 U19911 ( .A1(n18479), .A2(n16674), .B1(n18554), .B2(n16651), .ZN(
        n16652) );
  AOI211_X1 U19912 ( .C1(n18452), .C2(n16654), .A(n16653), .B(n16652), .ZN(
        n16655) );
  OAI211_X1 U19913 ( .C1(n17610), .C2(n16658), .A(n16656), .B(n16655), .ZN(
        P3_U2669) );
  AND2_X1 U19914 ( .A1(n18392), .A2(n16657), .ZN(n18565) );
  AOI22_X1 U19915 ( .A1(n16673), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n18565), .B2(
        n16670), .ZN(n16669) );
  OAI21_X1 U19916 ( .B1(n16660), .B2(n16659), .A(n16658), .ZN(n16667) );
  OAI22_X1 U19917 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16661), .B1(
        n16674), .B2(n18587), .ZN(n16666) );
  NAND2_X1 U19918 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16979) );
  NAND2_X1 U19919 ( .A1(n16662), .A2(n16979), .ZN(n16991) );
  OAI22_X1 U19920 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16664), .B1(n16663), 
        .B2(n16991), .ZN(n16665) );
  AOI211_X1 U19921 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16667), .A(
        n16666), .B(n16665), .ZN(n16668) );
  NAND2_X1 U19922 ( .A1(n16669), .A2(n16668), .ZN(P3_U2670) );
  AOI22_X1 U19923 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16671), .B1(n16670), 
        .B2(n18575), .ZN(n16677) );
  OAI21_X1 U19924 ( .B1(n16673), .B2(n16672), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16676) );
  NAND3_X1 U19925 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18556), .A3(
        n16674), .ZN(n16675) );
  NAND3_X1 U19926 ( .A1(n16677), .A2(n16676), .A3(n16675), .ZN(P3_U2671) );
  INV_X1 U19927 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16679) );
  NOR4_X1 U19928 ( .A1(n16679), .A2(n16678), .A3(n16759), .A4(n16796), .ZN(
        n16680) );
  NAND4_X1 U19929 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16715), .A4(n16680), .ZN(n16681) );
  NOR4_X1 U19930 ( .A1(n16714), .A2(n16727), .A3(n16724), .A4(n16681), .ZN(
        n16708) );
  NAND2_X1 U19931 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16708), .ZN(n16707) );
  NAND2_X1 U19932 ( .A1(n16707), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16684) );
  NAND2_X1 U19933 ( .A1(n17144), .A2(n16682), .ZN(n16683) );
  OAI22_X1 U19934 ( .A1(n16993), .A2(n16684), .B1(n16707), .B2(n16683), .ZN(
        P3_U2672) );
  AOI22_X1 U19935 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16688) );
  AOI22_X1 U19936 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16687) );
  AOI22_X1 U19937 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16686) );
  AOI22_X1 U19938 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16685) );
  NAND4_X1 U19939 ( .A1(n16688), .A2(n16687), .A3(n16686), .A4(n16685), .ZN(
        n16694) );
  AOI22_X1 U19940 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16692) );
  AOI22_X1 U19941 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16691) );
  AOI22_X1 U19942 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16690) );
  AOI22_X1 U19943 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16689) );
  NAND4_X1 U19944 ( .A1(n16692), .A2(n16691), .A3(n16690), .A4(n16689), .ZN(
        n16693) );
  NOR2_X1 U19945 ( .A1(n16694), .A2(n16693), .ZN(n16706) );
  AOI22_X1 U19946 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16705) );
  AOI22_X1 U19947 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16704) );
  AOI22_X1 U19948 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16695) );
  OAI21_X1 U19949 ( .B1(n16696), .B2(n20819), .A(n16695), .ZN(n16702) );
  AOI22_X1 U19950 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16700) );
  AOI22_X1 U19951 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16699) );
  AOI22_X1 U19952 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16698) );
  AOI22_X1 U19953 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16697) );
  NAND4_X1 U19954 ( .A1(n16700), .A2(n16699), .A3(n16698), .A4(n16697), .ZN(
        n16701) );
  AOI211_X1 U19955 ( .C1(n16934), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n16702), .B(n16701), .ZN(n16703) );
  NAND3_X1 U19956 ( .A1(n16705), .A2(n16704), .A3(n16703), .ZN(n16711) );
  NAND2_X1 U19957 ( .A1(n16712), .A2(n16711), .ZN(n16710) );
  XNOR2_X1 U19958 ( .A(n16706), .B(n16710), .ZN(n17006) );
  OAI211_X1 U19959 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16708), .A(n16707), .B(
        n16984), .ZN(n16709) );
  OAI21_X1 U19960 ( .B1(n17006), .B2(n16984), .A(n16709), .ZN(P3_U2673) );
  OAI21_X1 U19961 ( .B1(n16712), .B2(n16711), .A(n16710), .ZN(n17011) );
  OAI222_X1 U19962 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16716), .B1(
        P3_EBX_REG_29__SCAN_IN), .B2(n16715), .C1(n16714), .C2(n16713), .ZN(
        n16717) );
  OAI21_X1 U19963 ( .B1(n17011), .B2(n16984), .A(n16717), .ZN(P3_U2674) );
  OAI21_X1 U19964 ( .B1(n16722), .B2(n16719), .A(n16718), .ZN(n17020) );
  NAND3_X1 U19965 ( .A1(n16721), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n16984), 
        .ZN(n16720) );
  OAI221_X1 U19966 ( .B1(n16721), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n16984), 
        .C2(n17020), .A(n16720), .ZN(P3_U2676) );
  AOI21_X1 U19967 ( .B1(n16723), .B2(n16729), .A(n16722), .ZN(n17021) );
  NOR2_X1 U19968 ( .A1(n16724), .A2(n16728), .ZN(n16732) );
  AOI22_X1 U19969 ( .A1(n16993), .A2(n17021), .B1(n16732), .B2(n16727), .ZN(
        n16725) );
  OAI21_X1 U19970 ( .B1(n16727), .B2(n16726), .A(n16725), .ZN(P3_U2677) );
  INV_X1 U19971 ( .A(n16728), .ZN(n16737) );
  AOI21_X1 U19972 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16984), .A(n16737), .ZN(
        n16731) );
  OAI21_X1 U19973 ( .B1(n16733), .B2(n16730), .A(n16729), .ZN(n17030) );
  OAI22_X1 U19974 ( .A1(n16732), .A2(n16731), .B1(n17030), .B2(n16984), .ZN(
        P3_U2678) );
  AOI21_X1 U19975 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16984), .A(n16743), .ZN(
        n16736) );
  AOI21_X1 U19976 ( .B1(n16734), .B2(n16739), .A(n16733), .ZN(n17031) );
  INV_X1 U19977 ( .A(n17031), .ZN(n16735) );
  OAI22_X1 U19978 ( .A1(n16737), .A2(n16736), .B1(n16735), .B2(n16984), .ZN(
        P3_U2679) );
  INV_X1 U19979 ( .A(n16738), .ZN(n16758) );
  AOI21_X1 U19980 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n16984), .A(n16758), .ZN(
        n16742) );
  OAI21_X1 U19981 ( .B1(n16741), .B2(n16740), .A(n16739), .ZN(n17040) );
  OAI22_X1 U19982 ( .A1(n16743), .A2(n16742), .B1(n17040), .B2(n16984), .ZN(
        P3_U2680) );
  AOI21_X1 U19983 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n16984), .A(n16744), .ZN(
        n16757) );
  AOI22_X1 U19984 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16755) );
  AOI22_X1 U19985 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16754) );
  AOI22_X1 U19986 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16745) );
  OAI21_X1 U19987 ( .B1(n16746), .B2(n20819), .A(n16745), .ZN(n16752) );
  AOI22_X1 U19988 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16750) );
  AOI22_X1 U19989 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16749) );
  AOI22_X1 U19990 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16748) );
  AOI22_X1 U19991 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16747) );
  NAND4_X1 U19992 ( .A1(n16750), .A2(n16749), .A3(n16748), .A4(n16747), .ZN(
        n16751) );
  AOI211_X1 U19993 ( .C1(n16943), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n16752), .B(n16751), .ZN(n16753) );
  NAND3_X1 U19994 ( .A1(n16755), .A2(n16754), .A3(n16753), .ZN(n17041) );
  INV_X1 U19995 ( .A(n17041), .ZN(n16756) );
  OAI22_X1 U19996 ( .A1(n16758), .A2(n16757), .B1(n16756), .B2(n16984), .ZN(
        P3_U2681) );
  OAI21_X1 U19997 ( .B1(n16759), .B2(n16796), .A(n16984), .ZN(n16784) );
  AOI22_X1 U19998 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16763) );
  AOI22_X1 U19999 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16762) );
  AOI22_X1 U20000 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16761) );
  AOI22_X1 U20001 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16760) );
  NAND4_X1 U20002 ( .A1(n16763), .A2(n16762), .A3(n16761), .A4(n16760), .ZN(
        n16769) );
  AOI22_X1 U20003 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16767) );
  AOI22_X1 U20004 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16766) );
  AOI22_X1 U20005 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16765) );
  AOI22_X1 U20006 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16764) );
  NAND4_X1 U20007 ( .A1(n16767), .A2(n16766), .A3(n16765), .A4(n16764), .ZN(
        n16768) );
  NOR2_X1 U20008 ( .A1(n16769), .A2(n16768), .ZN(n17050) );
  OR2_X1 U20009 ( .A1(n17050), .A2(n16984), .ZN(n16770) );
  OAI221_X1 U20010 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16772), .C1(n16771), 
        .C2(n16784), .A(n16770), .ZN(P3_U2682) );
  AOI22_X1 U20011 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16776) );
  AOI22_X1 U20012 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16775) );
  AOI22_X1 U20013 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16774) );
  AOI22_X1 U20014 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16773) );
  NAND4_X1 U20015 ( .A1(n16776), .A2(n16775), .A3(n16774), .A4(n16773), .ZN(
        n16782) );
  AOI22_X1 U20016 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16780) );
  AOI22_X1 U20017 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16779) );
  AOI22_X1 U20018 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16778) );
  AOI22_X1 U20019 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16777) );
  NAND4_X1 U20020 ( .A1(n16780), .A2(n16779), .A3(n16778), .A4(n16777), .ZN(
        n16781) );
  NOR2_X1 U20021 ( .A1(n16782), .A2(n16781), .ZN(n17057) );
  NOR2_X1 U20022 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16783), .ZN(n16785) );
  OAI22_X1 U20023 ( .A1(n17057), .A2(n16984), .B1(n16785), .B2(n16784), .ZN(
        P3_U2683) );
  AOI22_X1 U20024 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16789) );
  AOI22_X1 U20025 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16788) );
  AOI22_X1 U20026 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16787) );
  AOI22_X1 U20027 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16786) );
  NAND4_X1 U20028 ( .A1(n16789), .A2(n16788), .A3(n16787), .A4(n16786), .ZN(
        n16795) );
  AOI22_X1 U20029 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16793) );
  AOI22_X1 U20030 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16792) );
  AOI22_X1 U20031 ( .A1(n11269), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16791) );
  AOI22_X1 U20032 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16790) );
  NAND4_X1 U20033 ( .A1(n16793), .A2(n16792), .A3(n16791), .A4(n16790), .ZN(
        n16794) );
  NOR2_X1 U20034 ( .A1(n16795), .A2(n16794), .ZN(n17063) );
  OAI21_X1 U20035 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16797), .A(n16796), .ZN(
        n16798) );
  AOI22_X1 U20036 ( .A1(n16993), .A2(n17063), .B1(n16798), .B2(n16984), .ZN(
        P3_U2684) );
  AOI22_X1 U20037 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16803) );
  AOI22_X1 U20038 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16932), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16802) );
  AOI22_X1 U20039 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16801) );
  AOI22_X1 U20040 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16800) );
  NAND4_X1 U20041 ( .A1(n16803), .A2(n16802), .A3(n16801), .A4(n16800), .ZN(
        n16809) );
  AOI22_X1 U20042 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16807) );
  AOI22_X1 U20043 ( .A1(n11269), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16806) );
  AOI22_X1 U20044 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16805) );
  AOI22_X1 U20045 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16804) );
  NAND4_X1 U20046 ( .A1(n16807), .A2(n16806), .A3(n16805), .A4(n16804), .ZN(
        n16808) );
  NOR2_X1 U20047 ( .A1(n16809), .A2(n16808), .ZN(n17067) );
  NAND2_X1 U20048 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16974), .ZN(n16813) );
  INV_X1 U20049 ( .A(n16990), .ZN(n16992) );
  OAI211_X1 U20050 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16811), .A(n16992), .B(
        n16810), .ZN(n16812) );
  OAI211_X1 U20051 ( .C1(n17067), .C2(n16984), .A(n16813), .B(n16812), .ZN(
        P3_U2685) );
  AOI22_X1 U20052 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9575), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n11393), .ZN(n16817) );
  AOI22_X1 U20053 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n16952), .ZN(n16816) );
  AOI22_X1 U20054 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n16926), .ZN(n16815) );
  AOI22_X1 U20055 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n16945), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n16951), .ZN(n16814) );
  NAND4_X1 U20056 ( .A1(n16817), .A2(n16816), .A3(n16815), .A4(n16814), .ZN(
        n16823) );
  AOI22_X1 U20057 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n16932), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n15502), .ZN(n16821) );
  AOI22_X1 U20058 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16927), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16820) );
  AOI22_X1 U20059 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n16881), .ZN(n16819) );
  AOI22_X1 U20060 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16818) );
  NAND4_X1 U20061 ( .A1(n16821), .A2(n16820), .A3(n16819), .A4(n16818), .ZN(
        n16822) );
  NOR2_X1 U20062 ( .A1(n16823), .A2(n16822), .ZN(n17073) );
  INV_X1 U20063 ( .A(n16824), .ZN(n16826) );
  NOR2_X1 U20064 ( .A1(n16826), .A2(n17991), .ZN(n16840) );
  OAI21_X1 U20065 ( .B1(n16840), .B2(n16974), .A(P3_EBX_REG_17__SCAN_IN), .ZN(
        n16828) );
  NAND3_X1 U20066 ( .A1(n16826), .A2(n16992), .A3(n16825), .ZN(n16827) );
  OAI211_X1 U20067 ( .C1(n17073), .C2(n16984), .A(n16828), .B(n16827), .ZN(
        P3_U2686) );
  AOI22_X1 U20068 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16832) );
  AOI22_X1 U20069 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16831) );
  AOI22_X1 U20070 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16830) );
  AOI22_X1 U20071 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16829) );
  NAND4_X1 U20072 ( .A1(n16832), .A2(n16831), .A3(n16830), .A4(n16829), .ZN(
        n16838) );
  AOI22_X1 U20073 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16836) );
  AOI22_X1 U20074 ( .A1(n16862), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16835) );
  AOI22_X1 U20075 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U20076 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16833) );
  NAND4_X1 U20077 ( .A1(n16836), .A2(n16835), .A3(n16834), .A4(n16833), .ZN(
        n16837) );
  NOR2_X1 U20078 ( .A1(n16838), .A2(n16837), .ZN(n17080) );
  OAI21_X1 U20079 ( .B1(n16839), .B2(n17991), .A(n16995), .ZN(n16860) );
  AND2_X1 U20080 ( .A1(n16995), .A2(n16839), .ZN(n16841) );
  AOI22_X1 U20081 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16860), .B1(n16841), 
        .B2(n16840), .ZN(n16842) );
  OAI21_X1 U20082 ( .B1(n17080), .B2(n16984), .A(n16842), .ZN(P3_U2687) );
  AOI22_X1 U20083 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16854) );
  AOI22_X1 U20084 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16853) );
  AOI22_X1 U20085 ( .A1(n16862), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16843) );
  OAI21_X1 U20086 ( .B1(n16844), .B2(n16966), .A(n16843), .ZN(n16851) );
  AOI22_X1 U20087 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16849) );
  AOI22_X1 U20088 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16848) );
  AOI22_X1 U20089 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16847) );
  AOI22_X1 U20090 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16846) );
  NAND4_X1 U20091 ( .A1(n16849), .A2(n16848), .A3(n16847), .A4(n16846), .ZN(
        n16850) );
  AOI211_X1 U20092 ( .C1(n16952), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n16851), .B(n16850), .ZN(n16852) );
  NAND3_X1 U20093 ( .A1(n16854), .A2(n16853), .A3(n16852), .ZN(n17082) );
  INV_X1 U20094 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20684) );
  NAND2_X1 U20095 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16978), .ZN(n16971) );
  NAND2_X1 U20096 ( .A1(n16856), .A2(n16970), .ZN(n16908) );
  OAI21_X1 U20097 ( .B1(n16858), .B2(n16908), .A(n16857), .ZN(n16859) );
  AOI22_X1 U20098 ( .A1(n16993), .A2(n17082), .B1(n16860), .B2(n16859), .ZN(
        n16861) );
  INV_X1 U20099 ( .A(n16861), .ZN(P3_U2688) );
  AOI21_X1 U20100 ( .B1(n16992), .B2(n16876), .A(n16892), .ZN(n16880) );
  INV_X1 U20101 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20102 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16873) );
  AOI22_X1 U20103 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16872) );
  AOI22_X1 U20104 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16863) );
  OAI21_X1 U20105 ( .B1(n16864), .B2(n20819), .A(n16863), .ZN(n16870) );
  AOI22_X1 U20106 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16868) );
  AOI22_X1 U20107 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20108 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16866) );
  AOI22_X1 U20109 ( .A1(n15502), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16865) );
  NAND4_X1 U20110 ( .A1(n16868), .A2(n16867), .A3(n16866), .A4(n16865), .ZN(
        n16869) );
  AOI211_X1 U20111 ( .C1(n9591), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n16870), .B(n16869), .ZN(n16871) );
  NAND3_X1 U20112 ( .A1(n16873), .A2(n16872), .A3(n16871), .ZN(n17085) );
  NOR4_X1 U20113 ( .A1(n16876), .A2(n16875), .A3(n16874), .A4(n16990), .ZN(
        n16877) );
  AOI22_X1 U20114 ( .A1(n16993), .A2(n17085), .B1(n16877), .B2(n16879), .ZN(
        n16878) );
  OAI21_X1 U20115 ( .B1(n16880), .B2(n16879), .A(n16878), .ZN(P3_U2689) );
  AOI22_X1 U20116 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16885) );
  AOI22_X1 U20117 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16884) );
  AOI22_X1 U20118 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16883) );
  AOI22_X1 U20119 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16882) );
  NAND4_X1 U20120 ( .A1(n16885), .A2(n16884), .A3(n16883), .A4(n16882), .ZN(
        n16891) );
  AOI22_X1 U20121 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11393), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U20122 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16888) );
  AOI22_X1 U20123 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20124 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16862), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16886) );
  NAND4_X1 U20125 ( .A1(n16889), .A2(n16888), .A3(n16887), .A4(n16886), .ZN(
        n16890) );
  NOR2_X1 U20126 ( .A1(n16891), .A2(n16890), .ZN(n17094) );
  INV_X1 U20127 ( .A(n16908), .ZN(n16893) );
  OAI21_X1 U20128 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16893), .A(n16892), .ZN(
        n16894) );
  OAI21_X1 U20129 ( .B1(n17094), .B2(n16984), .A(n16894), .ZN(P3_U2691) );
  AOI22_X1 U20130 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U20131 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16897) );
  AOI22_X1 U20132 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11393), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16896) );
  AOI22_X1 U20133 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16895) );
  NAND4_X1 U20134 ( .A1(n16898), .A2(n16897), .A3(n16896), .A4(n16895), .ZN(
        n16905) );
  AOI22_X1 U20135 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20136 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16899), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20137 ( .A1(n9575), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16901) );
  AOI22_X1 U20138 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16900) );
  NAND4_X1 U20139 ( .A1(n16903), .A2(n16902), .A3(n16901), .A4(n16900), .ZN(
        n16904) );
  NOR2_X1 U20140 ( .A1(n16905), .A2(n16904), .ZN(n17098) );
  NAND2_X1 U20141 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16970), .ZN(n16964) );
  OAI21_X1 U20142 ( .B1(n16907), .B2(n16964), .A(n16906), .ZN(n16909) );
  NAND3_X1 U20143 ( .A1(n16909), .A2(n16908), .A3(n16984), .ZN(n16910) );
  OAI21_X1 U20144 ( .B1(n17098), .B2(n16984), .A(n16910), .ZN(P3_U2692) );
  AOI22_X1 U20145 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11393), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16914) );
  AOI22_X1 U20146 ( .A1(n16862), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20147 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20148 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16911) );
  NAND4_X1 U20149 ( .A1(n16914), .A2(n16913), .A3(n16912), .A4(n16911), .ZN(
        n16920) );
  AOI22_X1 U20150 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20151 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16917) );
  AOI22_X1 U20152 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16916) );
  AOI22_X1 U20153 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16881), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16915) );
  NAND4_X1 U20154 ( .A1(n16918), .A2(n16917), .A3(n16916), .A4(n16915), .ZN(
        n16919) );
  NOR2_X1 U20155 ( .A1(n16920), .A2(n16919), .ZN(n17105) );
  INV_X1 U20156 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16922) );
  NOR2_X1 U20157 ( .A1(n16922), .A2(n16964), .ZN(n16963) );
  AOI21_X1 U20158 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n16963), .A(n16993), .ZN(
        n16941) );
  NOR2_X1 U20159 ( .A1(n17991), .A2(n16964), .ZN(n16961) );
  INV_X1 U20160 ( .A(n16961), .ZN(n16921) );
  NOR4_X1 U20161 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16923), .A3(n16922), .A4(
        n16921), .ZN(n16924) );
  AOI21_X1 U20162 ( .B1(n16941), .B2(P3_EBX_REG_10__SCAN_IN), .A(n16924), .ZN(
        n16925) );
  OAI21_X1 U20163 ( .B1(n17105), .B2(n16984), .A(n16925), .ZN(P3_U2693) );
  AOI22_X1 U20164 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n16899), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16931) );
  AOI22_X1 U20165 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16930) );
  AOI22_X1 U20166 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16945), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n16926), .ZN(n16929) );
  AOI22_X1 U20167 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16862), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n15502), .ZN(n16928) );
  NAND4_X1 U20168 ( .A1(n16931), .A2(n16930), .A3(n16929), .A4(n16928), .ZN(
        n16940) );
  AOI22_X1 U20169 ( .A1(n16932), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n11393), .ZN(n16938) );
  AOI22_X1 U20170 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16937) );
  AOI22_X1 U20171 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n16951), .ZN(n16936) );
  AOI22_X1 U20172 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n16933), .ZN(n16935) );
  NAND4_X1 U20173 ( .A1(n16938), .A2(n16937), .A3(n16936), .A4(n16935), .ZN(
        n16939) );
  NOR2_X1 U20174 ( .A1(n16940), .A2(n16939), .ZN(n17107) );
  OAI21_X1 U20175 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n16963), .A(n16941), .ZN(
        n16942) );
  OAI21_X1 U20176 ( .B1(n17107), .B2(n16984), .A(n16942), .ZN(P3_U2694) );
  AOI22_X1 U20177 ( .A1(n16899), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U20178 ( .A1(n16881), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9575), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20179 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16947) );
  AOI22_X1 U20180 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16946) );
  NAND4_X1 U20181 ( .A1(n16949), .A2(n16948), .A3(n16947), .A4(n16946), .ZN(
        n16960) );
  AOI22_X1 U20182 ( .A1(n16862), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16950), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U20183 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20184 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16956) );
  AOI22_X1 U20185 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15501), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16955) );
  NAND4_X1 U20186 ( .A1(n16958), .A2(n16957), .A3(n16956), .A4(n16955), .ZN(
        n16959) );
  NOR2_X1 U20187 ( .A1(n16960), .A2(n16959), .ZN(n17112) );
  OAI21_X1 U20188 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16961), .A(n16984), .ZN(
        n16962) );
  OAI22_X1 U20189 ( .A1(n17112), .A2(n16984), .B1(n16963), .B2(n16962), .ZN(
        P3_U2695) );
  OAI21_X1 U20190 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n16970), .A(n16964), .ZN(
        n16965) );
  AOI22_X1 U20191 ( .A1(n16993), .A2(n16966), .B1(n16965), .B2(n16984), .ZN(
        P3_U2696) );
  INV_X1 U20192 ( .A(n16971), .ZN(n16967) );
  OAI21_X1 U20193 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n16967), .A(n16984), .ZN(
        n16969) );
  INV_X1 U20194 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16968) );
  OAI22_X1 U20195 ( .A1(n16970), .A2(n16969), .B1(n16968), .B2(n16984), .ZN(
        P3_U2697) );
  OAI21_X1 U20196 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n16978), .A(n16971), .ZN(
        n16972) );
  AOI22_X1 U20197 ( .A1(n16993), .A2(n20785), .B1(n16972), .B2(n16984), .ZN(
        P3_U2698) );
  NOR2_X1 U20198 ( .A1(n16974), .A2(n16973), .ZN(n16975) );
  OAI21_X1 U20199 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n16975), .A(n16984), .ZN(
        n16977) );
  INV_X1 U20200 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16976) );
  OAI22_X1 U20201 ( .A1(n16978), .A2(n16977), .B1(n16976), .B2(n16984), .ZN(
        P3_U2699) );
  INV_X1 U20202 ( .A(n16979), .ZN(n16982) );
  NAND3_X1 U20203 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n16982), .A3(n16992), .ZN(
        n16983) );
  INV_X1 U20204 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16981) );
  NAND3_X1 U20205 ( .A1(n16983), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n16984), .ZN(
        n16980) );
  OAI221_X1 U20206 ( .B1(n16983), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n16984), 
        .C2(n16981), .A(n16980), .ZN(P3_U2700) );
  AOI21_X1 U20207 ( .B1(n16995), .B2(n16982), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n16987) );
  NAND2_X1 U20208 ( .A1(n16984), .A2(n16983), .ZN(n16986) );
  OAI22_X1 U20209 ( .A1(n16987), .A2(n16986), .B1(n16985), .B2(n16984), .ZN(
        P3_U2701) );
  INV_X1 U20210 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16988) );
  OAI222_X1 U20211 ( .A1(n16991), .A2(n16990), .B1(n16989), .B2(n16995), .C1(
        n16988), .C2(n16984), .ZN(P3_U2702) );
  AOI22_X1 U20212 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n16993), .B1(
        n16992), .B2(n20703), .ZN(n16994) );
  OAI21_X1 U20213 ( .B1(n16995), .B2(n20703), .A(n16994), .ZN(P3_U2703) );
  INV_X1 U20214 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17220) );
  INV_X1 U20215 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17214) );
  INV_X1 U20216 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17256) );
  NAND2_X1 U20217 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n17116) );
  NAND2_X1 U20218 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n17117) );
  INV_X1 U20219 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17226) );
  INV_X1 U20220 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17224) );
  NOR4_X1 U20221 ( .A1(n17116), .A2(n17117), .A3(n17226), .A4(n17224), .ZN(
        n16996) );
  NAND3_X1 U20222 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(n16996), .ZN(n17111) );
  NAND4_X1 U20223 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n16997)
         );
  NAND4_X1 U20224 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n16998), .ZN(n17081) );
  NAND2_X1 U20225 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .ZN(n17043) );
  NAND4_X1 U20226 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n16999)
         );
  NAND2_X1 U20227 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17037), .ZN(n17036) );
  NAND2_X1 U20228 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17033), .ZN(n17032) );
  NAND2_X1 U20229 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17022), .ZN(n17017) );
  NAND2_X1 U20230 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17007), .ZN(n17003) );
  NAND3_X1 U20231 ( .A1(n17136), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17003), 
        .ZN(n17002) );
  NAND2_X1 U20232 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17074), .ZN(n17001) );
  OAI211_X1 U20233 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17003), .A(n17002), .B(
        n17001), .ZN(P3_U2704) );
  NOR2_X2 U20234 ( .A1(n17981), .A2(n17136), .ZN(n17075) );
  AOI22_X1 U20235 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17074), .ZN(n17005) );
  OAI211_X1 U20236 ( .C1(n17007), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17136), .B(
        n17003), .ZN(n17004) );
  OAI211_X1 U20237 ( .C1(n17006), .C2(n17138), .A(n17005), .B(n17004), .ZN(
        P3_U2705) );
  AOI22_X1 U20238 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17074), .ZN(n17010) );
  AOI211_X1 U20239 ( .C1(n17220), .C2(n17013), .A(n17007), .B(n17058), .ZN(
        n17008) );
  INV_X1 U20240 ( .A(n17008), .ZN(n17009) );
  OAI211_X1 U20241 ( .C1(n17011), .C2(n17138), .A(n17010), .B(n17009), .ZN(
        P3_U2706) );
  AOI22_X1 U20242 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17075), .B1(n17146), .B2(
        n17012), .ZN(n17016) );
  OAI211_X1 U20243 ( .C1(n17014), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17136), .B(
        n17013), .ZN(n17015) );
  OAI211_X1 U20244 ( .C1(n17049), .C2(n17977), .A(n17016), .B(n17015), .ZN(
        P3_U2707) );
  AOI22_X1 U20245 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17074), .ZN(n17019) );
  OAI211_X1 U20246 ( .C1(n17022), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17136), .B(
        n17017), .ZN(n17018) );
  OAI211_X1 U20247 ( .C1(n17020), .C2(n17138), .A(n17019), .B(n17018), .ZN(
        P3_U2708) );
  AOI22_X1 U20248 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17075), .B1(n17146), .B2(
        n17021), .ZN(n17025) );
  AOI211_X1 U20249 ( .C1(n17214), .C2(n17026), .A(n17022), .B(n17058), .ZN(
        n17023) );
  INV_X1 U20250 ( .A(n17023), .ZN(n17024) );
  OAI211_X1 U20251 ( .C1(n17049), .C2(n14959), .A(n17025), .B(n17024), .ZN(
        P3_U2709) );
  AOI22_X1 U20252 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17074), .ZN(n17029) );
  OAI211_X1 U20253 ( .C1(n17027), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17136), .B(
        n17026), .ZN(n17028) );
  OAI211_X1 U20254 ( .C1(n17030), .C2(n17138), .A(n17029), .B(n17028), .ZN(
        P3_U2710) );
  AOI22_X1 U20255 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17075), .B1(n17146), .B2(
        n17031), .ZN(n17035) );
  OAI211_X1 U20256 ( .C1(n17033), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17136), .B(
        n17032), .ZN(n17034) );
  OAI211_X1 U20257 ( .C1(n17049), .C2(n17963), .A(n17035), .B(n17034), .ZN(
        P3_U2711) );
  AOI22_X1 U20258 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17074), .ZN(n17039) );
  OAI211_X1 U20259 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17037), .A(n17136), .B(
        n17036), .ZN(n17038) );
  OAI211_X1 U20260 ( .C1(n17040), .C2(n17138), .A(n17039), .B(n17038), .ZN(
        P3_U2712) );
  INV_X1 U20261 ( .A(n17075), .ZN(n17048) );
  AOI22_X1 U20262 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17074), .B1(n17146), .B2(
        n17041), .ZN(n17047) );
  INV_X1 U20263 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17200) );
  INV_X1 U20264 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17196) );
  NAND2_X1 U20265 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17068), .ZN(n17064) );
  NAND2_X1 U20266 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17059), .ZN(n17054) );
  NAND2_X1 U20267 ( .A1(n17136), .A2(n17054), .ZN(n17053) );
  OAI21_X1 U20268 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17142), .A(n17053), .ZN(
        n17045) );
  INV_X1 U20269 ( .A(n17059), .ZN(n17042) );
  NOR3_X1 U20270 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17043), .A3(n17042), .ZN(
        n17044) );
  AOI21_X1 U20271 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n17045), .A(n17044), .ZN(
        n17046) );
  OAI211_X1 U20272 ( .C1(n17987), .C2(n17048), .A(n17047), .B(n17046), .ZN(
        P3_U2713) );
  INV_X1 U20273 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17204) );
  OAI22_X1 U20274 ( .A1(n17050), .A2(n17138), .B1(n14995), .B2(n17049), .ZN(
        n17051) );
  AOI21_X1 U20275 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17075), .A(n17051), .ZN(
        n17052) );
  OAI221_X1 U20276 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17054), .C1(n17204), 
        .C2(n17053), .A(n17052), .ZN(P3_U2714) );
  AOI22_X1 U20277 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17074), .ZN(n17056) );
  OAI211_X1 U20278 ( .C1(n17059), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17136), .B(
        n17054), .ZN(n17055) );
  OAI211_X1 U20279 ( .C1(n17057), .C2(n17138), .A(n17056), .B(n17055), .ZN(
        P3_U2715) );
  AOI22_X1 U20280 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17074), .ZN(n17062) );
  AOI211_X1 U20281 ( .C1(n17200), .C2(n17064), .A(n17059), .B(n17058), .ZN(
        n17060) );
  INV_X1 U20282 ( .A(n17060), .ZN(n17061) );
  OAI211_X1 U20283 ( .C1(n17063), .C2(n17138), .A(n17062), .B(n17061), .ZN(
        P3_U2716) );
  AOI22_X1 U20284 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17074), .ZN(n17066) );
  OAI211_X1 U20285 ( .C1(n17068), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17136), .B(
        n17064), .ZN(n17065) );
  OAI211_X1 U20286 ( .C1(n17067), .C2(n17138), .A(n17066), .B(n17065), .ZN(
        P3_U2717) );
  AOI22_X1 U20287 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17074), .ZN(n17072) );
  INV_X1 U20288 ( .A(n17076), .ZN(n17070) );
  INV_X1 U20289 ( .A(n17068), .ZN(n17069) );
  OAI211_X1 U20290 ( .C1(n17070), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17136), .B(
        n17069), .ZN(n17071) );
  OAI211_X1 U20291 ( .C1(n17073), .C2(n17138), .A(n17072), .B(n17071), .ZN(
        P3_U2718) );
  AOI22_X1 U20292 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17075), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17074), .ZN(n17079) );
  OAI211_X1 U20293 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17077), .A(n17136), .B(
        n17076), .ZN(n17078) );
  OAI211_X1 U20294 ( .C1(n17080), .C2(n17138), .A(n17079), .B(n17078), .ZN(
        P3_U2719) );
  OR2_X1 U20295 ( .A1(n17991), .A2(n17081), .ZN(n17084) );
  NAND2_X1 U20296 ( .A1(n17136), .A2(n17081), .ZN(n17087) );
  AOI22_X1 U20297 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17147), .B1(n17146), .B2(
        n17082), .ZN(n17083) );
  OAI221_X1 U20298 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17084), .C1(n17256), 
        .C2(n17087), .A(n17083), .ZN(P3_U2720) );
  INV_X1 U20299 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17250) );
  INV_X1 U20300 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17245) );
  INV_X1 U20301 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17240) );
  NAND2_X1 U20302 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17114), .ZN(n17106) );
  NAND2_X1 U20303 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17102), .ZN(n17093) );
  NOR2_X1 U20304 ( .A1(n17250), .A2(n17093), .ZN(n17096) );
  NAND2_X1 U20305 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17096), .ZN(n17088) );
  INV_X1 U20306 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20307 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17147), .B1(n17146), .B2(
        n17085), .ZN(n17086) );
  OAI221_X1 U20308 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17088), .C1(n17254), 
        .C2(n17087), .A(n17086), .ZN(P3_U2721) );
  INV_X1 U20309 ( .A(n17088), .ZN(n17091) );
  AOI21_X1 U20310 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17136), .A(n17096), .ZN(
        n17090) );
  OAI222_X1 U20311 ( .A1(n17141), .A2(n17092), .B1(n17091), .B2(n17090), .C1(
        n17138), .C2(n17089), .ZN(P3_U2722) );
  INV_X1 U20312 ( .A(n17093), .ZN(n17100) );
  AOI21_X1 U20313 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17136), .A(n17100), .ZN(
        n17095) );
  OAI222_X1 U20314 ( .A1(n17141), .A2(n17097), .B1(n17096), .B2(n17095), .C1(
        n17138), .C2(n17094), .ZN(P3_U2723) );
  AOI21_X1 U20315 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17136), .A(n17102), .ZN(
        n17099) );
  OAI222_X1 U20316 ( .A1(n17141), .A2(n17101), .B1(n17100), .B2(n17099), .C1(
        n17138), .C2(n17098), .ZN(P3_U2724) );
  AOI21_X1 U20317 ( .B1(n17245), .B2(n17106), .A(n17102), .ZN(n17103) );
  AOI22_X1 U20318 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17147), .B1(n17103), .B2(
        n17136), .ZN(n17104) );
  OAI21_X1 U20319 ( .B1(n17105), .B2(n17138), .A(n17104), .ZN(P3_U2725) );
  INV_X1 U20320 ( .A(n17106), .ZN(n17109) );
  AOI21_X1 U20321 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17136), .A(n17114), .ZN(
        n17108) );
  OAI222_X1 U20322 ( .A1(n17141), .A2(n17110), .B1(n17109), .B2(n17108), .C1(
        n17138), .C2(n17107), .ZN(P3_U2726) );
  NOR2_X1 U20323 ( .A1(n17111), .A2(n17142), .ZN(n17120) );
  AOI21_X1 U20324 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17136), .A(n17120), .ZN(
        n17113) );
  OAI222_X1 U20325 ( .A1(n17141), .A2(n17115), .B1(n17114), .B2(n17113), .C1(
        n17138), .C2(n17112), .ZN(P3_U2727) );
  NOR3_X1 U20326 ( .A1(n20802), .A2(n17224), .A3(n17142), .ZN(n17135) );
  NAND2_X1 U20327 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17135), .ZN(n17134) );
  NOR2_X1 U20328 ( .A1(n17116), .A2(n17134), .ZN(n17130) );
  INV_X1 U20329 ( .A(n17130), .ZN(n17127) );
  NOR2_X1 U20330 ( .A1(n17117), .A2(n17127), .ZN(n17123) );
  AOI21_X1 U20331 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17136), .A(n17123), .ZN(
        n17119) );
  OAI222_X1 U20332 ( .A1(n17992), .A2(n17141), .B1(n17120), .B2(n17119), .C1(
        n17138), .C2(n17118), .ZN(P3_U2728) );
  AOI22_X1 U20333 ( .A1(n17130), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17136), .ZN(n17122) );
  OAI222_X1 U20334 ( .A1(n17987), .A2(n17141), .B1(n17123), .B2(n17122), .C1(
        n17138), .C2(n17121), .ZN(P3_U2729) );
  NAND3_X1 U20335 ( .A1(n17136), .A2(P3_EAX_REG_5__SCAN_IN), .A3(n17127), .ZN(
        n17126) );
  AOI22_X1 U20336 ( .A1(n17147), .A2(BUF2_REG_5__SCAN_IN), .B1(n17146), .B2(
        n17124), .ZN(n17125) );
  OAI211_X1 U20337 ( .C1(P3_EAX_REG_5__SCAN_IN), .C2(n17127), .A(n17126), .B(
        n17125), .ZN(P3_U2730) );
  INV_X1 U20338 ( .A(n17134), .ZN(n17140) );
  AOI22_X1 U20339 ( .A1(n17140), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n17136), .ZN(n17129) );
  OAI222_X1 U20340 ( .A1(n17978), .A2(n17141), .B1(n17130), .B2(n17129), .C1(
        n17138), .C2(n17128), .ZN(P3_U2731) );
  NAND3_X1 U20341 ( .A1(n17136), .A2(P3_EAX_REG_3__SCAN_IN), .A3(n17134), .ZN(
        n17133) );
  AOI22_X1 U20342 ( .A1(n17147), .A2(BUF2_REG_3__SCAN_IN), .B1(n17146), .B2(
        n17131), .ZN(n17132) );
  OAI211_X1 U20343 ( .C1(P3_EAX_REG_3__SCAN_IN), .C2(n17134), .A(n17133), .B(
        n17132), .ZN(P3_U2732) );
  AOI21_X1 U20344 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17136), .A(n17135), .ZN(
        n17139) );
  OAI222_X1 U20345 ( .A1(n20714), .A2(n17141), .B1(n17140), .B2(n17139), .C1(
        n17138), .C2(n17137), .ZN(P3_U2733) );
  OR2_X1 U20346 ( .A1(n20802), .A2(n17142), .ZN(n17150) );
  AOI21_X1 U20347 ( .B1(n17144), .B2(n20802), .A(n17143), .ZN(n17149) );
  AOI22_X1 U20348 ( .A1(n17147), .A2(BUF2_REG_1__SCAN_IN), .B1(n17146), .B2(
        n17145), .ZN(n17148) );
  OAI221_X1 U20349 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17150), .C1(n17224), 
        .C2(n17149), .A(n17148), .ZN(P3_U2734) );
  INV_X2 U20350 ( .A(n17179), .ZN(n18609) );
  NOR2_X4 U20351 ( .A1(n18609), .A2(n17177), .ZN(n17182) );
  AND2_X1 U20352 ( .A1(n17182), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20353 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20354 ( .A1(n18609), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17153) );
  OAI21_X1 U20355 ( .B1(n17222), .B2(n17168), .A(n17153), .ZN(P3_U2737) );
  AOI22_X1 U20356 ( .A1(n18609), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17154) );
  OAI21_X1 U20357 ( .B1(n17220), .B2(n17168), .A(n17154), .ZN(P3_U2738) );
  INV_X1 U20358 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20359 ( .A1(n18609), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17155) );
  OAI21_X1 U20360 ( .B1(n17218), .B2(n17168), .A(n17155), .ZN(P3_U2739) );
  INV_X1 U20361 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20362 ( .A1(n18609), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17156) );
  OAI21_X1 U20363 ( .B1(n17216), .B2(n17168), .A(n17156), .ZN(P3_U2740) );
  AOI22_X1 U20364 ( .A1(n18609), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17157) );
  OAI21_X1 U20365 ( .B1(n17214), .B2(n17168), .A(n17157), .ZN(P3_U2741) );
  INV_X1 U20366 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20367 ( .A1(n18609), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17158) );
  OAI21_X1 U20368 ( .B1(n17212), .B2(n17168), .A(n17158), .ZN(P3_U2742) );
  INV_X1 U20369 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20370 ( .A1(n18609), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17159) );
  OAI21_X1 U20371 ( .B1(n17210), .B2(n17168), .A(n17159), .ZN(P3_U2743) );
  INV_X1 U20372 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20373 ( .A1(n18609), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17160) );
  OAI21_X1 U20374 ( .B1(n17208), .B2(n17168), .A(n17160), .ZN(P3_U2744) );
  INV_X1 U20375 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U20376 ( .A1(n18609), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17161) );
  OAI21_X1 U20377 ( .B1(n17206), .B2(n17168), .A(n17161), .ZN(P3_U2745) );
  AOI22_X1 U20378 ( .A1(n18609), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17162) );
  OAI21_X1 U20379 ( .B1(n17204), .B2(n17168), .A(n17162), .ZN(P3_U2746) );
  INV_X1 U20380 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20381 ( .A1(n18609), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17163) );
  OAI21_X1 U20382 ( .B1(n17202), .B2(n17168), .A(n17163), .ZN(P3_U2747) );
  AOI22_X1 U20383 ( .A1(n18609), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17164) );
  OAI21_X1 U20384 ( .B1(n17200), .B2(n17168), .A(n17164), .ZN(P3_U2748) );
  INV_X1 U20385 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U20386 ( .A1(n18609), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17165) );
  OAI21_X1 U20387 ( .B1(n17198), .B2(n17168), .A(n17165), .ZN(P3_U2749) );
  AOI22_X1 U20388 ( .A1(n18609), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17166) );
  OAI21_X1 U20389 ( .B1(n17196), .B2(n17168), .A(n17166), .ZN(P3_U2750) );
  INV_X1 U20390 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20391 ( .A1(n18609), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17167) );
  OAI21_X1 U20392 ( .B1(n17194), .B2(n17168), .A(n17167), .ZN(P3_U2751) );
  AOI22_X1 U20393 ( .A1(n18609), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17169) );
  OAI21_X1 U20394 ( .B1(n17256), .B2(n17188), .A(n17169), .ZN(P3_U2752) );
  AOI22_X1 U20395 ( .A1(n18609), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17170) );
  OAI21_X1 U20396 ( .B1(n17254), .B2(n17188), .A(n17170), .ZN(P3_U2753) );
  INV_X1 U20397 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20398 ( .A1(n18609), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17171) );
  OAI21_X1 U20399 ( .B1(n17252), .B2(n17188), .A(n17171), .ZN(P3_U2754) );
  AOI22_X1 U20400 ( .A1(n18609), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17172) );
  OAI21_X1 U20401 ( .B1(n17250), .B2(n17188), .A(n17172), .ZN(P3_U2755) );
  INV_X1 U20402 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20403 ( .A1(n18609), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17173) );
  OAI21_X1 U20404 ( .B1(n17248), .B2(n17188), .A(n17173), .ZN(P3_U2756) );
  AOI22_X1 U20405 ( .A1(n18609), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17174) );
  OAI21_X1 U20406 ( .B1(n17245), .B2(n17188), .A(n17174), .ZN(P3_U2757) );
  INV_X1 U20407 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20408 ( .A1(n18609), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17175) );
  OAI21_X1 U20409 ( .B1(n17242), .B2(n17188), .A(n17175), .ZN(P3_U2758) );
  AOI22_X1 U20410 ( .A1(n18609), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17176) );
  OAI21_X1 U20411 ( .B1(n17240), .B2(n17188), .A(n17176), .ZN(P3_U2759) );
  INV_X1 U20412 ( .A(P3_LWORD_REG_7__SCAN_IN), .ZN(n20742) );
  AOI22_X1 U20413 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17177), .B1(n17182), .B2(
        P3_DATAO_REG_7__SCAN_IN), .ZN(n17178) );
  OAI21_X1 U20414 ( .B1(n17179), .B2(n20742), .A(n17178), .ZN(P3_U2760) );
  INV_X1 U20415 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20416 ( .A1(n18609), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17180) );
  OAI21_X1 U20417 ( .B1(n17236), .B2(n17188), .A(n17180), .ZN(P3_U2761) );
  INV_X1 U20418 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20419 ( .A1(n18609), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17181) );
  OAI21_X1 U20420 ( .B1(n17233), .B2(n17188), .A(n17181), .ZN(P3_U2762) );
  INV_X1 U20421 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20422 ( .A1(n18609), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17183) );
  OAI21_X1 U20423 ( .B1(n17230), .B2(n17188), .A(n17183), .ZN(P3_U2763) );
  INV_X1 U20424 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20425 ( .A1(n18609), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17184) );
  OAI21_X1 U20426 ( .B1(n17228), .B2(n17188), .A(n17184), .ZN(P3_U2764) );
  AOI22_X1 U20427 ( .A1(n18609), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17185) );
  OAI21_X1 U20428 ( .B1(n17226), .B2(n17188), .A(n17185), .ZN(P3_U2765) );
  AOI22_X1 U20429 ( .A1(n18609), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17186) );
  OAI21_X1 U20430 ( .B1(n17224), .B2(n17188), .A(n17186), .ZN(P3_U2766) );
  AOI22_X1 U20431 ( .A1(n18609), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17182), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17187) );
  OAI21_X1 U20432 ( .B1(n20802), .B2(n17188), .A(n17187), .ZN(P3_U2767) );
  OAI21_X4 U20433 ( .B1(n17191), .B2(n18443), .A(n17190), .ZN(n17234) );
  AOI22_X1 U20434 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17234), .ZN(n17193) );
  OAI21_X1 U20435 ( .B1(n17194), .B2(n17244), .A(n17193), .ZN(P3_U2768) );
  AOI22_X1 U20436 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17234), .ZN(n17195) );
  OAI21_X1 U20437 ( .B1(n17196), .B2(n17244), .A(n17195), .ZN(P3_U2769) );
  AOI22_X1 U20438 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17234), .ZN(n17197) );
  OAI21_X1 U20439 ( .B1(n17198), .B2(n17244), .A(n17197), .ZN(P3_U2770) );
  AOI22_X1 U20440 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17234), .ZN(n17199) );
  OAI21_X1 U20441 ( .B1(n17200), .B2(n17244), .A(n17199), .ZN(P3_U2771) );
  AOI22_X1 U20442 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17234), .ZN(n17201) );
  OAI21_X1 U20443 ( .B1(n17202), .B2(n17244), .A(n17201), .ZN(P3_U2772) );
  AOI22_X1 U20444 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17234), .ZN(n17203) );
  OAI21_X1 U20445 ( .B1(n17204), .B2(n17244), .A(n17203), .ZN(P3_U2773) );
  AOI22_X1 U20446 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17234), .ZN(n17205) );
  OAI21_X1 U20447 ( .B1(n17206), .B2(n17244), .A(n17205), .ZN(P3_U2774) );
  AOI22_X1 U20448 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17234), .ZN(n17207) );
  OAI21_X1 U20449 ( .B1(n17208), .B2(n17244), .A(n17207), .ZN(P3_U2775) );
  AOI22_X1 U20450 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17234), .ZN(n17209) );
  OAI21_X1 U20451 ( .B1(n17210), .B2(n17244), .A(n17209), .ZN(P3_U2776) );
  AOI22_X1 U20452 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17231), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17234), .ZN(n17211) );
  OAI21_X1 U20453 ( .B1(n17212), .B2(n17244), .A(n17211), .ZN(P3_U2777) );
  AOI22_X1 U20454 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17231), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17234), .ZN(n17213) );
  OAI21_X1 U20455 ( .B1(n17214), .B2(n17244), .A(n17213), .ZN(P3_U2778) );
  AOI22_X1 U20456 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20800), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17234), .ZN(n17215) );
  OAI21_X1 U20457 ( .B1(n17216), .B2(n17244), .A(n17215), .ZN(P3_U2779) );
  AOI22_X1 U20458 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17231), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17234), .ZN(n17217) );
  OAI21_X1 U20459 ( .B1(n17218), .B2(n17244), .A(n17217), .ZN(P3_U2780) );
  AOI22_X1 U20460 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17231), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17234), .ZN(n17219) );
  OAI21_X1 U20461 ( .B1(n17220), .B2(n17244), .A(n17219), .ZN(P3_U2781) );
  AOI22_X1 U20462 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17231), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17234), .ZN(n17221) );
  OAI21_X1 U20463 ( .B1(n17222), .B2(n17244), .A(n17221), .ZN(P3_U2782) );
  AOI22_X1 U20464 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17231), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17234), .ZN(n17223) );
  OAI21_X1 U20465 ( .B1(n17224), .B2(n17244), .A(n17223), .ZN(P3_U2784) );
  AOI22_X1 U20466 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17231), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17234), .ZN(n17225) );
  OAI21_X1 U20467 ( .B1(n17226), .B2(n17244), .A(n17225), .ZN(P3_U2785) );
  AOI22_X1 U20468 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17231), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17234), .ZN(n17227) );
  OAI21_X1 U20469 ( .B1(n17228), .B2(n17244), .A(n17227), .ZN(P3_U2786) );
  AOI22_X1 U20470 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17231), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17234), .ZN(n17229) );
  OAI21_X1 U20471 ( .B1(n17230), .B2(n17244), .A(n17229), .ZN(P3_U2787) );
  AOI22_X1 U20472 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17231), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17234), .ZN(n17232) );
  OAI21_X1 U20473 ( .B1(n17233), .B2(n17244), .A(n17232), .ZN(P3_U2788) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17234), .ZN(n17235) );
  OAI21_X1 U20475 ( .B1(n17236), .B2(n17244), .A(n17235), .ZN(P3_U2789) );
  AOI22_X1 U20476 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20800), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17246), .ZN(n17237) );
  OAI21_X1 U20477 ( .B1(n17238), .B2(n20742), .A(n17237), .ZN(P3_U2790) );
  AOI22_X1 U20478 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17234), .ZN(n17239) );
  OAI21_X1 U20479 ( .B1(n17240), .B2(n17244), .A(n17239), .ZN(P3_U2791) );
  AOI22_X1 U20480 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17234), .ZN(n17241) );
  OAI21_X1 U20481 ( .B1(n17242), .B2(n17244), .A(n17241), .ZN(P3_U2792) );
  AOI22_X1 U20482 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17234), .ZN(n17243) );
  OAI21_X1 U20483 ( .B1(n17245), .B2(n17244), .A(n17243), .ZN(P3_U2793) );
  AOI22_X1 U20484 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17234), .ZN(n17247) );
  OAI21_X1 U20485 ( .B1(n17248), .B2(n17244), .A(n17247), .ZN(P3_U2794) );
  AOI22_X1 U20486 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17234), .ZN(n17249) );
  OAI21_X1 U20487 ( .B1(n17250), .B2(n17244), .A(n17249), .ZN(P3_U2795) );
  AOI22_X1 U20488 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17234), .ZN(n17251) );
  OAI21_X1 U20489 ( .B1(n17252), .B2(n17244), .A(n17251), .ZN(P3_U2796) );
  AOI22_X1 U20490 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17234), .ZN(n17253) );
  OAI21_X1 U20491 ( .B1(n17254), .B2(n17244), .A(n17253), .ZN(P3_U2797) );
  AOI22_X1 U20492 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17234), .ZN(n17255) );
  OAI21_X1 U20493 ( .B1(n17256), .B2(n17244), .A(n17255), .ZN(P3_U2798) );
  OAI21_X1 U20494 ( .B1(n17257), .B2(n17624), .A(n9597), .ZN(n17258) );
  AOI21_X1 U20495 ( .B1(n17584), .B2(n16333), .A(n17258), .ZN(n17287) );
  OAI21_X1 U20496 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17399), .A(
        n17287), .ZN(n17277) );
  AOI22_X1 U20497 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17277), .B1(
        n17473), .B2(n17259), .ZN(n17273) );
  INV_X1 U20498 ( .A(n17260), .ZN(n17636) );
  NOR2_X1 U20499 ( .A1(n17638), .A2(n17292), .ZN(n17261) );
  AOI211_X1 U20500 ( .C1(n17628), .C2(n17482), .A(n17261), .B(n16215), .ZN(
        n17264) );
  INV_X1 U20501 ( .A(n17265), .ZN(n17268) );
  NAND2_X1 U20502 ( .A1(n17268), .A2(n17267), .ZN(n17269) );
  NAND2_X1 U20503 ( .A1(n9578), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17272) );
  NOR2_X1 U20504 ( .A1(n17383), .A2(n16333), .ZN(n17279) );
  OAI211_X1 U20505 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17279), .B(n17270), .ZN(n17271) );
  NAND4_X1 U20506 ( .A1(n17273), .A2(n9647), .A3(n17272), .A4(n17271), .ZN(
        P3_U2802) );
  AOI21_X1 U20507 ( .B1(n17528), .B2(n17274), .A(n9645), .ZN(n17642) );
  INV_X1 U20508 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17278) );
  OAI22_X1 U20509 ( .A1(n17852), .A2(n18526), .B1(n17460), .B2(n17275), .ZN(
        n17276) );
  AOI221_X1 U20510 ( .B1(n17279), .B2(n17278), .C1(n17277), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17276), .ZN(n17282) );
  AOI22_X1 U20511 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17292), .B1(
        n17280), .B2(n17638), .ZN(n17281) );
  OAI211_X1 U20512 ( .C1(n17642), .C2(n17529), .A(n17282), .B(n17281), .ZN(
        P3_U2803) );
  AOI21_X1 U20513 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17284), .A(
        n17283), .ZN(n17646) );
  INV_X1 U20514 ( .A(n17399), .ZN(n17289) );
  AOI21_X1 U20515 ( .B1(n17285), .B2(n18273), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17286) );
  OAI22_X1 U20516 ( .A1(n17287), .A2(n17286), .B1(n17852), .B2(n18524), .ZN(
        n17288) );
  AOI221_X1 U20517 ( .B1(n17473), .B2(n17290), .C1(n17289), .C2(n17290), .A(
        n17288), .ZN(n17294) );
  NOR2_X1 U20518 ( .A1(n17652), .A2(n17424), .ZN(n17291) );
  NOR2_X1 U20519 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17653), .ZN(
        n17643) );
  AOI22_X1 U20520 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17292), .B1(
        n17291), .B2(n17643), .ZN(n17293) );
  OAI211_X1 U20521 ( .C1(n17646), .C2(n17529), .A(n17294), .B(n17293), .ZN(
        P3_U2804) );
  AND2_X1 U20522 ( .A1(n16337), .A2(n18273), .ZN(n17329) );
  AOI211_X1 U20523 ( .C1(n17296), .C2(n17295), .A(n17582), .B(n17329), .ZN(
        n17326) );
  OAI21_X1 U20524 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17399), .A(
        n17326), .ZN(n17312) );
  AOI22_X1 U20525 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17312), .B1(
        n17473), .B2(n17297), .ZN(n17307) );
  XNOR2_X1 U20526 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17298), .ZN(
        n17661) );
  XNOR2_X1 U20527 ( .A(n17299), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17663) );
  OAI21_X1 U20528 ( .B1(n17528), .B2(n17301), .A(n17300), .ZN(n17302) );
  XNOR2_X1 U20529 ( .A(n17302), .B(n17653), .ZN(n17659) );
  OAI22_X1 U20530 ( .A1(n17628), .A2(n17663), .B1(n17529), .B2(n17659), .ZN(
        n17303) );
  AOI21_X1 U20531 ( .B1(n9600), .B2(n17661), .A(n17303), .ZN(n17306) );
  NAND2_X1 U20532 ( .A1(n9578), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17657) );
  NOR2_X1 U20533 ( .A1(n17383), .A2(n16337), .ZN(n17314) );
  OAI211_X1 U20534 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17314), .B(n17304), .ZN(n17305) );
  NAND4_X1 U20535 ( .A1(n17307), .A2(n17306), .A3(n17657), .A4(n17305), .ZN(
        P3_U2805) );
  AOI21_X1 U20536 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17309), .A(
        n17308), .ZN(n17679) );
  OAI22_X1 U20537 ( .A1(n17852), .A2(n18520), .B1(n17460), .B2(n17310), .ZN(
        n17311) );
  AOI221_X1 U20538 ( .B1(n17314), .B2(n17313), .C1(n17312), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17311), .ZN(n17317) );
  NAND2_X1 U20539 ( .A1(n17668), .A2(n17612), .ZN(n17318) );
  OAI21_X1 U20540 ( .B1(n17665), .B2(n17482), .A(n17318), .ZN(n17334) );
  NOR2_X1 U20541 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17315), .ZN(
        n17677) );
  AOI22_X1 U20542 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17334), .B1(
        n17372), .B2(n17677), .ZN(n17316) );
  OAI211_X1 U20543 ( .C1(n17679), .C2(n17529), .A(n17317), .B(n17316), .ZN(
        P3_U2806) );
  INV_X1 U20544 ( .A(n17318), .ZN(n17320) );
  NOR3_X1 U20545 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17482), .A3(
        n17767), .ZN(n17319) );
  AOI21_X1 U20546 ( .B1(n17320), .B2(n17688), .A(n17319), .ZN(n17337) );
  NOR2_X1 U20547 ( .A1(n17852), .A2(n18518), .ZN(n17683) );
  NOR2_X1 U20548 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17399), .ZN(
        n17321) );
  AOI22_X1 U20549 ( .A1(n17473), .A2(n17323), .B1(n17322), .B2(n17321), .ZN(
        n17324) );
  OAI21_X1 U20550 ( .B1(n17326), .B2(n17325), .A(n17324), .ZN(n17327) );
  AOI211_X1 U20551 ( .C1(n17329), .C2(n17328), .A(n17683), .B(n17327), .ZN(
        n17336) );
  AOI22_X1 U20552 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17528), .B1(
        n17331), .B2(n17339), .ZN(n17332) );
  NAND2_X1 U20553 ( .A1(n17330), .A2(n17332), .ZN(n17333) );
  XNOR2_X1 U20554 ( .A(n17333), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17684) );
  AOI22_X1 U20555 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17334), .B1(
        n17516), .B2(n17684), .ZN(n17335) );
  OAI211_X1 U20556 ( .C1(n17337), .C2(n17664), .A(n17336), .B(n17335), .ZN(
        P3_U2807) );
  INV_X1 U20557 ( .A(n17693), .ZN(n17680) );
  INV_X1 U20558 ( .A(n17330), .ZN(n17338) );
  AOI221_X1 U20559 ( .B1(n17340), .B2(n17339), .C1(n17680), .C2(n17339), .A(
        n17338), .ZN(n17341) );
  XNOR2_X1 U20560 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17341), .ZN(
        n17702) );
  NOR2_X1 U20561 ( .A1(n17680), .A2(n17424), .ZN(n17350) );
  NOR2_X1 U20562 ( .A1(n17612), .A2(n9600), .ZN(n17371) );
  NOR2_X1 U20563 ( .A1(n17688), .A2(n17628), .ZN(n17436) );
  AOI21_X1 U20564 ( .B1(n9600), .B2(n17767), .A(n17436), .ZN(n17422) );
  OAI21_X1 U20565 ( .B1(n17693), .B2(n17371), .A(n17422), .ZN(n17362) );
  OAI21_X1 U20566 ( .B1(n17342), .B2(n17624), .A(n9597), .ZN(n17343) );
  AOI21_X1 U20567 ( .B1(n17584), .B2(n17345), .A(n17343), .ZN(n17368) );
  OAI21_X1 U20568 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17399), .A(
        n17368), .ZN(n17356) );
  AOI22_X1 U20569 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17356), .B1(
        n17473), .B2(n17344), .ZN(n17348) );
  NOR2_X1 U20570 ( .A1(n17383), .A2(n17345), .ZN(n17357) );
  OAI211_X1 U20571 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17357), .B(n17346), .ZN(n17347) );
  OAI211_X1 U20572 ( .C1(n18516), .C2(n17852), .A(n17348), .B(n17347), .ZN(
        n17349) );
  AOI221_X1 U20573 ( .B1(n17350), .B2(n20760), .C1(n17362), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17349), .ZN(n17351) );
  OAI21_X1 U20574 ( .B1(n17529), .B2(n17702), .A(n17351), .ZN(P3_U2808) );
  NAND2_X1 U20575 ( .A1(n17708), .A2(n17352), .ZN(n17712) );
  INV_X1 U20576 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17388) );
  NOR2_X1 U20577 ( .A1(n17669), .A2(n17388), .ZN(n17703) );
  NAND2_X1 U20578 ( .A1(n17372), .A2(n17703), .ZN(n17380) );
  INV_X1 U20579 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20682) );
  AOI22_X1 U20580 ( .A1(n9578), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17473), 
        .B2(n17353), .ZN(n17354) );
  INV_X1 U20581 ( .A(n17354), .ZN(n17355) );
  AOI221_X1 U20582 ( .B1(n17357), .B2(n20682), .C1(n17356), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17355), .ZN(n17364) );
  NOR3_X1 U20583 ( .A1(n17388), .A2(n17528), .A3(n17358), .ZN(n17377) );
  INV_X1 U20584 ( .A(n17359), .ZN(n17378) );
  AOI22_X1 U20585 ( .A1(n17708), .A2(n17377), .B1(n17378), .B2(n17360), .ZN(
        n17361) );
  XNOR2_X1 U20586 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17361), .ZN(
        n17704) );
  AOI22_X1 U20587 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17362), .B1(
        n17516), .B2(n17704), .ZN(n17363) );
  OAI211_X1 U20588 ( .C1(n17712), .C2(n17380), .A(n17364), .B(n17363), .ZN(
        P3_U2809) );
  OAI221_X1 U20589 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17395), 
        .C1(n17713), .C2(n17377), .A(n17330), .ZN(n17365) );
  XNOR2_X1 U20590 ( .A(n17695), .B(n17365), .ZN(n17724) );
  AOI21_X1 U20591 ( .B1(n17366), .B2(n18273), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17367) );
  OAI22_X1 U20592 ( .A1(n17368), .A2(n17367), .B1(n17852), .B2(n18512), .ZN(
        n17369) );
  AOI221_X1 U20593 ( .B1(n17473), .B2(n17370), .C1(n17289), .C2(n17370), .A(
        n17369), .ZN(n17374) );
  INV_X1 U20594 ( .A(n17703), .ZN(n17691) );
  NOR2_X1 U20595 ( .A1(n17713), .A2(n17691), .ZN(n17716) );
  OAI21_X1 U20596 ( .B1(n17371), .B2(n17716), .A(n17422), .ZN(n17382) );
  AND2_X1 U20597 ( .A1(n17695), .A2(n17716), .ZN(n17719) );
  AOI22_X1 U20598 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17382), .B1(
        n17372), .B2(n17719), .ZN(n17373) );
  OAI211_X1 U20599 ( .C1(n17529), .C2(n17724), .A(n17374), .B(n17373), .ZN(
        P3_U2810) );
  AOI21_X1 U20600 ( .B1(n17584), .B2(n12168), .A(n17582), .ZN(n17402) );
  OAI21_X1 U20601 ( .B1(n17375), .B2(n17624), .A(n17402), .ZN(n17392) );
  AOI22_X1 U20602 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17392), .B1(
        n17473), .B2(n17376), .ZN(n17387) );
  AOI21_X1 U20603 ( .B1(n17378), .B2(n17395), .A(n17377), .ZN(n17379) );
  XNOR2_X1 U20604 ( .A(n17379), .B(n17713), .ZN(n17729) );
  OAI22_X1 U20605 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17380), .B1(
        n17729), .B2(n17529), .ZN(n17381) );
  AOI21_X1 U20606 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17382), .A(
        n17381), .ZN(n17386) );
  NAND2_X1 U20607 ( .A1(n9578), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17727) );
  NOR2_X1 U20608 ( .A1(n17383), .A2(n12168), .ZN(n17394) );
  OAI211_X1 U20609 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17394), .B(n17384), .ZN(n17385) );
  NAND4_X1 U20610 ( .A1(n17387), .A2(n17386), .A3(n17727), .A4(n17385), .ZN(
        P3_U2811) );
  NAND2_X1 U20611 ( .A1(n17737), .A2(n17388), .ZN(n17744) );
  AOI22_X1 U20612 ( .A1(n9578), .A2(P3_REIP_REG_18__SCAN_IN), .B1(n17473), 
        .B2(n17389), .ZN(n17390) );
  INV_X1 U20613 ( .A(n17390), .ZN(n17391) );
  AOI221_X1 U20614 ( .B1(n17394), .B2(n17393), .C1(n17392), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17391), .ZN(n17398) );
  OAI21_X1 U20615 ( .B1(n17737), .B2(n17424), .A(n17422), .ZN(n17407) );
  AOI21_X1 U20616 ( .B1(n17454), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17395), .ZN(n17396) );
  XNOR2_X1 U20617 ( .A(n17396), .B(n17359), .ZN(n17740) );
  AOI22_X1 U20618 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17407), .B1(
        n17516), .B2(n17740), .ZN(n17397) );
  OAI211_X1 U20619 ( .C1(n17424), .C2(n17744), .A(n17398), .B(n17397), .ZN(
        P3_U2812) );
  NAND2_X1 U20620 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17745), .ZN(
        n17751) );
  AOI21_X1 U20621 ( .B1(n18273), .B2(n17400), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17401) );
  OAI22_X1 U20622 ( .A1(n17402), .A2(n17401), .B1(n17852), .B2(n18507), .ZN(
        n17403) );
  AOI21_X1 U20623 ( .B1(n17404), .B2(n17614), .A(n17403), .ZN(n17409) );
  OAI21_X1 U20624 ( .B1(n17406), .B2(n17745), .A(n17405), .ZN(n17749) );
  AOI22_X1 U20625 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17407), .B1(
        n17516), .B2(n17749), .ZN(n17408) );
  OAI211_X1 U20626 ( .C1(n17424), .C2(n17751), .A(n17409), .B(n17408), .ZN(
        P3_U2813) );
  NAND2_X1 U20627 ( .A1(n17454), .A2(n17430), .ZN(n17514) );
  OAI22_X1 U20628 ( .A1(n17454), .A2(n17411), .B1(n17514), .B2(n17410), .ZN(
        n17412) );
  XNOR2_X1 U20629 ( .A(n17423), .B(n17412), .ZN(n17759) );
  NAND3_X1 U20630 ( .A1(n17413), .A2(n16492), .A3(n17471), .ZN(n17426) );
  OAI21_X1 U20631 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17414), .ZN(n17419) );
  AOI21_X1 U20632 ( .B1(n17584), .B2(n17415), .A(n17582), .ZN(n17441) );
  OAI21_X1 U20633 ( .B1(n17416), .B2(n17624), .A(n17441), .ZN(n17429) );
  AOI22_X1 U20634 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17429), .B1(
        n17473), .B2(n17417), .ZN(n17418) );
  NAND2_X1 U20635 ( .A1(n9578), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17761) );
  OAI211_X1 U20636 ( .C1(n17426), .C2(n17419), .A(n17418), .B(n17761), .ZN(
        n17420) );
  AOI21_X1 U20637 ( .B1(n17516), .B2(n17759), .A(n17420), .ZN(n17421) );
  OAI221_X1 U20638 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17424), 
        .C1(n17423), .C2(n17422), .A(n17421), .ZN(P3_U2814) );
  NOR2_X1 U20639 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17446), .ZN(
        n17770) );
  NAND2_X1 U20640 ( .A1(n9600), .A2(n17767), .ZN(n17439) );
  NOR2_X1 U20641 ( .A1(n17852), .A2(n18502), .ZN(n17428) );
  OAI22_X1 U20642 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17426), .B1(
        n17425), .B2(n17460), .ZN(n17427) );
  AOI211_X1 U20643 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17429), .A(
        n17428), .B(n17427), .ZN(n17438) );
  INV_X1 U20644 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17790) );
  NAND4_X1 U20645 ( .A1(n17810), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n17430), .ZN(n17431) );
  AOI22_X1 U20646 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17528), .B1(
        n17432), .B2(n17431), .ZN(n17433) );
  OAI21_X1 U20647 ( .B1(n17790), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17433), .ZN(n17434) );
  XOR2_X1 U20648 ( .A(n17434), .B(n17435), .Z(n17764) );
  NAND2_X1 U20649 ( .A1(n17440), .A2(n17435), .ZN(n17773) );
  AOI22_X1 U20650 ( .A1(n17516), .A2(n17764), .B1(n17436), .B2(n17773), .ZN(
        n17437) );
  OAI211_X1 U20651 ( .C1(n17770), .C2(n17439), .A(n17438), .B(n17437), .ZN(
        P3_U2815) );
  OAI221_X1 U20652 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17800), .A(n17440), .ZN(
        n17797) );
  NAND2_X1 U20653 ( .A1(n18273), .A2(n16492), .ZN(n17487) );
  AOI221_X1 U20654 ( .B1(n17443), .B2(n17442), .C1(n17487), .C2(n17442), .A(
        n17441), .ZN(n17444) );
  NOR2_X1 U20655 ( .A1(n17852), .A2(n18501), .ZN(n17792) );
  AOI211_X1 U20656 ( .C1(n17445), .C2(n17614), .A(n17444), .B(n17792), .ZN(
        n17450) );
  NOR2_X1 U20657 ( .A1(n17807), .A2(n17455), .ZN(n17765) );
  INV_X1 U20658 ( .A(n17765), .ZN(n17782) );
  AOI221_X1 U20659 ( .B1(n17466), .B2(n17790), .C1(n17782), .C2(n17790), .A(
        n17446), .ZN(n17794) );
  INV_X1 U20660 ( .A(n17514), .ZN(n17494) );
  AOI21_X1 U20661 ( .B1(n17494), .B2(n17765), .A(n17447), .ZN(n17448) );
  XNOR2_X1 U20662 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17448), .ZN(
        n17793) );
  AOI22_X1 U20663 ( .A1(n9600), .A2(n17794), .B1(n17516), .B2(n17793), .ZN(
        n17449) );
  OAI211_X1 U20664 ( .C1(n17628), .C2(n17797), .A(n17450), .B(n17449), .ZN(
        P3_U2816) );
  AND2_X1 U20665 ( .A1(n17492), .A2(n17451), .ZN(n17469) );
  OAI22_X1 U20666 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17454), .B1(
        n17452), .B2(n17807), .ZN(n17453) );
  OAI21_X1 U20667 ( .B1(n17454), .B2(n17469), .A(n17453), .ZN(n17456) );
  XNOR2_X1 U20668 ( .A(n17456), .B(n17455), .ZN(n17806) );
  AOI21_X1 U20669 ( .B1(n17584), .B2(n17457), .A(n17582), .ZN(n17458) );
  OAI21_X1 U20670 ( .B1(n17459), .B2(n17624), .A(n17458), .ZN(n17474) );
  INV_X1 U20671 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20814) );
  NOR2_X1 U20672 ( .A1(n17852), .A2(n20814), .ZN(n17465) );
  OAI211_X1 U20673 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n16492), .B(n17471), .ZN(n17462) );
  OAI22_X1 U20674 ( .A1(n17463), .A2(n17462), .B1(n17461), .B2(n17460), .ZN(
        n17464) );
  AOI211_X1 U20675 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17474), .A(
        n17465), .B(n17464), .ZN(n17468) );
  NOR2_X1 U20676 ( .A1(n17807), .A2(n17466), .ZN(n17799) );
  OAI22_X1 U20677 ( .A1(n17800), .A2(n17628), .B1(n17799), .B2(n17482), .ZN(
        n17478) );
  NOR2_X1 U20678 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17807), .ZN(
        n17798) );
  AOI22_X1 U20679 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17478), .B1(
        n17798), .B2(n17498), .ZN(n17467) );
  OAI211_X1 U20680 ( .C1(n17529), .C2(n17806), .A(n17468), .B(n17467), .ZN(
        P3_U2817) );
  AOI21_X1 U20681 ( .B1(n17494), .B2(n17810), .A(n17469), .ZN(n17470) );
  XOR2_X1 U20682 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17470), .Z(
        n17817) );
  NAND2_X1 U20683 ( .A1(n16492), .A2(n17471), .ZN(n17476) );
  AOI22_X1 U20684 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17474), .B1(
        n17473), .B2(n17472), .ZN(n17475) );
  NAND2_X1 U20685 ( .A1(n9578), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17815) );
  OAI211_X1 U20686 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17476), .A(
        n17475), .B(n17815), .ZN(n17477) );
  AOI21_X1 U20687 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17478), .A(
        n17477), .ZN(n17480) );
  NAND3_X1 U20688 ( .A1(n17810), .A2(n9954), .A3(n17498), .ZN(n17479) );
  OAI211_X1 U20689 ( .C1(n17817), .C2(n17529), .A(n17480), .B(n17479), .ZN(
        P3_U2818) );
  OAI22_X1 U20690 ( .A1(n17824), .A2(n17482), .B1(n17628), .B2(n17481), .ZN(
        n17517) );
  AOI21_X1 U20691 ( .B1(n17827), .B2(n17498), .A(n17517), .ZN(n17501) );
  NAND3_X1 U20692 ( .A1(n18273), .A2(n17535), .A3(n16551), .ZN(n17509) );
  NOR2_X1 U20693 ( .A1(n17508), .A2(n17509), .ZN(n17507) );
  NAND2_X1 U20694 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17507), .ZN(
        n17505) );
  OAI21_X1 U20695 ( .B1(n17619), .B2(n17483), .A(n17505), .ZN(n17486) );
  OAI22_X1 U20696 ( .A1(n17607), .A2(n17484), .B1(n17852), .B2(n18497), .ZN(
        n17485) );
  AOI21_X1 U20697 ( .B1(n17487), .B2(n17486), .A(n17485), .ZN(n17491) );
  OAI21_X1 U20698 ( .B1(n17827), .B2(n17514), .A(n17488), .ZN(n17489) );
  XNOR2_X1 U20699 ( .A(n17489), .B(n17492), .ZN(n17831) );
  NOR2_X1 U20700 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17827), .ZN(
        n17830) );
  AOI22_X1 U20701 ( .A1(n17516), .A2(n17831), .B1(n17830), .B2(n17498), .ZN(
        n17490) );
  OAI211_X1 U20702 ( .C1(n17501), .C2(n17492), .A(n17491), .B(n17490), .ZN(
        P3_U2819) );
  AOI21_X1 U20703 ( .B1(n17494), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17493), .ZN(n17495) );
  XNOR2_X1 U20704 ( .A(n17495), .B(n17838), .ZN(n17841) );
  INV_X1 U20705 ( .A(n17507), .ZN(n17496) );
  OAI21_X1 U20706 ( .B1(n17619), .B2(n17497), .A(n17496), .ZN(n17504) );
  NOR2_X1 U20707 ( .A1(n17852), .A2(n18495), .ZN(n17503) );
  AOI21_X1 U20708 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17498), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17500) );
  OAI22_X1 U20709 ( .A1(n17501), .A2(n17500), .B1(n17607), .B2(n17499), .ZN(
        n17502) );
  AOI211_X1 U20710 ( .C1(n17505), .C2(n17504), .A(n17503), .B(n17502), .ZN(
        n17506) );
  OAI21_X1 U20711 ( .B1(n17841), .B2(n17529), .A(n17506), .ZN(P3_U2820) );
  AOI211_X1 U20712 ( .C1(n17509), .C2(n17508), .A(n17619), .B(n17507), .ZN(
        n17511) );
  NOR2_X1 U20713 ( .A1(n17852), .A2(n18493), .ZN(n17510) );
  AOI211_X1 U20714 ( .C1(n17512), .C2(n17614), .A(n17511), .B(n17510), .ZN(
        n17519) );
  NAND2_X1 U20715 ( .A1(n17514), .A2(n17513), .ZN(n17515) );
  XOR2_X1 U20716 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n17515), .Z(
        n17849) );
  AOI22_X1 U20717 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17517), .B1(
        n17516), .B2(n17849), .ZN(n17518) );
  OAI211_X1 U20718 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17520), .A(
        n17519), .B(n17518), .ZN(P3_U2821) );
  AOI21_X1 U20719 ( .B1(n17584), .B2(n17521), .A(n17582), .ZN(n17547) );
  INV_X1 U20720 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18491) );
  NOR2_X1 U20721 ( .A1(n17852), .A2(n18491), .ZN(n17860) );
  NAND2_X1 U20722 ( .A1(n17535), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17522) );
  AOI211_X1 U20723 ( .C1(n17534), .C2(n17522), .A(n16551), .B(n17995), .ZN(
        n17523) );
  AOI211_X1 U20724 ( .C1(n17866), .C2(n9600), .A(n17860), .B(n17523), .ZN(
        n17533) );
  AOI21_X1 U20725 ( .B1(n17526), .B2(n17862), .A(n17525), .ZN(n17864) );
  OAI21_X1 U20726 ( .B1(n17866), .B2(n17528), .A(n17527), .ZN(n17869) );
  OAI22_X1 U20727 ( .A1(n17607), .A2(n17530), .B1(n17529), .B2(n17869), .ZN(
        n17531) );
  AOI21_X1 U20728 ( .B1(n17612), .B2(n17864), .A(n17531), .ZN(n17532) );
  OAI211_X1 U20729 ( .C1(n17547), .C2(n17534), .A(n17533), .B(n17532), .ZN(
        P3_U2822) );
  NAND2_X1 U20730 ( .A1(n18273), .A2(n17535), .ZN(n17539) );
  NAND2_X1 U20731 ( .A1(n17537), .A2(n17536), .ZN(n17538) );
  XNOR2_X1 U20732 ( .A(n17538), .B(n17874), .ZN(n17879) );
  OAI22_X1 U20733 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17539), .B1(
        n17628), .B2(n17879), .ZN(n17540) );
  AOI21_X1 U20734 ( .B1(n9578), .B2(P3_REIP_REG_7__SCAN_IN), .A(n17540), .ZN(
        n17545) );
  AOI21_X1 U20735 ( .B1(n17874), .B2(n17542), .A(n17541), .ZN(n17877) );
  AOI22_X1 U20736 ( .A1(n9599), .A2(n17877), .B1(n17543), .B2(n17614), .ZN(
        n17544) );
  OAI211_X1 U20737 ( .C1(n17547), .C2(n17546), .A(n17545), .B(n17544), .ZN(
        P3_U2823) );
  AOI21_X1 U20738 ( .B1(n17858), .B2(n17549), .A(n17548), .ZN(n17883) );
  NOR2_X1 U20739 ( .A1(n17995), .A2(n16599), .ZN(n17550) );
  AOI22_X1 U20740 ( .A1(n17612), .A2(n17883), .B1(n17550), .B2(n17555), .ZN(
        n17559) );
  AOI21_X1 U20741 ( .B1(n17553), .B2(n17552), .A(n17551), .ZN(n17880) );
  OAI21_X1 U20742 ( .B1(n16599), .B2(n17995), .A(n17554), .ZN(n17571) );
  OAI22_X1 U20743 ( .A1(n17607), .A2(n17556), .B1(n17555), .B2(n17571), .ZN(
        n17557) );
  AOI21_X1 U20744 ( .B1(n9599), .B2(n17880), .A(n17557), .ZN(n17558) );
  OAI211_X1 U20745 ( .C1(n17852), .C2(n18487), .A(n17559), .B(n17558), .ZN(
        P3_U2824) );
  AOI21_X1 U20746 ( .B1(n17560), .B2(n9597), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17572) );
  AOI21_X1 U20747 ( .B1(n17563), .B2(n17562), .A(n17561), .ZN(n17888) );
  AOI22_X1 U20748 ( .A1(n17612), .A2(n17888), .B1(n9578), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17570) );
  AOI21_X1 U20749 ( .B1(n17564), .B2(n17566), .A(n17565), .ZN(n17567) );
  XNOR2_X1 U20750 ( .A(n17567), .B(n17890), .ZN(n17887) );
  AOI22_X1 U20751 ( .A1(n9599), .A2(n17887), .B1(n17568), .B2(n17614), .ZN(
        n17569) );
  OAI211_X1 U20752 ( .C1(n17572), .C2(n17571), .A(n17570), .B(n17569), .ZN(
        P3_U2825) );
  OAI21_X1 U20753 ( .B1(n17575), .B2(n17574), .A(n17573), .ZN(n17576) );
  XNOR2_X1 U20754 ( .A(n17576), .B(n11288), .ZN(n17905) );
  AOI22_X1 U20755 ( .A1(n9578), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18273), .B2(
        n17577), .ZN(n17589) );
  OAI21_X1 U20756 ( .B1(n17580), .B2(n17579), .A(n17578), .ZN(n17581) );
  XNOR2_X1 U20757 ( .A(n17581), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17894) );
  AOI21_X1 U20758 ( .B1(n17584), .B2(n17583), .A(n17582), .ZN(n17599) );
  OAI22_X1 U20759 ( .A1(n17607), .A2(n17586), .B1(n17585), .B2(n17599), .ZN(
        n17587) );
  AOI21_X1 U20760 ( .B1(n9599), .B2(n17894), .A(n17587), .ZN(n17588) );
  OAI211_X1 U20761 ( .C1(n17628), .C2(n17905), .A(n17589), .B(n17588), .ZN(
        P3_U2826) );
  AOI21_X1 U20762 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n9597), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17600) );
  AOI21_X1 U20763 ( .B1(n17592), .B2(n17591), .A(n17590), .ZN(n17907) );
  AOI22_X1 U20764 ( .A1(n9599), .A2(n17907), .B1(n9578), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17598) );
  AOI21_X1 U20765 ( .B1(n17595), .B2(n17594), .A(n17593), .ZN(n17908) );
  AOI22_X1 U20766 ( .A1(n17612), .A2(n17908), .B1(n17596), .B2(n17614), .ZN(
        n17597) );
  OAI211_X1 U20767 ( .C1(n17600), .C2(n17599), .A(n17598), .B(n17597), .ZN(
        P3_U2827) );
  AOI21_X1 U20768 ( .B1(n17603), .B2(n17602), .A(n17601), .ZN(n17917) );
  NOR2_X1 U20769 ( .A1(n17852), .A2(n18479), .ZN(n17925) );
  XNOR2_X1 U20770 ( .A(n17605), .B(n17604), .ZN(n17927) );
  OAI22_X1 U20771 ( .A1(n17607), .A2(n17606), .B1(n17627), .B2(n17927), .ZN(
        n17608) );
  AOI211_X1 U20772 ( .C1(n17612), .C2(n17917), .A(n17925), .B(n17608), .ZN(
        n17609) );
  OAI221_X1 U20773 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17995), .C1(
        n17610), .C2(n9597), .A(n17609), .ZN(P3_U2828) );
  OAI21_X1 U20774 ( .B1(n17622), .B2(n11452), .A(n17611), .ZN(n17928) );
  AOI22_X1 U20775 ( .A1(n17612), .A2(n17928), .B1(n9578), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17617) );
  AOI21_X1 U20776 ( .B1(n11452), .B2(n17620), .A(n17613), .ZN(n17933) );
  AOI22_X1 U20777 ( .A1(n9599), .A2(n17933), .B1(n17618), .B2(n17614), .ZN(
        n17616) );
  OAI211_X1 U20778 ( .C1(n17619), .C2(n17618), .A(n17617), .B(n17616), .ZN(
        P3_U2829) );
  INV_X1 U20779 ( .A(n17620), .ZN(n17621) );
  NOR2_X1 U20780 ( .A1(n17622), .A2(n17621), .ZN(n17629) );
  INV_X1 U20781 ( .A(n17629), .ZN(n17948) );
  NAND3_X1 U20782 ( .A1(n18553), .A2(n17624), .A3(n9597), .ZN(n17625) );
  AOI22_X1 U20783 ( .A1(n9578), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17625), .ZN(n17626) );
  OAI221_X1 U20784 ( .B1(n17629), .B2(n17628), .C1(n17948), .C2(n17627), .A(
        n17626), .ZN(P3_U2830) );
  AOI22_X1 U20785 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17936), .B1(
        n9578), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n17641) );
  NOR3_X1 U20786 ( .A1(n17681), .A2(n17652), .A3(n17630), .ZN(n17639) );
  NOR2_X1 U20787 ( .A1(n18403), .A2(n18395), .ZN(n17919) );
  NOR2_X1 U20788 ( .A1(n9569), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17921) );
  NOR2_X1 U20789 ( .A1(n17921), .A2(n17631), .ZN(n17633) );
  OAI211_X1 U20790 ( .C1(n17919), .C2(n17633), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17632), .ZN(n17655) );
  NOR2_X1 U20791 ( .A1(n17634), .A2(n17655), .ZN(n17635) );
  INV_X1 U20792 ( .A(n17859), .ZN(n17758) );
  OAI222_X1 U20793 ( .A1(n17823), .A2(n17637), .B1(n9776), .B2(n17636), .C1(
        n17635), .C2(n17758), .ZN(n17645) );
  OAI221_X1 U20794 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17639), 
        .C1(n17638), .C2(n17645), .A(n9564), .ZN(n17640) );
  OAI211_X1 U20795 ( .C1(n17642), .C2(n17870), .A(n17641), .B(n17640), .ZN(
        P3_U2835) );
  NOR2_X1 U20796 ( .A1(n17681), .A2(n17652), .ZN(n17644) );
  AOI22_X1 U20797 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17645), .B1(
        n17644), .B2(n17643), .ZN(n17650) );
  INV_X1 U20798 ( .A(n17646), .ZN(n17647) );
  AOI22_X1 U20799 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17936), .B1(
        n17850), .B2(n17647), .ZN(n17649) );
  NAND2_X1 U20800 ( .A1(n9578), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17648) );
  OAI211_X1 U20801 ( .C1(n17650), .C2(n9563), .A(n17649), .B(n17648), .ZN(
        P3_U2836) );
  INV_X1 U20802 ( .A(n17651), .ZN(n17654) );
  AOI221_X1 U20803 ( .B1(n17654), .B2(n17653), .C1(n17652), .C2(n17653), .A(
        n9563), .ZN(n17656) );
  AOI22_X1 U20804 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17936), .B1(
        n17656), .B2(n17655), .ZN(n17658) );
  OAI211_X1 U20805 ( .C1(n17659), .C2(n17870), .A(n17658), .B(n17657), .ZN(
        n17660) );
  AOI21_X1 U20806 ( .B1(n17865), .B2(n17661), .A(n17660), .ZN(n17662) );
  OAI21_X1 U20807 ( .B1(n17939), .B2(n17663), .A(n17662), .ZN(P3_U2837) );
  NOR2_X1 U20808 ( .A1(n17852), .A2(n18520), .ZN(n17676) );
  NOR3_X1 U20809 ( .A1(n17921), .A2(n17734), .A3(n17664), .ZN(n17666) );
  OAI22_X1 U20810 ( .A1(n17919), .A2(n17666), .B1(n17665), .B2(n17823), .ZN(
        n17667) );
  AOI211_X1 U20811 ( .C1(n18439), .C2(n17668), .A(n17936), .B(n17667), .ZN(
        n17674) );
  NOR2_X1 U20812 ( .A1(n17669), .A2(n17692), .ZN(n17736) );
  OAI221_X1 U20813 ( .B1(n18429), .B2(n17670), .C1(n18429), .C2(n17736), .A(
        n17674), .ZN(n17671) );
  OAI21_X1 U20814 ( .B1(n17672), .B2(n17671), .A(n17852), .ZN(n17687) );
  AOI211_X1 U20815 ( .C1(n17758), .C2(n17674), .A(n17673), .B(n17687), .ZN(
        n17675) );
  AOI211_X1 U20816 ( .C1(n17677), .C2(n17720), .A(n17676), .B(n17675), .ZN(
        n17678) );
  OAI21_X1 U20817 ( .B1(n17679), .B2(n17870), .A(n17678), .ZN(P3_U2838) );
  NOR2_X1 U20818 ( .A1(n17681), .A2(n17680), .ZN(n17699) );
  OAI221_X1 U20819 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17699), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17900), .A(n17682), .ZN(
        n17686) );
  AOI21_X1 U20820 ( .B1(n17684), .B2(n17850), .A(n17683), .ZN(n17685) );
  OAI21_X1 U20821 ( .B1(n17687), .B2(n17686), .A(n17685), .ZN(P3_U2839) );
  AOI22_X1 U20822 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17936), .B1(
        n9578), .B2(P3_REIP_REG_22__SCAN_IN), .ZN(n17701) );
  NOR2_X1 U20823 ( .A1(n17688), .A2(n9776), .ZN(n17774) );
  AOI21_X1 U20824 ( .B1(n17768), .B2(n17767), .A(n17774), .ZN(n17705) );
  NOR2_X1 U20825 ( .A1(n18439), .A2(n17768), .ZN(n17818) );
  AOI21_X1 U20826 ( .B1(n17689), .B2(n17716), .A(n17942), .ZN(n17690) );
  AOI221_X1 U20827 ( .B1(n17692), .B2(n18411), .C1(n17691), .C2(n18411), .A(
        n17690), .ZN(n17714) );
  OAI21_X1 U20828 ( .B1(n17693), .B2(n17818), .A(n17714), .ZN(n17694) );
  AOI21_X1 U20829 ( .B1(n18403), .B2(n17695), .A(n17694), .ZN(n17707) );
  NAND2_X1 U20830 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17708), .ZN(
        n17696) );
  AOI21_X1 U20831 ( .B1(n17753), .B2(n17703), .A(n9569), .ZN(n17706) );
  AOI211_X1 U20832 ( .C1(n17859), .C2(n17696), .A(n17706), .B(n20760), .ZN(
        n17697) );
  NAND3_X1 U20833 ( .A1(n17705), .A2(n17707), .A3(n17697), .ZN(n17698) );
  OAI211_X1 U20834 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17699), .A(
        n9564), .B(n17698), .ZN(n17700) );
  OAI211_X1 U20835 ( .C1(n17702), .C2(n17870), .A(n17701), .B(n17700), .ZN(
        P3_U2840) );
  NAND2_X1 U20836 ( .A1(n17720), .A2(n17703), .ZN(n17726) );
  AOI22_X1 U20837 ( .A1(n9578), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17850), 
        .B2(n17704), .ZN(n17711) );
  NOR2_X1 U20838 ( .A1(n18411), .A2(n18395), .ZN(n17935) );
  NAND2_X1 U20839 ( .A1(n9564), .A2(n17705), .ZN(n17752) );
  NOR2_X1 U20840 ( .A1(n17706), .A2(n17752), .ZN(n17715) );
  OAI211_X1 U20841 ( .C1(n17708), .C2(n17935), .A(n17715), .B(n17707), .ZN(
        n17709) );
  NAND3_X1 U20842 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17852), .A3(
        n17709), .ZN(n17710) );
  OAI211_X1 U20843 ( .C1(n17726), .C2(n17712), .A(n17711), .B(n17710), .ZN(
        P3_U2841) );
  NAND2_X1 U20844 ( .A1(n17713), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17718) );
  OAI211_X1 U20845 ( .C1(n17716), .C2(n17818), .A(n17715), .B(n17714), .ZN(
        n17717) );
  NAND2_X1 U20846 ( .A1(n17852), .A2(n17717), .ZN(n17725) );
  OAI21_X1 U20847 ( .B1(n17935), .B2(n17718), .A(n17725), .ZN(n17721) );
  AOI22_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17721), .B1(
        n17720), .B2(n17719), .ZN(n17723) );
  NAND2_X1 U20849 ( .A1(n9578), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17722) );
  OAI211_X1 U20850 ( .C1(n17724), .C2(n17870), .A(n17723), .B(n17722), .ZN(
        P3_U2842) );
  MUX2_X1 U20851 ( .A(n17726), .B(n17725), .S(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(n17728) );
  OAI211_X1 U20852 ( .C1(n17729), .C2(n17870), .A(n17728), .B(n17727), .ZN(
        P3_U2843) );
  INV_X1 U20853 ( .A(n17730), .ZN(n17898) );
  OAI22_X1 U20854 ( .A1(n18429), .A2(n17913), .B1(n17914), .B2(n17898), .ZN(
        n17906) );
  INV_X1 U20855 ( .A(n17906), .ZN(n17854) );
  NOR2_X1 U20856 ( .A1(n17854), .A2(n17731), .ZN(n17766) );
  NOR2_X1 U20857 ( .A1(n17766), .A2(n17732), .ZN(n17812) );
  NAND2_X1 U20858 ( .A1(n17733), .A2(n17848), .ZN(n17763) );
  NOR2_X1 U20859 ( .A1(n17921), .A2(n17734), .ZN(n17735) );
  AOI21_X1 U20860 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17735), .A(
        n17919), .ZN(n17739) );
  OAI22_X1 U20861 ( .A1(n17737), .A2(n17818), .B1(n17736), .B2(n18429), .ZN(
        n17738) );
  NOR3_X1 U20862 ( .A1(n17739), .A2(n17752), .A3(n17738), .ZN(n17746) );
  AOI221_X1 U20863 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17746), 
        .C1(n17919), .C2(n17746), .A(n9578), .ZN(n17741) );
  AOI22_X1 U20864 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17741), .B1(
        n17850), .B2(n17740), .ZN(n17743) );
  NAND2_X1 U20865 ( .A1(n9578), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17742) );
  OAI211_X1 U20866 ( .C1(n17744), .C2(n17763), .A(n17743), .B(n17742), .ZN(
        P3_U2844) );
  NOR2_X1 U20867 ( .A1(n17852), .A2(n18507), .ZN(n17748) );
  NOR3_X1 U20868 ( .A1(n9578), .A2(n17746), .A3(n17745), .ZN(n17747) );
  AOI211_X1 U20869 ( .C1(n17850), .C2(n17749), .A(n17748), .B(n17747), .ZN(
        n17750) );
  OAI21_X1 U20870 ( .B1(n17763), .B2(n17751), .A(n17750), .ZN(P3_U2845) );
  INV_X1 U20871 ( .A(n17752), .ZN(n17757) );
  NOR2_X1 U20872 ( .A1(n17780), .A2(n18429), .ZN(n17820) );
  NAND2_X1 U20873 ( .A1(n18403), .A2(n17783), .ZN(n17834) );
  OAI211_X1 U20874 ( .C1(n17753), .C2(n9569), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17834), .ZN(n17754) );
  AOI211_X1 U20875 ( .C1(n17756), .C2(n17755), .A(n17820), .B(n17754), .ZN(
        n17772) );
  AOI221_X1 U20876 ( .B1(n17758), .B2(n17757), .C1(n17772), .C2(n17757), .A(
        n9578), .ZN(n17760) );
  AOI22_X1 U20877 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17760), .B1(
        n17850), .B2(n17759), .ZN(n17762) );
  OAI211_X1 U20878 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17763), .A(
        n17762), .B(n17761), .ZN(P3_U2846) );
  INV_X1 U20879 ( .A(n17764), .ZN(n17778) );
  AOI22_X1 U20880 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17936), .B1(
        n9578), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n17777) );
  AND2_X1 U20881 ( .A1(n17766), .A2(n17765), .ZN(n17779) );
  AOI21_X1 U20882 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17779), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17771) );
  NAND2_X1 U20883 ( .A1(n17768), .A2(n17767), .ZN(n17769) );
  OAI22_X1 U20884 ( .A1(n17772), .A2(n17771), .B1(n17770), .B2(n17769), .ZN(
        n17775) );
  OAI221_X1 U20885 ( .B1(n17775), .B2(n17774), .C1(n17775), .C2(n17773), .A(
        n9564), .ZN(n17776) );
  OAI211_X1 U20886 ( .C1(n17870), .C2(n17778), .A(n17777), .B(n17776), .ZN(
        P3_U2847) );
  INV_X1 U20887 ( .A(n17779), .ZN(n17788) );
  AOI21_X1 U20888 ( .B1(n17781), .B2(n17780), .A(n18429), .ZN(n17786) );
  OAI21_X1 U20889 ( .B1(n17783), .B2(n17782), .A(n18403), .ZN(n17784) );
  OAI21_X1 U20890 ( .B1(n17807), .B2(n17842), .A(n18395), .ZN(n17802) );
  OAI211_X1 U20891 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n17935), .A(
        n17784), .B(n17802), .ZN(n17785) );
  NOR2_X1 U20892 ( .A1(n17786), .A2(n17785), .ZN(n17787) );
  MUX2_X1 U20893 ( .A(n17788), .B(n17787), .S(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n17789) );
  OAI22_X1 U20894 ( .A1(n17790), .A2(n17900), .B1(n9563), .B2(n17789), .ZN(
        n17791) );
  AOI211_X1 U20895 ( .C1(n17850), .C2(n17793), .A(n17792), .B(n17791), .ZN(
        n17796) );
  NAND2_X1 U20896 ( .A1(n17865), .A2(n17794), .ZN(n17795) );
  OAI211_X1 U20897 ( .C1(n17797), .C2(n17939), .A(n17796), .B(n17795), .ZN(
        P3_U2848) );
  AOI22_X1 U20898 ( .A1(n9578), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n17848), 
        .B2(n17798), .ZN(n17805) );
  OAI21_X1 U20899 ( .B1(n17836), .B2(n17810), .A(n17834), .ZN(n17829) );
  OAI22_X1 U20900 ( .A1(n17800), .A2(n9776), .B1(n17799), .B2(n17823), .ZN(
        n17801) );
  NOR3_X1 U20901 ( .A1(n17820), .A2(n17829), .A3(n17801), .ZN(n17809) );
  OAI211_X1 U20902 ( .C1(n17836), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17809), .B(n17802), .ZN(n17803) );
  OAI211_X1 U20903 ( .C1(n9563), .C2(n17803), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17852), .ZN(n17804) );
  OAI211_X1 U20904 ( .C1(n17870), .C2(n17806), .A(n17805), .B(n17804), .ZN(
        P3_U2849) );
  OAI22_X1 U20905 ( .A1(n18395), .A2(n9954), .B1(n17807), .B2(n17842), .ZN(
        n17808) );
  AOI21_X1 U20906 ( .B1(n17809), .B2(n17808), .A(n9563), .ZN(n17814) );
  INV_X1 U20907 ( .A(n17810), .ZN(n17811) );
  OAI21_X1 U20908 ( .B1(n17812), .B2(n17811), .A(n9954), .ZN(n17813) );
  AOI22_X1 U20909 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17936), .B1(
        n17814), .B2(n17813), .ZN(n17816) );
  OAI211_X1 U20910 ( .C1(n17817), .C2(n17870), .A(n17816), .B(n17815), .ZN(
        P3_U2850) );
  INV_X1 U20911 ( .A(n17818), .ZN(n17826) );
  AOI21_X1 U20912 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17819), .A(
        n9569), .ZN(n17825) );
  AOI211_X1 U20913 ( .C1(n17821), .C2(n18439), .A(n17820), .B(n9563), .ZN(
        n17822) );
  OAI21_X1 U20914 ( .B1(n17824), .B2(n17823), .A(n17822), .ZN(n17846) );
  AOI211_X1 U20915 ( .C1(n17827), .C2(n17826), .A(n17825), .B(n17846), .ZN(
        n17835) );
  OAI21_X1 U20916 ( .B1(n9569), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17835), .ZN(n17828) );
  OAI21_X1 U20917 ( .B1(n17829), .B2(n17828), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U20918 ( .A1(n17850), .A2(n17831), .B1(n17848), .B2(n17830), .ZN(
        n17832) );
  OAI221_X1 U20919 ( .B1(n9578), .B2(n17833), .C1(n17852), .C2(n18497), .A(
        n17832), .ZN(P3_U2851) );
  OAI211_X1 U20920 ( .C1(n17836), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17835), .B(n17834), .ZN(n17837) );
  OAI221_X1 U20921 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n17852), .C1(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n9578), .A(n17837), .ZN(
        n17840) );
  NAND3_X1 U20922 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17848), .A3(
        n17838), .ZN(n17839) );
  OAI211_X1 U20923 ( .C1(n17841), .C2(n17870), .A(n17840), .B(n17839), .ZN(
        P3_U2852) );
  OAI21_X1 U20924 ( .B1(n17862), .B2(n18395), .A(n17842), .ZN(n17844) );
  OAI22_X1 U20925 ( .A1(n17919), .A2(n17844), .B1(n17942), .B2(n17843), .ZN(
        n17845) );
  OAI21_X1 U20926 ( .B1(n17846), .B2(n17845), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17853) );
  INV_X1 U20927 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17847) );
  AOI22_X1 U20928 ( .A1(n17850), .A2(n17849), .B1(n17848), .B2(n17847), .ZN(
        n17851) );
  OAI221_X1 U20929 ( .B1(n9578), .B2(n17853), .C1(n17852), .C2(n18493), .A(
        n17851), .ZN(P3_U2853) );
  NOR3_X1 U20930 ( .A1(n17854), .A2(n9563), .A3(n17897), .ZN(n17901) );
  NAND3_X1 U20931 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n17901), .ZN(n17886) );
  NOR2_X1 U20932 ( .A1(n17855), .A2(n17886), .ZN(n17863) );
  AOI21_X1 U20933 ( .B1(n17913), .B2(n18411), .A(n17921), .ZN(n17895) );
  INV_X1 U20934 ( .A(n17919), .ZN(n17899) );
  NAND2_X1 U20935 ( .A1(n17899), .A2(n17856), .ZN(n17857) );
  OAI211_X1 U20936 ( .C1(n17871), .C2(n18429), .A(n17895), .B(n17857), .ZN(
        n17881) );
  AOI211_X1 U20937 ( .C1(n17859), .C2(n17858), .A(n17874), .B(n17881), .ZN(
        n17872) );
  OAI21_X1 U20938 ( .B1(n17872), .B2(n17929), .A(n17900), .ZN(n17861) );
  AOI221_X1 U20939 ( .B1(n17863), .B2(n17862), .C1(n17861), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n17860), .ZN(n17868) );
  AOI22_X1 U20940 ( .A1(n17866), .A2(n17865), .B1(n17945), .B2(n17864), .ZN(
        n17867) );
  OAI211_X1 U20941 ( .C1(n17870), .C2(n17869), .A(n17868), .B(n17867), .ZN(
        P3_U2854) );
  NAND3_X1 U20942 ( .A1(n17871), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n17906), .ZN(n17873) );
  AOI211_X1 U20943 ( .C1(n17874), .C2(n17873), .A(n17872), .B(n9563), .ZN(
        n17876) );
  OAI22_X1 U20944 ( .A1(n17874), .A2(n17900), .B1(n17852), .B2(n18489), .ZN(
        n17875) );
  AOI211_X1 U20945 ( .C1(n17877), .C2(n17932), .A(n17876), .B(n17875), .ZN(
        n17878) );
  OAI21_X1 U20946 ( .B1(n17939), .B2(n17879), .A(n17878), .ZN(P3_U2855) );
  AOI22_X1 U20947 ( .A1(n9578), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17932), .B2(
        n17880), .ZN(n17885) );
  INV_X1 U20948 ( .A(n17881), .ZN(n17882) );
  AOI21_X1 U20949 ( .B1(n9564), .B2(n17882), .A(n9578), .ZN(n17889) );
  AOI22_X1 U20950 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17889), .B1(
        n17945), .B2(n17883), .ZN(n17884) );
  OAI211_X1 U20951 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n17886), .A(
        n17885), .B(n17884), .ZN(P3_U2856) );
  AOI22_X1 U20952 ( .A1(n9578), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17932), .B2(
        n17887), .ZN(n17893) );
  AOI22_X1 U20953 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17889), .B1(
        n17945), .B2(n17888), .ZN(n17892) );
  NAND3_X1 U20954 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17901), .A3(
        n17890), .ZN(n17891) );
  NAND3_X1 U20955 ( .A1(n17893), .A2(n17892), .A3(n17891), .ZN(P3_U2857) );
  AOI22_X1 U20956 ( .A1(n9578), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n17932), .B2(
        n17894), .ZN(n17904) );
  INV_X1 U20957 ( .A(n17895), .ZN(n17896) );
  AOI211_X1 U20958 ( .C1(n17899), .C2(n17898), .A(n17897), .B(n17896), .ZN(
        n17912) );
  OAI21_X1 U20959 ( .B1(n17912), .B2(n17929), .A(n17900), .ZN(n17902) );
  AOI22_X1 U20960 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17902), .B1(
        n17901), .B2(n11288), .ZN(n17903) );
  OAI211_X1 U20961 ( .C1(n17939), .C2(n17905), .A(n17904), .B(n17903), .ZN(
        P3_U2858) );
  OAI21_X1 U20962 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17906), .A(
        n9564), .ZN(n17911) );
  AOI22_X1 U20963 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17936), .B1(
        n9578), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n17910) );
  AOI22_X1 U20964 ( .A1(n17945), .A2(n17908), .B1(n17932), .B2(n17907), .ZN(
        n17909) );
  OAI211_X1 U20965 ( .C1(n17912), .C2(n17911), .A(n17910), .B(n17909), .ZN(
        P3_U2859) );
  INV_X1 U20966 ( .A(n17932), .ZN(n17949) );
  AND2_X1 U20967 ( .A1(n18411), .A2(n17913), .ZN(n17916) );
  NOR3_X1 U20968 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20679), .A3(
        n17914), .ZN(n17915) );
  AOI211_X1 U20969 ( .C1(n18439), .C2(n17917), .A(n17916), .B(n17915), .ZN(
        n17923) );
  NAND2_X1 U20970 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17918) );
  OAI22_X1 U20971 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17919), .B1(
        n18429), .B2(n17918), .ZN(n17920) );
  OAI21_X1 U20972 ( .B1(n17921), .B2(n17920), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17922) );
  AOI21_X1 U20973 ( .B1(n17923), .B2(n17922), .A(n9563), .ZN(n17924) );
  AOI211_X1 U20974 ( .C1(n17936), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n17925), .B(n17924), .ZN(n17926) );
  OAI21_X1 U20975 ( .B1(n17949), .B2(n17927), .A(n17926), .ZN(P3_U2860) );
  INV_X1 U20976 ( .A(n17928), .ZN(n17940) );
  NOR2_X1 U20977 ( .A1(n17852), .A2(n18587), .ZN(n17931) );
  AOI211_X1 U20978 ( .C1(n17942), .C2(n18572), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n17929), .ZN(n17930) );
  AOI211_X1 U20979 ( .C1(n17933), .C2(n17932), .A(n17931), .B(n17930), .ZN(
        n17938) );
  NOR3_X1 U20980 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17935), .A3(
        n9563), .ZN(n17944) );
  OAI21_X1 U20981 ( .B1(n17936), .B2(n17944), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17937) );
  OAI211_X1 U20982 ( .C1(n17940), .C2(n17939), .A(n17938), .B(n17937), .ZN(
        P3_U2861) );
  AOI211_X1 U20983 ( .C1(n17942), .C2(n9564), .A(n9578), .B(n18572), .ZN(
        n17943) );
  AOI211_X1 U20984 ( .C1(n17945), .C2(n17948), .A(n17944), .B(n17943), .ZN(
        n17947) );
  NAND2_X1 U20985 ( .A1(n9578), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n17946) );
  OAI211_X1 U20986 ( .C1(n17949), .C2(n17948), .A(n17947), .B(n17946), .ZN(
        P3_U2862) );
  AOI21_X1 U20987 ( .B1(n17952), .B2(n17951), .A(n17950), .ZN(n18447) );
  OAI21_X1 U20988 ( .B1(n18447), .B2(n17999), .A(n17957), .ZN(n17953) );
  OAI221_X1 U20989 ( .B1(n18404), .B2(n18605), .C1(n18404), .C2(n17957), .A(
        n17953), .ZN(P3_U2863) );
  NOR2_X1 U20990 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20820), .ZN(
        n18086) );
  NOR2_X1 U20991 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18425), .ZN(
        n18200) );
  NOR2_X1 U20992 ( .A1(n18086), .A2(n18200), .ZN(n17955) );
  OAI22_X1 U20993 ( .A1(n17956), .A2(n18425), .B1(n17955), .B2(n17954), .ZN(
        P3_U2866) );
  NOR2_X1 U20994 ( .A1(n18426), .A2(n17957), .ZN(P3_U2867) );
  NOR2_X1 U20995 ( .A1(n17959), .A2(n17958), .ZN(n17990) );
  NAND2_X1 U20996 ( .A1(n17960), .A2(n17990), .ZN(n18338) );
  NOR2_X1 U20997 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18408) );
  NAND2_X1 U20998 ( .A1(n20820), .A2(n18425), .ZN(n18042) );
  INV_X1 U20999 ( .A(n18042), .ZN(n18001) );
  NAND2_X1 U21000 ( .A1(n18408), .A2(n18001), .ZN(n18041) );
  NAND2_X1 U21001 ( .A1(n18273), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18303) );
  INV_X1 U21002 ( .A(n18303), .ZN(n18331) );
  NOR2_X1 U21003 ( .A1(n18425), .A2(n18109), .ZN(n18333) );
  INV_X1 U21004 ( .A(n18333), .ZN(n18328) );
  NOR2_X2 U21005 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18328), .ZN(
        n18321) );
  NOR2_X2 U21006 ( .A1(n18000), .A2(n17961), .ZN(n18330) );
  NOR2_X2 U21007 ( .A1(n18404), .A2(n18328), .ZN(n18341) );
  NOR2_X1 U21008 ( .A1(n18341), .A2(n18059), .ZN(n18021) );
  NOR2_X1 U21009 ( .A1(n18329), .A2(n18021), .ZN(n17993) );
  AOI22_X1 U21010 ( .A1(n18331), .A2(n18321), .B1(n18330), .B2(n17993), .ZN(
        n17965) );
  NAND2_X1 U21011 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18405), .ZN(
        n18177) );
  INV_X1 U21012 ( .A(n18177), .ZN(n18085) );
  NOR2_X1 U21013 ( .A1(n20820), .A2(n18425), .ZN(n18271) );
  NAND2_X1 U21014 ( .A1(n18085), .A2(n18271), .ZN(n18345) );
  NAND2_X1 U21015 ( .A1(n18345), .A2(n18318), .ZN(n18299) );
  AOI21_X1 U21016 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18000), .ZN(n18296) );
  INV_X1 U21017 ( .A(n18021), .ZN(n17962) );
  AOI22_X1 U21018 ( .A1(n18273), .A2(n18299), .B1(n18296), .B2(n17962), .ZN(
        n17996) );
  NOR2_X2 U21019 ( .A1(n17963), .A2(n17995), .ZN(n18335) );
  INV_X1 U21020 ( .A(n18345), .ZN(n18379) );
  AOI22_X1 U21021 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17996), .B1(
        n18335), .B2(n18379), .ZN(n17964) );
  OAI211_X1 U21022 ( .C1(n18338), .C2(n18041), .A(n17965), .B(n17964), .ZN(
        P3_U2868) );
  NAND2_X1 U21023 ( .A1(n18273), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18346) );
  NOR2_X2 U21024 ( .A1(n18000), .A2(n17966), .ZN(n18340) );
  AND2_X1 U21025 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18273), .ZN(n18339) );
  AOI22_X1 U21026 ( .A1(n18340), .A2(n17993), .B1(n18339), .B2(n18379), .ZN(
        n17968) );
  NAND2_X1 U21027 ( .A1(n18598), .A2(n17990), .ZN(n18307) );
  INV_X1 U21028 ( .A(n18307), .ZN(n18342) );
  AOI22_X1 U21029 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17996), .B1(
        n18342), .B2(n18059), .ZN(n17967) );
  OAI211_X1 U21030 ( .C1(n18346), .C2(n18318), .A(n17968), .B(n17967), .ZN(
        P3_U2869) );
  NAND2_X1 U21031 ( .A1(n17990), .A2(n17969), .ZN(n18352) );
  NOR2_X2 U21032 ( .A1(n18000), .A2(n20714), .ZN(n18347) );
  AOI22_X1 U21033 ( .A1(n18348), .A2(n18321), .B1(n18347), .B2(n17993), .ZN(
        n17971) );
  NOR2_X2 U21034 ( .A1(n14959), .A2(n17995), .ZN(n18349) );
  AOI22_X1 U21035 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n17996), .B1(
        n18349), .B2(n18379), .ZN(n17970) );
  OAI211_X1 U21036 ( .C1(n18352), .C2(n18041), .A(n17971), .B(n17970), .ZN(
        P3_U2870) );
  NAND2_X1 U21037 ( .A1(n18273), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18283) );
  NOR2_X2 U21038 ( .A1(n18000), .A2(n17972), .ZN(n18353) );
  AND2_X1 U21039 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18273), .ZN(n18355) );
  AOI22_X1 U21040 ( .A1(n18353), .A2(n17993), .B1(n18355), .B2(n18379), .ZN(
        n17975) );
  NAND2_X1 U21041 ( .A1(n17973), .A2(n17990), .ZN(n18358) );
  AOI22_X1 U21042 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n17996), .B1(
        n18280), .B2(n18059), .ZN(n17974) );
  OAI211_X1 U21043 ( .C1(n18283), .C2(n18318), .A(n17975), .B(n17974), .ZN(
        P3_U2871) );
  NAND2_X1 U21044 ( .A1(n17990), .A2(n17976), .ZN(n18364) );
  NOR2_X2 U21045 ( .A1(n17977), .A2(n17995), .ZN(n18360) );
  NOR2_X2 U21046 ( .A1(n18000), .A2(n17978), .ZN(n18359) );
  AOI22_X1 U21047 ( .A1(n18360), .A2(n18379), .B1(n18359), .B2(n17993), .ZN(
        n17980) );
  AND2_X1 U21048 ( .A1(n18273), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18361) );
  AOI22_X1 U21049 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n17996), .B1(
        n18361), .B2(n18321), .ZN(n17979) );
  OAI211_X1 U21050 ( .C1(n18364), .C2(n18041), .A(n17980), .B(n17979), .ZN(
        P3_U2872) );
  NAND2_X1 U21051 ( .A1(n17990), .A2(n17981), .ZN(n18370) );
  AND2_X1 U21052 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18273), .ZN(n18367) );
  NOR2_X2 U21053 ( .A1(n18000), .A2(n17982), .ZN(n18365) );
  AOI22_X1 U21054 ( .A1(n18367), .A2(n18379), .B1(n18365), .B2(n17993), .ZN(
        n17984) );
  NOR2_X2 U21055 ( .A1(n17995), .A2(n14995), .ZN(n18366) );
  AOI22_X1 U21056 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n17996), .B1(
        n18366), .B2(n18321), .ZN(n17983) );
  OAI211_X1 U21057 ( .C1(n18370), .C2(n18041), .A(n17984), .B(n17983), .ZN(
        P3_U2873) );
  NAND2_X1 U21058 ( .A1(n17990), .A2(n17985), .ZN(n18376) );
  NOR2_X2 U21059 ( .A1(n17986), .A2(n17995), .ZN(n18372) );
  NOR2_X2 U21060 ( .A1(n18000), .A2(n17987), .ZN(n18371) );
  AOI22_X1 U21061 ( .A1(n18372), .A2(n18379), .B1(n18371), .B2(n17993), .ZN(
        n17989) );
  AND2_X1 U21062 ( .A1(n18273), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U21063 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17996), .B1(
        n18373), .B2(n18321), .ZN(n17988) );
  OAI211_X1 U21064 ( .C1(n18376), .C2(n18041), .A(n17989), .B(n17988), .ZN(
        P3_U2874) );
  NAND2_X1 U21065 ( .A1(n17991), .A2(n17990), .ZN(n18387) );
  NAND2_X1 U21066 ( .A1(n18273), .A2(BUF2_REG_23__SCAN_IN), .ZN(n18327) );
  INV_X1 U21067 ( .A(n18327), .ZN(n18380) );
  NOR2_X2 U21068 ( .A1(n18000), .A2(n17992), .ZN(n18378) );
  AOI22_X1 U21069 ( .A1(n18380), .A2(n18321), .B1(n18378), .B2(n17993), .ZN(
        n17998) );
  NOR2_X2 U21070 ( .A1(n17995), .A2(n17994), .ZN(n18382) );
  AOI22_X1 U21071 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17996), .B1(
        n18382), .B2(n18379), .ZN(n17997) );
  OAI211_X1 U21072 ( .C1(n18387), .C2(n18041), .A(n17998), .B(n17997), .ZN(
        P3_U2875) );
  INV_X1 U21073 ( .A(n18329), .ZN(n18294) );
  NAND2_X1 U21074 ( .A1(n18405), .A2(n18294), .ZN(n18268) );
  NOR2_X1 U21075 ( .A1(n18042), .A2(n18268), .ZN(n18016) );
  AOI22_X1 U21076 ( .A1(n18330), .A2(n18016), .B1(n18335), .B2(n18321), .ZN(
        n18003) );
  NOR2_X1 U21077 ( .A1(n18000), .A2(n17999), .ZN(n18332) );
  INV_X1 U21078 ( .A(n18332), .ZN(n18087) );
  NOR2_X1 U21079 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18087), .ZN(
        n18270) );
  AOI22_X1 U21080 ( .A1(n18273), .A2(n18333), .B1(n18001), .B2(n18270), .ZN(
        n18017) );
  NOR2_X2 U21081 ( .A1(n18042), .A2(n18177), .ZN(n18080) );
  INV_X1 U21082 ( .A(n18338), .ZN(n18300) );
  AOI22_X1 U21083 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18017), .B1(
        n18080), .B2(n18300), .ZN(n18002) );
  OAI211_X1 U21084 ( .C1(n18303), .C2(n18386), .A(n18003), .B(n18002), .ZN(
        P3_U2876) );
  AOI22_X1 U21085 ( .A1(n18340), .A2(n18016), .B1(n18339), .B2(n18321), .ZN(
        n18005) );
  AOI22_X1 U21086 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18017), .B1(
        n18080), .B2(n18342), .ZN(n18004) );
  OAI211_X1 U21087 ( .C1(n18346), .C2(n18386), .A(n18005), .B(n18004), .ZN(
        P3_U2877) );
  INV_X1 U21088 ( .A(n18080), .ZN(n18020) );
  AOI22_X1 U21089 ( .A1(n18348), .A2(n18341), .B1(n18347), .B2(n18016), .ZN(
        n18007) );
  AOI22_X1 U21090 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18017), .B1(
        n18349), .B2(n18321), .ZN(n18006) );
  OAI211_X1 U21091 ( .C1(n18020), .C2(n18352), .A(n18007), .B(n18006), .ZN(
        P3_U2878) );
  INV_X1 U21092 ( .A(n18283), .ZN(n18354) );
  AOI22_X1 U21093 ( .A1(n18354), .A2(n18341), .B1(n18353), .B2(n18016), .ZN(
        n18009) );
  AOI22_X1 U21094 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18017), .B1(
        n18355), .B2(n18321), .ZN(n18008) );
  OAI211_X1 U21095 ( .C1(n18020), .C2(n18358), .A(n18009), .B(n18008), .ZN(
        P3_U2879) );
  AOI22_X1 U21096 ( .A1(n18360), .A2(n18321), .B1(n18359), .B2(n18016), .ZN(
        n18011) );
  AOI22_X1 U21097 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18017), .B1(
        n18361), .B2(n18341), .ZN(n18010) );
  OAI211_X1 U21098 ( .C1(n18020), .C2(n18364), .A(n18011), .B(n18010), .ZN(
        P3_U2880) );
  AOI22_X1 U21099 ( .A1(n18366), .A2(n18341), .B1(n18365), .B2(n18016), .ZN(
        n18013) );
  AOI22_X1 U21100 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18017), .B1(
        n18367), .B2(n18321), .ZN(n18012) );
  OAI211_X1 U21101 ( .C1(n18020), .C2(n18370), .A(n18013), .B(n18012), .ZN(
        P3_U2881) );
  AOI22_X1 U21102 ( .A1(n18373), .A2(n18341), .B1(n18371), .B2(n18016), .ZN(
        n18015) );
  AOI22_X1 U21103 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18017), .B1(
        n18372), .B2(n18321), .ZN(n18014) );
  OAI211_X1 U21104 ( .C1(n18020), .C2(n18376), .A(n18015), .B(n18014), .ZN(
        P3_U2882) );
  AOI22_X1 U21105 ( .A1(n18380), .A2(n18341), .B1(n18378), .B2(n18016), .ZN(
        n18019) );
  AOI22_X1 U21106 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18017), .B1(
        n18382), .B2(n18321), .ZN(n18018) );
  OAI211_X1 U21107 ( .C1(n18020), .C2(n18387), .A(n18019), .B(n18018), .ZN(
        P3_U2883) );
  NOR2_X1 U21108 ( .A1(n18405), .A2(n18042), .ZN(n18089) );
  NAND2_X1 U21109 ( .A1(n18089), .A2(n18404), .ZN(n18084) );
  NOR2_X1 U21110 ( .A1(n18105), .A2(n18080), .ZN(n18063) );
  NOR2_X1 U21111 ( .A1(n18329), .A2(n18063), .ZN(n18037) );
  AOI22_X1 U21112 ( .A1(n18330), .A2(n18037), .B1(n18335), .B2(n18341), .ZN(
        n18024) );
  OAI21_X1 U21113 ( .B1(n18021), .B2(n18245), .A(n18063), .ZN(n18022) );
  OAI211_X1 U21114 ( .C1(n18105), .C2(n18543), .A(n18247), .B(n18022), .ZN(
        n18038) );
  AOI22_X1 U21115 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18038), .B1(
        n18105), .B2(n18300), .ZN(n18023) );
  OAI211_X1 U21116 ( .C1(n18303), .C2(n18041), .A(n18024), .B(n18023), .ZN(
        P3_U2884) );
  AOI22_X1 U21117 ( .A1(n18304), .A2(n18059), .B1(n18340), .B2(n18037), .ZN(
        n18026) );
  AOI22_X1 U21118 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18038), .B1(
        n18339), .B2(n18341), .ZN(n18025) );
  OAI211_X1 U21119 ( .C1(n18084), .C2(n18307), .A(n18026), .B(n18025), .ZN(
        P3_U2885) );
  AOI22_X1 U21120 ( .A1(n18348), .A2(n18059), .B1(n18347), .B2(n18037), .ZN(
        n18028) );
  AOI22_X1 U21121 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18038), .B1(
        n18349), .B2(n18341), .ZN(n18027) );
  OAI211_X1 U21122 ( .C1(n18084), .C2(n18352), .A(n18028), .B(n18027), .ZN(
        P3_U2886) );
  AOI22_X1 U21123 ( .A1(n18353), .A2(n18037), .B1(n18355), .B2(n18341), .ZN(
        n18030) );
  AOI22_X1 U21124 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18038), .B1(
        n18105), .B2(n18280), .ZN(n18029) );
  OAI211_X1 U21125 ( .C1(n18283), .C2(n18041), .A(n18030), .B(n18029), .ZN(
        P3_U2887) );
  AOI22_X1 U21126 ( .A1(n18359), .A2(n18037), .B1(n18361), .B2(n18059), .ZN(
        n18032) );
  AOI22_X1 U21127 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18038), .B1(
        n18360), .B2(n18341), .ZN(n18031) );
  OAI211_X1 U21128 ( .C1(n18084), .C2(n18364), .A(n18032), .B(n18031), .ZN(
        P3_U2888) );
  AOI22_X1 U21129 ( .A1(n18366), .A2(n18059), .B1(n18365), .B2(n18037), .ZN(
        n18034) );
  AOI22_X1 U21130 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18038), .B1(
        n18367), .B2(n18341), .ZN(n18033) );
  OAI211_X1 U21131 ( .C1(n18084), .C2(n18370), .A(n18034), .B(n18033), .ZN(
        P3_U2889) );
  AOI22_X1 U21132 ( .A1(n18372), .A2(n18341), .B1(n18371), .B2(n18037), .ZN(
        n18036) );
  AOI22_X1 U21133 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18038), .B1(
        n18373), .B2(n18059), .ZN(n18035) );
  OAI211_X1 U21134 ( .C1(n18084), .C2(n18376), .A(n18036), .B(n18035), .ZN(
        P3_U2890) );
  AOI22_X1 U21135 ( .A1(n18382), .A2(n18341), .B1(n18378), .B2(n18037), .ZN(
        n18040) );
  INV_X1 U21136 ( .A(n18387), .ZN(n18322) );
  AOI22_X1 U21137 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18038), .B1(
        n18105), .B2(n18322), .ZN(n18039) );
  OAI211_X1 U21138 ( .C1(n18327), .C2(n18041), .A(n18040), .B(n18039), .ZN(
        P3_U2891) );
  NAND2_X1 U21139 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18089), .ZN(
        n18110) );
  AND2_X1 U21140 ( .A1(n18294), .A2(n18089), .ZN(n18058) );
  AOI22_X1 U21141 ( .A1(n18330), .A2(n18058), .B1(n18335), .B2(n18059), .ZN(
        n18045) );
  OAI21_X1 U21142 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18042), .A(n18110), 
        .ZN(n18043) );
  NAND3_X1 U21143 ( .A1(n18247), .A2(n18133), .A3(n18043), .ZN(n18060) );
  AOI22_X1 U21144 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18060), .B1(
        n18331), .B2(n18080), .ZN(n18044) );
  OAI211_X1 U21145 ( .C1(n18110), .C2(n18338), .A(n18045), .B(n18044), .ZN(
        P3_U2892) );
  AOI22_X1 U21146 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18060), .B1(
        n18340), .B2(n18058), .ZN(n18047) );
  AOI22_X1 U21147 ( .A1(n18080), .A2(n18304), .B1(n18339), .B2(n18059), .ZN(
        n18046) );
  OAI211_X1 U21148 ( .C1(n18110), .C2(n18307), .A(n18047), .B(n18046), .ZN(
        P3_U2893) );
  AOI22_X1 U21149 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18060), .B1(
        n18347), .B2(n18058), .ZN(n18049) );
  AOI22_X1 U21150 ( .A1(n18080), .A2(n18348), .B1(n18349), .B2(n18059), .ZN(
        n18048) );
  OAI211_X1 U21151 ( .C1(n18110), .C2(n18352), .A(n18049), .B(n18048), .ZN(
        P3_U2894) );
  AOI22_X1 U21152 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18060), .B1(
        n18353), .B2(n18058), .ZN(n18051) );
  AOI22_X1 U21153 ( .A1(n18080), .A2(n18354), .B1(n18355), .B2(n18059), .ZN(
        n18050) );
  OAI211_X1 U21154 ( .C1(n18110), .C2(n18358), .A(n18051), .B(n18050), .ZN(
        P3_U2895) );
  AOI22_X1 U21155 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18060), .B1(
        n18359), .B2(n18058), .ZN(n18053) );
  AOI22_X1 U21156 ( .A1(n18080), .A2(n18361), .B1(n18360), .B2(n18059), .ZN(
        n18052) );
  OAI211_X1 U21157 ( .C1(n18110), .C2(n18364), .A(n18053), .B(n18052), .ZN(
        P3_U2896) );
  AOI22_X1 U21158 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18060), .B1(
        n18365), .B2(n18058), .ZN(n18055) );
  AOI22_X1 U21159 ( .A1(n18080), .A2(n18366), .B1(n18367), .B2(n18059), .ZN(
        n18054) );
  OAI211_X1 U21160 ( .C1(n18110), .C2(n18370), .A(n18055), .B(n18054), .ZN(
        P3_U2897) );
  AOI22_X1 U21161 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18060), .B1(
        n18371), .B2(n18058), .ZN(n18057) );
  AOI22_X1 U21162 ( .A1(n18080), .A2(n18373), .B1(n18372), .B2(n18059), .ZN(
        n18056) );
  OAI211_X1 U21163 ( .C1(n18110), .C2(n18376), .A(n18057), .B(n18056), .ZN(
        P3_U2898) );
  AOI22_X1 U21164 ( .A1(n18080), .A2(n18380), .B1(n18378), .B2(n18058), .ZN(
        n18062) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18060), .B1(
        n18382), .B2(n18059), .ZN(n18061) );
  OAI211_X1 U21166 ( .C1(n18110), .C2(n18387), .A(n18062), .B(n18061), .ZN(
        P3_U2899) );
  NAND2_X1 U21167 ( .A1(n18408), .A2(n18086), .ZN(n18117) );
  AOI21_X1 U21168 ( .B1(n18117), .B2(n18110), .A(n18329), .ZN(n18079) );
  AOI22_X1 U21169 ( .A1(n18080), .A2(n18335), .B1(n18330), .B2(n18079), .ZN(
        n18066) );
  AOI221_X1 U21170 ( .B1(n18063), .B2(n18110), .C1(n18245), .C2(n18110), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18064) );
  OAI21_X1 U21171 ( .B1(n18151), .B2(n18064), .A(n18247), .ZN(n18081) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18081), .B1(
        n18151), .B2(n18300), .ZN(n18065) );
  OAI211_X1 U21173 ( .C1(n18303), .C2(n18084), .A(n18066), .B(n18065), .ZN(
        P3_U2900) );
  AOI22_X1 U21174 ( .A1(n18080), .A2(n18339), .B1(n18079), .B2(n18340), .ZN(
        n18068) );
  AOI22_X1 U21175 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18081), .B1(
        n18151), .B2(n18342), .ZN(n18067) );
  OAI211_X1 U21176 ( .C1(n18084), .C2(n18346), .A(n18068), .B(n18067), .ZN(
        P3_U2901) );
  AOI22_X1 U21177 ( .A1(n18105), .A2(n18348), .B1(n18079), .B2(n18347), .ZN(
        n18070) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18081), .B1(
        n18080), .B2(n18349), .ZN(n18069) );
  OAI211_X1 U21179 ( .C1(n18117), .C2(n18352), .A(n18070), .B(n18069), .ZN(
        P3_U2902) );
  AOI22_X1 U21180 ( .A1(n18080), .A2(n18355), .B1(n18079), .B2(n18353), .ZN(
        n18072) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18081), .B1(
        n18151), .B2(n18280), .ZN(n18071) );
  OAI211_X1 U21182 ( .C1(n18084), .C2(n18283), .A(n18072), .B(n18071), .ZN(
        P3_U2903) );
  AOI22_X1 U21183 ( .A1(n18105), .A2(n18361), .B1(n18079), .B2(n18359), .ZN(
        n18074) );
  AOI22_X1 U21184 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18081), .B1(
        n18080), .B2(n18360), .ZN(n18073) );
  OAI211_X1 U21185 ( .C1(n18117), .C2(n18364), .A(n18074), .B(n18073), .ZN(
        P3_U2904) );
  AOI22_X1 U21186 ( .A1(n18105), .A2(n18366), .B1(n18079), .B2(n18365), .ZN(
        n18076) );
  AOI22_X1 U21187 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18081), .B1(
        n18080), .B2(n18367), .ZN(n18075) );
  OAI211_X1 U21188 ( .C1(n18117), .C2(n18370), .A(n18076), .B(n18075), .ZN(
        P3_U2905) );
  AOI22_X1 U21189 ( .A1(n18105), .A2(n18373), .B1(n18079), .B2(n18371), .ZN(
        n18078) );
  AOI22_X1 U21190 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18081), .B1(
        n18080), .B2(n18372), .ZN(n18077) );
  OAI211_X1 U21191 ( .C1(n18117), .C2(n18376), .A(n18078), .B(n18077), .ZN(
        P3_U2906) );
  AOI22_X1 U21192 ( .A1(n18080), .A2(n18382), .B1(n18079), .B2(n18378), .ZN(
        n18083) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18081), .B1(
        n18151), .B2(n18322), .ZN(n18082) );
  OAI211_X1 U21194 ( .C1(n18084), .C2(n18327), .A(n18083), .B(n18082), .ZN(
        P3_U2907) );
  NAND2_X1 U21195 ( .A1(n18086), .A2(n18085), .ZN(n18143) );
  INV_X1 U21196 ( .A(n18110), .ZN(n18129) );
  INV_X1 U21197 ( .A(n18086), .ZN(n18088) );
  NOR2_X1 U21198 ( .A1(n18088), .A2(n18268), .ZN(n18104) );
  AOI22_X1 U21199 ( .A1(n18331), .A2(n18129), .B1(n18330), .B2(n18104), .ZN(
        n18091) );
  NOR2_X1 U21200 ( .A1(n18088), .A2(n18087), .ZN(n18134) );
  AOI22_X1 U21201 ( .A1(n18089), .A2(n18273), .B1(n18134), .B2(n18405), .ZN(
        n18106) );
  AOI22_X1 U21202 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18106), .B1(
        n18105), .B2(n18335), .ZN(n18090) );
  OAI211_X1 U21203 ( .C1(n18338), .C2(n18143), .A(n18091), .B(n18090), .ZN(
        P3_U2908) );
  AOI22_X1 U21204 ( .A1(n18129), .A2(n18304), .B1(n18340), .B2(n18104), .ZN(
        n18093) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18106), .B1(
        n18105), .B2(n18339), .ZN(n18092) );
  OAI211_X1 U21206 ( .C1(n18307), .C2(n18143), .A(n18093), .B(n18092), .ZN(
        P3_U2909) );
  AOI22_X1 U21207 ( .A1(n18105), .A2(n18349), .B1(n18347), .B2(n18104), .ZN(
        n18095) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18106), .B1(
        n18129), .B2(n18348), .ZN(n18094) );
  OAI211_X1 U21209 ( .C1(n18352), .C2(n18143), .A(n18095), .B(n18094), .ZN(
        P3_U2910) );
  AOI22_X1 U21210 ( .A1(n18105), .A2(n18355), .B1(n18353), .B2(n18104), .ZN(
        n18097) );
  AOI22_X1 U21211 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18106), .B1(
        n18129), .B2(n18354), .ZN(n18096) );
  OAI211_X1 U21212 ( .C1(n18358), .C2(n18143), .A(n18097), .B(n18096), .ZN(
        P3_U2911) );
  AOI22_X1 U21213 ( .A1(n18105), .A2(n18360), .B1(n18359), .B2(n18104), .ZN(
        n18099) );
  AOI22_X1 U21214 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18106), .B1(
        n18129), .B2(n18361), .ZN(n18098) );
  OAI211_X1 U21215 ( .C1(n18364), .C2(n18143), .A(n18099), .B(n18098), .ZN(
        P3_U2912) );
  AOI22_X1 U21216 ( .A1(n18105), .A2(n18367), .B1(n18365), .B2(n18104), .ZN(
        n18101) );
  AOI22_X1 U21217 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18106), .B1(
        n18129), .B2(n18366), .ZN(n18100) );
  OAI211_X1 U21218 ( .C1(n18370), .C2(n18143), .A(n18101), .B(n18100), .ZN(
        P3_U2913) );
  AOI22_X1 U21219 ( .A1(n18129), .A2(n18373), .B1(n18371), .B2(n18104), .ZN(
        n18103) );
  AOI22_X1 U21220 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18106), .B1(
        n18105), .B2(n18372), .ZN(n18102) );
  OAI211_X1 U21221 ( .C1(n18376), .C2(n18143), .A(n18103), .B(n18102), .ZN(
        P3_U2914) );
  AOI22_X1 U21222 ( .A1(n18129), .A2(n18380), .B1(n18378), .B2(n18104), .ZN(
        n18108) );
  AOI22_X1 U21223 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18106), .B1(
        n18105), .B2(n18382), .ZN(n18107) );
  OAI211_X1 U21224 ( .C1(n18387), .C2(n18143), .A(n18108), .B(n18107), .ZN(
        P3_U2915) );
  NOR2_X1 U21225 ( .A1(n18109), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18179) );
  NAND2_X1 U21226 ( .A1(n18404), .A2(n18179), .ZN(n18176) );
  NOR2_X1 U21227 ( .A1(n18172), .A2(n18195), .ZN(n18155) );
  NOR2_X1 U21228 ( .A1(n18329), .A2(n18155), .ZN(n18128) );
  AOI22_X1 U21229 ( .A1(n18129), .A2(n18335), .B1(n18330), .B2(n18128), .ZN(
        n18114) );
  INV_X1 U21230 ( .A(n18155), .ZN(n18112) );
  NAND2_X1 U21231 ( .A1(n18117), .A2(n18110), .ZN(n18111) );
  OAI221_X1 U21232 ( .B1(n18112), .B2(n18298), .C1(n18112), .C2(n18111), .A(
        n18296), .ZN(n18130) );
  AOI22_X1 U21233 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18130), .B1(
        n18300), .B2(n18195), .ZN(n18113) );
  OAI211_X1 U21234 ( .C1(n18303), .C2(n18117), .A(n18114), .B(n18113), .ZN(
        P3_U2916) );
  AOI22_X1 U21235 ( .A1(n18129), .A2(n18339), .B1(n18340), .B2(n18128), .ZN(
        n18116) );
  AOI22_X1 U21236 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18130), .B1(
        n18342), .B2(n18195), .ZN(n18115) );
  OAI211_X1 U21237 ( .C1(n18117), .C2(n18346), .A(n18116), .B(n18115), .ZN(
        P3_U2917) );
  AOI22_X1 U21238 ( .A1(n18129), .A2(n18349), .B1(n18347), .B2(n18128), .ZN(
        n18119) );
  AOI22_X1 U21239 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18130), .B1(
        n18151), .B2(n18348), .ZN(n18118) );
  OAI211_X1 U21240 ( .C1(n18352), .C2(n18176), .A(n18119), .B(n18118), .ZN(
        P3_U2918) );
  AOI22_X1 U21241 ( .A1(n18151), .A2(n18354), .B1(n18353), .B2(n18128), .ZN(
        n18121) );
  AOI22_X1 U21242 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18130), .B1(
        n18129), .B2(n18355), .ZN(n18120) );
  OAI211_X1 U21243 ( .C1(n18358), .C2(n18176), .A(n18121), .B(n18120), .ZN(
        P3_U2919) );
  AOI22_X1 U21244 ( .A1(n18151), .A2(n18361), .B1(n18359), .B2(n18128), .ZN(
        n18123) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18130), .B1(
        n18129), .B2(n18360), .ZN(n18122) );
  OAI211_X1 U21246 ( .C1(n18364), .C2(n18176), .A(n18123), .B(n18122), .ZN(
        P3_U2920) );
  AOI22_X1 U21247 ( .A1(n18151), .A2(n18366), .B1(n18365), .B2(n18128), .ZN(
        n18125) );
  AOI22_X1 U21248 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18130), .B1(
        n18129), .B2(n18367), .ZN(n18124) );
  OAI211_X1 U21249 ( .C1(n18370), .C2(n18176), .A(n18125), .B(n18124), .ZN(
        P3_U2921) );
  AOI22_X1 U21250 ( .A1(n18129), .A2(n18372), .B1(n18371), .B2(n18128), .ZN(
        n18127) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18130), .B1(
        n18151), .B2(n18373), .ZN(n18126) );
  OAI211_X1 U21252 ( .C1(n18376), .C2(n18176), .A(n18127), .B(n18126), .ZN(
        P3_U2922) );
  AOI22_X1 U21253 ( .A1(n18151), .A2(n18380), .B1(n18378), .B2(n18128), .ZN(
        n18132) );
  AOI22_X1 U21254 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18130), .B1(
        n18129), .B2(n18382), .ZN(n18131) );
  OAI211_X1 U21255 ( .C1(n18387), .C2(n18176), .A(n18132), .B(n18131), .ZN(
        P3_U2923) );
  AND2_X1 U21256 ( .A1(n18294), .A2(n18179), .ZN(n18150) );
  AOI22_X1 U21257 ( .A1(n18151), .A2(n18335), .B1(n18330), .B2(n18150), .ZN(
        n18136) );
  NAND2_X1 U21258 ( .A1(n18134), .A2(n18133), .ZN(n18152) );
  NAND2_X1 U21259 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18179), .ZN(
        n18199) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18152), .B1(
        n18300), .B2(n18219), .ZN(n18135) );
  OAI211_X1 U21261 ( .C1(n18303), .C2(n18143), .A(n18136), .B(n18135), .ZN(
        P3_U2924) );
  AOI22_X1 U21262 ( .A1(n18151), .A2(n18339), .B1(n18340), .B2(n18150), .ZN(
        n18138) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18152), .B1(
        n18342), .B2(n18219), .ZN(n18137) );
  OAI211_X1 U21264 ( .C1(n18346), .C2(n18143), .A(n18138), .B(n18137), .ZN(
        P3_U2925) );
  AOI22_X1 U21265 ( .A1(n18151), .A2(n18349), .B1(n18347), .B2(n18150), .ZN(
        n18140) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18152), .B1(
        n18348), .B2(n18172), .ZN(n18139) );
  OAI211_X1 U21267 ( .C1(n18352), .C2(n18199), .A(n18140), .B(n18139), .ZN(
        P3_U2926) );
  AOI22_X1 U21268 ( .A1(n18151), .A2(n18355), .B1(n18353), .B2(n18150), .ZN(
        n18142) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18152), .B1(
        n18280), .B2(n18219), .ZN(n18141) );
  OAI211_X1 U21270 ( .C1(n18283), .C2(n18143), .A(n18142), .B(n18141), .ZN(
        P3_U2927) );
  AOI22_X1 U21271 ( .A1(n18151), .A2(n18360), .B1(n18359), .B2(n18150), .ZN(
        n18145) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18152), .B1(
        n18361), .B2(n18172), .ZN(n18144) );
  OAI211_X1 U21273 ( .C1(n18364), .C2(n18199), .A(n18145), .B(n18144), .ZN(
        P3_U2928) );
  AOI22_X1 U21274 ( .A1(n18151), .A2(n18367), .B1(n18365), .B2(n18150), .ZN(
        n18147) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18152), .B1(
        n18366), .B2(n18172), .ZN(n18146) );
  OAI211_X1 U21276 ( .C1(n18370), .C2(n18199), .A(n18147), .B(n18146), .ZN(
        P3_U2929) );
  AOI22_X1 U21277 ( .A1(n18151), .A2(n18372), .B1(n18371), .B2(n18150), .ZN(
        n18149) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18152), .B1(
        n18373), .B2(n18172), .ZN(n18148) );
  OAI211_X1 U21279 ( .C1(n18376), .C2(n18199), .A(n18149), .B(n18148), .ZN(
        P3_U2930) );
  AOI22_X1 U21280 ( .A1(n18380), .A2(n18172), .B1(n18378), .B2(n18150), .ZN(
        n18154) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18152), .B1(
        n18151), .B2(n18382), .ZN(n18153) );
  OAI211_X1 U21282 ( .C1(n18387), .C2(n18199), .A(n18154), .B(n18153), .ZN(
        P3_U2931) );
  NAND2_X1 U21283 ( .A1(n18408), .A2(n18200), .ZN(n18223) );
  INV_X1 U21284 ( .A(n18223), .ZN(n18241) );
  NOR2_X1 U21285 ( .A1(n18219), .A2(n18241), .ZN(n18201) );
  NOR2_X1 U21286 ( .A1(n18329), .A2(n18201), .ZN(n18171) );
  AOI22_X1 U21287 ( .A1(n18330), .A2(n18171), .B1(n18335), .B2(n18172), .ZN(
        n18158) );
  OAI21_X1 U21288 ( .B1(n18155), .B2(n18245), .A(n18201), .ZN(n18156) );
  OAI211_X1 U21289 ( .C1(n18241), .C2(n18543), .A(n18247), .B(n18156), .ZN(
        n18173) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18173), .B1(
        n18331), .B2(n18195), .ZN(n18157) );
  OAI211_X1 U21291 ( .C1(n18338), .C2(n18223), .A(n18158), .B(n18157), .ZN(
        P3_U2932) );
  AOI22_X1 U21292 ( .A1(n18304), .A2(n18195), .B1(n18340), .B2(n18171), .ZN(
        n18160) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18173), .B1(
        n18339), .B2(n18172), .ZN(n18159) );
  OAI211_X1 U21294 ( .C1(n18307), .C2(n18223), .A(n18160), .B(n18159), .ZN(
        P3_U2933) );
  AOI22_X1 U21295 ( .A1(n18348), .A2(n18195), .B1(n18347), .B2(n18171), .ZN(
        n18162) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18173), .B1(
        n18349), .B2(n18172), .ZN(n18161) );
  OAI211_X1 U21297 ( .C1(n18352), .C2(n18223), .A(n18162), .B(n18161), .ZN(
        P3_U2934) );
  AOI22_X1 U21298 ( .A1(n18353), .A2(n18171), .B1(n18355), .B2(n18172), .ZN(
        n18164) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18173), .B1(
        n18280), .B2(n18241), .ZN(n18163) );
  OAI211_X1 U21300 ( .C1(n18283), .C2(n18176), .A(n18164), .B(n18163), .ZN(
        P3_U2935) );
  AOI22_X1 U21301 ( .A1(n18360), .A2(n18172), .B1(n18359), .B2(n18171), .ZN(
        n18166) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18173), .B1(
        n18361), .B2(n18195), .ZN(n18165) );
  OAI211_X1 U21303 ( .C1(n18364), .C2(n18223), .A(n18166), .B(n18165), .ZN(
        P3_U2936) );
  AOI22_X1 U21304 ( .A1(n18367), .A2(n18172), .B1(n18365), .B2(n18171), .ZN(
        n18168) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18173), .B1(
        n18366), .B2(n18195), .ZN(n18167) );
  OAI211_X1 U21306 ( .C1(n18370), .C2(n18223), .A(n18168), .B(n18167), .ZN(
        P3_U2937) );
  AOI22_X1 U21307 ( .A1(n18372), .A2(n18172), .B1(n18371), .B2(n18171), .ZN(
        n18170) );
  AOI22_X1 U21308 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18173), .B1(
        n18373), .B2(n18195), .ZN(n18169) );
  OAI211_X1 U21309 ( .C1(n18376), .C2(n18223), .A(n18170), .B(n18169), .ZN(
        P3_U2938) );
  AOI22_X1 U21310 ( .A1(n18382), .A2(n18172), .B1(n18378), .B2(n18171), .ZN(
        n18175) );
  AOI22_X1 U21311 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18173), .B1(
        n18322), .B2(n18241), .ZN(n18174) );
  OAI211_X1 U21312 ( .C1(n18327), .C2(n18176), .A(n18175), .B(n18174), .ZN(
        P3_U2939) );
  INV_X1 U21313 ( .A(n18200), .ZN(n18178) );
  NOR2_X2 U21314 ( .A1(n18177), .A2(n18178), .ZN(n18264) );
  INV_X1 U21315 ( .A(n18264), .ZN(n18194) );
  NOR2_X1 U21316 ( .A1(n18178), .A2(n18268), .ZN(n18225) );
  AOI22_X1 U21317 ( .A1(n18331), .A2(n18219), .B1(n18330), .B2(n18225), .ZN(
        n18181) );
  AOI22_X1 U21318 ( .A1(n18273), .A2(n18179), .B1(n18200), .B2(n18270), .ZN(
        n18196) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18196), .B1(
        n18335), .B2(n18195), .ZN(n18180) );
  OAI211_X1 U21320 ( .C1(n18338), .C2(n18194), .A(n18181), .B(n18180), .ZN(
        P3_U2940) );
  AOI22_X1 U21321 ( .A1(n18304), .A2(n18219), .B1(n18340), .B2(n18225), .ZN(
        n18183) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18196), .B1(
        n18339), .B2(n18195), .ZN(n18182) );
  OAI211_X1 U21323 ( .C1(n18307), .C2(n18194), .A(n18183), .B(n18182), .ZN(
        P3_U2941) );
  AOI22_X1 U21324 ( .A1(n18349), .A2(n18195), .B1(n18347), .B2(n18225), .ZN(
        n18185) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18196), .B1(
        n18348), .B2(n18219), .ZN(n18184) );
  OAI211_X1 U21326 ( .C1(n18352), .C2(n18194), .A(n18185), .B(n18184), .ZN(
        P3_U2942) );
  AOI22_X1 U21327 ( .A1(n18353), .A2(n18225), .B1(n18355), .B2(n18195), .ZN(
        n18187) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18196), .B1(
        n18280), .B2(n18264), .ZN(n18186) );
  OAI211_X1 U21329 ( .C1(n18283), .C2(n18199), .A(n18187), .B(n18186), .ZN(
        P3_U2943) );
  AOI22_X1 U21330 ( .A1(n18359), .A2(n18225), .B1(n18361), .B2(n18219), .ZN(
        n18189) );
  AOI22_X1 U21331 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18196), .B1(
        n18360), .B2(n18195), .ZN(n18188) );
  OAI211_X1 U21332 ( .C1(n18364), .C2(n18194), .A(n18189), .B(n18188), .ZN(
        P3_U2944) );
  AOI22_X1 U21333 ( .A1(n18366), .A2(n18219), .B1(n18365), .B2(n18225), .ZN(
        n18191) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18196), .B1(
        n18367), .B2(n18195), .ZN(n18190) );
  OAI211_X1 U21335 ( .C1(n18370), .C2(n18194), .A(n18191), .B(n18190), .ZN(
        P3_U2945) );
  AOI22_X1 U21336 ( .A1(n18372), .A2(n18195), .B1(n18371), .B2(n18225), .ZN(
        n18193) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18196), .B1(
        n18373), .B2(n18219), .ZN(n18192) );
  OAI211_X1 U21338 ( .C1(n18376), .C2(n18194), .A(n18193), .B(n18192), .ZN(
        P3_U2946) );
  AOI22_X1 U21339 ( .A1(n18382), .A2(n18195), .B1(n18378), .B2(n18225), .ZN(
        n18198) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18196), .B1(
        n18322), .B2(n18264), .ZN(n18197) );
  OAI211_X1 U21341 ( .C1(n18327), .C2(n18199), .A(n18198), .B(n18197), .ZN(
        P3_U2947) );
  NAND2_X1 U21342 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18200), .ZN(
        n18224) );
  NOR2_X1 U21343 ( .A1(n18264), .A2(n9562), .ZN(n18246) );
  NOR2_X1 U21344 ( .A1(n18329), .A2(n18246), .ZN(n18218) );
  AOI22_X1 U21345 ( .A1(n18330), .A2(n18218), .B1(n18335), .B2(n18219), .ZN(
        n18204) );
  OAI21_X1 U21346 ( .B1(n18201), .B2(n18245), .A(n18246), .ZN(n18202) );
  OAI211_X1 U21347 ( .C1(n9562), .C2(n18543), .A(n18247), .B(n18202), .ZN(
        n18220) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18220), .B1(
        n18300), .B2(n9562), .ZN(n18203) );
  OAI211_X1 U21349 ( .C1(n18303), .C2(n18223), .A(n18204), .B(n18203), .ZN(
        P3_U2948) );
  INV_X1 U21350 ( .A(n9562), .ZN(n18217) );
  AOI22_X1 U21351 ( .A1(n18304), .A2(n18241), .B1(n18340), .B2(n18218), .ZN(
        n18206) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18220), .B1(
        n18339), .B2(n18219), .ZN(n18205) );
  OAI211_X1 U21353 ( .C1(n18307), .C2(n18217), .A(n18206), .B(n18205), .ZN(
        P3_U2949) );
  AOI22_X1 U21354 ( .A1(n18349), .A2(n18219), .B1(n18347), .B2(n18218), .ZN(
        n18208) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18220), .B1(
        n18348), .B2(n18241), .ZN(n18207) );
  OAI211_X1 U21356 ( .C1(n18352), .C2(n18217), .A(n18208), .B(n18207), .ZN(
        P3_U2950) );
  AOI22_X1 U21357 ( .A1(n18353), .A2(n18218), .B1(n18355), .B2(n18219), .ZN(
        n18210) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18220), .B1(
        n18280), .B2(n9562), .ZN(n18209) );
  OAI211_X1 U21359 ( .C1(n18283), .C2(n18223), .A(n18210), .B(n18209), .ZN(
        P3_U2951) );
  AOI22_X1 U21360 ( .A1(n18359), .A2(n18218), .B1(n18361), .B2(n18241), .ZN(
        n18212) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18220), .B1(
        n18360), .B2(n18219), .ZN(n18211) );
  OAI211_X1 U21362 ( .C1(n18364), .C2(n18217), .A(n18212), .B(n18211), .ZN(
        P3_U2952) );
  AOI22_X1 U21363 ( .A1(n18367), .A2(n18219), .B1(n18365), .B2(n18218), .ZN(
        n18214) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18220), .B1(
        n18366), .B2(n18241), .ZN(n18213) );
  OAI211_X1 U21365 ( .C1(n18370), .C2(n18217), .A(n18214), .B(n18213), .ZN(
        P3_U2953) );
  AOI22_X1 U21366 ( .A1(n18373), .A2(n18241), .B1(n18371), .B2(n18218), .ZN(
        n18216) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18220), .B1(
        n18372), .B2(n18219), .ZN(n18215) );
  OAI211_X1 U21368 ( .C1(n18376), .C2(n18217), .A(n18216), .B(n18215), .ZN(
        P3_U2954) );
  AOI22_X1 U21369 ( .A1(n18382), .A2(n18219), .B1(n18378), .B2(n18218), .ZN(
        n18222) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18220), .B1(
        n18322), .B2(n9562), .ZN(n18221) );
  OAI211_X1 U21371 ( .C1(n18327), .C2(n18223), .A(n18222), .B(n18221), .ZN(
        P3_U2955) );
  INV_X1 U21372 ( .A(n18224), .ZN(n18272) );
  NAND2_X1 U21373 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18272), .ZN(
        n18295) );
  NOR2_X1 U21374 ( .A1(n18329), .A2(n18224), .ZN(n18240) );
  AOI22_X1 U21375 ( .A1(n18330), .A2(n18240), .B1(n18335), .B2(n18241), .ZN(
        n18227) );
  AOI22_X1 U21376 ( .A1(n18273), .A2(n18225), .B1(n18272), .B2(n18332), .ZN(
        n18242) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18242), .B1(
        n18331), .B2(n18264), .ZN(n18226) );
  OAI211_X1 U21378 ( .C1(n18338), .C2(n18295), .A(n18227), .B(n18226), .ZN(
        P3_U2956) );
  AOI22_X1 U21379 ( .A1(n18304), .A2(n18264), .B1(n18340), .B2(n18240), .ZN(
        n18229) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18242), .B1(
        n18339), .B2(n18241), .ZN(n18228) );
  OAI211_X1 U21381 ( .C1(n18307), .C2(n18295), .A(n18229), .B(n18228), .ZN(
        P3_U2957) );
  AOI22_X1 U21382 ( .A1(n18349), .A2(n18241), .B1(n18347), .B2(n18240), .ZN(
        n18231) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18242), .B1(
        n18348), .B2(n18264), .ZN(n18230) );
  OAI211_X1 U21384 ( .C1(n18352), .C2(n18295), .A(n18231), .B(n18230), .ZN(
        P3_U2958) );
  AOI22_X1 U21385 ( .A1(n18353), .A2(n18240), .B1(n18355), .B2(n18241), .ZN(
        n18233) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18242), .B1(
        n18354), .B2(n18264), .ZN(n18232) );
  OAI211_X1 U21387 ( .C1(n18358), .C2(n18295), .A(n18233), .B(n18232), .ZN(
        P3_U2959) );
  AOI22_X1 U21388 ( .A1(n18359), .A2(n18240), .B1(n18361), .B2(n18264), .ZN(
        n18235) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18242), .B1(
        n18360), .B2(n18241), .ZN(n18234) );
  OAI211_X1 U21390 ( .C1(n18364), .C2(n18295), .A(n18235), .B(n18234), .ZN(
        P3_U2960) );
  AOI22_X1 U21391 ( .A1(n18367), .A2(n18241), .B1(n18365), .B2(n18240), .ZN(
        n18237) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18242), .B1(
        n18366), .B2(n18264), .ZN(n18236) );
  OAI211_X1 U21393 ( .C1(n18370), .C2(n18295), .A(n18237), .B(n18236), .ZN(
        P3_U2961) );
  AOI22_X1 U21394 ( .A1(n18373), .A2(n18264), .B1(n18371), .B2(n18240), .ZN(
        n18239) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18242), .B1(
        n18372), .B2(n18241), .ZN(n18238) );
  OAI211_X1 U21396 ( .C1(n18376), .C2(n18295), .A(n18239), .B(n18238), .ZN(
        P3_U2962) );
  AOI22_X1 U21397 ( .A1(n18380), .A2(n18264), .B1(n18378), .B2(n18240), .ZN(
        n18244) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18242), .B1(
        n18382), .B2(n18241), .ZN(n18243) );
  OAI211_X1 U21399 ( .C1(n18387), .C2(n18295), .A(n18244), .B(n18243), .ZN(
        P3_U2963) );
  NAND2_X1 U21400 ( .A1(n18408), .A2(n18271), .ZN(n18326) );
  AOI21_X1 U21401 ( .B1(n18326), .B2(n18295), .A(n18329), .ZN(n18263) );
  AOI22_X1 U21402 ( .A1(n18331), .A2(n9562), .B1(n18330), .B2(n18263), .ZN(
        n18250) );
  INV_X1 U21403 ( .A(n18326), .ZN(n18381) );
  AOI221_X1 U21404 ( .B1(n18246), .B2(n18295), .C1(n18245), .C2(n18295), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18248) );
  OAI21_X1 U21405 ( .B1(n18381), .B2(n18248), .A(n18247), .ZN(n18265) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18265), .B1(
        n18335), .B2(n18264), .ZN(n18249) );
  OAI211_X1 U21407 ( .C1(n18338), .C2(n18326), .A(n18250), .B(n18249), .ZN(
        P3_U2964) );
  AOI22_X1 U21408 ( .A1(n18304), .A2(n9562), .B1(n18340), .B2(n18263), .ZN(
        n18252) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18265), .B1(
        n18339), .B2(n18264), .ZN(n18251) );
  OAI211_X1 U21410 ( .C1(n18307), .C2(n18326), .A(n18252), .B(n18251), .ZN(
        P3_U2965) );
  AOI22_X1 U21411 ( .A1(n18349), .A2(n18264), .B1(n18347), .B2(n18263), .ZN(
        n18254) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18265), .B1(
        n18348), .B2(n9562), .ZN(n18253) );
  OAI211_X1 U21413 ( .C1(n18352), .C2(n18326), .A(n18254), .B(n18253), .ZN(
        P3_U2966) );
  AOI22_X1 U21414 ( .A1(n18354), .A2(n9562), .B1(n18353), .B2(n18263), .ZN(
        n18256) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18265), .B1(
        n18355), .B2(n18264), .ZN(n18255) );
  OAI211_X1 U21416 ( .C1(n18358), .C2(n18326), .A(n18256), .B(n18255), .ZN(
        P3_U2967) );
  AOI22_X1 U21417 ( .A1(n18360), .A2(n18264), .B1(n18359), .B2(n18263), .ZN(
        n18258) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18265), .B1(
        n18361), .B2(n9562), .ZN(n18257) );
  OAI211_X1 U21419 ( .C1(n18364), .C2(n18326), .A(n18258), .B(n18257), .ZN(
        P3_U2968) );
  AOI22_X1 U21420 ( .A1(n18366), .A2(n9562), .B1(n18365), .B2(n18263), .ZN(
        n18260) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18265), .B1(
        n18367), .B2(n18264), .ZN(n18259) );
  OAI211_X1 U21422 ( .C1(n18370), .C2(n18326), .A(n18260), .B(n18259), .ZN(
        P3_U2969) );
  AOI22_X1 U21423 ( .A1(n18373), .A2(n9562), .B1(n18371), .B2(n18263), .ZN(
        n18262) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18265), .B1(
        n18372), .B2(n18264), .ZN(n18261) );
  OAI211_X1 U21425 ( .C1(n18376), .C2(n18326), .A(n18262), .B(n18261), .ZN(
        P3_U2970) );
  AOI22_X1 U21426 ( .A1(n18380), .A2(n9562), .B1(n18378), .B2(n18263), .ZN(
        n18267) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18265), .B1(
        n18382), .B2(n18264), .ZN(n18266) );
  OAI211_X1 U21428 ( .C1(n18387), .C2(n18326), .A(n18267), .B(n18266), .ZN(
        P3_U2971) );
  INV_X1 U21429 ( .A(n18295), .ZN(n18320) );
  INV_X1 U21430 ( .A(n18271), .ZN(n18269) );
  NOR2_X1 U21431 ( .A1(n18269), .A2(n18268), .ZN(n18334) );
  AOI22_X1 U21432 ( .A1(n18331), .A2(n18320), .B1(n18330), .B2(n18334), .ZN(
        n18275) );
  AOI22_X1 U21433 ( .A1(n18273), .A2(n18272), .B1(n18271), .B2(n18270), .ZN(
        n18291) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18291), .B1(
        n18335), .B2(n9562), .ZN(n18274) );
  OAI211_X1 U21435 ( .C1(n18338), .C2(n18345), .A(n18275), .B(n18274), .ZN(
        P3_U2972) );
  AOI22_X1 U21436 ( .A1(n18304), .A2(n18320), .B1(n18340), .B2(n18334), .ZN(
        n18277) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18291), .B1(
        n18339), .B2(n9562), .ZN(n18276) );
  OAI211_X1 U21438 ( .C1(n18307), .C2(n18345), .A(n18277), .B(n18276), .ZN(
        P3_U2973) );
  AOI22_X1 U21439 ( .A1(n18349), .A2(n9562), .B1(n18347), .B2(n18334), .ZN(
        n18279) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18291), .B1(
        n18348), .B2(n18320), .ZN(n18278) );
  OAI211_X1 U21441 ( .C1(n18352), .C2(n18345), .A(n18279), .B(n18278), .ZN(
        P3_U2974) );
  AOI22_X1 U21442 ( .A1(n18353), .A2(n18334), .B1(n18355), .B2(n9562), .ZN(
        n18282) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18291), .B1(
        n18280), .B2(n18379), .ZN(n18281) );
  OAI211_X1 U21444 ( .C1(n18283), .C2(n18295), .A(n18282), .B(n18281), .ZN(
        P3_U2975) );
  AOI22_X1 U21445 ( .A1(n18359), .A2(n18334), .B1(n18361), .B2(n18320), .ZN(
        n18285) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18291), .B1(
        n18360), .B2(n9562), .ZN(n18284) );
  OAI211_X1 U21447 ( .C1(n18364), .C2(n18345), .A(n18285), .B(n18284), .ZN(
        P3_U2976) );
  AOI22_X1 U21448 ( .A1(n18367), .A2(n9562), .B1(n18365), .B2(n18334), .ZN(
        n18287) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18291), .B1(
        n18366), .B2(n18320), .ZN(n18286) );
  OAI211_X1 U21450 ( .C1(n18370), .C2(n18345), .A(n18287), .B(n18286), .ZN(
        P3_U2977) );
  AOI22_X1 U21451 ( .A1(n18373), .A2(n18320), .B1(n18371), .B2(n18334), .ZN(
        n18290) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18291), .B1(
        n18372), .B2(n9562), .ZN(n18289) );
  OAI211_X1 U21453 ( .C1(n18376), .C2(n18345), .A(n18290), .B(n18289), .ZN(
        P3_U2978) );
  AOI22_X1 U21454 ( .A1(n18380), .A2(n18320), .B1(n18378), .B2(n18334), .ZN(
        n18293) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18291), .B1(
        n18382), .B2(n9562), .ZN(n18292) );
  OAI211_X1 U21456 ( .C1(n18387), .C2(n18345), .A(n18293), .B(n18292), .ZN(
        P3_U2979) );
  AND2_X1 U21457 ( .A1(n18294), .A2(n18299), .ZN(n18319) );
  AOI22_X1 U21458 ( .A1(n18330), .A2(n18319), .B1(n18335), .B2(n18320), .ZN(
        n18302) );
  NAND2_X1 U21459 ( .A1(n18326), .A2(n18295), .ZN(n18297) );
  OAI221_X1 U21460 ( .B1(n18299), .B2(n18298), .C1(n18299), .C2(n18297), .A(
        n18296), .ZN(n18323) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18323), .B1(
        n18300), .B2(n18321), .ZN(n18301) );
  OAI211_X1 U21462 ( .C1(n18303), .C2(n18326), .A(n18302), .B(n18301), .ZN(
        P3_U2980) );
  AOI22_X1 U21463 ( .A1(n18304), .A2(n18381), .B1(n18340), .B2(n18319), .ZN(
        n18306) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18323), .B1(
        n18339), .B2(n18320), .ZN(n18305) );
  OAI211_X1 U21465 ( .C1(n18307), .C2(n18318), .A(n18306), .B(n18305), .ZN(
        P3_U2981) );
  AOI22_X1 U21466 ( .A1(n18349), .A2(n18320), .B1(n18347), .B2(n18319), .ZN(
        n18309) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18323), .B1(
        n18348), .B2(n18381), .ZN(n18308) );
  OAI211_X1 U21468 ( .C1(n18352), .C2(n18318), .A(n18309), .B(n18308), .ZN(
        P3_U2982) );
  AOI22_X1 U21469 ( .A1(n18354), .A2(n18381), .B1(n18353), .B2(n18319), .ZN(
        n18311) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18323), .B1(
        n18355), .B2(n18320), .ZN(n18310) );
  OAI211_X1 U21471 ( .C1(n18358), .C2(n18318), .A(n18311), .B(n18310), .ZN(
        P3_U2983) );
  AOI22_X1 U21472 ( .A1(n18359), .A2(n18319), .B1(n18361), .B2(n18381), .ZN(
        n18313) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18323), .B1(
        n18360), .B2(n18320), .ZN(n18312) );
  OAI211_X1 U21474 ( .C1(n18364), .C2(n18318), .A(n18313), .B(n18312), .ZN(
        P3_U2984) );
  AOI22_X1 U21475 ( .A1(n18367), .A2(n18320), .B1(n18365), .B2(n18319), .ZN(
        n18315) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18323), .B1(
        n18366), .B2(n18381), .ZN(n18314) );
  OAI211_X1 U21477 ( .C1(n18370), .C2(n18318), .A(n18315), .B(n18314), .ZN(
        P3_U2985) );
  AOI22_X1 U21478 ( .A1(n18372), .A2(n18320), .B1(n18371), .B2(n18319), .ZN(
        n18317) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18323), .B1(
        n18373), .B2(n18381), .ZN(n18316) );
  OAI211_X1 U21480 ( .C1(n18376), .C2(n18318), .A(n18317), .B(n18316), .ZN(
        P3_U2986) );
  AOI22_X1 U21481 ( .A1(n18382), .A2(n18320), .B1(n18378), .B2(n18319), .ZN(
        n18325) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18323), .B1(
        n18322), .B2(n18321), .ZN(n18324) );
  OAI211_X1 U21483 ( .C1(n18327), .C2(n18326), .A(n18325), .B(n18324), .ZN(
        P3_U2987) );
  NOR2_X1 U21484 ( .A1(n18329), .A2(n18328), .ZN(n18377) );
  AOI22_X1 U21485 ( .A1(n18331), .A2(n18379), .B1(n18330), .B2(n18377), .ZN(
        n18337) );
  AOI22_X1 U21486 ( .A1(n18273), .A2(n18334), .B1(n18333), .B2(n18332), .ZN(
        n18383) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18383), .B1(
        n18335), .B2(n18381), .ZN(n18336) );
  OAI211_X1 U21488 ( .C1(n18338), .C2(n18386), .A(n18337), .B(n18336), .ZN(
        P3_U2988) );
  AOI22_X1 U21489 ( .A1(n18340), .A2(n18377), .B1(n18339), .B2(n18381), .ZN(
        n18344) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18383), .B1(
        n18342), .B2(n18341), .ZN(n18343) );
  OAI211_X1 U21491 ( .C1(n18346), .C2(n18345), .A(n18344), .B(n18343), .ZN(
        P3_U2989) );
  AOI22_X1 U21492 ( .A1(n18348), .A2(n18379), .B1(n18347), .B2(n18377), .ZN(
        n18351) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18383), .B1(
        n18349), .B2(n18381), .ZN(n18350) );
  OAI211_X1 U21494 ( .C1(n18352), .C2(n18386), .A(n18351), .B(n18350), .ZN(
        P3_U2990) );
  AOI22_X1 U21495 ( .A1(n18354), .A2(n18379), .B1(n18353), .B2(n18377), .ZN(
        n18357) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18383), .B1(
        n18355), .B2(n18381), .ZN(n18356) );
  OAI211_X1 U21497 ( .C1(n18358), .C2(n18386), .A(n18357), .B(n18356), .ZN(
        P3_U2991) );
  AOI22_X1 U21498 ( .A1(n18360), .A2(n18381), .B1(n18359), .B2(n18377), .ZN(
        n18363) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18383), .B1(
        n18361), .B2(n18379), .ZN(n18362) );
  OAI211_X1 U21500 ( .C1(n18364), .C2(n18386), .A(n18363), .B(n18362), .ZN(
        P3_U2992) );
  AOI22_X1 U21501 ( .A1(n18366), .A2(n18379), .B1(n18365), .B2(n18377), .ZN(
        n18369) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18383), .B1(
        n18367), .B2(n18381), .ZN(n18368) );
  OAI211_X1 U21503 ( .C1(n18370), .C2(n18386), .A(n18369), .B(n18368), .ZN(
        P3_U2993) );
  AOI22_X1 U21504 ( .A1(n18372), .A2(n18381), .B1(n18371), .B2(n18377), .ZN(
        n18375) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18383), .B1(
        n18373), .B2(n18379), .ZN(n18374) );
  OAI211_X1 U21506 ( .C1(n18376), .C2(n18386), .A(n18375), .B(n18374), .ZN(
        P3_U2994) );
  AOI22_X1 U21507 ( .A1(n18380), .A2(n18379), .B1(n18378), .B2(n18377), .ZN(
        n18385) );
  AOI22_X1 U21508 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18383), .B1(
        n18382), .B2(n18381), .ZN(n18384) );
  OAI211_X1 U21509 ( .C1(n18387), .C2(n18386), .A(n18385), .B(n18384), .ZN(
        P3_U2995) );
  NOR2_X1 U21510 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18441) );
  AOI21_X1 U21511 ( .B1(n18390), .B2(n18389), .A(n18388), .ZN(n18391) );
  INV_X1 U21512 ( .A(n18391), .ZN(n18419) );
  AND3_X1 U21513 ( .A1(n18392), .A2(n18419), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18398) );
  INV_X1 U21514 ( .A(n18415), .ZN(n18393) );
  AOI211_X1 U21515 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18395), .A(
        n18394), .B(n18393), .ZN(n18401) );
  AOI211_X1 U21516 ( .C1(n18560), .C2(n18568), .A(n18401), .B(n18396), .ZN(
        n18397) );
  AOI211_X1 U21517 ( .C1(n18411), .C2(n18554), .A(n18398), .B(n18397), .ZN(
        n18557) );
  MUX2_X1 U21518 ( .A(n18560), .B(n18557), .S(n18422), .Z(n18423) );
  NAND2_X1 U21519 ( .A1(n9569), .A2(n18399), .ZN(n18402) );
  INV_X1 U21520 ( .A(n18401), .ZN(n18412) );
  AOI22_X1 U21521 ( .A1(n18565), .A2(n18402), .B1(n18568), .B2(n18412), .ZN(
        n18561) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18403), .B1(
        n18402), .B2(n18575), .ZN(n18406) );
  INV_X1 U21523 ( .A(n18406), .ZN(n18570) );
  NOR3_X1 U21524 ( .A1(n18405), .A2(n18404), .A3(n18570), .ZN(n18407) );
  OAI22_X1 U21525 ( .A1(n18561), .A2(n18407), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18406), .ZN(n18409) );
  AOI21_X1 U21526 ( .B1(n18409), .B2(n18422), .A(n18408), .ZN(n18410) );
  AOI222_X1 U21527 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18423), 
        .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18410), .C1(n18423), 
        .C2(n18410), .ZN(n18440) );
  AOI22_X1 U21528 ( .A1(n18396), .A2(n18412), .B1(n18411), .B2(n18416), .ZN(
        n18413) );
  NOR2_X1 U21529 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18413), .ZN(
        n18548) );
  AOI21_X1 U21530 ( .B1(n18415), .B2(n18414), .A(n18396), .ZN(n18418) );
  INV_X1 U21531 ( .A(n18416), .ZN(n18417) );
  AOI211_X1 U21532 ( .C1(n18420), .C2(n18419), .A(n18418), .B(n18417), .ZN(
        n18545) );
  AOI21_X1 U21533 ( .B1(n18545), .B2(n18422), .A(n18551), .ZN(n18421) );
  AOI21_X1 U21534 ( .B1(n18422), .B2(n18548), .A(n18421), .ZN(n18437) );
  INV_X1 U21535 ( .A(n18423), .ZN(n18424) );
  AOI221_X1 U21536 ( .B1(n18440), .B2(n18426), .C1(n18425), .C2(n18426), .A(
        n18424), .ZN(n18436) );
  AOI221_X1 U21537 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n18428), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n18428), .A(n18427), .ZN(n18435) );
  OAI22_X1 U21538 ( .A1(n18431), .A2(n18430), .B1(n18591), .B2(n18429), .ZN(
        n18592) );
  AOI211_X1 U21539 ( .C1(n18433), .C2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18432), .B(n18592), .ZN(n18434) );
  OAI211_X1 U21540 ( .C1(n18437), .C2(n18436), .A(n18435), .B(n18434), .ZN(
        n18438) );
  AOI211_X1 U21541 ( .C1(n18441), .C2(n18440), .A(n18439), .B(n18438), .ZN(
        n18451) );
  INV_X1 U21542 ( .A(n18602), .ZN(n18458) );
  AOI22_X1 U21543 ( .A1(n18569), .A2(n18458), .B1(n18600), .B2(n18609), .ZN(
        n18448) );
  INV_X1 U21544 ( .A(n18451), .ZN(n18442) );
  AOI211_X1 U21545 ( .C1(n18444), .C2(n18443), .A(n18450), .B(n18442), .ZN(
        n18445) );
  NOR2_X1 U21546 ( .A1(n18445), .A2(n18603), .ZN(n18544) );
  OAI211_X1 U21547 ( .C1(P3_STATE2_REG_2__SCAN_IN), .C2(n18608), .A(n18544), 
        .B(n18446), .ZN(n18454) );
  OAI22_X1 U21548 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18448), .B1(n18447), 
        .B2(n18454), .ZN(n18449) );
  OAI21_X1 U21549 ( .B1(n18451), .B2(n18450), .A(n18449), .ZN(P3_U2996) );
  NOR4_X1 U21550 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18553), .A3(n18603), 
        .A4(n18608), .ZN(n18456) );
  AOI211_X1 U21551 ( .C1(n18600), .C2(n18609), .A(n18452), .B(n18456), .ZN(
        n18453) );
  OAI21_X1 U21552 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18454), .A(n18453), 
        .ZN(P3_U2997) );
  NOR4_X1 U21553 ( .A1(n18458), .A2(n18457), .A3(n18456), .A4(n18455), .ZN(
        P3_U2998) );
  AND2_X1 U21554 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18459), .ZN(
        P3_U2999) );
  AND2_X1 U21555 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18459), .ZN(
        P3_U3000) );
  AND2_X1 U21556 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18459), .ZN(
        P3_U3001) );
  AND2_X1 U21557 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18459), .ZN(
        P3_U3002) );
  AND2_X1 U21558 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18459), .ZN(
        P3_U3003) );
  AND2_X1 U21559 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18459), .ZN(
        P3_U3004) );
  AND2_X1 U21560 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18459), .ZN(
        P3_U3005) );
  AND2_X1 U21561 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18459), .ZN(
        P3_U3006) );
  AND2_X1 U21562 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18459), .ZN(
        P3_U3007) );
  AND2_X1 U21563 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18459), .ZN(
        P3_U3008) );
  AND2_X1 U21564 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18459), .ZN(
        P3_U3009) );
  AND2_X1 U21565 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18459), .ZN(
        P3_U3010) );
  AND2_X1 U21566 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18459), .ZN(
        P3_U3011) );
  NOR2_X1 U21567 ( .A1(n20780), .A2(n18541), .ZN(P3_U3012) );
  AND2_X1 U21568 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18459), .ZN(
        P3_U3013) );
  AND2_X1 U21569 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18459), .ZN(
        P3_U3014) );
  AND2_X1 U21570 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18459), .ZN(
        P3_U3015) );
  AND2_X1 U21571 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18459), .ZN(
        P3_U3016) );
  AND2_X1 U21572 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18459), .ZN(
        P3_U3017) );
  NOR2_X1 U21573 ( .A1(n20678), .A2(n18541), .ZN(P3_U3018) );
  AND2_X1 U21574 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18459), .ZN(
        P3_U3019) );
  AND2_X1 U21575 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18459), .ZN(
        P3_U3020) );
  AND2_X1 U21576 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18459), .ZN(P3_U3021) );
  AND2_X1 U21577 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18459), .ZN(P3_U3022) );
  AND2_X1 U21578 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18459), .ZN(P3_U3023) );
  AND2_X1 U21579 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18459), .ZN(P3_U3024) );
  AND2_X1 U21580 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18459), .ZN(P3_U3025) );
  AND2_X1 U21581 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18459), .ZN(P3_U3026) );
  AND2_X1 U21582 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18459), .ZN(P3_U3027) );
  AND2_X1 U21583 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18459), .ZN(P3_U3028) );
  INV_X1 U21584 ( .A(n18460), .ZN(n18461) );
  INV_X1 U21585 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18465) );
  AOI21_X1 U21586 ( .B1(HOLD), .B2(n18461), .A(n18465), .ZN(n18464) );
  NAND2_X1 U21587 ( .A1(n18600), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18471) );
  INV_X1 U21588 ( .A(n18471), .ZN(n18466) );
  NOR2_X1 U21589 ( .A1(n18466), .A2(n18475), .ZN(n18477) );
  INV_X1 U21590 ( .A(NA), .ZN(n20587) );
  OAI21_X1 U21591 ( .B1(n20587), .B2(n18462), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18476) );
  INV_X1 U21592 ( .A(n18476), .ZN(n18463) );
  OAI22_X1 U21593 ( .A1(n18532), .A2(n18464), .B1(n18477), .B2(n18463), .ZN(
        P3_U3029) );
  NOR2_X1 U21594 ( .A1(n18478), .A2(n20581), .ZN(n18473) );
  NOR3_X1 U21595 ( .A1(n18473), .A2(n18465), .A3(n18475), .ZN(n18467) );
  NOR2_X1 U21596 ( .A1(n18467), .A2(n18466), .ZN(n18469) );
  OAI211_X1 U21597 ( .C1(n20581), .C2(n18470), .A(n18469), .B(n18468), .ZN(
        P3_U3030) );
  OAI22_X1 U21598 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18471), .ZN(n18472) );
  OAI22_X1 U21599 ( .A1(n18473), .A2(n18472), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18474) );
  OAI22_X1 U21600 ( .A1(n18477), .A2(n18476), .B1(n18475), .B2(n18474), .ZN(
        P3_U3031) );
  NAND2_X1 U21601 ( .A1(n18532), .A2(n18478), .ZN(n18528) );
  CLKBUF_X1 U21602 ( .A(n18528), .Z(n18533) );
  OAI222_X1 U21603 ( .A1(n18587), .A2(n18537), .B1(n20727), .B2(n18532), .C1(
        n18479), .C2(n18533), .ZN(P3_U3032) );
  OAI222_X1 U21604 ( .A1(n18533), .A2(n18482), .B1(n18480), .B2(n18532), .C1(
        n18479), .C2(n18537), .ZN(P3_U3033) );
  OAI222_X1 U21605 ( .A1(n18482), .A2(n18537), .B1(n18481), .B2(n18532), .C1(
        n18483), .C2(n18533), .ZN(P3_U3034) );
  INV_X1 U21606 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18485) );
  OAI222_X1 U21607 ( .A1(n18528), .A2(n18485), .B1(n18484), .B2(n18532), .C1(
        n18483), .C2(n18537), .ZN(P3_U3035) );
  OAI222_X1 U21608 ( .A1(n18528), .A2(n18487), .B1(n18486), .B2(n18532), .C1(
        n18485), .C2(n18537), .ZN(P3_U3036) );
  OAI222_X1 U21609 ( .A1(n18528), .A2(n18489), .B1(n18488), .B2(n18532), .C1(
        n18487), .C2(n18537), .ZN(P3_U3037) );
  OAI222_X1 U21610 ( .A1(n18528), .A2(n18491), .B1(n18490), .B2(n18532), .C1(
        n18489), .C2(n18537), .ZN(P3_U3038) );
  OAI222_X1 U21611 ( .A1(n18528), .A2(n18493), .B1(n18492), .B2(n18532), .C1(
        n18491), .C2(n18537), .ZN(P3_U3039) );
  OAI222_X1 U21612 ( .A1(n18533), .A2(n18495), .B1(n18494), .B2(n18532), .C1(
        n18493), .C2(n18537), .ZN(P3_U3040) );
  OAI222_X1 U21613 ( .A1(n18533), .A2(n18497), .B1(n18496), .B2(n18532), .C1(
        n18495), .C2(n18537), .ZN(P3_U3041) );
  INV_X1 U21614 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20712) );
  OAI222_X1 U21615 ( .A1(n18533), .A2(n20712), .B1(n18498), .B2(n18532), .C1(
        n18497), .C2(n18537), .ZN(P3_U3042) );
  OAI222_X1 U21616 ( .A1(n20712), .A2(n18537), .B1(n20700), .B2(n18532), .C1(
        n20814), .C2(n18533), .ZN(P3_U3043) );
  OAI222_X1 U21617 ( .A1(n20814), .A2(n18537), .B1(n18499), .B2(n18532), .C1(
        n18501), .C2(n18533), .ZN(P3_U3044) );
  OAI222_X1 U21618 ( .A1(n18501), .A2(n18537), .B1(n18500), .B2(n18532), .C1(
        n18502), .C2(n18533), .ZN(P3_U3045) );
  OAI222_X1 U21619 ( .A1(n18533), .A2(n18504), .B1(n18503), .B2(n18532), .C1(
        n18502), .C2(n18537), .ZN(P3_U3046) );
  OAI222_X1 U21620 ( .A1(n18533), .A2(n18507), .B1(n18505), .B2(n18532), .C1(
        n18504), .C2(n18537), .ZN(P3_U3047) );
  OAI222_X1 U21621 ( .A1(n18507), .A2(n18537), .B1(n18506), .B2(n18532), .C1(
        n18508), .C2(n18533), .ZN(P3_U3048) );
  OAI222_X1 U21622 ( .A1(n18533), .A2(n18510), .B1(n18509), .B2(n18532), .C1(
        n18508), .C2(n18537), .ZN(P3_U3049) );
  OAI222_X1 U21623 ( .A1(n18528), .A2(n18512), .B1(n18511), .B2(n18532), .C1(
        n18510), .C2(n18537), .ZN(P3_U3050) );
  OAI222_X1 U21624 ( .A1(n18528), .A2(n18514), .B1(n18513), .B2(n18532), .C1(
        n18512), .C2(n18537), .ZN(P3_U3051) );
  OAI222_X1 U21625 ( .A1(n18528), .A2(n18516), .B1(n18515), .B2(n18532), .C1(
        n18514), .C2(n18537), .ZN(P3_U3052) );
  OAI222_X1 U21626 ( .A1(n18528), .A2(n18518), .B1(n18517), .B2(n18532), .C1(
        n18516), .C2(n18537), .ZN(P3_U3053) );
  OAI222_X1 U21627 ( .A1(n18528), .A2(n18520), .B1(n18519), .B2(n18532), .C1(
        n18518), .C2(n18537), .ZN(P3_U3054) );
  OAI222_X1 U21628 ( .A1(n18528), .A2(n18522), .B1(n18521), .B2(n18532), .C1(
        n18520), .C2(n18537), .ZN(P3_U3055) );
  OAI222_X1 U21629 ( .A1(n18533), .A2(n18524), .B1(n18523), .B2(n18532), .C1(
        n18522), .C2(n18537), .ZN(P3_U3056) );
  OAI222_X1 U21630 ( .A1(n18533), .A2(n18526), .B1(n18525), .B2(n18532), .C1(
        n18524), .C2(n18537), .ZN(P3_U3057) );
  INV_X1 U21631 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18530) );
  OAI222_X1 U21632 ( .A1(n18528), .A2(n18530), .B1(n18527), .B2(n18532), .C1(
        n18526), .C2(n18537), .ZN(P3_U3058) );
  OAI222_X1 U21633 ( .A1(n18530), .A2(n18537), .B1(n18529), .B2(n18532), .C1(
        n18531), .C2(n18533), .ZN(P3_U3059) );
  OAI222_X1 U21634 ( .A1(n18533), .A2(n18536), .B1(n20722), .B2(n18532), .C1(
        n18531), .C2(n18537), .ZN(P3_U3060) );
  OAI222_X1 U21635 ( .A1(n18537), .A2(n18536), .B1(n18535), .B2(n18532), .C1(
        n18534), .C2(n18533), .ZN(P3_U3061) );
  MUX2_X1 U21636 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n18532), .Z(P3_U3274) );
  MUX2_X1 U21637 ( .A(P3_BE_N_REG_2__SCAN_IN), .B(P3_BYTEENABLE_REG_2__SCAN_IN), .S(n18532), .Z(P3_U3275) );
  MUX2_X1 U21638 ( .A(P3_BE_N_REG_1__SCAN_IN), .B(P3_BYTEENABLE_REG_1__SCAN_IN), .S(n18532), .Z(P3_U3276) );
  MUX2_X1 U21639 ( .A(P3_BE_N_REG_0__SCAN_IN), .B(P3_BYTEENABLE_REG_0__SCAN_IN), .S(n18532), .Z(P3_U3277) );
  OAI21_X1 U21640 ( .B1(n18541), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18539), 
        .ZN(n18538) );
  INV_X1 U21641 ( .A(n18538), .ZN(P3_U3280) );
  INV_X1 U21642 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18540) );
  OAI21_X1 U21643 ( .B1(n18541), .B2(n18540), .A(n18539), .ZN(P3_U3281) );
  OAI21_X1 U21644 ( .B1(n18544), .B2(n18543), .A(n18542), .ZN(P3_U3282) );
  NOR2_X1 U21645 ( .A1(n18545), .A2(n18556), .ZN(n18546) );
  INV_X1 U21646 ( .A(n18573), .ZN(n18576) );
  NOR2_X1 U21647 ( .A1(n18546), .A2(n18576), .ZN(n18550) );
  AOI22_X1 U21648 ( .A1(n18571), .A2(n18548), .B1(n18569), .B2(n18547), .ZN(
        n18549) );
  OAI22_X1 U21649 ( .A1(n18551), .A2(n18550), .B1(n18576), .B2(n18549), .ZN(
        P3_U3285) );
  AOI22_X1 U21650 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n18552), .B2(n20679), .ZN(
        n18562) );
  NOR2_X1 U21651 ( .A1(n18553), .A2(n18572), .ZN(n18563) );
  INV_X1 U21652 ( .A(n18569), .ZN(n18555) );
  OAI22_X1 U21653 ( .A1(n18557), .A2(n18556), .B1(n18555), .B2(n18554), .ZN(
        n18558) );
  AOI21_X1 U21654 ( .B1(n18562), .B2(n18563), .A(n18558), .ZN(n18559) );
  AOI22_X1 U21655 ( .A1(n18576), .A2(n18560), .B1(n18559), .B2(n18573), .ZN(
        P3_U3288) );
  INV_X1 U21656 ( .A(n18561), .ZN(n18566) );
  INV_X1 U21657 ( .A(n18562), .ZN(n18564) );
  AOI222_X1 U21658 ( .A1(n18566), .A2(n18571), .B1(n18569), .B2(n18565), .C1(
        n18564), .C2(n18563), .ZN(n18567) );
  AOI22_X1 U21659 ( .A1(n18576), .A2(n18568), .B1(n18567), .B2(n18573), .ZN(
        P3_U3289) );
  AOI222_X1 U21660 ( .A1(n18572), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18571), 
        .B2(n18570), .C1(n18575), .C2(n18569), .ZN(n18574) );
  AOI22_X1 U21661 ( .A1(n18576), .A2(n18575), .B1(n18574), .B2(n18573), .ZN(
        P3_U3290) );
  NOR2_X1 U21662 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18578) );
  AOI211_X1 U21663 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(n20741), .A(n18578), 
        .B(n18577), .ZN(n18582) );
  NOR2_X1 U21664 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n18587), .ZN(n18580) );
  INV_X1 U21665 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18579) );
  MUX2_X1 U21666 ( .A(n18580), .B(n18579), .S(n18586), .Z(n18581) );
  NOR2_X1 U21667 ( .A1(n18582), .A2(n18581), .ZN(P3_U3292) );
  OAI21_X1 U21668 ( .B1(n18584), .B2(P3_BYTEENABLE_REG_0__SCAN_IN), .A(n18583), 
        .ZN(n18585) );
  OAI21_X1 U21669 ( .B1(n18587), .B2(n18586), .A(n18585), .ZN(P3_U3293) );
  INV_X1 U21670 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18588) );
  AOI22_X1 U21671 ( .A1(n18532), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18588), 
        .B2(n18612), .ZN(P3_U3294) );
  INV_X1 U21672 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n18596) );
  OAI22_X1 U21673 ( .A1(n18591), .A2(n9776), .B1(n18590), .B2(n18589), .ZN(
        n18593) );
  OAI21_X1 U21674 ( .B1(n18593), .B2(n18592), .A(n18595), .ZN(n18594) );
  OAI21_X1 U21675 ( .B1(n18596), .B2(n18595), .A(n18594), .ZN(P3_U3295) );
  OAI21_X1 U21676 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18598), .A(n18597), 
        .ZN(n18601) );
  AOI211_X1 U21677 ( .C1(n18615), .C2(n18601), .A(n18600), .B(n18599), .ZN(
        n18604) );
  OAI21_X1 U21678 ( .B1(n18604), .B2(n18603), .A(n18602), .ZN(n18611) );
  OAI21_X1 U21679 ( .B1(n18606), .B2(n18605), .A(n18616), .ZN(n18607) );
  AOI21_X1 U21680 ( .B1(n18609), .B2(n18608), .A(n18607), .ZN(n18610) );
  MUX2_X1 U21681 ( .A(n18611), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18610), 
        .Z(P3_U3296) );
  INV_X1 U21682 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18613) );
  AOI22_X1 U21683 ( .A1(n18532), .A2(n18613), .B1(n20699), .B2(n18612), .ZN(
        P3_U3297) );
  OAI21_X1 U21684 ( .B1(n18617), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n18616), 
        .ZN(n18614) );
  OAI21_X1 U21685 ( .B1(n18616), .B2(n18615), .A(n18614), .ZN(P3_U3298) );
  NOR2_X1 U21686 ( .A1(n18617), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18619)
         );
  OAI21_X1 U21687 ( .B1(n18620), .B2(n18619), .A(n18618), .ZN(P3_U3299) );
  INV_X1 U21688 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19560) );
  INV_X1 U21689 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18621) );
  NAND2_X1 U21690 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19578), .ZN(n19568) );
  NAND2_X1 U21691 ( .A1(n19560), .A2(n20696), .ZN(n19564) );
  OAI21_X1 U21692 ( .B1(n19560), .B2(n19568), .A(n19564), .ZN(n19631) );
  OAI21_X1 U21693 ( .B1(n19560), .B2(n18621), .A(n19559), .ZN(P2_U2815) );
  INV_X1 U21694 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18624) );
  OAI22_X1 U21695 ( .A1(n18623), .A2(n18624), .B1(n12317), .B2(n18622), .ZN(
        P2_U2816) );
  AOI21_X1 U21696 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n18624), .A(n19572), 
        .ZN(n18626) );
  INV_X1 U21697 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n18625) );
  OAI22_X1 U21698 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n18626), .B1(n19613), 
        .B2(n18625), .ZN(P2_U2817) );
  OAI21_X1 U21699 ( .B1(n19572), .B2(BS16), .A(n19631), .ZN(n19629) );
  OAI21_X1 U21700 ( .B1(n19631), .B2(n19633), .A(n19629), .ZN(P2_U2818) );
  NOR4_X1 U21701 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18630) );
  NOR4_X1 U21702 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18629) );
  NOR4_X1 U21703 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18628) );
  NOR4_X1 U21704 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18627) );
  NAND4_X1 U21705 ( .A1(n18630), .A2(n18629), .A3(n18628), .A4(n18627), .ZN(
        n18636) );
  NOR4_X1 U21706 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18634) );
  AOI211_X1 U21707 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18633) );
  NOR4_X1 U21708 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18632) );
  NOR4_X1 U21709 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18631) );
  NAND4_X1 U21710 ( .A1(n18634), .A2(n18633), .A3(n18632), .A4(n18631), .ZN(
        n18635) );
  NOR2_X1 U21711 ( .A1(n18636), .A2(n18635), .ZN(n18643) );
  INV_X1 U21712 ( .A(n18643), .ZN(n18642) );
  NOR2_X1 U21713 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18642), .ZN(n18637) );
  INV_X1 U21714 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19627) );
  AOI22_X1 U21715 ( .A1(n18637), .A2(n10804), .B1(n18642), .B2(n19627), .ZN(
        P2_U2820) );
  OR3_X1 U21716 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18641) );
  INV_X1 U21717 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19625) );
  AOI22_X1 U21718 ( .A1(n18637), .A2(n18641), .B1(n18642), .B2(n19625), .ZN(
        P2_U2821) );
  INV_X1 U21719 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19630) );
  NAND2_X1 U21720 ( .A1(n18637), .A2(n19630), .ZN(n18640) );
  OAI21_X1 U21721 ( .B1(n10804), .B2(n10240), .A(n18643), .ZN(n18638) );
  OAI21_X1 U21722 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18643), .A(n18638), 
        .ZN(n18639) );
  OAI221_X1 U21723 ( .B1(n18640), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18640), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18639), .ZN(P2_U2822) );
  INV_X1 U21724 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20739) );
  OAI221_X1 U21725 ( .B1(n18643), .B2(n20739), .C1(n18642), .C2(n18641), .A(
        n18640), .ZN(P2_U2823) );
  NOR2_X1 U21726 ( .A1(n18657), .A2(n18656), .ZN(n18655) );
  NOR2_X1 U21727 ( .A1(n18830), .A2(n18655), .ZN(n18645) );
  AOI211_X1 U21728 ( .C1(n18646), .C2(n18645), .A(n18644), .B(n19555), .ZN(
        n18652) );
  AOI22_X1 U21729 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n18853), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n18856), .ZN(n18649) );
  AOI22_X1 U21730 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18838), .B1(
        n18647), .B2(n18852), .ZN(n18648) );
  OAI211_X1 U21731 ( .C1(n18650), .C2(n18842), .A(n18649), .B(n18648), .ZN(
        n18651) );
  AOI211_X1 U21732 ( .C1(n18854), .C2(n18653), .A(n18652), .B(n18651), .ZN(
        n18654) );
  INV_X1 U21733 ( .A(n18654), .ZN(P2_U2835) );
  AOI211_X1 U21734 ( .C1(n18657), .C2(n18656), .A(n18655), .B(n19555), .ZN(
        n18662) );
  AOI21_X1 U21735 ( .B1(P2_REIP_REG_19__SCAN_IN), .B2(n18853), .A(n18980), 
        .ZN(n18659) );
  AOI22_X1 U21736 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18859), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n18856), .ZN(n18658) );
  OAI211_X1 U21737 ( .C1(n18660), .C2(n18810), .A(n18659), .B(n18658), .ZN(
        n18661) );
  AOI211_X1 U21738 ( .C1(n18854), .C2(n18663), .A(n18662), .B(n18661), .ZN(
        n18664) );
  OAI21_X1 U21739 ( .B1(n18665), .B2(n18842), .A(n18664), .ZN(P2_U2836) );
  OAI21_X1 U21740 ( .B1(n19598), .B2(n18792), .A(n19016), .ZN(n18669) );
  OAI22_X1 U21741 ( .A1(n18826), .A2(n18667), .B1(n18666), .B2(n18810), .ZN(
        n18668) );
  AOI211_X1 U21742 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18838), .A(
        n18669), .B(n18668), .ZN(n18675) );
  NOR2_X1 U21743 ( .A1(n18830), .A2(n18670), .ZN(n18683) );
  XNOR2_X1 U21744 ( .A(n18683), .B(n18671), .ZN(n18672) );
  AOI22_X1 U21745 ( .A1(n18673), .A2(n18854), .B1(n18818), .B2(n18672), .ZN(
        n18674) );
  OAI211_X1 U21746 ( .C1(n18676), .C2(n18842), .A(n18675), .B(n18674), .ZN(
        P2_U2837) );
  AOI22_X1 U21747 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18859), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n18856), .ZN(n18677) );
  OAI211_X1 U21748 ( .C1(n10984), .C2(n18792), .A(n18677), .B(n19016), .ZN(
        n18680) );
  NAND2_X1 U21749 ( .A1(n18818), .A2(n18830), .ZN(n18749) );
  OAI22_X1 U21750 ( .A1(n18678), .A2(n18810), .B1(n18684), .B2(n18749), .ZN(
        n18679) );
  AOI211_X1 U21751 ( .C1(n18681), .C2(n18855), .A(n18680), .B(n18679), .ZN(
        n18687) );
  INV_X1 U21752 ( .A(n18682), .ZN(n18685) );
  OAI211_X1 U21753 ( .C1(n18685), .C2(n18684), .A(n18818), .B(n18683), .ZN(
        n18686) );
  OAI211_X1 U21754 ( .C1(n18822), .C2(n18688), .A(n18687), .B(n18686), .ZN(
        P2_U2838) );
  INV_X1 U21755 ( .A(n18689), .ZN(n18690) );
  OAI22_X1 U21756 ( .A1(n18690), .A2(n18810), .B1(n11094), .B2(n18826), .ZN(
        n18691) );
  AOI211_X1 U21757 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18853), .A(n18980), 
        .B(n18691), .ZN(n18700) );
  NOR2_X1 U21758 ( .A1(n18830), .A2(n18692), .ZN(n18693) );
  XNOR2_X1 U21759 ( .A(n18694), .B(n18693), .ZN(n18698) );
  OAI22_X1 U21760 ( .A1(n18696), .A2(n18842), .B1(n18695), .B2(n18822), .ZN(
        n18697) );
  AOI21_X1 U21761 ( .B1(n18698), .B2(n18818), .A(n18697), .ZN(n18699) );
  OAI211_X1 U21762 ( .C1(n18701), .C2(n18742), .A(n18700), .B(n18699), .ZN(
        P2_U2839) );
  NAND2_X1 U21763 ( .A1(n18814), .A2(n18702), .ZN(n18704) );
  XOR2_X1 U21764 ( .A(n18704), .B(n18703), .Z(n18711) );
  AOI22_X1 U21765 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n18856), .B1(n18705), 
        .B2(n18852), .ZN(n18706) );
  OAI211_X1 U21766 ( .C1(n11091), .C2(n18792), .A(n18706), .B(n19016), .ZN(
        n18709) );
  OAI22_X1 U21767 ( .A1(n18707), .A2(n18822), .B1(n18871), .B2(n18842), .ZN(
        n18708) );
  AOI211_X1 U21768 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18838), .A(
        n18709), .B(n18708), .ZN(n18710) );
  OAI21_X1 U21769 ( .B1(n18711), .B2(n19555), .A(n18710), .ZN(P2_U2840) );
  AOI22_X1 U21770 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18859), .B1(
        n18712), .B2(n18852), .ZN(n18713) );
  OAI211_X1 U21771 ( .C1(n10962), .C2(n18792), .A(n18713), .B(n19016), .ZN(
        n18714) );
  AOI21_X1 U21772 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n18856), .A(n18714), .ZN(
        n18721) );
  NOR2_X1 U21773 ( .A1(n18830), .A2(n18715), .ZN(n18717) );
  XNOR2_X1 U21774 ( .A(n18717), .B(n18716), .ZN(n18718) );
  AOI22_X1 U21775 ( .A1(n18719), .A2(n18854), .B1(n18818), .B2(n18718), .ZN(
        n18720) );
  OAI211_X1 U21776 ( .C1(n18873), .C2(n18842), .A(n18721), .B(n18720), .ZN(
        P2_U2841) );
  NAND2_X1 U21777 ( .A1(n18814), .A2(n18722), .ZN(n18723) );
  XOR2_X1 U21778 ( .A(n18724), .B(n18723), .Z(n18731) );
  AOI22_X1 U21779 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18859), .B1(
        n18725), .B2(n18852), .ZN(n18726) );
  OAI211_X1 U21780 ( .C1(n10936), .C2(n18792), .A(n18726), .B(n19016), .ZN(
        n18727) );
  AOI21_X1 U21781 ( .B1(P2_EBX_REG_13__SCAN_IN), .B2(n18856), .A(n18727), .ZN(
        n18730) );
  AOI22_X1 U21782 ( .A1(n18728), .A2(n18854), .B1(n18876), .B2(n18855), .ZN(
        n18729) );
  OAI211_X1 U21783 ( .C1(n19555), .C2(n18731), .A(n18730), .B(n18729), .ZN(
        P2_U2842) );
  INV_X1 U21784 ( .A(n18737), .ZN(n18732) );
  AOI211_X1 U21785 ( .C1(n18814), .C2(n18732), .A(n19555), .B(n18738), .ZN(
        n18735) );
  AOI22_X1 U21786 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18859), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n18856), .ZN(n18733) );
  OAI211_X1 U21787 ( .C1(n10932), .C2(n18792), .A(n18733), .B(n19016), .ZN(
        n18734) );
  AOI211_X1 U21788 ( .C1(n18852), .C2(n18736), .A(n18735), .B(n18734), .ZN(
        n18741) );
  NOR3_X1 U21789 ( .A1(n18830), .A2(n18737), .A3(n19555), .ZN(n18752) );
  AOI22_X1 U21790 ( .A1(n18739), .A2(n18854), .B1(n18752), .B2(n18738), .ZN(
        n18740) );
  OAI211_X1 U21791 ( .C1(n18879), .C2(n18842), .A(n18741), .B(n18740), .ZN(
        P2_U2843) );
  OAI22_X1 U21792 ( .A1(n18826), .A2(n18744), .B1(n18743), .B2(n18742), .ZN(
        n18745) );
  AOI211_X1 U21793 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n18853), .A(n18980), 
        .B(n18745), .ZN(n18746) );
  OAI21_X1 U21794 ( .B1(n18747), .B2(n18810), .A(n18746), .ZN(n18748) );
  AOI21_X1 U21795 ( .B1(n18880), .B2(n18855), .A(n18748), .ZN(n18755) );
  INV_X1 U21796 ( .A(n18749), .ZN(n18845) );
  NAND2_X1 U21797 ( .A1(n18753), .A2(n18750), .ZN(n18751) );
  AOI22_X1 U21798 ( .A1(n18753), .A2(n18845), .B1(n18752), .B2(n18751), .ZN(
        n18754) );
  OAI211_X1 U21799 ( .C1(n18756), .C2(n18822), .A(n18755), .B(n18754), .ZN(
        P2_U2844) );
  AOI22_X1 U21800 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18859), .B1(
        n18757), .B2(n18852), .ZN(n18758) );
  OAI211_X1 U21801 ( .C1(n10905), .C2(n18792), .A(n18758), .B(n19016), .ZN(
        n18759) );
  AOI21_X1 U21802 ( .B1(P2_EBX_REG_10__SCAN_IN), .B2(n18856), .A(n18759), .ZN(
        n18766) );
  NOR2_X1 U21803 ( .A1(n18830), .A2(n18760), .ZN(n18762) );
  XNOR2_X1 U21804 ( .A(n18762), .B(n18761), .ZN(n18763) );
  AOI22_X1 U21805 ( .A1(n18764), .A2(n18854), .B1(n18818), .B2(n18763), .ZN(
        n18765) );
  OAI211_X1 U21806 ( .C1(n18884), .C2(n18842), .A(n18766), .B(n18765), .ZN(
        P2_U2845) );
  AOI22_X1 U21807 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18859), .B1(
        n18852), .B2(n18767), .ZN(n18768) );
  OAI21_X1 U21808 ( .B1(n18826), .B2(n11066), .A(n18768), .ZN(n18769) );
  AOI211_X1 U21809 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18853), .A(n18980), .B(
        n18769), .ZN(n18775) );
  NAND2_X1 U21810 ( .A1(n18814), .A2(n18770), .ZN(n18771) );
  XNOR2_X1 U21811 ( .A(n18772), .B(n18771), .ZN(n18773) );
  AOI22_X1 U21812 ( .A1(n18885), .A2(n18855), .B1(n18818), .B2(n18773), .ZN(
        n18774) );
  OAI211_X1 U21813 ( .C1(n18776), .C2(n18822), .A(n18775), .B(n18774), .ZN(
        P2_U2846) );
  AOI22_X1 U21814 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18859), .B1(
        n18777), .B2(n18852), .ZN(n18778) );
  OAI211_X1 U21815 ( .C1(n10875), .C2(n18792), .A(n18778), .B(n19016), .ZN(
        n18779) );
  AOI21_X1 U21816 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n18856), .A(n18779), .ZN(
        n18786) );
  NOR2_X1 U21817 ( .A1(n18830), .A2(n18780), .ZN(n18782) );
  XNOR2_X1 U21818 ( .A(n18782), .B(n18781), .ZN(n18784) );
  AOI22_X1 U21819 ( .A1(n18818), .A2(n18784), .B1(n18854), .B2(n18783), .ZN(
        n18785) );
  OAI211_X1 U21820 ( .C1(n18842), .C2(n18889), .A(n18786), .B(n18785), .ZN(
        P2_U2847) );
  NAND2_X1 U21821 ( .A1(n18814), .A2(n18787), .ZN(n18789) );
  XOR2_X1 U21822 ( .A(n18789), .B(n18788), .Z(n18797) );
  AOI22_X1 U21823 ( .A1(P2_EBX_REG_7__SCAN_IN), .A2(n18856), .B1(n18790), .B2(
        n18852), .ZN(n18791) );
  OAI211_X1 U21824 ( .C1(n10861), .C2(n18792), .A(n18791), .B(n19016), .ZN(
        n18795) );
  OAI22_X1 U21825 ( .A1(n18842), .A2(n18891), .B1(n18822), .B2(n18793), .ZN(
        n18794) );
  AOI211_X1 U21826 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18838), .A(
        n18795), .B(n18794), .ZN(n18796) );
  OAI21_X1 U21827 ( .B1(n18797), .B2(n19555), .A(n18796), .ZN(P2_U2848) );
  NOR2_X1 U21828 ( .A1(n18830), .A2(n18798), .ZN(n18800) );
  XOR2_X1 U21829 ( .A(n18800), .B(n18799), .Z(n18808) );
  AOI22_X1 U21830 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18859), .B1(
        P2_EBX_REG_6__SCAN_IN), .B2(n18856), .ZN(n18801) );
  OAI21_X1 U21831 ( .B1(n18802), .B2(n18810), .A(n18801), .ZN(n18803) );
  AOI211_X1 U21832 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n18853), .A(n18980), .B(
        n18803), .ZN(n18807) );
  INV_X1 U21833 ( .A(n18804), .ZN(n18893) );
  AOI22_X1 U21834 ( .A1(n18855), .A2(n18893), .B1(n18854), .B2(n18805), .ZN(
        n18806) );
  OAI211_X1 U21835 ( .C1(n19555), .C2(n18808), .A(n18807), .B(n18806), .ZN(
        P2_U2849) );
  AOI22_X1 U21836 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n18859), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n18856), .ZN(n18809) );
  OAI21_X1 U21837 ( .B1(n18811), .B2(n18810), .A(n18809), .ZN(n18812) );
  AOI211_X1 U21838 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18853), .A(n18980), .B(
        n18812), .ZN(n18820) );
  NAND2_X1 U21839 ( .A1(n18814), .A2(n18813), .ZN(n18815) );
  XNOR2_X1 U21840 ( .A(n18816), .B(n18815), .ZN(n18817) );
  AOI22_X1 U21841 ( .A1(n18855), .A2(n18896), .B1(n18818), .B2(n18817), .ZN(
        n18819) );
  OAI211_X1 U21842 ( .C1(n18822), .C2(n18821), .A(n18820), .B(n18819), .ZN(
        P2_U2850) );
  AOI22_X1 U21843 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18859), .B1(
        n18823), .B2(n18852), .ZN(n18837) );
  OAI22_X1 U21844 ( .A1(n18826), .A2(n18825), .B1(n18842), .B2(n18824), .ZN(
        n18827) );
  AOI211_X1 U21845 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n18853), .A(n18980), .B(
        n18827), .ZN(n18836) );
  INV_X1 U21846 ( .A(n18828), .ZN(n18897) );
  AOI22_X1 U21847 ( .A1(n18897), .A2(n18857), .B1(n18987), .B2(n18854), .ZN(
        n18835) );
  INV_X1 U21848 ( .A(n18991), .ZN(n18833) );
  NOR2_X1 U21849 ( .A1(n18830), .A2(n18829), .ZN(n18832) );
  AOI21_X1 U21850 ( .B1(n18833), .B2(n18832), .A(n19555), .ZN(n18831) );
  OAI21_X1 U21851 ( .B1(n18833), .B2(n18832), .A(n18831), .ZN(n18834) );
  NAND4_X1 U21852 ( .A1(n18837), .A2(n18836), .A3(n18835), .A4(n18834), .ZN(
        P2_U2851) );
  INV_X1 U21853 ( .A(n19658), .ZN(n18843) );
  AOI22_X1 U21854 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18838), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n18856), .ZN(n18841) );
  AOI22_X1 U21855 ( .A1(n18853), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n18839), 
        .B2(n18852), .ZN(n18840) );
  OAI211_X1 U21856 ( .C1(n18843), .C2(n18842), .A(n18841), .B(n18840), .ZN(
        n18844) );
  AOI21_X1 U21857 ( .B1(n9598), .B2(n18854), .A(n18844), .ZN(n18849) );
  AOI22_X1 U21858 ( .A1(n18847), .A2(n18857), .B1(n18846), .B2(n18845), .ZN(
        n18848) );
  OAI211_X1 U21859 ( .C1(n19555), .C2(n18850), .A(n18849), .B(n18848), .ZN(
        P2_U2854) );
  AOI22_X1 U21860 ( .A1(n18853), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n18852), 
        .B2(n18851), .ZN(n18863) );
  AOI222_X1 U21861 ( .A1(n18856), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n18924), 
        .B2(n18855), .C1(n12340), .C2(n18854), .ZN(n18862) );
  AOI22_X1 U21862 ( .A1(n18818), .A2(n18858), .B1(n19663), .B2(n18857), .ZN(
        n18861) );
  NAND2_X1 U21863 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18859), .ZN(
        n18860) );
  NAND4_X1 U21864 ( .A1(n18863), .A2(n18862), .A3(n18861), .A4(n18860), .ZN(
        P2_U2855) );
  AOI22_X1 U21865 ( .A1(n15930), .A2(n18921), .B1(n18864), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18867) );
  AOI22_X1 U21866 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n18865), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n18920), .ZN(n18866) );
  NAND2_X1 U21867 ( .A1(n18867), .A2(n18866), .ZN(P2_U2888) );
  INV_X1 U21868 ( .A(n18921), .ZN(n18869) );
  OAI222_X1 U21869 ( .A1(n18937), .A2(n18892), .B1(n18871), .B2(n18890), .C1(
        n18870), .C2(n18927), .ZN(P2_U2904) );
  AOI22_X1 U21870 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n18920), .B1(n18972), 
        .B2(n18874), .ZN(n18872) );
  OAI21_X1 U21871 ( .B1(n18890), .B2(n18873), .A(n18872), .ZN(P2_U2905) );
  INV_X1 U21872 ( .A(n18890), .ZN(n18895) );
  AOI22_X1 U21873 ( .A1(n18876), .A2(n18895), .B1(n18875), .B2(n18874), .ZN(
        n18877) );
  OAI21_X1 U21874 ( .B1(n18892), .B2(n18941), .A(n18877), .ZN(P2_U2906) );
  INV_X1 U21875 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18943) );
  OAI222_X1 U21876 ( .A1(n18943), .A2(n18892), .B1(n18879), .B2(n18890), .C1(
        n18927), .C2(n18878), .ZN(P2_U2907) );
  AOI22_X1 U21877 ( .A1(n18880), .A2(n18895), .B1(P2_EAX_REG_11__SCAN_IN), 
        .B2(n18920), .ZN(n18881) );
  OAI21_X1 U21878 ( .B1(n18882), .B2(n18927), .A(n18881), .ZN(P2_U2908) );
  INV_X1 U21879 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20788) );
  OAI222_X1 U21880 ( .A1(n20788), .A2(n18892), .B1(n18884), .B2(n18890), .C1(
        n18927), .C2(n18883), .ZN(P2_U2909) );
  AOI22_X1 U21881 ( .A1(n18885), .A2(n18895), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n18920), .ZN(n18886) );
  OAI21_X1 U21882 ( .B1(n18887), .B2(n18927), .A(n18886), .ZN(P2_U2910) );
  INV_X1 U21883 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n18950) );
  OAI222_X1 U21884 ( .A1(n18950), .A2(n18892), .B1(n18889), .B2(n18890), .C1(
        n18927), .C2(n18888), .ZN(P2_U2911) );
  INV_X1 U21885 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18952) );
  OAI222_X1 U21886 ( .A1(n18952), .A2(n18892), .B1(n18891), .B2(n18890), .C1(
        n18927), .C2(n19053), .ZN(P2_U2912) );
  AOI22_X1 U21887 ( .A1(n18893), .A2(n18895), .B1(P2_EAX_REG_6__SCAN_IN), .B2(
        n18920), .ZN(n18894) );
  OAI21_X1 U21888 ( .B1(n19044), .B2(n18927), .A(n18894), .ZN(P2_U2913) );
  AOI22_X1 U21889 ( .A1(n18896), .A2(n18895), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n18920), .ZN(n18900) );
  NAND3_X1 U21890 ( .A1(n18898), .A2(n18897), .A3(n18922), .ZN(n18899) );
  OAI211_X1 U21891 ( .C1(n19040), .C2(n18927), .A(n18900), .B(n18899), .ZN(
        P2_U2914) );
  AOI22_X1 U21892 ( .A1(n18921), .A2(n18901), .B1(n18920), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n18907) );
  OAI21_X1 U21893 ( .B1(n18904), .B2(n18903), .A(n18902), .ZN(n18905) );
  NAND2_X1 U21894 ( .A1(n18905), .A2(n18922), .ZN(n18906) );
  OAI211_X1 U21895 ( .C1(n19034), .C2(n18927), .A(n18907), .B(n18906), .ZN(
        P2_U2916) );
  AOI22_X1 U21896 ( .A1(n18921), .A2(n19649), .B1(n18920), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n18913) );
  OAI21_X1 U21897 ( .B1(n18910), .B2(n18909), .A(n18908), .ZN(n18911) );
  NAND2_X1 U21898 ( .A1(n18911), .A2(n18922), .ZN(n18912) );
  OAI211_X1 U21899 ( .C1(n19029), .C2(n18927), .A(n18913), .B(n18912), .ZN(
        P2_U2917) );
  AOI22_X1 U21900 ( .A1(n18921), .A2(n19658), .B1(n18920), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n18918) );
  OAI21_X1 U21901 ( .B1(n18915), .B2(n18923), .A(n18914), .ZN(n18916) );
  NAND2_X1 U21902 ( .A1(n18916), .A2(n18922), .ZN(n18917) );
  OAI211_X1 U21903 ( .C1(n18919), .C2(n18927), .A(n18918), .B(n18917), .ZN(
        P2_U2918) );
  AOI22_X1 U21904 ( .A1(n18921), .A2(n18924), .B1(n18920), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n18926) );
  OAI211_X1 U21905 ( .C1(n19663), .C2(n18924), .A(n18923), .B(n18922), .ZN(
        n18925) );
  OAI211_X1 U21906 ( .C1(n18928), .C2(n18927), .A(n18926), .B(n18925), .ZN(
        P2_U2919) );
  INV_X1 U21907 ( .A(n18966), .ZN(n18933) );
  NOR2_X1 U21908 ( .A1(n18933), .A2(n18929), .ZN(P2_U2920) );
  INV_X1 U21909 ( .A(n18930), .ZN(n18934) );
  AOI22_X1 U21910 ( .A1(n18934), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n18963), .ZN(n18931) );
  OAI21_X1 U21911 ( .B1(n18933), .B2(n18932), .A(n18931), .ZN(P2_U2921) );
  INV_X1 U21912 ( .A(P2_UWORD_REG_13__SCAN_IN), .ZN(n20709) );
  AOI22_X1 U21913 ( .A1(n18934), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n18935) );
  OAI21_X1 U21914 ( .B1(n19679), .B2(n20709), .A(n18935), .ZN(P2_U2922) );
  AOI22_X1 U21915 ( .A1(n18963), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18936) );
  OAI21_X1 U21916 ( .B1(n18937), .B2(n18968), .A(n18936), .ZN(P2_U2936) );
  INV_X1 U21917 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18939) );
  AOI22_X1 U21918 ( .A1(n18963), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18938) );
  OAI21_X1 U21919 ( .B1(n18939), .B2(n18968), .A(n18938), .ZN(P2_U2937) );
  AOI22_X1 U21920 ( .A1(n18963), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18940) );
  OAI21_X1 U21921 ( .B1(n18941), .B2(n18968), .A(n18940), .ZN(P2_U2938) );
  AOI22_X1 U21922 ( .A1(n18963), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18942) );
  OAI21_X1 U21923 ( .B1(n18943), .B2(n18968), .A(n18942), .ZN(P2_U2939) );
  INV_X1 U21924 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18945) );
  AOI22_X1 U21925 ( .A1(n18963), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18944) );
  OAI21_X1 U21926 ( .B1(n18945), .B2(n18968), .A(n18944), .ZN(P2_U2940) );
  AOI22_X1 U21927 ( .A1(n18963), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18946) );
  OAI21_X1 U21928 ( .B1(n20788), .B2(n18968), .A(n18946), .ZN(P2_U2941) );
  INV_X1 U21929 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18948) );
  AOI22_X1 U21930 ( .A1(n18963), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18947) );
  OAI21_X1 U21931 ( .B1(n18948), .B2(n18968), .A(n18947), .ZN(P2_U2942) );
  AOI22_X1 U21932 ( .A1(n18963), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18949) );
  OAI21_X1 U21933 ( .B1(n18950), .B2(n18968), .A(n18949), .ZN(P2_U2943) );
  AOI22_X1 U21934 ( .A1(n18963), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18951) );
  OAI21_X1 U21935 ( .B1(n18952), .B2(n18968), .A(n18951), .ZN(P2_U2944) );
  INV_X1 U21936 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18954) );
  AOI22_X1 U21937 ( .A1(n18963), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18953) );
  OAI21_X1 U21938 ( .B1(n18954), .B2(n18968), .A(n18953), .ZN(P2_U2945) );
  INV_X1 U21939 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18956) );
  AOI22_X1 U21940 ( .A1(n18963), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18955) );
  OAI21_X1 U21941 ( .B1(n18956), .B2(n18968), .A(n18955), .ZN(P2_U2946) );
  INV_X1 U21942 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n18958) );
  AOI22_X1 U21943 ( .A1(n18963), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18957) );
  OAI21_X1 U21944 ( .B1(n18958), .B2(n18968), .A(n18957), .ZN(P2_U2947) );
  INV_X1 U21945 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18960) );
  AOI22_X1 U21946 ( .A1(n18963), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n18959) );
  OAI21_X1 U21947 ( .B1(n18960), .B2(n18968), .A(n18959), .ZN(P2_U2948) );
  INV_X1 U21948 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18962) );
  AOI22_X1 U21949 ( .A1(n18963), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18961) );
  OAI21_X1 U21950 ( .B1(n18962), .B2(n18968), .A(n18961), .ZN(P2_U2949) );
  INV_X1 U21951 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18965) );
  AOI22_X1 U21952 ( .A1(n18963), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18964) );
  OAI21_X1 U21953 ( .B1(n18965), .B2(n18968), .A(n18964), .ZN(P2_U2950) );
  AOI22_X1 U21954 ( .A1(n18963), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18966), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18967) );
  OAI21_X1 U21955 ( .B1(n10806), .B2(n18968), .A(n18967), .ZN(P2_U2951) );
  INV_X1 U21956 ( .A(n18969), .ZN(n18970) );
  AOI21_X1 U21957 ( .B1(n18975), .B2(P2_EAX_REG_29__SCAN_IN), .A(n18970), .ZN(
        n18971) );
  OAI21_X1 U21958 ( .B1(n20709), .B2(n12392), .A(n18971), .ZN(P2_U2965) );
  AOI22_X1 U21959 ( .A1(n18976), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n18975), .ZN(n18974) );
  NAND2_X1 U21960 ( .A1(n18973), .A2(n18972), .ZN(n18977) );
  NAND2_X1 U21961 ( .A1(n18974), .A2(n18977), .ZN(P2_U2966) );
  AOI22_X1 U21962 ( .A1(n18976), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n18975), .ZN(n18978) );
  NAND2_X1 U21963 ( .A1(n18978), .A2(n18977), .ZN(P2_U2981) );
  AOI22_X1 U21964 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n18980), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18979), .ZN(n18990) );
  INV_X1 U21965 ( .A(n18981), .ZN(n18985) );
  OAI22_X1 U21966 ( .A1(n18985), .A2(n18984), .B1(n18983), .B2(n18982), .ZN(
        n18986) );
  AOI21_X1 U21967 ( .B1(n18988), .B2(n18987), .A(n18986), .ZN(n18989) );
  OAI211_X1 U21968 ( .C1(n18992), .C2(n18991), .A(n18990), .B(n18989), .ZN(
        P2_U3010) );
  INV_X1 U21969 ( .A(n19649), .ZN(n18996) );
  OAI22_X1 U21970 ( .A1(n18996), .A2(n18995), .B1(n18994), .B2(n18993), .ZN(
        n18997) );
  AOI21_X1 U21971 ( .B1(n18999), .B2(n18998), .A(n18997), .ZN(n19015) );
  NAND2_X1 U21972 ( .A1(n19000), .A2(n19008), .ZN(n19002) );
  OAI211_X1 U21973 ( .C1(n19006), .C2(n19008), .A(n19002), .B(n19001), .ZN(
        n19003) );
  NAND2_X1 U21974 ( .A1(n19003), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19013) );
  NAND2_X1 U21975 ( .A1(n19005), .A2(n19004), .ZN(n19011) );
  INV_X1 U21976 ( .A(n19006), .ZN(n19009) );
  NAND3_X1 U21977 ( .A1(n19009), .A2(n19008), .A3(n19007), .ZN(n19010) );
  AND4_X1 U21978 ( .A1(n19013), .A2(n19012), .A3(n19011), .A4(n19010), .ZN(
        n19014) );
  OAI211_X1 U21979 ( .C1(n10269), .C2(n19016), .A(n19015), .B(n19014), .ZN(
        P2_U3044) );
  INV_X1 U21980 ( .A(n19395), .ZN(n19017) );
  NAND2_X1 U21981 ( .A1(n12670), .A2(n19651), .ZN(n19117) );
  NOR2_X1 U21982 ( .A1(n19250), .A2(n19117), .ZN(n19051) );
  AOI22_X1 U21983 ( .A1(n19502), .A2(n19052), .B1(n19494), .B2(n19051), .ZN(
        n19026) );
  AOI21_X1 U21984 ( .B1(n19548), .B2(n19086), .A(n19633), .ZN(n19018) );
  INV_X1 U21985 ( .A(n19642), .ZN(n19449) );
  NOR2_X1 U21986 ( .A1(n19018), .A2(n19449), .ZN(n19021) );
  AOI21_X1 U21987 ( .B1(n19022), .B2(n19639), .A(n19642), .ZN(n19019) );
  AOI21_X1 U21988 ( .B1(n19021), .B2(n19497), .A(n19019), .ZN(n19020) );
  OAI21_X1 U21989 ( .B1(n19020), .B2(n19051), .A(n19392), .ZN(n19055) );
  INV_X1 U21990 ( .A(n19497), .ZN(n19540) );
  OAI21_X1 U21991 ( .B1(n19540), .B2(n19051), .A(n19021), .ZN(n19024) );
  OAI21_X1 U21992 ( .B1(n19022), .B2(n19051), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19023) );
  NAND2_X1 U21993 ( .A1(n19024), .A2(n19023), .ZN(n19054) );
  AOI22_X1 U21994 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19055), .B1(
        n13025), .B2(n19054), .ZN(n19025) );
  OAI211_X1 U21995 ( .C1(n19505), .C2(n19086), .A(n19026), .B(n19025), .ZN(
        P2_U3048) );
  AOI22_X1 U21996 ( .A1(n19507), .A2(n19052), .B1(n19506), .B2(n19051), .ZN(
        n19028) );
  AOI22_X1 U21997 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19055), .B1(
        n13050), .B2(n19054), .ZN(n19027) );
  OAI211_X1 U21998 ( .C1(n19510), .C2(n19086), .A(n19028), .B(n19027), .ZN(
        P2_U3049) );
  AOI22_X1 U21999 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19047), .ZN(n19515) );
  AOI22_X1 U22000 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19047), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19048), .ZN(n19410) );
  AOI22_X1 U22001 ( .A1(n19512), .A2(n19052), .B1(n19511), .B2(n19051), .ZN(
        n19032) );
  AOI22_X1 U22002 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19055), .B1(
        n19030), .B2(n19054), .ZN(n19031) );
  OAI211_X1 U22003 ( .C1(n19515), .C2(n19086), .A(n19032), .B(n19031), .ZN(
        P2_U3050) );
  AOI22_X1 U22004 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19047), .ZN(n19520) );
  AOI22_X1 U22005 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19047), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19048), .ZN(n19416) );
  NOR2_X2 U22006 ( .A1(n10221), .A2(n19033), .ZN(n19516) );
  AOI22_X1 U22007 ( .A1(n19517), .A2(n19052), .B1(n19516), .B2(n19051), .ZN(
        n19037) );
  AOI22_X1 U22008 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19055), .B1(
        n19035), .B2(n19054), .ZN(n19036) );
  OAI211_X1 U22009 ( .C1(n19520), .C2(n19086), .A(n19037), .B(n19036), .ZN(
        P2_U3051) );
  AOI22_X1 U22010 ( .A1(n19523), .A2(n19052), .B1(n19521), .B2(n19051), .ZN(
        n19039) );
  AOI22_X1 U22011 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19055), .B1(
        n19522), .B2(n19054), .ZN(n19038) );
  OAI211_X1 U22012 ( .C1(n19526), .C2(n19086), .A(n19039), .B(n19038), .ZN(
        P2_U3052) );
  AOI22_X1 U22013 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19047), .ZN(n19532) );
  AOI22_X1 U22014 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19047), .ZN(n19428) );
  AOI22_X1 U22015 ( .A1(n19529), .A2(n19052), .B1(n19527), .B2(n19051), .ZN(
        n19042) );
  NOR2_X2 U22016 ( .A1(n19040), .A2(n19496), .ZN(n19528) );
  AOI22_X1 U22017 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19055), .B1(
        n19528), .B2(n19054), .ZN(n19041) );
  OAI211_X1 U22018 ( .C1(n19532), .C2(n19086), .A(n19042), .B(n19041), .ZN(
        P2_U3053) );
  AOI22_X1 U22019 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19047), .ZN(n19538) );
  AOI22_X1 U22020 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19047), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19048), .ZN(n19434) );
  AOI22_X1 U22021 ( .A1(n19535), .A2(n19052), .B1(n19533), .B2(n19051), .ZN(
        n19046) );
  NOR2_X2 U22022 ( .A1(n19044), .A2(n19496), .ZN(n19534) );
  AOI22_X1 U22023 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19055), .B1(
        n19534), .B2(n19054), .ZN(n19045) );
  OAI211_X1 U22024 ( .C1(n19538), .C2(n19086), .A(n19046), .B(n19045), .ZN(
        P2_U3054) );
  AOI22_X1 U22025 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19047), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19048), .ZN(n19549) );
  AOI22_X1 U22026 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19048), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19047), .ZN(n19444) );
  AOI22_X1 U22027 ( .A1(n19543), .A2(n19052), .B1(n19539), .B2(n19051), .ZN(
        n19057) );
  NOR2_X2 U22028 ( .A1(n19053), .A2(n19496), .ZN(n19541) );
  AOI22_X1 U22029 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19055), .B1(
        n19541), .B2(n19054), .ZN(n19056) );
  OAI211_X1 U22030 ( .C1(n19549), .C2(n19086), .A(n19057), .B(n19056), .ZN(
        P2_U3055) );
  NOR2_X1 U22031 ( .A1(n19117), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19065) );
  INV_X1 U22032 ( .A(n19065), .ZN(n19060) );
  INV_X1 U22033 ( .A(n19551), .ZN(n19059) );
  NOR2_X1 U22034 ( .A1(n19666), .A2(n19060), .ZN(n19081) );
  NOR3_X1 U22035 ( .A1(n19058), .A2(n19081), .A3(n19493), .ZN(n19061) );
  AOI211_X2 U22036 ( .C1(n19060), .C2(n19493), .A(n19059), .B(n19061), .ZN(
        n19082) );
  AOI22_X1 U22037 ( .A1(n19082), .A2(n13025), .B1(n19494), .B2(n19081), .ZN(
        n19068) );
  INV_X1 U22038 ( .A(n19081), .ZN(n19062) );
  AOI211_X1 U22039 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19062), .A(n19496), 
        .B(n19061), .ZN(n19063) );
  OAI221_X1 U22040 ( .B1(n19065), .B2(n19064), .C1(n19065), .C2(n19225), .A(
        n19063), .ZN(n19083) );
  AOI22_X1 U22041 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19083), .B1(
        n19112), .B2(n19453), .ZN(n19067) );
  OAI211_X1 U22042 ( .C1(n19398), .C2(n19086), .A(n19068), .B(n19067), .ZN(
        P2_U3056) );
  AOI22_X1 U22043 ( .A1(n19082), .A2(n13050), .B1(n19506), .B2(n19081), .ZN(
        n19070) );
  AOI22_X1 U22044 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19083), .B1(
        n19112), .B2(n19461), .ZN(n19069) );
  OAI211_X1 U22045 ( .C1(n19404), .C2(n19086), .A(n19070), .B(n19069), .ZN(
        P2_U3057) );
  AOI22_X1 U22046 ( .A1(n19082), .A2(n19030), .B1(n19511), .B2(n19081), .ZN(
        n19072) );
  AOI22_X1 U22047 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19083), .B1(
        n19112), .B2(n19464), .ZN(n19071) );
  OAI211_X1 U22048 ( .C1(n19410), .C2(n19086), .A(n19072), .B(n19071), .ZN(
        P2_U3058) );
  AOI22_X1 U22049 ( .A1(n19082), .A2(n19035), .B1(n19516), .B2(n19081), .ZN(
        n19074) );
  AOI22_X1 U22050 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19083), .B1(
        n19112), .B2(n19467), .ZN(n19073) );
  OAI211_X1 U22051 ( .C1(n19416), .C2(n19086), .A(n19074), .B(n19073), .ZN(
        P2_U3059) );
  AOI22_X1 U22052 ( .A1(n19082), .A2(n19522), .B1(n19081), .B2(n19521), .ZN(
        n19076) );
  AOI22_X1 U22053 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19083), .B1(
        n19112), .B2(n19470), .ZN(n19075) );
  OAI211_X1 U22054 ( .C1(n19422), .C2(n19086), .A(n19076), .B(n19075), .ZN(
        P2_U3060) );
  AOI22_X1 U22055 ( .A1(n19082), .A2(n19528), .B1(n19527), .B2(n19081), .ZN(
        n19078) );
  AOI22_X1 U22056 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19083), .B1(
        n19112), .B2(n19474), .ZN(n19077) );
  OAI211_X1 U22057 ( .C1(n19428), .C2(n19086), .A(n19078), .B(n19077), .ZN(
        P2_U3061) );
  AOI22_X1 U22058 ( .A1(n19082), .A2(n19534), .B1(n19533), .B2(n19081), .ZN(
        n19080) );
  AOI22_X1 U22059 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19083), .B1(
        n19112), .B2(n19477), .ZN(n19079) );
  OAI211_X1 U22060 ( .C1(n19434), .C2(n19086), .A(n19080), .B(n19079), .ZN(
        P2_U3062) );
  AOI22_X1 U22061 ( .A1(n19082), .A2(n19541), .B1(n19539), .B2(n19081), .ZN(
        n19085) );
  AOI22_X1 U22062 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19083), .B1(
        n19112), .B2(n19482), .ZN(n19084) );
  OAI211_X1 U22063 ( .C1(n19444), .C2(n19086), .A(n19085), .B(n19084), .ZN(
        P2_U3063) );
  NOR3_X2 U22064 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10817), .A3(
        n19117), .ZN(n19110) );
  OAI21_X1 U22065 ( .B1(n19088), .B2(n19110), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19091) );
  INV_X1 U22066 ( .A(n19305), .ZN(n19090) );
  INV_X1 U22067 ( .A(n19117), .ZN(n19089) );
  NAND2_X1 U22068 ( .A1(n19090), .A2(n19089), .ZN(n19092) );
  NAND2_X1 U22069 ( .A1(n19091), .A2(n19092), .ZN(n19111) );
  AOI22_X1 U22070 ( .A1(n19111), .A2(n13025), .B1(n19494), .B2(n19110), .ZN(
        n19097) );
  AOI21_X1 U22071 ( .B1(n10423), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19095) );
  OAI21_X1 U22072 ( .B1(n19112), .B2(n19142), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19093) );
  NAND3_X1 U22073 ( .A1(n19093), .A2(n19642), .A3(n19092), .ZN(n19094) );
  OAI211_X1 U22074 ( .C1(n19110), .C2(n19095), .A(n19094), .B(n19392), .ZN(
        n19113) );
  AOI22_X1 U22075 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19502), .ZN(n19096) );
  OAI211_X1 U22076 ( .C1(n19505), .C2(n19116), .A(n19097), .B(n19096), .ZN(
        P2_U3064) );
  AOI22_X1 U22077 ( .A1(n19111), .A2(n13050), .B1(n19506), .B2(n19110), .ZN(
        n19099) );
  AOI22_X1 U22078 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19507), .ZN(n19098) );
  OAI211_X1 U22079 ( .C1(n19510), .C2(n19116), .A(n19099), .B(n19098), .ZN(
        P2_U3065) );
  AOI22_X1 U22080 ( .A1(n19111), .A2(n19030), .B1(n19511), .B2(n19110), .ZN(
        n19101) );
  AOI22_X1 U22081 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19512), .ZN(n19100) );
  OAI211_X1 U22082 ( .C1(n19515), .C2(n19116), .A(n19101), .B(n19100), .ZN(
        P2_U3066) );
  AOI22_X1 U22083 ( .A1(n19111), .A2(n19035), .B1(n19516), .B2(n19110), .ZN(
        n19103) );
  AOI22_X1 U22084 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19517), .ZN(n19102) );
  OAI211_X1 U22085 ( .C1(n19520), .C2(n19116), .A(n19103), .B(n19102), .ZN(
        P2_U3067) );
  AOI22_X1 U22086 ( .A1(n19111), .A2(n19522), .B1(n19110), .B2(n19521), .ZN(
        n19105) );
  AOI22_X1 U22087 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19523), .ZN(n19104) );
  OAI211_X1 U22088 ( .C1(n19526), .C2(n19116), .A(n19105), .B(n19104), .ZN(
        P2_U3068) );
  AOI22_X1 U22089 ( .A1(n19111), .A2(n19528), .B1(n19527), .B2(n19110), .ZN(
        n19107) );
  AOI22_X1 U22090 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19529), .ZN(n19106) );
  OAI211_X1 U22091 ( .C1(n19532), .C2(n19116), .A(n19107), .B(n19106), .ZN(
        P2_U3069) );
  AOI22_X1 U22092 ( .A1(n19111), .A2(n19534), .B1(n19533), .B2(n19110), .ZN(
        n19109) );
  AOI22_X1 U22093 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19535), .ZN(n19108) );
  OAI211_X1 U22094 ( .C1(n19538), .C2(n19116), .A(n19109), .B(n19108), .ZN(
        P2_U3070) );
  AOI22_X1 U22095 ( .A1(n19111), .A2(n19541), .B1(n19539), .B2(n19110), .ZN(
        n19115) );
  AOI22_X1 U22096 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19543), .ZN(n19114) );
  OAI211_X1 U22097 ( .C1(n19549), .C2(n19116), .A(n19115), .B(n19114), .ZN(
        P2_U3071) );
  OR2_X1 U22098 ( .A1(n10817), .A2(n19117), .ZN(n19120) );
  NOR2_X1 U22099 ( .A1(n19449), .A2(n19120), .ZN(n19119) );
  NOR2_X1 U22100 ( .A1(n19335), .A2(n19117), .ZN(n19141) );
  INV_X1 U22101 ( .A(n19141), .ZN(n19122) );
  AOI21_X1 U22102 ( .B1(n19123), .B2(n19122), .A(n19493), .ZN(n19118) );
  NOR2_X1 U22103 ( .A1(n19119), .A2(n19118), .ZN(n19146) );
  INV_X1 U22104 ( .A(n13025), .ZN(n19386) );
  NOR2_X2 U22105 ( .A1(n19229), .A2(n19303), .ZN(n19171) );
  AOI22_X1 U22106 ( .A1(n19453), .A2(n19171), .B1(n19494), .B2(n19141), .ZN(
        n19128) );
  NAND2_X1 U22107 ( .A1(n19225), .A2(n19632), .ZN(n19121) );
  NAND2_X1 U22108 ( .A1(n19121), .A2(n19120), .ZN(n19125) );
  OAI21_X1 U22109 ( .B1(n19123), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19122), 
        .ZN(n19124) );
  MUX2_X1 U22110 ( .A(n19125), .B(n19124), .S(n19449), .Z(n19126) );
  NAND2_X1 U22111 ( .A1(n19126), .A2(n19392), .ZN(n19143) );
  AOI22_X1 U22112 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19143), .B1(
        n19142), .B2(n19502), .ZN(n19127) );
  OAI211_X1 U22113 ( .C1(n19146), .C2(n19386), .A(n19128), .B(n19127), .ZN(
        P2_U3072) );
  INV_X1 U22114 ( .A(n13050), .ZN(n19400) );
  AOI22_X1 U22115 ( .A1(n19507), .A2(n19142), .B1(n19506), .B2(n19141), .ZN(
        n19130) );
  AOI22_X1 U22116 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19143), .B1(
        n19171), .B2(n19461), .ZN(n19129) );
  OAI211_X1 U22117 ( .C1(n19146), .C2(n19400), .A(n19130), .B(n19129), .ZN(
        P2_U3073) );
  INV_X1 U22118 ( .A(n19030), .ZN(n19406) );
  AOI22_X1 U22119 ( .A1(n19464), .A2(n19171), .B1(n19141), .B2(n19511), .ZN(
        n19132) );
  AOI22_X1 U22120 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19143), .B1(
        n19142), .B2(n19512), .ZN(n19131) );
  OAI211_X1 U22121 ( .C1(n19146), .C2(n19406), .A(n19132), .B(n19131), .ZN(
        P2_U3074) );
  INV_X1 U22122 ( .A(n19035), .ZN(n19412) );
  AOI22_X1 U22123 ( .A1(n19517), .A2(n19142), .B1(n19141), .B2(n19516), .ZN(
        n19134) );
  AOI22_X1 U22124 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19143), .B1(
        n19171), .B2(n19467), .ZN(n19133) );
  OAI211_X1 U22125 ( .C1(n19146), .C2(n19412), .A(n19134), .B(n19133), .ZN(
        P2_U3075) );
  AOI22_X1 U22126 ( .A1(n19470), .A2(n19171), .B1(n19141), .B2(n19521), .ZN(
        n19136) );
  AOI22_X1 U22127 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19143), .B1(
        n19142), .B2(n19523), .ZN(n19135) );
  OAI211_X1 U22128 ( .C1(n19146), .C2(n19418), .A(n19136), .B(n19135), .ZN(
        P2_U3076) );
  INV_X1 U22129 ( .A(n19528), .ZN(n19424) );
  AOI22_X1 U22130 ( .A1(n19529), .A2(n19142), .B1(n19141), .B2(n19527), .ZN(
        n19138) );
  AOI22_X1 U22131 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19143), .B1(
        n19171), .B2(n19474), .ZN(n19137) );
  OAI211_X1 U22132 ( .C1(n19146), .C2(n19424), .A(n19138), .B(n19137), .ZN(
        P2_U3077) );
  INV_X1 U22133 ( .A(n19534), .ZN(n19430) );
  AOI22_X1 U22134 ( .A1(n19535), .A2(n19142), .B1(n19141), .B2(n19533), .ZN(
        n19140) );
  AOI22_X1 U22135 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19143), .B1(
        n19171), .B2(n19477), .ZN(n19139) );
  OAI211_X1 U22136 ( .C1(n19146), .C2(n19430), .A(n19140), .B(n19139), .ZN(
        P2_U3078) );
  INV_X1 U22137 ( .A(n19541), .ZN(n19437) );
  AOI22_X1 U22138 ( .A1(n19482), .A2(n19171), .B1(n19141), .B2(n19539), .ZN(
        n19145) );
  AOI22_X1 U22139 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19143), .B1(
        n19142), .B2(n19543), .ZN(n19144) );
  OAI211_X1 U22140 ( .C1(n19146), .C2(n19437), .A(n19145), .B(n19144), .ZN(
        P2_U3079) );
  OR2_X1 U22141 ( .A1(n19148), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19153) );
  NOR2_X1 U22142 ( .A1(n19250), .A2(n19221), .ZN(n19169) );
  OAI21_X1 U22143 ( .B1(n19149), .B2(n19169), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19150) );
  OAI21_X1 U22144 ( .B1(n19153), .B2(n19449), .A(n19150), .ZN(n19170) );
  AOI22_X1 U22145 ( .A1(n19170), .A2(n13025), .B1(n19494), .B2(n19169), .ZN(
        n19156) );
  OAI21_X1 U22146 ( .B1(n19171), .B2(n19197), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19152) );
  AOI211_X1 U22147 ( .C1(n19149), .C2(n19639), .A(n19642), .B(n19169), .ZN(
        n19151) );
  AOI211_X1 U22148 ( .C1(n19153), .C2(n19152), .A(n19496), .B(n19151), .ZN(
        n19154) );
  AOI22_X1 U22149 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19172), .B1(
        n19171), .B2(n19502), .ZN(n19155) );
  OAI211_X1 U22150 ( .C1(n19505), .C2(n19175), .A(n19156), .B(n19155), .ZN(
        P2_U3080) );
  AOI22_X1 U22151 ( .A1(n19170), .A2(n13050), .B1(n19506), .B2(n19169), .ZN(
        n19158) );
  AOI22_X1 U22152 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19172), .B1(
        n19171), .B2(n19507), .ZN(n19157) );
  OAI211_X1 U22153 ( .C1(n19510), .C2(n19175), .A(n19158), .B(n19157), .ZN(
        P2_U3081) );
  AOI22_X1 U22154 ( .A1(n19170), .A2(n19030), .B1(n19511), .B2(n19169), .ZN(
        n19160) );
  AOI22_X1 U22155 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19172), .B1(
        n19171), .B2(n19512), .ZN(n19159) );
  OAI211_X1 U22156 ( .C1(n19515), .C2(n19175), .A(n19160), .B(n19159), .ZN(
        P2_U3082) );
  AOI22_X1 U22157 ( .A1(n19170), .A2(n19035), .B1(n19516), .B2(n19169), .ZN(
        n19162) );
  AOI22_X1 U22158 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19172), .B1(
        n19171), .B2(n19517), .ZN(n19161) );
  OAI211_X1 U22159 ( .C1(n19520), .C2(n19175), .A(n19162), .B(n19161), .ZN(
        P2_U3083) );
  AOI22_X1 U22160 ( .A1(n19170), .A2(n19522), .B1(n19169), .B2(n19521), .ZN(
        n19164) );
  AOI22_X1 U22161 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19172), .B1(
        n19171), .B2(n19523), .ZN(n19163) );
  OAI211_X1 U22162 ( .C1(n19526), .C2(n19175), .A(n19164), .B(n19163), .ZN(
        P2_U3084) );
  AOI22_X1 U22163 ( .A1(n19170), .A2(n19528), .B1(n19527), .B2(n19169), .ZN(
        n19166) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19172), .B1(
        n19171), .B2(n19529), .ZN(n19165) );
  OAI211_X1 U22165 ( .C1(n19532), .C2(n19175), .A(n19166), .B(n19165), .ZN(
        P2_U3085) );
  AOI22_X1 U22166 ( .A1(n19170), .A2(n19534), .B1(n19533), .B2(n19169), .ZN(
        n19168) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19172), .B1(
        n19171), .B2(n19535), .ZN(n19167) );
  OAI211_X1 U22168 ( .C1(n19538), .C2(n19175), .A(n19168), .B(n19167), .ZN(
        P2_U3086) );
  AOI22_X1 U22169 ( .A1(n19170), .A2(n19541), .B1(n19539), .B2(n19169), .ZN(
        n19174) );
  AOI22_X1 U22170 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19172), .B1(
        n19171), .B2(n19543), .ZN(n19173) );
  OAI211_X1 U22171 ( .C1(n19549), .C2(n19175), .A(n19174), .B(n19173), .ZN(
        P2_U3087) );
  INV_X1 U22172 ( .A(n19394), .ZN(n19388) );
  AOI21_X1 U22173 ( .B1(n19225), .B2(n19388), .A(n19449), .ZN(n19177) );
  NOR2_X1 U22174 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19221), .ZN(
        n19180) );
  NAND2_X1 U22175 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19180), .ZN(
        n19178) );
  AOI21_X1 U22176 ( .B1(n10426), .B2(n19178), .A(n19493), .ZN(n19176) );
  INV_X1 U22177 ( .A(n19178), .ZN(n19196) );
  AOI22_X1 U22178 ( .A1(n19197), .A2(n19502), .B1(n19494), .B2(n19196), .ZN(
        n19183) );
  INV_X1 U22179 ( .A(n19177), .ZN(n19181) );
  OAI211_X1 U22180 ( .C1(n10426), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19178), 
        .B(n19449), .ZN(n19179) );
  OAI211_X1 U22181 ( .C1(n19181), .C2(n19180), .A(n19392), .B(n19179), .ZN(
        n19198) );
  AOI22_X1 U22182 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19198), .B1(
        n19216), .B2(n19453), .ZN(n19182) );
  OAI211_X1 U22183 ( .C1(n19201), .C2(n19386), .A(n19183), .B(n19182), .ZN(
        P2_U3088) );
  AOI22_X1 U22184 ( .A1(n19197), .A2(n19507), .B1(n19506), .B2(n19196), .ZN(
        n19185) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19198), .B1(
        n19216), .B2(n19461), .ZN(n19184) );
  OAI211_X1 U22186 ( .C1(n19201), .C2(n19400), .A(n19185), .B(n19184), .ZN(
        P2_U3089) );
  AOI22_X1 U22187 ( .A1(n19197), .A2(n19512), .B1(n19511), .B2(n19196), .ZN(
        n19187) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19198), .B1(
        n19216), .B2(n19464), .ZN(n19186) );
  OAI211_X1 U22189 ( .C1(n19201), .C2(n19406), .A(n19187), .B(n19186), .ZN(
        P2_U3090) );
  AOI22_X1 U22190 ( .A1(n19467), .A2(n19216), .B1(n19196), .B2(n19516), .ZN(
        n19189) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19198), .B1(
        n19197), .B2(n19517), .ZN(n19188) );
  OAI211_X1 U22192 ( .C1(n19201), .C2(n19412), .A(n19189), .B(n19188), .ZN(
        P2_U3091) );
  AOI22_X1 U22193 ( .A1(n19470), .A2(n19216), .B1(n19521), .B2(n19196), .ZN(
        n19191) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19198), .B1(
        n19197), .B2(n19523), .ZN(n19190) );
  OAI211_X1 U22195 ( .C1(n19201), .C2(n19418), .A(n19191), .B(n19190), .ZN(
        P2_U3092) );
  AOI22_X1 U22196 ( .A1(n19474), .A2(n19216), .B1(n19196), .B2(n19527), .ZN(
        n19193) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19198), .B1(
        n19197), .B2(n19529), .ZN(n19192) );
  OAI211_X1 U22198 ( .C1(n19201), .C2(n19424), .A(n19193), .B(n19192), .ZN(
        P2_U3093) );
  AOI22_X1 U22199 ( .A1(n19477), .A2(n19216), .B1(n19196), .B2(n19533), .ZN(
        n19195) );
  AOI22_X1 U22200 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19198), .B1(
        n19197), .B2(n19535), .ZN(n19194) );
  OAI211_X1 U22201 ( .C1(n19201), .C2(n19430), .A(n19195), .B(n19194), .ZN(
        P2_U3094) );
  AOI22_X1 U22202 ( .A1(n19482), .A2(n19216), .B1(n19539), .B2(n19196), .ZN(
        n19200) );
  AOI22_X1 U22203 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19198), .B1(
        n19197), .B2(n19543), .ZN(n19199) );
  OAI211_X1 U22204 ( .C1(n19201), .C2(n19437), .A(n19200), .B(n19199), .ZN(
        P2_U3095) );
  AOI22_X1 U22205 ( .A1(n19215), .A2(n13050), .B1(n19506), .B2(n19214), .ZN(
        n19203) );
  AOI22_X1 U22206 ( .A1(n19216), .A2(n19507), .B1(n19220), .B2(n19461), .ZN(
        n19202) );
  OAI211_X1 U22207 ( .C1(n19219), .C2(n10309), .A(n19203), .B(n19202), .ZN(
        P2_U3097) );
  AOI22_X1 U22208 ( .A1(n19215), .A2(n19030), .B1(n19214), .B2(n19511), .ZN(
        n19205) );
  AOI22_X1 U22209 ( .A1(n19216), .A2(n19512), .B1(n19220), .B2(n19464), .ZN(
        n19204) );
  OAI211_X1 U22210 ( .C1(n19219), .C2(n14161), .A(n19205), .B(n19204), .ZN(
        P2_U3098) );
  AOI22_X1 U22211 ( .A1(n19215), .A2(n19035), .B1(n19214), .B2(n19516), .ZN(
        n19207) );
  AOI22_X1 U22212 ( .A1(n19216), .A2(n19517), .B1(n19220), .B2(n19467), .ZN(
        n19206) );
  OAI211_X1 U22213 ( .C1(n19219), .C2(n14185), .A(n19207), .B(n19206), .ZN(
        P2_U3099) );
  AOI22_X1 U22214 ( .A1(n19215), .A2(n19522), .B1(n19214), .B2(n19521), .ZN(
        n19209) );
  AOI22_X1 U22215 ( .A1(n19216), .A2(n19523), .B1(n19220), .B2(n19470), .ZN(
        n19208) );
  OAI211_X1 U22216 ( .C1(n19219), .C2(n14217), .A(n19209), .B(n19208), .ZN(
        P2_U3100) );
  AOI22_X1 U22217 ( .A1(n19215), .A2(n19528), .B1(n19214), .B2(n19527), .ZN(
        n19211) );
  AOI22_X1 U22218 ( .A1(n19216), .A2(n19529), .B1(n19220), .B2(n19474), .ZN(
        n19210) );
  OAI211_X1 U22219 ( .C1(n19219), .C2(n14237), .A(n19211), .B(n19210), .ZN(
        P2_U3101) );
  AOI22_X1 U22220 ( .A1(n19215), .A2(n19534), .B1(n19214), .B2(n19533), .ZN(
        n19213) );
  AOI22_X1 U22221 ( .A1(n19216), .A2(n19535), .B1(n19220), .B2(n19477), .ZN(
        n19212) );
  OAI211_X1 U22222 ( .C1(n19219), .C2(n10512), .A(n19213), .B(n19212), .ZN(
        P2_U3102) );
  AOI22_X1 U22223 ( .A1(n19215), .A2(n19541), .B1(n19214), .B2(n19539), .ZN(
        n19218) );
  AOI22_X1 U22224 ( .A1(n19216), .A2(n19543), .B1(n19220), .B2(n19482), .ZN(
        n19217) );
  OAI211_X1 U22225 ( .C1(n19219), .C2(n14291), .A(n19218), .B(n19217), .ZN(
        P2_U3103) );
  NOR2_X1 U22226 ( .A1(n19489), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19228) );
  INV_X1 U22227 ( .A(n19228), .ZN(n19224) );
  NOR2_X1 U22228 ( .A1(n19335), .A2(n19221), .ZN(n19251) );
  OAI21_X1 U22229 ( .B1(n19222), .B2(n19251), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19223) );
  OAI21_X1 U22230 ( .B1(n19224), .B2(n19449), .A(n19223), .ZN(n19244) );
  AOI22_X1 U22231 ( .A1(n19244), .A2(n13025), .B1(n19494), .B2(n19251), .ZN(
        n19231) );
  AND2_X1 U22232 ( .A1(n19225), .A2(n19500), .ZN(n19643) );
  INV_X1 U22233 ( .A(n19251), .ZN(n19226) );
  OAI211_X1 U22234 ( .C1(n10418), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19449), 
        .B(n19226), .ZN(n19227) );
  OAI211_X1 U22235 ( .C1(n19643), .C2(n19228), .A(n19392), .B(n19227), .ZN(
        n19245) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19245), .B1(
        n19279), .B2(n19453), .ZN(n19230) );
  OAI211_X1 U22237 ( .C1(n19398), .C2(n19248), .A(n19231), .B(n19230), .ZN(
        P2_U3104) );
  AOI22_X1 U22238 ( .A1(n19244), .A2(n13050), .B1(n19506), .B2(n19251), .ZN(
        n19233) );
  AOI22_X1 U22239 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19245), .B1(
        n19279), .B2(n19461), .ZN(n19232) );
  OAI211_X1 U22240 ( .C1(n19404), .C2(n19248), .A(n19233), .B(n19232), .ZN(
        P2_U3105) );
  AOI22_X1 U22241 ( .A1(n19244), .A2(n19030), .B1(n19251), .B2(n19511), .ZN(
        n19235) );
  AOI22_X1 U22242 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19245), .B1(
        n19279), .B2(n19464), .ZN(n19234) );
  OAI211_X1 U22243 ( .C1(n19410), .C2(n19248), .A(n19235), .B(n19234), .ZN(
        P2_U3106) );
  AOI22_X1 U22244 ( .A1(n19244), .A2(n19035), .B1(n19251), .B2(n19516), .ZN(
        n19237) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19245), .B1(
        n19279), .B2(n19467), .ZN(n19236) );
  OAI211_X1 U22246 ( .C1(n19416), .C2(n19248), .A(n19237), .B(n19236), .ZN(
        P2_U3107) );
  AOI22_X1 U22247 ( .A1(n19244), .A2(n19522), .B1(n19251), .B2(n19521), .ZN(
        n19239) );
  AOI22_X1 U22248 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19245), .B1(
        n19279), .B2(n19470), .ZN(n19238) );
  OAI211_X1 U22249 ( .C1(n19422), .C2(n19248), .A(n19239), .B(n19238), .ZN(
        P2_U3108) );
  AOI22_X1 U22250 ( .A1(n19244), .A2(n19528), .B1(n19251), .B2(n19527), .ZN(
        n19241) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19245), .B1(
        n19279), .B2(n19474), .ZN(n19240) );
  OAI211_X1 U22252 ( .C1(n19428), .C2(n19248), .A(n19241), .B(n19240), .ZN(
        P2_U3109) );
  AOI22_X1 U22253 ( .A1(n19244), .A2(n19534), .B1(n19251), .B2(n19533), .ZN(
        n19243) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19245), .B1(
        n19279), .B2(n19477), .ZN(n19242) );
  OAI211_X1 U22255 ( .C1(n19434), .C2(n19248), .A(n19243), .B(n19242), .ZN(
        P2_U3110) );
  AOI22_X1 U22256 ( .A1(n19244), .A2(n19541), .B1(n19251), .B2(n19539), .ZN(
        n19247) );
  AOI22_X1 U22257 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19245), .B1(
        n19279), .B2(n19482), .ZN(n19246) );
  OAI211_X1 U22258 ( .C1(n19444), .C2(n19248), .A(n19247), .B(n19246), .ZN(
        P2_U3111) );
  OAI21_X1 U22259 ( .B1(n19297), .B2(n19279), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19249) );
  NAND2_X1 U22260 ( .A1(n19249), .A2(n19642), .ZN(n19256) );
  INV_X1 U22261 ( .A(n19256), .ZN(n19253) );
  NOR2_X1 U22262 ( .A1(n19250), .A2(n19334), .ZN(n19278) );
  NOR2_X1 U22263 ( .A1(n19278), .A2(n19251), .ZN(n19254) );
  INV_X1 U22264 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n19259) );
  AOI22_X1 U22265 ( .A1(n19453), .A2(n19297), .B1(n19494), .B2(n19278), .ZN(
        n19258) );
  OAI21_X1 U22266 ( .B1(n10407), .B2(n19278), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19255) );
  AOI22_X1 U22267 ( .A1(n19256), .A2(n19255), .B1(n19254), .B2(n19493), .ZN(
        n19280) );
  AOI22_X1 U22268 ( .A1(n13025), .A2(n19280), .B1(n19279), .B2(n19502), .ZN(
        n19257) );
  OAI211_X1 U22269 ( .C1(n19284), .C2(n19259), .A(n19258), .B(n19257), .ZN(
        P2_U3112) );
  INV_X1 U22270 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n19262) );
  AOI22_X1 U22271 ( .A1(n19461), .A2(n19297), .B1(n19506), .B2(n19278), .ZN(
        n19261) );
  AOI22_X1 U22272 ( .A1(n13050), .A2(n19280), .B1(n19279), .B2(n19507), .ZN(
        n19260) );
  OAI211_X1 U22273 ( .C1(n19284), .C2(n19262), .A(n19261), .B(n19260), .ZN(
        P2_U3113) );
  AOI22_X1 U22274 ( .A1(n19464), .A2(n19297), .B1(n19511), .B2(n19278), .ZN(
        n19264) );
  AOI22_X1 U22275 ( .A1(n19030), .A2(n19280), .B1(n19279), .B2(n19512), .ZN(
        n19263) );
  OAI211_X1 U22276 ( .C1(n19284), .C2(n19265), .A(n19264), .B(n19263), .ZN(
        P2_U3114) );
  INV_X1 U22277 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n19268) );
  AOI22_X1 U22278 ( .A1(n19467), .A2(n19297), .B1(n19516), .B2(n19278), .ZN(
        n19267) );
  AOI22_X1 U22279 ( .A1(n19035), .A2(n19280), .B1(n19279), .B2(n19517), .ZN(
        n19266) );
  OAI211_X1 U22280 ( .C1(n19284), .C2(n19268), .A(n19267), .B(n19266), .ZN(
        P2_U3115) );
  INV_X1 U22281 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n19271) );
  AOI22_X1 U22282 ( .A1(n19470), .A2(n19297), .B1(n19521), .B2(n19278), .ZN(
        n19270) );
  AOI22_X1 U22283 ( .A1(n19522), .A2(n19280), .B1(n19279), .B2(n19523), .ZN(
        n19269) );
  OAI211_X1 U22284 ( .C1(n19284), .C2(n19271), .A(n19270), .B(n19269), .ZN(
        P2_U3116) );
  INV_X1 U22285 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n19274) );
  AOI22_X1 U22286 ( .A1(n19474), .A2(n19297), .B1(n19527), .B2(n19278), .ZN(
        n19273) );
  AOI22_X1 U22287 ( .A1(n19528), .A2(n19280), .B1(n19279), .B2(n19529), .ZN(
        n19272) );
  OAI211_X1 U22288 ( .C1(n19284), .C2(n19274), .A(n19273), .B(n19272), .ZN(
        P2_U3117) );
  AOI22_X1 U22289 ( .A1(n19477), .A2(n19297), .B1(n19533), .B2(n19278), .ZN(
        n19276) );
  AOI22_X1 U22290 ( .A1(n19534), .A2(n19280), .B1(n19279), .B2(n19535), .ZN(
        n19275) );
  OAI211_X1 U22291 ( .C1(n19284), .C2(n19277), .A(n19276), .B(n19275), .ZN(
        P2_U3118) );
  INV_X1 U22292 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n19283) );
  AOI22_X1 U22293 ( .A1(n19482), .A2(n19297), .B1(n19539), .B2(n19278), .ZN(
        n19282) );
  AOI22_X1 U22294 ( .A1(n19541), .A2(n19280), .B1(n19279), .B2(n19543), .ZN(
        n19281) );
  OAI211_X1 U22295 ( .C1(n19284), .C2(n19283), .A(n19282), .B(n19281), .ZN(
        P2_U3119) );
  INV_X1 U22296 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n19287) );
  AOI22_X1 U22297 ( .A1(n19512), .A2(n19297), .B1(n19306), .B2(n19511), .ZN(
        n19286) );
  AOI22_X1 U22298 ( .A1(n19030), .A2(n19298), .B1(n19329), .B2(n19464), .ZN(
        n19285) );
  OAI211_X1 U22299 ( .C1(n19302), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P2_U3122) );
  INV_X1 U22300 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n19290) );
  AOI22_X1 U22301 ( .A1(n19467), .A2(n19329), .B1(n19306), .B2(n19516), .ZN(
        n19289) );
  AOI22_X1 U22302 ( .A1(n19035), .A2(n19298), .B1(n19297), .B2(n19517), .ZN(
        n19288) );
  OAI211_X1 U22303 ( .C1(n19302), .C2(n19290), .A(n19289), .B(n19288), .ZN(
        P2_U3123) );
  INV_X1 U22304 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n19293) );
  AOI22_X1 U22305 ( .A1(n19474), .A2(n19329), .B1(n19306), .B2(n19527), .ZN(
        n19292) );
  AOI22_X1 U22306 ( .A1(n19528), .A2(n19298), .B1(n19297), .B2(n19529), .ZN(
        n19291) );
  OAI211_X1 U22307 ( .C1(n19302), .C2(n19293), .A(n19292), .B(n19291), .ZN(
        P2_U3125) );
  AOI22_X1 U22308 ( .A1(n19477), .A2(n19329), .B1(n19306), .B2(n19533), .ZN(
        n19295) );
  AOI22_X1 U22309 ( .A1(n19534), .A2(n19298), .B1(n19297), .B2(n19535), .ZN(
        n19294) );
  OAI211_X1 U22310 ( .C1(n19302), .C2(n19296), .A(n19295), .B(n19294), .ZN(
        P2_U3126) );
  INV_X1 U22311 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n19301) );
  AOI22_X1 U22312 ( .A1(n19482), .A2(n19329), .B1(n19306), .B2(n19539), .ZN(
        n19300) );
  AOI22_X1 U22313 ( .A1(n19541), .A2(n19298), .B1(n19297), .B2(n19543), .ZN(
        n19299) );
  OAI211_X1 U22314 ( .C1(n19302), .C2(n19301), .A(n19300), .B(n19299), .ZN(
        P2_U3127) );
  NOR3_X2 U22315 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10817), .A3(
        n19334), .ZN(n19327) );
  OAI21_X1 U22316 ( .B1(n19308), .B2(n19327), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19304) );
  OAI21_X1 U22317 ( .B1(n19334), .B2(n19305), .A(n19304), .ZN(n19328) );
  AOI22_X1 U22318 ( .A1(n19328), .A2(n13025), .B1(n19494), .B2(n19327), .ZN(
        n19314) );
  AOI221_X1 U22319 ( .B1(n19329), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19307), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19306), .ZN(n19310) );
  INV_X1 U22320 ( .A(n19308), .ZN(n19309) );
  MUX2_X1 U22321 ( .A(n19310), .B(n19309), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19311) );
  NOR2_X1 U22322 ( .A1(n19311), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19312) );
  OAI21_X1 U22323 ( .B1(n19312), .B2(n19327), .A(n19392), .ZN(n19330) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19502), .ZN(n19313) );
  OAI211_X1 U22325 ( .C1(n19505), .C2(n19361), .A(n19314), .B(n19313), .ZN(
        P2_U3128) );
  AOI22_X1 U22326 ( .A1(n19328), .A2(n13050), .B1(n19506), .B2(n19327), .ZN(
        n19316) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19507), .ZN(n19315) );
  OAI211_X1 U22328 ( .C1(n19510), .C2(n19361), .A(n19316), .B(n19315), .ZN(
        P2_U3129) );
  AOI22_X1 U22329 ( .A1(n19328), .A2(n19030), .B1(n19511), .B2(n19327), .ZN(
        n19318) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19512), .ZN(n19317) );
  OAI211_X1 U22331 ( .C1(n19515), .C2(n19361), .A(n19318), .B(n19317), .ZN(
        P2_U3130) );
  AOI22_X1 U22332 ( .A1(n19328), .A2(n19035), .B1(n19516), .B2(n19327), .ZN(
        n19320) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19517), .ZN(n19319) );
  OAI211_X1 U22334 ( .C1(n19520), .C2(n19361), .A(n19320), .B(n19319), .ZN(
        P2_U3131) );
  AOI22_X1 U22335 ( .A1(n19328), .A2(n19522), .B1(n19327), .B2(n19521), .ZN(
        n19322) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19523), .ZN(n19321) );
  OAI211_X1 U22337 ( .C1(n19526), .C2(n19361), .A(n19322), .B(n19321), .ZN(
        P2_U3132) );
  AOI22_X1 U22338 ( .A1(n19328), .A2(n19528), .B1(n19527), .B2(n19327), .ZN(
        n19324) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19529), .ZN(n19323) );
  OAI211_X1 U22340 ( .C1(n19532), .C2(n19361), .A(n19324), .B(n19323), .ZN(
        P2_U3133) );
  AOI22_X1 U22341 ( .A1(n19328), .A2(n19534), .B1(n19533), .B2(n19327), .ZN(
        n19326) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19535), .ZN(n19325) );
  OAI211_X1 U22343 ( .C1(n19538), .C2(n19361), .A(n19326), .B(n19325), .ZN(
        P2_U3134) );
  AOI22_X1 U22344 ( .A1(n19328), .A2(n19541), .B1(n19539), .B2(n19327), .ZN(
        n19332) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19543), .ZN(n19331) );
  OAI211_X1 U22346 ( .C1(n19549), .C2(n19361), .A(n19332), .B(n19331), .ZN(
        P2_U3135) );
  NAND2_X1 U22347 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19333), .ZN(
        n19337) );
  OR2_X1 U22348 ( .A1(n19337), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19336) );
  NOR2_X1 U22349 ( .A1(n19335), .A2(n19334), .ZN(n19356) );
  NOR3_X1 U22350 ( .A1(n10415), .A2(n19356), .A3(n19493), .ZN(n19338) );
  AOI21_X1 U22351 ( .B1(n19493), .B2(n19336), .A(n19338), .ZN(n19357) );
  AOI22_X1 U22352 ( .A1(n19357), .A2(n13025), .B1(n19494), .B2(n19356), .ZN(
        n19343) );
  INV_X1 U22353 ( .A(n19337), .ZN(n19341) );
  INV_X1 U22354 ( .A(n19356), .ZN(n19339) );
  AOI211_X1 U22355 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19339), .A(n19496), 
        .B(n19338), .ZN(n19340) );
  OAI221_X1 U22356 ( .B1(n19341), .B2(n19632), .C1(n19341), .C2(n19499), .A(
        n19340), .ZN(n19358) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19358), .B1(
        n19375), .B2(n19453), .ZN(n19342) );
  OAI211_X1 U22358 ( .C1(n19398), .C2(n19361), .A(n19343), .B(n19342), .ZN(
        P2_U3136) );
  AOI22_X1 U22359 ( .A1(n19357), .A2(n13050), .B1(n19506), .B2(n19356), .ZN(
        n19345) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19358), .B1(
        n19375), .B2(n19461), .ZN(n19344) );
  OAI211_X1 U22361 ( .C1(n19404), .C2(n19361), .A(n19345), .B(n19344), .ZN(
        P2_U3137) );
  AOI22_X1 U22362 ( .A1(n19357), .A2(n19030), .B1(n19511), .B2(n19356), .ZN(
        n19347) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19358), .B1(
        n19375), .B2(n19464), .ZN(n19346) );
  OAI211_X1 U22364 ( .C1(n19410), .C2(n19361), .A(n19347), .B(n19346), .ZN(
        P2_U3138) );
  AOI22_X1 U22365 ( .A1(n19357), .A2(n19035), .B1(n19516), .B2(n19356), .ZN(
        n19349) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19358), .B1(
        n19375), .B2(n19467), .ZN(n19348) );
  OAI211_X1 U22367 ( .C1(n19416), .C2(n19361), .A(n19349), .B(n19348), .ZN(
        P2_U3139) );
  AOI22_X1 U22368 ( .A1(n19357), .A2(n19522), .B1(n19356), .B2(n19521), .ZN(
        n19351) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19358), .B1(
        n19375), .B2(n19470), .ZN(n19350) );
  OAI211_X1 U22370 ( .C1(n19422), .C2(n19361), .A(n19351), .B(n19350), .ZN(
        P2_U3140) );
  AOI22_X1 U22371 ( .A1(n19357), .A2(n19528), .B1(n19527), .B2(n19356), .ZN(
        n19353) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19358), .B1(
        n19375), .B2(n19474), .ZN(n19352) );
  OAI211_X1 U22373 ( .C1(n19428), .C2(n19361), .A(n19353), .B(n19352), .ZN(
        P2_U3141) );
  AOI22_X1 U22374 ( .A1(n19357), .A2(n19534), .B1(n19533), .B2(n19356), .ZN(
        n19355) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19358), .B1(
        n19375), .B2(n19477), .ZN(n19354) );
  OAI211_X1 U22376 ( .C1(n19434), .C2(n19361), .A(n19355), .B(n19354), .ZN(
        P2_U3142) );
  AOI22_X1 U22377 ( .A1(n19357), .A2(n19541), .B1(n19539), .B2(n19356), .ZN(
        n19360) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19358), .B1(
        n19375), .B2(n19482), .ZN(n19359) );
  OAI211_X1 U22379 ( .C1(n19444), .C2(n19361), .A(n19360), .B(n19359), .ZN(
        P2_U3143) );
  AOI22_X1 U22380 ( .A1(n19374), .A2(n19030), .B1(n19373), .B2(n19511), .ZN(
        n19363) );
  AOI22_X1 U22381 ( .A1(n19375), .A2(n19512), .B1(n19380), .B2(n19464), .ZN(
        n19362) );
  OAI211_X1 U22382 ( .C1(n19379), .C2(n19364), .A(n19363), .B(n19362), .ZN(
        P2_U3146) );
  AOI22_X1 U22383 ( .A1(n19374), .A2(n19035), .B1(n19373), .B2(n19516), .ZN(
        n19366) );
  AOI22_X1 U22384 ( .A1(n19375), .A2(n19517), .B1(n19380), .B2(n19467), .ZN(
        n19365) );
  OAI211_X1 U22385 ( .C1(n19379), .C2(n14191), .A(n19366), .B(n19365), .ZN(
        P2_U3147) );
  AOI22_X1 U22386 ( .A1(n19374), .A2(n19522), .B1(n19373), .B2(n19521), .ZN(
        n19368) );
  AOI22_X1 U22387 ( .A1(n19375), .A2(n19523), .B1(n19380), .B2(n19470), .ZN(
        n19367) );
  OAI211_X1 U22388 ( .C1(n19379), .C2(n14208), .A(n19368), .B(n19367), .ZN(
        P2_U3148) );
  AOI22_X1 U22389 ( .A1(n19374), .A2(n19528), .B1(n19373), .B2(n19527), .ZN(
        n19370) );
  AOI22_X1 U22390 ( .A1(n19375), .A2(n19529), .B1(n19380), .B2(n19474), .ZN(
        n19369) );
  OAI211_X1 U22391 ( .C1(n19379), .C2(n14243), .A(n19370), .B(n19369), .ZN(
        P2_U3149) );
  AOI22_X1 U22392 ( .A1(n19374), .A2(n19534), .B1(n19373), .B2(n19533), .ZN(
        n19372) );
  AOI22_X1 U22393 ( .A1(n19375), .A2(n19535), .B1(n19380), .B2(n19477), .ZN(
        n19371) );
  OAI211_X1 U22394 ( .C1(n19379), .C2(n14266), .A(n19372), .B(n19371), .ZN(
        P2_U3150) );
  INV_X1 U22395 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n19378) );
  AOI22_X1 U22396 ( .A1(n19374), .A2(n19541), .B1(n19373), .B2(n19539), .ZN(
        n19377) );
  AOI22_X1 U22397 ( .A1(n19375), .A2(n19543), .B1(n19380), .B2(n19482), .ZN(
        n19376) );
  OAI211_X1 U22398 ( .C1(n19379), .C2(n19378), .A(n19377), .B(n19376), .ZN(
        P2_U3151) );
  NOR2_X1 U22399 ( .A1(n19666), .A2(n19390), .ZN(n19451) );
  INV_X1 U22400 ( .A(n19451), .ZN(n19435) );
  NAND2_X1 U22401 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19435), .ZN(n19381) );
  NOR2_X1 U22402 ( .A1(n19382), .A2(n19381), .ZN(n19389) );
  INV_X1 U22403 ( .A(n19390), .ZN(n19383) );
  AOI21_X1 U22404 ( .B1(n19639), .B2(n19383), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19384) );
  OAI22_X1 U22405 ( .A1(n19438), .A2(n19386), .B1(n19385), .B2(n19435), .ZN(
        n19387) );
  INV_X1 U22406 ( .A(n19387), .ZN(n19397) );
  NAND2_X1 U22407 ( .A1(n19499), .A2(n19388), .ZN(n19391) );
  AOI21_X1 U22408 ( .B1(n19391), .B2(n19390), .A(n19389), .ZN(n19393) );
  OAI211_X1 U22409 ( .C1(n19451), .C2(n19639), .A(n19393), .B(n19392), .ZN(
        n19440) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19440), .B1(
        n19483), .B2(n19453), .ZN(n19396) );
  OAI211_X1 U22411 ( .C1(n19398), .C2(n19443), .A(n19397), .B(n19396), .ZN(
        P2_U3152) );
  OAI22_X1 U22412 ( .A1(n19438), .A2(n19400), .B1(n19399), .B2(n19435), .ZN(
        n19401) );
  INV_X1 U22413 ( .A(n19401), .ZN(n19403) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19440), .B1(
        n19483), .B2(n19461), .ZN(n19402) );
  OAI211_X1 U22415 ( .C1(n19404), .C2(n19443), .A(n19403), .B(n19402), .ZN(
        P2_U3153) );
  INV_X1 U22416 ( .A(n19511), .ZN(n19405) );
  OAI22_X1 U22417 ( .A1(n19438), .A2(n19406), .B1(n19405), .B2(n19435), .ZN(
        n19407) );
  INV_X1 U22418 ( .A(n19407), .ZN(n19409) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19440), .B1(
        n19483), .B2(n19464), .ZN(n19408) );
  OAI211_X1 U22420 ( .C1(n19410), .C2(n19443), .A(n19409), .B(n19408), .ZN(
        P2_U3154) );
  INV_X1 U22421 ( .A(n19516), .ZN(n19411) );
  OAI22_X1 U22422 ( .A1(n19438), .A2(n19412), .B1(n19411), .B2(n19435), .ZN(
        n19413) );
  INV_X1 U22423 ( .A(n19413), .ZN(n19415) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19440), .B1(
        n19483), .B2(n19467), .ZN(n19414) );
  OAI211_X1 U22425 ( .C1(n19416), .C2(n19443), .A(n19415), .B(n19414), .ZN(
        P2_U3155) );
  OAI22_X1 U22426 ( .A1(n19438), .A2(n19418), .B1(n19435), .B2(n19417), .ZN(
        n19419) );
  INV_X1 U22427 ( .A(n19419), .ZN(n19421) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19440), .B1(
        n19483), .B2(n19470), .ZN(n19420) );
  OAI211_X1 U22429 ( .C1(n19422), .C2(n19443), .A(n19421), .B(n19420), .ZN(
        P2_U3156) );
  INV_X1 U22430 ( .A(n19527), .ZN(n19423) );
  OAI22_X1 U22431 ( .A1(n19438), .A2(n19424), .B1(n19423), .B2(n19435), .ZN(
        n19425) );
  INV_X1 U22432 ( .A(n19425), .ZN(n19427) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19440), .B1(
        n19483), .B2(n19474), .ZN(n19426) );
  OAI211_X1 U22434 ( .C1(n19428), .C2(n19443), .A(n19427), .B(n19426), .ZN(
        P2_U3157) );
  INV_X1 U22435 ( .A(n19533), .ZN(n19429) );
  OAI22_X1 U22436 ( .A1(n19438), .A2(n19430), .B1(n19429), .B2(n19435), .ZN(
        n19431) );
  INV_X1 U22437 ( .A(n19431), .ZN(n19433) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19440), .B1(
        n19483), .B2(n19477), .ZN(n19432) );
  OAI211_X1 U22439 ( .C1(n19434), .C2(n19443), .A(n19433), .B(n19432), .ZN(
        P2_U3158) );
  INV_X1 U22440 ( .A(n19539), .ZN(n19436) );
  OAI22_X1 U22441 ( .A1(n19438), .A2(n19437), .B1(n19436), .B2(n19435), .ZN(
        n19439) );
  INV_X1 U22442 ( .A(n19439), .ZN(n19442) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19440), .B1(
        n19483), .B2(n19482), .ZN(n19441) );
  OAI211_X1 U22444 ( .C1(n19444), .C2(n19443), .A(n19442), .B(n19441), .ZN(
        P2_U3159) );
  INV_X1 U22445 ( .A(n19544), .ZN(n19448) );
  INV_X1 U22446 ( .A(n19483), .ZN(n19447) );
  NAND2_X1 U22447 ( .A1(n19448), .A2(n19447), .ZN(n19450) );
  AOI21_X1 U22448 ( .B1(n19450), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19449), 
        .ZN(n19454) );
  NOR3_X2 U22449 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12670), .A3(
        n19489), .ZN(n19481) );
  NOR2_X1 U22450 ( .A1(n19481), .A2(n19451), .ZN(n19456) );
  AOI22_X1 U22451 ( .A1(n19453), .A2(n19544), .B1(n19494), .B2(n19481), .ZN(
        n19459) );
  INV_X1 U22452 ( .A(n19454), .ZN(n19457) );
  OAI21_X1 U22453 ( .B1(n10524), .B2(n19481), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19455) );
  AOI22_X1 U22454 ( .A1(n13025), .A2(n19484), .B1(n19483), .B2(n19502), .ZN(
        n19458) );
  OAI211_X1 U22455 ( .C1(n19488), .C2(n19460), .A(n19459), .B(n19458), .ZN(
        P2_U3160) );
  AOI22_X1 U22456 ( .A1(n19461), .A2(n19544), .B1(n19506), .B2(n19481), .ZN(
        n19463) );
  AOI22_X1 U22457 ( .A1(n13050), .A2(n19484), .B1(n19483), .B2(n19507), .ZN(
        n19462) );
  OAI211_X1 U22458 ( .C1(n19488), .C2(n14142), .A(n19463), .B(n19462), .ZN(
        P2_U3161) );
  AOI22_X1 U22459 ( .A1(n19512), .A2(n19483), .B1(n19511), .B2(n19481), .ZN(
        n19466) );
  AOI22_X1 U22460 ( .A1(n19030), .A2(n19484), .B1(n19544), .B2(n19464), .ZN(
        n19465) );
  OAI211_X1 U22461 ( .C1(n19488), .C2(n14168), .A(n19466), .B(n19465), .ZN(
        P2_U3162) );
  AOI22_X1 U22462 ( .A1(n19517), .A2(n19483), .B1(n19516), .B2(n19481), .ZN(
        n19469) );
  AOI22_X1 U22463 ( .A1(n19035), .A2(n19484), .B1(n19544), .B2(n19467), .ZN(
        n19468) );
  OAI211_X1 U22464 ( .C1(n19488), .C2(n14193), .A(n19469), .B(n19468), .ZN(
        P2_U3163) );
  INV_X1 U22465 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19473) );
  AOI22_X1 U22466 ( .A1(n19470), .A2(n19544), .B1(n19521), .B2(n19481), .ZN(
        n19472) );
  AOI22_X1 U22467 ( .A1(n19522), .A2(n19484), .B1(n19483), .B2(n19523), .ZN(
        n19471) );
  OAI211_X1 U22468 ( .C1(n19488), .C2(n19473), .A(n19472), .B(n19471), .ZN(
        P2_U3164) );
  AOI22_X1 U22469 ( .A1(n19529), .A2(n19483), .B1(n19527), .B2(n19481), .ZN(
        n19476) );
  AOI22_X1 U22470 ( .A1(n19528), .A2(n19484), .B1(n19544), .B2(n19474), .ZN(
        n19475) );
  OAI211_X1 U22471 ( .C1(n19488), .C2(n14245), .A(n19476), .B(n19475), .ZN(
        P2_U3165) );
  INV_X1 U22472 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n19480) );
  AOI22_X1 U22473 ( .A1(n19535), .A2(n19483), .B1(n19533), .B2(n19481), .ZN(
        n19479) );
  AOI22_X1 U22474 ( .A1(n19534), .A2(n19484), .B1(n19544), .B2(n19477), .ZN(
        n19478) );
  OAI211_X1 U22475 ( .C1(n19488), .C2(n19480), .A(n19479), .B(n19478), .ZN(
        P2_U3166) );
  INV_X1 U22476 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19487) );
  AOI22_X1 U22477 ( .A1(n19482), .A2(n19544), .B1(n19539), .B2(n19481), .ZN(
        n19486) );
  AOI22_X1 U22478 ( .A1(n19541), .A2(n19484), .B1(n19483), .B2(n19543), .ZN(
        n19485) );
  OAI211_X1 U22479 ( .C1(n19488), .C2(n19487), .A(n19486), .B(n19485), .ZN(
        P2_U3167) );
  NOR2_X1 U22480 ( .A1(n12670), .A2(n19489), .ZN(n19501) );
  INV_X1 U22481 ( .A(n19501), .ZN(n19490) );
  OR2_X1 U22482 ( .A1(n19490), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19492) );
  NOR3_X1 U22483 ( .A1(n19491), .A2(n19540), .A3(n19493), .ZN(n19495) );
  AOI21_X1 U22484 ( .B1(n19493), .B2(n19492), .A(n19495), .ZN(n19542) );
  AOI22_X1 U22485 ( .A1(n19542), .A2(n13025), .B1(n19540), .B2(n19494), .ZN(
        n19504) );
  AOI211_X1 U22486 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19497), .A(n19496), 
        .B(n19495), .ZN(n19498) );
  OAI221_X1 U22487 ( .B1(n19501), .B2(n19500), .C1(n19501), .C2(n19499), .A(
        n19498), .ZN(n19545) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19502), .ZN(n19503) );
  OAI211_X1 U22489 ( .C1(n19505), .C2(n19548), .A(n19504), .B(n19503), .ZN(
        P2_U3168) );
  AOI22_X1 U22490 ( .A1(n19542), .A2(n13050), .B1(n19540), .B2(n19506), .ZN(
        n19509) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19507), .ZN(n19508) );
  OAI211_X1 U22492 ( .C1(n19510), .C2(n19548), .A(n19509), .B(n19508), .ZN(
        P2_U3169) );
  AOI22_X1 U22493 ( .A1(n19542), .A2(n19030), .B1(n19540), .B2(n19511), .ZN(
        n19514) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19512), .ZN(n19513) );
  OAI211_X1 U22495 ( .C1(n19515), .C2(n19548), .A(n19514), .B(n19513), .ZN(
        P2_U3170) );
  AOI22_X1 U22496 ( .A1(n19542), .A2(n19035), .B1(n19540), .B2(n19516), .ZN(
        n19519) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19517), .ZN(n19518) );
  OAI211_X1 U22498 ( .C1(n19520), .C2(n19548), .A(n19519), .B(n19518), .ZN(
        P2_U3171) );
  AOI22_X1 U22499 ( .A1(n19542), .A2(n19522), .B1(n19540), .B2(n19521), .ZN(
        n19525) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19523), .ZN(n19524) );
  OAI211_X1 U22501 ( .C1(n19526), .C2(n19548), .A(n19525), .B(n19524), .ZN(
        P2_U3172) );
  AOI22_X1 U22502 ( .A1(n19542), .A2(n19528), .B1(n19540), .B2(n19527), .ZN(
        n19531) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19529), .ZN(n19530) );
  OAI211_X1 U22504 ( .C1(n19532), .C2(n19548), .A(n19531), .B(n19530), .ZN(
        P2_U3173) );
  AOI22_X1 U22505 ( .A1(n19542), .A2(n19534), .B1(n19540), .B2(n19533), .ZN(
        n19537) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19535), .ZN(n19536) );
  OAI211_X1 U22507 ( .C1(n19538), .C2(n19548), .A(n19537), .B(n19536), .ZN(
        P2_U3174) );
  AOI22_X1 U22508 ( .A1(n19542), .A2(n19541), .B1(n19540), .B2(n19539), .ZN(
        n19547) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19543), .ZN(n19546) );
  OAI211_X1 U22510 ( .C1(n19549), .C2(n19548), .A(n19547), .B(n19546), .ZN(
        P2_U3175) );
  INV_X1 U22511 ( .A(n19550), .ZN(n19552) );
  OAI211_X1 U22512 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19685), .A(n19552), 
        .B(n19551), .ZN(n19557) );
  OAI21_X1 U22513 ( .B1(n19554), .B2(n19553), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n19556) );
  OAI211_X1 U22514 ( .C1(n19558), .C2(n19557), .A(n19556), .B(n19555), .ZN(
        P2_U3177) );
  AND2_X1 U22515 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19559), .ZN(
        P2_U3179) );
  AND2_X1 U22516 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19559), .ZN(
        P2_U3180) );
  AND2_X1 U22517 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19559), .ZN(
        P2_U3181) );
  AND2_X1 U22518 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19559), .ZN(
        P2_U3182) );
  AND2_X1 U22519 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19559), .ZN(
        P2_U3183) );
  AND2_X1 U22520 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19559), .ZN(
        P2_U3184) );
  AND2_X1 U22521 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19559), .ZN(
        P2_U3185) );
  AND2_X1 U22522 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19559), .ZN(
        P2_U3186) );
  AND2_X1 U22523 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19559), .ZN(
        P2_U3187) );
  AND2_X1 U22524 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19559), .ZN(
        P2_U3188) );
  AND2_X1 U22525 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19559), .ZN(
        P2_U3189) );
  AND2_X1 U22526 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19559), .ZN(
        P2_U3190) );
  AND2_X1 U22527 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19559), .ZN(
        P2_U3191) );
  AND2_X1 U22528 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19559), .ZN(
        P2_U3192) );
  AND2_X1 U22529 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19559), .ZN(
        P2_U3193) );
  AND2_X1 U22530 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19559), .ZN(
        P2_U3194) );
  AND2_X1 U22531 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19559), .ZN(
        P2_U3195) );
  AND2_X1 U22532 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19559), .ZN(
        P2_U3196) );
  AND2_X1 U22533 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19559), .ZN(
        P2_U3197) );
  AND2_X1 U22534 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19559), .ZN(
        P2_U3198) );
  AND2_X1 U22535 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19559), .ZN(
        P2_U3199) );
  AND2_X1 U22536 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19559), .ZN(
        P2_U3200) );
  AND2_X1 U22537 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19559), .ZN(P2_U3201) );
  AND2_X1 U22538 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19559), .ZN(P2_U3202) );
  AND2_X1 U22539 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19559), .ZN(P2_U3203) );
  AND2_X1 U22540 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19559), .ZN(P2_U3204) );
  AND2_X1 U22541 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19559), .ZN(P2_U3205) );
  AND2_X1 U22542 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19559), .ZN(P2_U3206) );
  AND2_X1 U22543 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19559), .ZN(P2_U3207) );
  AND2_X1 U22544 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19559), .ZN(P2_U3208) );
  NOR2_X1 U22545 ( .A1(n19685), .A2(n20696), .ZN(n19571) );
  INV_X1 U22546 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19694) );
  OR3_X1 U22547 ( .A1(n19571), .A2(n19694), .A3(n19560), .ZN(n19562) );
  AOI211_X1 U22548 ( .C1(n20581), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19572), .B(n19613), .ZN(n19561) );
  NOR2_X1 U22549 ( .A1(n20587), .A2(n19564), .ZN(n19577) );
  AOI211_X1 U22550 ( .C1(n19578), .C2(n19562), .A(n19561), .B(n19577), .ZN(
        n19563) );
  INV_X1 U22551 ( .A(n19563), .ZN(P2_U3209) );
  AOI21_X1 U22552 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20581), .A(n19578), 
        .ZN(n19569) );
  NOR2_X1 U22553 ( .A1(n19694), .A2(n19569), .ZN(n19565) );
  AOI21_X1 U22554 ( .B1(n19565), .B2(n19564), .A(n19571), .ZN(n19567) );
  OAI211_X1 U22555 ( .C1(n20581), .C2(n19568), .A(n19567), .B(n19566), .ZN(
        P2_U3210) );
  AOI21_X1 U22556 ( .B1(n19570), .B2(n19680), .A(n19569), .ZN(n19576) );
  AOI22_X1 U22557 ( .A1(n19694), .A2(n19572), .B1(n20587), .B2(n19571), .ZN(
        n19573) );
  INV_X1 U22558 ( .A(n19573), .ZN(n19574) );
  OAI211_X1 U22559 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19574), .ZN(n19575) );
  OAI21_X1 U22560 ( .B1(n19577), .B2(n19576), .A(n19575), .ZN(P2_U3211) );
  NAND2_X1 U22561 ( .A1(n19613), .A2(n19578), .ZN(n19622) );
  CLKBUF_X1 U22562 ( .A(n19622), .Z(n19619) );
  NAND2_X2 U22563 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19613), .ZN(n19620) );
  OAI222_X1 U22564 ( .A1(n19619), .A2(n10269), .B1(n19579), .B2(n19613), .C1(
        n10240), .C2(n19620), .ZN(P2_U3212) );
  OAI222_X1 U22565 ( .A1(n19620), .A2(n10269), .B1(n19580), .B2(n19613), .C1(
        n12737), .C2(n19619), .ZN(P2_U3213) );
  OAI222_X1 U22566 ( .A1(n19620), .A2(n12737), .B1(n19581), .B2(n19613), .C1(
        n10842), .C2(n19619), .ZN(P2_U3214) );
  OAI222_X1 U22567 ( .A1(n19622), .A2(n10845), .B1(n19582), .B2(n19613), .C1(
        n10842), .C2(n19620), .ZN(P2_U3215) );
  OAI222_X1 U22568 ( .A1(n19622), .A2(n10855), .B1(n19583), .B2(n19613), .C1(
        n10845), .C2(n19620), .ZN(P2_U3216) );
  OAI222_X1 U22569 ( .A1(n19622), .A2(n10861), .B1(n19584), .B2(n19613), .C1(
        n10855), .C2(n19620), .ZN(P2_U3217) );
  OAI222_X1 U22570 ( .A1(n19622), .A2(n10875), .B1(n19585), .B2(n19613), .C1(
        n10861), .C2(n19620), .ZN(P2_U3218) );
  OAI222_X1 U22571 ( .A1(n19622), .A2(n10879), .B1(n19586), .B2(n19613), .C1(
        n10875), .C2(n19620), .ZN(P2_U3219) );
  OAI222_X1 U22572 ( .A1(n19619), .A2(n10905), .B1(n19587), .B2(n19613), .C1(
        n10879), .C2(n19620), .ZN(P2_U3220) );
  INV_X1 U22573 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19589) );
  OAI222_X1 U22574 ( .A1(n19619), .A2(n19589), .B1(n19588), .B2(n19613), .C1(
        n10905), .C2(n19620), .ZN(P2_U3221) );
  OAI222_X1 U22575 ( .A1(n19619), .A2(n10932), .B1(n19590), .B2(n19613), .C1(
        n19589), .C2(n19620), .ZN(P2_U3222) );
  OAI222_X1 U22576 ( .A1(n19619), .A2(n10936), .B1(n19591), .B2(n19613), .C1(
        n10932), .C2(n19620), .ZN(P2_U3223) );
  OAI222_X1 U22577 ( .A1(n19619), .A2(n10962), .B1(n19592), .B2(n19613), .C1(
        n10936), .C2(n19620), .ZN(P2_U3224) );
  OAI222_X1 U22578 ( .A1(n19619), .A2(n11091), .B1(n19593), .B2(n19613), .C1(
        n10962), .C2(n19620), .ZN(P2_U3225) );
  OAI222_X1 U22579 ( .A1(n19622), .A2(n19595), .B1(n19594), .B2(n19613), .C1(
        n11091), .C2(n19620), .ZN(P2_U3226) );
  OAI222_X1 U22580 ( .A1(n19622), .A2(n10984), .B1(n19596), .B2(n19613), .C1(
        n19595), .C2(n19620), .ZN(P2_U3227) );
  OAI222_X1 U22581 ( .A1(n19622), .A2(n19598), .B1(n19597), .B2(n19613), .C1(
        n10984), .C2(n19620), .ZN(P2_U3228) );
  OAI222_X1 U22582 ( .A1(n19622), .A2(n15097), .B1(n19599), .B2(n19613), .C1(
        n19598), .C2(n19620), .ZN(P2_U3229) );
  OAI222_X1 U22583 ( .A1(n19622), .A2(n19601), .B1(n19600), .B2(n19613), .C1(
        n15097), .C2(n19620), .ZN(P2_U3230) );
  OAI222_X1 U22584 ( .A1(n19622), .A2(n19602), .B1(n20761), .B2(n19613), .C1(
        n19601), .C2(n19620), .ZN(P2_U3231) );
  OAI222_X1 U22585 ( .A1(n19619), .A2(n19604), .B1(n19603), .B2(n19613), .C1(
        n19602), .C2(n19620), .ZN(P2_U3232) );
  OAI222_X1 U22586 ( .A1(n19619), .A2(n10998), .B1(n19605), .B2(n19613), .C1(
        n19604), .C2(n19620), .ZN(P2_U3233) );
  OAI222_X1 U22587 ( .A1(n19619), .A2(n19607), .B1(n19606), .B2(n19613), .C1(
        n10998), .C2(n19620), .ZN(P2_U3234) );
  OAI222_X1 U22588 ( .A1(n19619), .A2(n19609), .B1(n19608), .B2(n19613), .C1(
        n19607), .C2(n19620), .ZN(P2_U3235) );
  OAI222_X1 U22589 ( .A1(n19619), .A2(n19611), .B1(n19610), .B2(n19613), .C1(
        n19609), .C2(n19620), .ZN(P2_U3236) );
  OAI222_X1 U22590 ( .A1(n19619), .A2(n19615), .B1(n19612), .B2(n19613), .C1(
        n19611), .C2(n19620), .ZN(P2_U3237) );
  OAI222_X1 U22591 ( .A1(n19620), .A2(n19615), .B1(n19614), .B2(n19613), .C1(
        n19616), .C2(n19619), .ZN(P2_U3238) );
  OAI222_X1 U22592 ( .A1(n19619), .A2(n14037), .B1(n19617), .B2(n19613), .C1(
        n19616), .C2(n19620), .ZN(P2_U3239) );
  OAI222_X1 U22593 ( .A1(n19619), .A2(n15022), .B1(n19618), .B2(n19613), .C1(
        n14037), .C2(n19620), .ZN(P2_U3240) );
  OAI222_X1 U22594 ( .A1(n19622), .A2(n14029), .B1(n19621), .B2(n19613), .C1(
        n15022), .C2(n19620), .ZN(P2_U3241) );
  INV_X1 U22595 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19623) );
  AOI22_X1 U22596 ( .A1(n19613), .A2(n20739), .B1(n19623), .B2(n19695), .ZN(
        P2_U3585) );
  MUX2_X1 U22597 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19613), .Z(P2_U3586) );
  INV_X1 U22598 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19624) );
  AOI22_X1 U22599 ( .A1(n19613), .A2(n19625), .B1(n19624), .B2(n19695), .ZN(
        P2_U3587) );
  INV_X1 U22600 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19626) );
  AOI22_X1 U22601 ( .A1(n19613), .A2(n19627), .B1(n19626), .B2(n19695), .ZN(
        P2_U3588) );
  OAI21_X1 U22602 ( .B1(n19631), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19629), 
        .ZN(n19628) );
  INV_X1 U22603 ( .A(n19628), .ZN(P2_U3591) );
  OAI21_X1 U22604 ( .B1(n19631), .B2(n19630), .A(n19629), .ZN(P2_U3592) );
  AND2_X1 U22605 ( .A1(n19642), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19655) );
  NAND2_X1 U22606 ( .A1(n19632), .A2(n19655), .ZN(n19645) );
  OR2_X1 U22607 ( .A1(n19634), .A2(n19633), .ZN(n19635) );
  OAI21_X1 U22608 ( .B1(n19654), .B2(n19635), .A(n19662), .ZN(n19646) );
  NAND2_X1 U22609 ( .A1(n19645), .A2(n19646), .ZN(n19637) );
  NAND2_X1 U22610 ( .A1(n19637), .A2(n19636), .ZN(n19638) );
  OAI21_X1 U22611 ( .B1(n19640), .B2(n19639), .A(n19638), .ZN(n19641) );
  AOI21_X1 U22612 ( .B1(n19643), .B2(n19642), .A(n19641), .ZN(n19644) );
  AOI22_X1 U22613 ( .A1(n19667), .A2(n12670), .B1(n19644), .B2(n19664), .ZN(
        P2_U3602) );
  OAI21_X1 U22614 ( .B1(n19647), .B2(n19646), .A(n19645), .ZN(n19648) );
  AOI21_X1 U22615 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19649), .A(n19648), 
        .ZN(n19650) );
  AOI22_X1 U22616 ( .A1(n19667), .A2(n19651), .B1(n19650), .B2(n19664), .ZN(
        P2_U3603) );
  INV_X1 U22617 ( .A(n19662), .ZN(n19653) );
  NOR2_X1 U22618 ( .A1(n19653), .A2(n19652), .ZN(n19656) );
  MUX2_X1 U22619 ( .A(n19656), .B(n19655), .S(n19654), .Z(n19657) );
  AOI21_X1 U22620 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19658), .A(n19657), 
        .ZN(n19659) );
  AOI22_X1 U22621 ( .A1(n19667), .A2(n10817), .B1(n19659), .B2(n19664), .ZN(
        P2_U3604) );
  NOR2_X1 U22622 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19639), .ZN(
        n19661) );
  AOI211_X1 U22623 ( .C1(n19663), .C2(n19662), .A(n19661), .B(n19660), .ZN(
        n19665) );
  AOI22_X1 U22624 ( .A1(n19667), .A2(n19666), .B1(n19665), .B2(n19664), .ZN(
        P2_U3605) );
  INV_X1 U22625 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19668) );
  AOI22_X1 U22626 ( .A1(n19613), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19668), 
        .B2(n19695), .ZN(P2_U3608) );
  INV_X1 U22627 ( .A(n19669), .ZN(n19674) );
  NAND2_X1 U22628 ( .A1(n19671), .A2(n19670), .ZN(n19672) );
  OAI211_X1 U22629 ( .C1(n19675), .C2(n19674), .A(n19673), .B(n19672), .ZN(
        n19677) );
  MUX2_X1 U22630 ( .A(P2_MORE_REG_SCAN_IN), .B(n19677), .S(n19676), .Z(
        P2_U3609) );
  OAI21_X1 U22631 ( .B1(n19680), .B2(n19679), .A(n19678), .ZN(n19681) );
  AOI21_X1 U22632 ( .B1(n19639), .B2(n19682), .A(n19681), .ZN(n19693) );
  NOR4_X1 U22633 ( .A1(n19688), .A2(n19683), .A3(n10217), .A4(n12317), .ZN(
        n19687) );
  AOI21_X1 U22634 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19685), .A(n19684), 
        .ZN(n19686) );
  NOR2_X1 U22635 ( .A1(n19687), .A2(n19686), .ZN(n19692) );
  AOI21_X1 U22636 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19688), .A(n9573), 
        .ZN(n19689) );
  AOI21_X1 U22637 ( .B1(n19690), .B2(n19689), .A(n19693), .ZN(n19691) );
  AOI22_X1 U22638 ( .A1(n19694), .A2(n19693), .B1(n19692), .B2(n19691), .ZN(
        P2_U3610) );
  INV_X1 U22639 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19696) );
  AOI22_X1 U22640 ( .A1(n19613), .A2(n19697), .B1(n19696), .B2(n19695), .ZN(
        P2_U3611) );
  OAI21_X1 U22641 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n19698), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20590) );
  OAI21_X1 U22642 ( .B1(n20590), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20675), .ZN(
        n19699) );
  INV_X1 U22643 ( .A(n19699), .ZN(P1_U2802) );
  NAND2_X1 U22644 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n19700), .ZN(n19705) );
  INV_X1 U22645 ( .A(n19701), .ZN(n19702) );
  OAI21_X1 U22646 ( .B1(n19703), .B2(n19702), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19704) );
  OAI21_X1 U22647 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19705), .A(n19704), 
        .ZN(P1_U2803) );
  NOR2_X1 U22648 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19707) );
  OAI21_X1 U22649 ( .B1(n19707), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20675), .ZN(
        n19706) );
  OAI21_X1 U22650 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20675), .A(n19706), 
        .ZN(P1_U2804) );
  INV_X1 U22651 ( .A(n20649), .ZN(n20653) );
  OAI21_X1 U22652 ( .B1(BS16), .B2(n19707), .A(n20653), .ZN(n20651) );
  OAI21_X1 U22653 ( .B1(n20653), .B2(n20055), .A(n20651), .ZN(P1_U2805) );
  OAI21_X1 U22654 ( .B1(n19710), .B2(n19709), .A(n19708), .ZN(P1_U2806) );
  NOR4_X1 U22655 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19714) );
  NOR4_X1 U22656 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19713) );
  NOR4_X1 U22657 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19712) );
  NOR4_X1 U22658 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19711) );
  NAND4_X1 U22659 ( .A1(n19714), .A2(n19713), .A3(n19712), .A4(n19711), .ZN(
        n19720) );
  NOR4_X1 U22660 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19718) );
  AOI211_X1 U22661 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_11__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19717) );
  NOR4_X1 U22662 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19716) );
  NOR4_X1 U22663 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19715) );
  NAND4_X1 U22664 ( .A1(n19718), .A2(n19717), .A3(n19716), .A4(n19715), .ZN(
        n19719) );
  NOR2_X1 U22665 ( .A1(n19720), .A2(n19719), .ZN(n20657) );
  INV_X1 U22666 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20646) );
  NOR3_X1 U22667 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19722) );
  OAI21_X1 U22668 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19722), .A(n20657), .ZN(
        n19721) );
  OAI21_X1 U22669 ( .B1(n20657), .B2(n20646), .A(n19721), .ZN(P1_U2807) );
  INV_X1 U22670 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20652) );
  AOI21_X1 U22671 ( .B1(n12892), .B2(n20652), .A(n19722), .ZN(n19723) );
  INV_X1 U22672 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20758) );
  INV_X1 U22673 ( .A(n20657), .ZN(n20660) );
  AOI22_X1 U22674 ( .A1(n20657), .A2(n19723), .B1(n20758), .B2(n20660), .ZN(
        P1_U2808) );
  NOR2_X1 U22675 ( .A1(n19724), .A2(n19747), .ZN(n19737) );
  NOR2_X1 U22676 ( .A1(n19725), .A2(n19737), .ZN(n19746) );
  AOI22_X1 U22677 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n19774), .B1(n19773), .B2(
        n19791), .ZN(n19732) );
  INV_X1 U22678 ( .A(n19726), .ZN(n19730) );
  OAI21_X1 U22679 ( .B1(n19728), .B2(n19727), .A(n19927), .ZN(n19729) );
  AOI21_X1 U22680 ( .B1(n19778), .B2(n19730), .A(n19729), .ZN(n19731) );
  OAI211_X1 U22681 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n19733), .A(n19732), .B(
        n19731), .ZN(n19734) );
  AOI21_X1 U22682 ( .B1(n19794), .B2(n19755), .A(n19734), .ZN(n19735) );
  OAI21_X1 U22683 ( .B1(n19746), .B2(n20605), .A(n19735), .ZN(P1_U2831) );
  INV_X1 U22684 ( .A(n19736), .ZN(n19738) );
  AOI22_X1 U22685 ( .A1(n19739), .A2(n19778), .B1(n19738), .B2(n19737), .ZN(
        n19745) );
  AOI22_X1 U22686 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(n19774), .ZN(n19740) );
  OAI211_X1 U22687 ( .C1(n19741), .C2(n19761), .A(n19927), .B(n19740), .ZN(
        n19742) );
  AOI21_X1 U22688 ( .B1(n19743), .B2(n19755), .A(n19742), .ZN(n19744) );
  OAI211_X1 U22689 ( .C1(n19746), .C2(n20603), .A(n19745), .B(n19744), .ZN(
        P1_U2832) );
  NOR2_X1 U22690 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19747), .ZN(n19748) );
  AOI22_X1 U22691 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n19774), .B1(n19749), .B2(
        n19748), .ZN(n19759) );
  OAI22_X1 U22692 ( .A1(n19752), .A2(n19751), .B1(n19761), .B2(n19750), .ZN(
        n19753) );
  AOI211_X1 U22693 ( .C1(n19779), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19913), .B(n19753), .ZN(n19758) );
  AOI22_X1 U22694 ( .A1(n19756), .A2(n19755), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n19754), .ZN(n19757) );
  NAND3_X1 U22695 ( .A1(n19759), .A2(n19758), .A3(n19757), .ZN(P1_U2833) );
  AOI22_X1 U22696 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19779), .B1(
        P1_EBX_REG_4__SCAN_IN), .B2(n19774), .ZN(n19771) );
  INV_X1 U22697 ( .A(n19911), .ZN(n19765) );
  INV_X1 U22698 ( .A(n19760), .ZN(n19763) );
  OAI22_X1 U22699 ( .A1(n19763), .A2(n19762), .B1(n19761), .B2(n19928), .ZN(
        n19764) );
  AOI21_X1 U22700 ( .B1(n19765), .B2(n19778), .A(n19764), .ZN(n19770) );
  NAND2_X1 U22701 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19772) );
  INV_X1 U22702 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20597) );
  OAI21_X1 U22703 ( .B1(n19772), .B2(n19790), .A(n20597), .ZN(n19768) );
  INV_X1 U22704 ( .A(n19766), .ZN(n19785) );
  AOI22_X1 U22705 ( .A1(n19768), .A2(n19767), .B1(n19907), .B2(n19785), .ZN(
        n19769) );
  NAND4_X1 U22706 ( .A1(n19771), .A2(n19770), .A3(n19769), .A4(n19927), .ZN(
        P1_U2836) );
  OAI21_X1 U22707 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .A(n19772), .ZN(n19789) );
  AOI22_X1 U22708 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(n19774), .B1(n19773), .B2(
        n19935), .ZN(n19788) );
  INV_X1 U22709 ( .A(n19775), .ZN(n19783) );
  INV_X1 U22710 ( .A(n19776), .ZN(n19777) );
  AOI22_X1 U22711 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n19779), .B1(
        n19778), .B2(n19777), .ZN(n19782) );
  NAND2_X1 U22712 ( .A1(n20255), .A2(n19780), .ZN(n19781) );
  OAI211_X1 U22713 ( .C1(n19783), .C2(n12905), .A(n19782), .B(n19781), .ZN(
        n19784) );
  AOI21_X1 U22714 ( .B1(n19786), .B2(n19785), .A(n19784), .ZN(n19787) );
  OAI211_X1 U22715 ( .C1(n19790), .C2(n19789), .A(n19788), .B(n19787), .ZN(
        P1_U2837) );
  INV_X1 U22716 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U22717 ( .A1(n19794), .A2(n19793), .B1(n19792), .B2(n19791), .ZN(
        n19795) );
  OAI21_X1 U22718 ( .B1(n19797), .B2(n19796), .A(n19795), .ZN(P1_U2863) );
  INV_X1 U22719 ( .A(n19798), .ZN(n19799) );
  AOI22_X1 U22720 ( .A1(n19799), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20667), .ZN(n19800) );
  OAI21_X1 U22721 ( .B1(n20782), .B2(n19801), .A(n19800), .ZN(P1_U2906) );
  AOI22_X1 U22722 ( .A1(n20667), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19803) );
  OAI21_X1 U22723 ( .B1(n19804), .B2(n19822), .A(n19803), .ZN(P1_U2921) );
  AOI22_X1 U22724 ( .A1(n20667), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19805) );
  OAI21_X1 U22725 ( .B1(n14600), .B2(n19822), .A(n19805), .ZN(P1_U2922) );
  INV_X1 U22726 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19892) );
  AOI22_X1 U22727 ( .A1(n20667), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19806) );
  OAI21_X1 U22728 ( .B1(n19892), .B2(n19822), .A(n19806), .ZN(P1_U2923) );
  AOI22_X1 U22729 ( .A1(n20667), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19807) );
  OAI21_X1 U22730 ( .B1(n20786), .B2(n19822), .A(n19807), .ZN(P1_U2924) );
  INV_X1 U22731 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U22732 ( .A1(n19817), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19808) );
  OAI21_X1 U22733 ( .B1(n19887), .B2(n19822), .A(n19808), .ZN(P1_U2925) );
  INV_X1 U22734 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U22735 ( .A1(n19817), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19809) );
  OAI21_X1 U22736 ( .B1(n19884), .B2(n19822), .A(n19809), .ZN(P1_U2926) );
  INV_X1 U22737 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U22738 ( .A1(n19817), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19810) );
  OAI21_X1 U22739 ( .B1(n19881), .B2(n19822), .A(n19810), .ZN(P1_U2927) );
  AOI22_X1 U22740 ( .A1(n19817), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19811) );
  OAI21_X1 U22741 ( .B1(n13305), .B2(n19822), .A(n19811), .ZN(P1_U2928) );
  AOI22_X1 U22742 ( .A1(n19817), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19812) );
  OAI21_X1 U22743 ( .B1(n19876), .B2(n19822), .A(n19812), .ZN(P1_U2929) );
  AOI22_X1 U22744 ( .A1(n19817), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19813) );
  OAI21_X1 U22745 ( .B1(n19873), .B2(n19822), .A(n19813), .ZN(P1_U2930) );
  AOI22_X1 U22746 ( .A1(n19817), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19814) );
  OAI21_X1 U22747 ( .B1(n13102), .B2(n19822), .A(n19814), .ZN(P1_U2931) );
  INV_X1 U22748 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U22749 ( .A1(n19817), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19815) );
  OAI21_X1 U22750 ( .B1(n19868), .B2(n19822), .A(n19815), .ZN(P1_U2932) );
  AOI22_X1 U22751 ( .A1(n19817), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19816) );
  OAI21_X1 U22752 ( .B1(n20744), .B2(n19822), .A(n19816), .ZN(P1_U2933) );
  AOI22_X1 U22753 ( .A1(n19817), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19818) );
  OAI21_X1 U22754 ( .B1(n19864), .B2(n19822), .A(n19818), .ZN(P1_U2934) );
  AOI22_X1 U22755 ( .A1(n20667), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19819) );
  OAI21_X1 U22756 ( .B1(n19861), .B2(n19822), .A(n19819), .ZN(P1_U2935) );
  AOI22_X1 U22757 ( .A1(n20667), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19820), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19821) );
  OAI21_X1 U22758 ( .B1(n19858), .B2(n19822), .A(n19821), .ZN(P1_U2936) );
  INV_X2 U22759 ( .A(n19899), .ZN(n19897) );
  OAI21_X1 U22760 ( .B1(n19826), .B2(n20666), .A(n19825), .ZN(n19898) );
  OR3_X1 U22761 ( .A1(n19828), .A2(n19827), .A3(n20585), .ZN(n19901) );
  AOI22_X1 U22762 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19856), .ZN(n19829) );
  OAI21_X1 U22763 ( .B1(n20815), .B2(n19897), .A(n19829), .ZN(P1_U2937) );
  AOI22_X1 U22764 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19859), .ZN(n19830) );
  OAI21_X1 U22765 ( .B1(n19831), .B2(n19897), .A(n19830), .ZN(P1_U2938) );
  AOI22_X1 U22766 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19862), .ZN(n19832) );
  OAI21_X1 U22767 ( .B1(n19833), .B2(n19897), .A(n19832), .ZN(P1_U2939) );
  AOI22_X1 U22768 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19865), .ZN(n19834) );
  OAI21_X1 U22769 ( .B1(n19835), .B2(n19897), .A(n19834), .ZN(P1_U2940) );
  AOI22_X1 U22770 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n20002), .ZN(n19836) );
  OAI21_X1 U22771 ( .B1(n19837), .B2(n19897), .A(n19836), .ZN(P1_U2941) );
  AOI22_X1 U22772 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19869), .ZN(n19838) );
  OAI21_X1 U22773 ( .B1(n19839), .B2(n19897), .A(n19838), .ZN(P1_U2942) );
  AOI22_X1 U22774 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19871), .ZN(n19840) );
  OAI21_X1 U22775 ( .B1(n19841), .B2(n19897), .A(n19840), .ZN(P1_U2943) );
  AOI22_X1 U22776 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19898), .B1(n19894), 
        .B2(n19874), .ZN(n19842) );
  OAI21_X1 U22777 ( .B1(n19843), .B2(n19897), .A(n19842), .ZN(P1_U2944) );
  AOI22_X1 U22778 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19898), .B1(n19894), 
        .B2(n19877), .ZN(n19844) );
  OAI21_X1 U22779 ( .B1(n14563), .B2(n19897), .A(n19844), .ZN(P1_U2945) );
  AOI22_X1 U22780 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19898), .B1(n19894), 
        .B2(n19879), .ZN(n19845) );
  OAI21_X1 U22781 ( .B1(n19846), .B2(n19897), .A(n19845), .ZN(P1_U2946) );
  AOI22_X1 U22782 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19898), .B1(n19894), 
        .B2(n19882), .ZN(n19847) );
  OAI21_X1 U22783 ( .B1(n19848), .B2(n19897), .A(n19847), .ZN(P1_U2947) );
  AOI22_X1 U22784 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19885), .ZN(n19849) );
  OAI21_X1 U22785 ( .B1(n19850), .B2(n19897), .A(n19849), .ZN(P1_U2948) );
  AOI22_X1 U22786 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19888), .ZN(n19851) );
  OAI21_X1 U22787 ( .B1(n19852), .B2(n19897), .A(n19851), .ZN(P1_U2949) );
  AOI22_X1 U22788 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19890), .ZN(n19853) );
  OAI21_X1 U22789 ( .B1(n19854), .B2(n19897), .A(n19853), .ZN(P1_U2950) );
  AOI22_X1 U22790 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19893), .ZN(n19855) );
  OAI21_X1 U22791 ( .B1(n14538), .B2(n19897), .A(n19855), .ZN(P1_U2951) );
  AOI22_X1 U22792 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19856), .ZN(n19857) );
  OAI21_X1 U22793 ( .B1(n19858), .B2(n19897), .A(n19857), .ZN(P1_U2952) );
  AOI22_X1 U22794 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19859), .ZN(n19860) );
  OAI21_X1 U22795 ( .B1(n19861), .B2(n19897), .A(n19860), .ZN(P1_U2953) );
  AOI22_X1 U22796 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19862), .ZN(n19863) );
  OAI21_X1 U22797 ( .B1(n19864), .B2(n19897), .A(n19863), .ZN(P1_U2954) );
  AOI22_X1 U22798 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19865), .ZN(n19866) );
  OAI21_X1 U22799 ( .B1(n20744), .B2(n19897), .A(n19866), .ZN(P1_U2955) );
  AOI22_X1 U22800 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n20002), .ZN(n19867) );
  OAI21_X1 U22801 ( .B1(n19868), .B2(n19897), .A(n19867), .ZN(P1_U2956) );
  AOI22_X1 U22802 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19869), .ZN(n19870) );
  OAI21_X1 U22803 ( .B1(n13102), .B2(n19897), .A(n19870), .ZN(P1_U2957) );
  AOI22_X1 U22804 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19871), .ZN(n19872) );
  OAI21_X1 U22805 ( .B1(n19873), .B2(n19897), .A(n19872), .ZN(P1_U2958) );
  AOI22_X1 U22806 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19874), .ZN(n19875) );
  OAI21_X1 U22807 ( .B1(n19876), .B2(n19897), .A(n19875), .ZN(P1_U2959) );
  AOI22_X1 U22808 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19877), .ZN(n19878) );
  OAI21_X1 U22809 ( .B1(n13305), .B2(n19897), .A(n19878), .ZN(P1_U2960) );
  AOI22_X1 U22810 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n19898), .B1(n19894), 
        .B2(n19879), .ZN(n19880) );
  OAI21_X1 U22811 ( .B1(n19881), .B2(n19897), .A(n19880), .ZN(P1_U2961) );
  AOI22_X1 U22812 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19898), .B1(n19894), 
        .B2(n19882), .ZN(n19883) );
  OAI21_X1 U22813 ( .B1(n19884), .B2(n19897), .A(n19883), .ZN(P1_U2962) );
  AOI22_X1 U22814 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19898), .B1(n19894), 
        .B2(n19885), .ZN(n19886) );
  OAI21_X1 U22815 ( .B1(n19887), .B2(n19897), .A(n19886), .ZN(P1_U2963) );
  AOI22_X1 U22816 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n19898), .B1(n19894), 
        .B2(n19888), .ZN(n19889) );
  OAI21_X1 U22817 ( .B1(n20786), .B2(n19897), .A(n19889), .ZN(P1_U2964) );
  AOI22_X1 U22818 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19898), .B1(n19894), 
        .B2(n19890), .ZN(n19891) );
  OAI21_X1 U22819 ( .B1(n19892), .B2(n19897), .A(n19891), .ZN(P1_U2965) );
  AOI22_X1 U22820 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19895), .B1(n19894), 
        .B2(n19893), .ZN(n19896) );
  OAI21_X1 U22821 ( .B1(n14600), .B2(n19897), .A(n19896), .ZN(P1_U2966) );
  AOI22_X1 U22822 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n19899), .B1(
        P1_LWORD_REG_15__SCAN_IN), .B2(n19898), .ZN(n19900) );
  OAI21_X1 U22823 ( .B1(n19902), .B2(n19901), .A(n19900), .ZN(P1_U2967) );
  AOI22_X1 U22824 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19910) );
  OR2_X1 U22825 ( .A1(n19904), .A2(n19903), .ZN(n19905) );
  NAND2_X1 U22826 ( .A1(n19906), .A2(n19905), .ZN(n19926) );
  INV_X1 U22827 ( .A(n19926), .ZN(n19908) );
  AOI22_X1 U22828 ( .A1(n19908), .A2(n19917), .B1(n15781), .B2(n19907), .ZN(
        n19909) );
  OAI211_X1 U22829 ( .C1(n19912), .C2(n19911), .A(n19910), .B(n19909), .ZN(
        P1_U2995) );
  AOI22_X1 U22830 ( .A1(n19914), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19913), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n19920) );
  INV_X1 U22831 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19915) );
  AOI22_X1 U22832 ( .A1(n19918), .A2(n19917), .B1(n19916), .B2(n19915), .ZN(
        n19919) );
  OAI211_X1 U22833 ( .C1(n19967), .C2(n19921), .A(n19920), .B(n19919), .ZN(
        P1_U2998) );
  NOR2_X1 U22834 ( .A1(n19946), .A2(n19922), .ZN(n19957) );
  NOR2_X1 U22835 ( .A1(n19957), .A2(n19923), .ZN(n19944) );
  AOI211_X1 U22836 ( .C1(n19933), .C2(n19943), .A(n19924), .B(n19938), .ZN(
        n19931) );
  NOR2_X1 U22837 ( .A1(n19926), .A2(n19925), .ZN(n19930) );
  OAI22_X1 U22838 ( .A1(n19955), .A2(n19928), .B1(n20597), .B2(n19927), .ZN(
        n19929) );
  NOR3_X1 U22839 ( .A1(n19931), .A2(n19930), .A3(n19929), .ZN(n19932) );
  OAI21_X1 U22840 ( .B1(n19944), .B2(n19933), .A(n19932), .ZN(P1_U3027) );
  AOI21_X1 U22841 ( .B1(n19936), .B2(n19935), .A(n19934), .ZN(n19942) );
  INV_X1 U22842 ( .A(n19937), .ZN(n19940) );
  INV_X1 U22843 ( .A(n19938), .ZN(n19939) );
  AOI22_X1 U22844 ( .A1(n19940), .A2(n19952), .B1(n19943), .B2(n19939), .ZN(
        n19941) );
  OAI211_X1 U22845 ( .C1(n19944), .C2(n19943), .A(n19942), .B(n19941), .ZN(
        P1_U3028) );
  NAND2_X1 U22846 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19945), .ZN(
        n19962) );
  NOR3_X1 U22847 ( .A1(n19947), .A2(n19951), .A3(n19946), .ZN(n19949) );
  AOI211_X1 U22848 ( .C1(n19951), .C2(n19950), .A(n19949), .B(n19948), .ZN(
        n19960) );
  AND3_X1 U22849 ( .A1(n12720), .A2(n19953), .A3(n19952), .ZN(n19958) );
  OAI22_X1 U22850 ( .A1(n19955), .A2(n19954), .B1(n12715), .B2(n19927), .ZN(
        n19956) );
  NOR3_X1 U22851 ( .A1(n19958), .A2(n19957), .A3(n19956), .ZN(n19959) );
  OAI221_X1 U22852 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19962), .C1(
        n19961), .C2(n19960), .A(n19959), .ZN(P1_U3029) );
  NOR2_X1 U22853 ( .A1(n19964), .A2(n19963), .ZN(P1_U3032) );
  NOR2_X2 U22854 ( .A1(n19967), .A2(n19966), .ZN(n20014) );
  AOI22_X1 U22855 ( .A1(DATAI_16_), .A2(n20013), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20014), .ZN(n20438) );
  NAND2_X1 U22856 ( .A1(n20053), .A2(n19970), .ZN(n20355) );
  AOI22_X2 U22857 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20014), .B1(DATAI_24_), 
        .B2(n20013), .ZN(n20522) );
  INV_X1 U22858 ( .A(n20522), .ZN(n20435) );
  NAND2_X1 U22859 ( .A1(n20016), .A2(n19972), .ZN(n20380) );
  NAND2_X1 U22860 ( .A1(n20058), .A2(n20256), .ZN(n20093) );
  OR2_X1 U22861 ( .A1(n20379), .A2(n20093), .ZN(n20017) );
  NOR2_X1 U22862 ( .A1(n20380), .A2(n20017), .ZN(n19973) );
  AOI21_X1 U22863 ( .B1(n20564), .B2(n20435), .A(n19973), .ZN(n19984) );
  OR2_X1 U22864 ( .A1(n20257), .A2(n20312), .ZN(n20136) );
  INV_X1 U22865 ( .A(n20136), .ZN(n19977) );
  NAND2_X1 U22866 ( .A1(n19980), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20473) );
  NAND2_X1 U22867 ( .A1(n20041), .A2(n20518), .ZN(n19974) );
  NAND2_X1 U22868 ( .A1(n20518), .A2(n20055), .ZN(n20382) );
  OAI21_X1 U22869 ( .B1(n19974), .B2(n20564), .A(n20382), .ZN(n19979) );
  OR2_X1 U22870 ( .A1(n20255), .A2(n19975), .ZN(n20057) );
  OR2_X1 U22871 ( .A1(n20057), .A2(n20471), .ZN(n19981) );
  AOI22_X1 U22872 ( .A1(n19979), .A2(n19981), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20017), .ZN(n19976) );
  OAI211_X1 U22873 ( .C1(n19977), .C2(n20573), .A(n20315), .B(n19976), .ZN(
        n20021) );
  NOR2_X2 U22874 ( .A1(n19978), .A2(n20140), .ZN(n20511) );
  INV_X1 U22875 ( .A(n19979), .ZN(n19982) );
  OR2_X1 U22876 ( .A1(n19980), .A2(n20573), .ZN(n20318) );
  AOI22_X1 U22877 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20021), .B1(
        n20511), .B2(n20020), .ZN(n19983) );
  OAI211_X1 U22878 ( .C1(n20438), .C2(n20041), .A(n19984), .B(n19983), .ZN(
        P1_U3033) );
  AOI22_X1 U22879 ( .A1(DATAI_17_), .A2(n20013), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20014), .ZN(n20442) );
  AOI22_X1 U22880 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20014), .B1(DATAI_25_), 
        .B2(n20013), .ZN(n20528) );
  INV_X1 U22881 ( .A(n20528), .ZN(n20439) );
  NAND2_X1 U22882 ( .A1(n20016), .A2(n19985), .ZN(n20394) );
  NOR2_X1 U22883 ( .A1(n20394), .A2(n20017), .ZN(n19986) );
  AOI21_X1 U22884 ( .B1(n20564), .B2(n20439), .A(n19986), .ZN(n19989) );
  NOR2_X2 U22885 ( .A1(n19987), .A2(n20140), .ZN(n20524) );
  AOI22_X1 U22886 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20021), .B1(
        n20524), .B2(n20020), .ZN(n19988) );
  OAI211_X1 U22887 ( .C1(n20442), .C2(n20041), .A(n19989), .B(n19988), .ZN(
        P1_U3034) );
  AOI22_X1 U22888 ( .A1(DATAI_18_), .A2(n20013), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20014), .ZN(n20446) );
  INV_X1 U22889 ( .A(n20534), .ZN(n20443) );
  NAND2_X1 U22890 ( .A1(n20016), .A2(n11974), .ZN(n20398) );
  NOR2_X1 U22891 ( .A1(n20398), .A2(n20017), .ZN(n19990) );
  AOI21_X1 U22892 ( .B1(n20564), .B2(n20443), .A(n19990), .ZN(n19993) );
  NOR2_X2 U22893 ( .A1(n19991), .A2(n20140), .ZN(n20530) );
  AOI22_X1 U22894 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20021), .B1(
        n20530), .B2(n20020), .ZN(n19992) );
  OAI211_X1 U22895 ( .C1(n20446), .C2(n20041), .A(n19993), .B(n19992), .ZN(
        P1_U3035) );
  AOI22_X1 U22896 ( .A1(DATAI_19_), .A2(n20013), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20014), .ZN(n20450) );
  AOI22_X1 U22897 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20014), .B1(DATAI_27_), 
        .B2(n20013), .ZN(n20540) );
  INV_X1 U22898 ( .A(n20540), .ZN(n20447) );
  NAND2_X1 U22899 ( .A1(n20016), .A2(n19994), .ZN(n20402) );
  NOR2_X1 U22900 ( .A1(n20402), .A2(n20017), .ZN(n19995) );
  AOI21_X1 U22901 ( .B1(n20564), .B2(n20447), .A(n19995), .ZN(n19998) );
  NOR2_X2 U22902 ( .A1(n19996), .A2(n20140), .ZN(n20536) );
  AOI22_X1 U22903 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20021), .B1(
        n20536), .B2(n20020), .ZN(n19997) );
  OAI211_X1 U22904 ( .C1(n20450), .C2(n20041), .A(n19998), .B(n19997), .ZN(
        P1_U3036) );
  AOI22_X1 U22905 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20014), .B1(DATAI_20_), 
        .B2(n20013), .ZN(n20454) );
  INV_X1 U22906 ( .A(n20546), .ZN(n20451) );
  NAND2_X1 U22907 ( .A1(n20016), .A2(n19999), .ZN(n20406) );
  NOR2_X1 U22908 ( .A1(n20406), .A2(n20017), .ZN(n20000) );
  AOI21_X1 U22909 ( .B1(n20564), .B2(n20451), .A(n20000), .ZN(n20004) );
  AOI22_X1 U22910 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20021), .B1(
        n20541), .B2(n20020), .ZN(n20003) );
  OAI211_X1 U22911 ( .C1(n20454), .C2(n20041), .A(n20004), .B(n20003), .ZN(
        P1_U3037) );
  AOI22_X1 U22912 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20014), .B1(DATAI_29_), 
        .B2(n20013), .ZN(n20552) );
  INV_X1 U22913 ( .A(n20552), .ZN(n20455) );
  NAND2_X1 U22914 ( .A1(n20016), .A2(n11767), .ZN(n20410) );
  NOR2_X1 U22915 ( .A1(n20410), .A2(n20017), .ZN(n20005) );
  AOI21_X1 U22916 ( .B1(n20564), .B2(n20455), .A(n20005), .ZN(n20008) );
  NOR2_X2 U22917 ( .A1(n20006), .A2(n20140), .ZN(n20548) );
  AOI22_X1 U22918 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20021), .B1(
        n20548), .B2(n20020), .ZN(n20007) );
  OAI211_X1 U22919 ( .C1(n20458), .C2(n20041), .A(n20008), .B(n20007), .ZN(
        P1_U3038) );
  AOI22_X1 U22920 ( .A1(DATAI_22_), .A2(n20013), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20014), .ZN(n20462) );
  AOI22_X1 U22921 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20014), .B1(DATAI_30_), 
        .B2(n20013), .ZN(n20558) );
  INV_X1 U22922 ( .A(n20558), .ZN(n20459) );
  NAND2_X1 U22923 ( .A1(n20016), .A2(n11655), .ZN(n20414) );
  NOR2_X1 U22924 ( .A1(n20414), .A2(n20017), .ZN(n20009) );
  AOI21_X1 U22925 ( .B1(n20564), .B2(n20459), .A(n20009), .ZN(n20012) );
  NOR2_X2 U22926 ( .A1(n20010), .A2(n20140), .ZN(n20554) );
  AOI22_X1 U22927 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20021), .B1(
        n20554), .B2(n20020), .ZN(n20011) );
  OAI211_X1 U22928 ( .C1(n20462), .C2(n20041), .A(n20012), .B(n20011), .ZN(
        P1_U3039) );
  AOI22_X1 U22929 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20014), .B1(DATAI_23_), 
        .B2(n20013), .ZN(n20470) );
  AOI22_X1 U22930 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20014), .B1(DATAI_31_), 
        .B2(n20013), .ZN(n20569) );
  INV_X1 U22931 ( .A(n20569), .ZN(n20465) );
  NAND2_X1 U22932 ( .A1(n20016), .A2(n20015), .ZN(n20419) );
  NOR2_X1 U22933 ( .A1(n20419), .A2(n20017), .ZN(n20018) );
  AOI21_X1 U22934 ( .B1(n20564), .B2(n20465), .A(n20018), .ZN(n20023) );
  NOR2_X2 U22935 ( .A1(n20019), .A2(n20140), .ZN(n20562) );
  AOI22_X1 U22936 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20021), .B1(
        n20562), .B2(n20020), .ZN(n20022) );
  OAI211_X1 U22937 ( .C1(n20470), .C2(n20041), .A(n20023), .B(n20022), .ZN(
        P1_U3040) );
  INV_X1 U22938 ( .A(n20057), .ZN(n20097) );
  INV_X1 U22939 ( .A(n20024), .ZN(n20429) );
  NOR3_X2 U22940 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20428), .A3(
        n20093), .ZN(n20046) );
  AOI21_X1 U22941 ( .B1(n20097), .B2(n20429), .A(n20046), .ZN(n20026) );
  NOR2_X1 U22942 ( .A1(n20093), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20029) );
  INV_X1 U22943 ( .A(n20029), .ZN(n20025) );
  OAI22_X1 U22944 ( .A1(n20026), .A2(n20509), .B1(n20025), .B2(n20573), .ZN(
        n20047) );
  AOI22_X1 U22945 ( .A1(n20511), .A2(n20047), .B1(n20510), .B2(n20046), .ZN(
        n20031) );
  INV_X1 U22946 ( .A(n20100), .ZN(n20027) );
  INV_X1 U22947 ( .A(n20382), .ZN(n20432) );
  OAI21_X1 U22948 ( .B1(n20027), .B2(n20432), .A(n20026), .ZN(n20028) );
  OAI211_X1 U22949 ( .C1(n20518), .C2(n20029), .A(n20516), .B(n20028), .ZN(
        n20049) );
  INV_X1 U22950 ( .A(n20084), .ZN(n20038) );
  INV_X1 U22951 ( .A(n20438), .ZN(n20519) );
  AOI22_X1 U22952 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20049), .B1(
        n20038), .B2(n20519), .ZN(n20030) );
  OAI211_X1 U22953 ( .C1(n20522), .C2(n20041), .A(n20031), .B(n20030), .ZN(
        P1_U3041) );
  AOI22_X1 U22954 ( .A1(n20524), .A2(n20047), .B1(n20523), .B2(n20046), .ZN(
        n20033) );
  INV_X1 U22955 ( .A(n20041), .ZN(n20048) );
  AOI22_X1 U22956 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20049), .B1(
        n20048), .B2(n20439), .ZN(n20032) );
  OAI211_X1 U22957 ( .C1(n20442), .C2(n20084), .A(n20033), .B(n20032), .ZN(
        P1_U3042) );
  AOI22_X1 U22958 ( .A1(n20530), .A2(n20047), .B1(n20529), .B2(n20046), .ZN(
        n20035) );
  INV_X1 U22959 ( .A(n20446), .ZN(n20531) );
  AOI22_X1 U22960 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20049), .B1(
        n20038), .B2(n20531), .ZN(n20034) );
  OAI211_X1 U22961 ( .C1(n20534), .C2(n20041), .A(n20035), .B(n20034), .ZN(
        P1_U3043) );
  AOI22_X1 U22962 ( .A1(n20536), .A2(n20047), .B1(n20535), .B2(n20046), .ZN(
        n20037) );
  AOI22_X1 U22963 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20049), .B1(
        n20048), .B2(n20447), .ZN(n20036) );
  OAI211_X1 U22964 ( .C1(n20450), .C2(n20084), .A(n20037), .B(n20036), .ZN(
        P1_U3044) );
  AOI22_X1 U22965 ( .A1(n20542), .A2(n20046), .B1(n20047), .B2(n20541), .ZN(
        n20040) );
  INV_X1 U22966 ( .A(n20454), .ZN(n20543) );
  AOI22_X1 U22967 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20049), .B1(
        n20038), .B2(n20543), .ZN(n20039) );
  OAI211_X1 U22968 ( .C1(n20546), .C2(n20041), .A(n20040), .B(n20039), .ZN(
        P1_U3045) );
  AOI22_X1 U22969 ( .A1(n20548), .A2(n20047), .B1(n20547), .B2(n20046), .ZN(
        n20043) );
  AOI22_X1 U22970 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20049), .B1(
        n20048), .B2(n20455), .ZN(n20042) );
  OAI211_X1 U22971 ( .C1(n20458), .C2(n20084), .A(n20043), .B(n20042), .ZN(
        P1_U3046) );
  AOI22_X1 U22972 ( .A1(n20554), .A2(n20047), .B1(n20553), .B2(n20046), .ZN(
        n20045) );
  AOI22_X1 U22973 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20049), .B1(
        n20048), .B2(n20459), .ZN(n20044) );
  OAI211_X1 U22974 ( .C1(n20462), .C2(n20084), .A(n20045), .B(n20044), .ZN(
        P1_U3047) );
  AOI22_X1 U22975 ( .A1(n20562), .A2(n20047), .B1(n20560), .B2(n20046), .ZN(
        n20051) );
  AOI22_X1 U22976 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20049), .B1(
        n20048), .B2(n20465), .ZN(n20050) );
  OAI211_X1 U22977 ( .C1(n20470), .C2(n20084), .A(n20051), .B(n20050), .ZN(
        P1_U3048) );
  OR3_X1 U22978 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20507), .A3(
        n20093), .ZN(n20083) );
  OAI22_X1 U22979 ( .A1(n20084), .A2(n20522), .B1(n20380), .B2(n20083), .ZN(
        n20054) );
  INV_X1 U22980 ( .A(n20054), .ZN(n20064) );
  AOI21_X1 U22981 ( .B1(n20128), .B2(n20084), .A(n20055), .ZN(n20056) );
  NOR2_X1 U22982 ( .A1(n20056), .A2(n20509), .ZN(n20060) );
  OR2_X1 U22983 ( .A1(n20057), .A2(n12955), .ZN(n20061) );
  AOI22_X1 U22984 ( .A1(n20060), .A2(n20061), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20083), .ZN(n20059) );
  NAND2_X1 U22985 ( .A1(n20312), .A2(n20058), .ZN(n20194) );
  NAND2_X1 U22986 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20194), .ZN(n20191) );
  NAND3_X1 U22987 ( .A1(n20315), .A2(n20059), .A3(n20191), .ZN(n20087) );
  INV_X1 U22988 ( .A(n20060), .ZN(n20062) );
  AOI22_X1 U22989 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20087), .B1(
        n20511), .B2(n20086), .ZN(n20063) );
  OAI211_X1 U22990 ( .C1(n20438), .C2(n20128), .A(n20064), .B(n20063), .ZN(
        P1_U3049) );
  OAI22_X1 U22991 ( .A1(n20128), .A2(n20442), .B1(n20394), .B2(n20083), .ZN(
        n20065) );
  INV_X1 U22992 ( .A(n20065), .ZN(n20067) );
  AOI22_X1 U22993 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20087), .B1(
        n20524), .B2(n20086), .ZN(n20066) );
  OAI211_X1 U22994 ( .C1(n20528), .C2(n20084), .A(n20067), .B(n20066), .ZN(
        P1_U3050) );
  OAI22_X1 U22995 ( .A1(n20128), .A2(n20446), .B1(n20398), .B2(n20083), .ZN(
        n20068) );
  INV_X1 U22996 ( .A(n20068), .ZN(n20070) );
  AOI22_X1 U22997 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20087), .B1(
        n20530), .B2(n20086), .ZN(n20069) );
  OAI211_X1 U22998 ( .C1(n20534), .C2(n20084), .A(n20070), .B(n20069), .ZN(
        P1_U3051) );
  OAI22_X1 U22999 ( .A1(n20084), .A2(n20540), .B1(n20402), .B2(n20083), .ZN(
        n20071) );
  INV_X1 U23000 ( .A(n20071), .ZN(n20073) );
  AOI22_X1 U23001 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20087), .B1(
        n20536), .B2(n20086), .ZN(n20072) );
  OAI211_X1 U23002 ( .C1(n20450), .C2(n20128), .A(n20073), .B(n20072), .ZN(
        P1_U3052) );
  OAI22_X1 U23003 ( .A1(n20084), .A2(n20546), .B1(n20406), .B2(n20083), .ZN(
        n20074) );
  INV_X1 U23004 ( .A(n20074), .ZN(n20076) );
  AOI22_X1 U23005 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20087), .B1(
        n20541), .B2(n20086), .ZN(n20075) );
  OAI211_X1 U23006 ( .C1(n20454), .C2(n20128), .A(n20076), .B(n20075), .ZN(
        P1_U3053) );
  OAI22_X1 U23007 ( .A1(n20128), .A2(n20458), .B1(n20410), .B2(n20083), .ZN(
        n20077) );
  INV_X1 U23008 ( .A(n20077), .ZN(n20079) );
  AOI22_X1 U23009 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20087), .B1(
        n20548), .B2(n20086), .ZN(n20078) );
  OAI211_X1 U23010 ( .C1(n20552), .C2(n20084), .A(n20079), .B(n20078), .ZN(
        P1_U3054) );
  OAI22_X1 U23011 ( .A1(n20128), .A2(n20462), .B1(n20414), .B2(n20083), .ZN(
        n20080) );
  INV_X1 U23012 ( .A(n20080), .ZN(n20082) );
  AOI22_X1 U23013 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20087), .B1(
        n20554), .B2(n20086), .ZN(n20081) );
  OAI211_X1 U23014 ( .C1(n20558), .C2(n20084), .A(n20082), .B(n20081), .ZN(
        P1_U3055) );
  OAI22_X1 U23015 ( .A1(n20084), .A2(n20569), .B1(n20419), .B2(n20083), .ZN(
        n20085) );
  INV_X1 U23016 ( .A(n20085), .ZN(n20089) );
  AOI22_X1 U23017 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20087), .B1(
        n20562), .B2(n20086), .ZN(n20088) );
  OAI211_X1 U23018 ( .C1(n20470), .C2(n20128), .A(n20089), .B(n20088), .ZN(
        P1_U3056) );
  INV_X1 U23019 ( .A(n20093), .ZN(n20090) );
  NAND2_X1 U23020 ( .A1(n20091), .A2(n20090), .ZN(n20127) );
  OAI22_X1 U23021 ( .A1(n20128), .A2(n20522), .B1(n20380), .B2(n20127), .ZN(
        n20092) );
  INV_X1 U23022 ( .A(n20092), .ZN(n20108) );
  NOR2_X1 U23023 ( .A1(n20507), .A2(n20093), .ZN(n20103) );
  INV_X1 U23024 ( .A(n20094), .ZN(n20095) );
  AND2_X1 U23025 ( .A1(n12253), .A2(n20095), .ZN(n20504) );
  INV_X1 U23026 ( .A(n20127), .ZN(n20096) );
  AOI21_X1 U23027 ( .B1(n20097), .B2(n20504), .A(n20096), .ZN(n20105) );
  INV_X1 U23028 ( .A(n20098), .ZN(n20099) );
  AOI21_X1 U23029 ( .B1(n20100), .B2(n20099), .A(n20509), .ZN(n20102) );
  NAND2_X1 U23030 ( .A1(n20105), .A2(n20102), .ZN(n20101) );
  OAI211_X1 U23031 ( .C1(n20518), .C2(n20103), .A(n20516), .B(n20101), .ZN(
        n20131) );
  INV_X1 U23032 ( .A(n20102), .ZN(n20106) );
  INV_X1 U23033 ( .A(n20103), .ZN(n20104) );
  OAI22_X1 U23034 ( .A1(n20106), .A2(n20105), .B1(n20573), .B2(n20104), .ZN(
        n20130) );
  AOI22_X1 U23035 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20131), .B1(
        n20511), .B2(n20130), .ZN(n20107) );
  OAI211_X1 U23036 ( .C1(n20438), .C2(n20137), .A(n20108), .B(n20107), .ZN(
        P1_U3057) );
  OAI22_X1 U23037 ( .A1(n20128), .A2(n20528), .B1(n20394), .B2(n20127), .ZN(
        n20109) );
  INV_X1 U23038 ( .A(n20109), .ZN(n20111) );
  AOI22_X1 U23039 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20131), .B1(
        n20524), .B2(n20130), .ZN(n20110) );
  OAI211_X1 U23040 ( .C1(n20442), .C2(n20137), .A(n20111), .B(n20110), .ZN(
        P1_U3058) );
  OAI22_X1 U23041 ( .A1(n20128), .A2(n20534), .B1(n20398), .B2(n20127), .ZN(
        n20112) );
  INV_X1 U23042 ( .A(n20112), .ZN(n20114) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20131), .B1(
        n20530), .B2(n20130), .ZN(n20113) );
  OAI211_X1 U23044 ( .C1(n20446), .C2(n20137), .A(n20114), .B(n20113), .ZN(
        P1_U3059) );
  OAI22_X1 U23045 ( .A1(n20128), .A2(n20540), .B1(n20402), .B2(n20127), .ZN(
        n20115) );
  INV_X1 U23046 ( .A(n20115), .ZN(n20117) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20131), .B1(
        n20536), .B2(n20130), .ZN(n20116) );
  OAI211_X1 U23048 ( .C1(n20450), .C2(n20137), .A(n20117), .B(n20116), .ZN(
        P1_U3060) );
  OAI22_X1 U23049 ( .A1(n20128), .A2(n20546), .B1(n20406), .B2(n20127), .ZN(
        n20118) );
  INV_X1 U23050 ( .A(n20118), .ZN(n20120) );
  AOI22_X1 U23051 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20131), .B1(
        n20541), .B2(n20130), .ZN(n20119) );
  OAI211_X1 U23052 ( .C1(n20454), .C2(n20137), .A(n20120), .B(n20119), .ZN(
        P1_U3061) );
  OAI22_X1 U23053 ( .A1(n20128), .A2(n20552), .B1(n20410), .B2(n20127), .ZN(
        n20121) );
  INV_X1 U23054 ( .A(n20121), .ZN(n20123) );
  AOI22_X1 U23055 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20131), .B1(
        n20548), .B2(n20130), .ZN(n20122) );
  OAI211_X1 U23056 ( .C1(n20458), .C2(n20137), .A(n20123), .B(n20122), .ZN(
        P1_U3062) );
  OAI22_X1 U23057 ( .A1(n20128), .A2(n20558), .B1(n20414), .B2(n20127), .ZN(
        n20124) );
  INV_X1 U23058 ( .A(n20124), .ZN(n20126) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20131), .B1(
        n20554), .B2(n20130), .ZN(n20125) );
  OAI211_X1 U23060 ( .C1(n20462), .C2(n20137), .A(n20126), .B(n20125), .ZN(
        P1_U3063) );
  OAI22_X1 U23061 ( .A1(n20128), .A2(n20569), .B1(n20419), .B2(n20127), .ZN(
        n20129) );
  INV_X1 U23062 ( .A(n20129), .ZN(n20133) );
  AOI22_X1 U23063 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20131), .B1(
        n20562), .B2(n20130), .ZN(n20132) );
  OAI211_X1 U23064 ( .C1(n20470), .C2(n20137), .A(n20133), .B(n20132), .ZN(
        P1_U3064) );
  OR2_X1 U23065 ( .A1(n12770), .A2(n20134), .ZN(n20190) );
  NAND3_X1 U23066 ( .A1(n20225), .A2(n20518), .A3(n12955), .ZN(n20135) );
  OAI21_X1 U23067 ( .B1(n20136), .B2(n20473), .A(n20135), .ZN(n20157) );
  AOI22_X1 U23068 ( .A1(n20511), .A2(n20157), .B1(n20510), .B2(n10092), .ZN(
        n20144) );
  INV_X1 U23069 ( .A(n20186), .ZN(n20138) );
  OAI21_X1 U23070 ( .B1(n20158), .B2(n20138), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20139) );
  OAI21_X1 U23071 ( .B1(n20471), .B2(n20190), .A(n20139), .ZN(n20142) );
  INV_X1 U23072 ( .A(n20318), .ZN(n20141) );
  AOI22_X1 U23073 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20159), .B1(
        n20158), .B2(n20435), .ZN(n20143) );
  OAI211_X1 U23074 ( .C1(n20438), .C2(n20186), .A(n20144), .B(n20143), .ZN(
        P1_U3065) );
  AOI22_X1 U23075 ( .A1(n20524), .A2(n20157), .B1(n20523), .B2(n10092), .ZN(
        n20146) );
  AOI22_X1 U23076 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20159), .B1(
        n20158), .B2(n20439), .ZN(n20145) );
  OAI211_X1 U23077 ( .C1(n20442), .C2(n20186), .A(n20146), .B(n20145), .ZN(
        P1_U3066) );
  AOI22_X1 U23078 ( .A1(n20530), .A2(n20157), .B1(n20529), .B2(n10092), .ZN(
        n20148) );
  AOI22_X1 U23079 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20159), .B1(
        n20158), .B2(n20443), .ZN(n20147) );
  OAI211_X1 U23080 ( .C1(n20446), .C2(n20186), .A(n20148), .B(n20147), .ZN(
        P1_U3067) );
  AOI22_X1 U23081 ( .A1(n20536), .A2(n20157), .B1(n20535), .B2(n10092), .ZN(
        n20150) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20159), .B1(
        n20158), .B2(n20447), .ZN(n20149) );
  OAI211_X1 U23083 ( .C1(n20450), .C2(n20186), .A(n20150), .B(n20149), .ZN(
        P1_U3068) );
  AOI22_X1 U23084 ( .A1(n20542), .A2(n10092), .B1(n20541), .B2(n20157), .ZN(
        n20152) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20159), .B1(
        n20158), .B2(n20451), .ZN(n20151) );
  OAI211_X1 U23086 ( .C1(n20454), .C2(n20186), .A(n20152), .B(n20151), .ZN(
        P1_U3069) );
  AOI22_X1 U23087 ( .A1(n20548), .A2(n20157), .B1(n20547), .B2(n10092), .ZN(
        n20154) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20159), .B1(
        n20158), .B2(n20455), .ZN(n20153) );
  OAI211_X1 U23089 ( .C1(n20458), .C2(n20186), .A(n20154), .B(n20153), .ZN(
        P1_U3070) );
  AOI22_X1 U23090 ( .A1(n20554), .A2(n20157), .B1(n20553), .B2(n10092), .ZN(
        n20156) );
  AOI22_X1 U23091 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20159), .B1(
        n20158), .B2(n20459), .ZN(n20155) );
  OAI211_X1 U23092 ( .C1(n20462), .C2(n20186), .A(n20156), .B(n20155), .ZN(
        P1_U3071) );
  AOI22_X1 U23093 ( .A1(n20562), .A2(n20157), .B1(n20560), .B2(n10092), .ZN(
        n20161) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20159), .B1(
        n20158), .B2(n20465), .ZN(n20160) );
  OAI211_X1 U23095 ( .C1(n20470), .C2(n20186), .A(n20161), .B(n20160), .ZN(
        P1_U3072) );
  NOR2_X1 U23096 ( .A1(n20187), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20165) );
  INV_X1 U23097 ( .A(n20165), .ZN(n20162) );
  NOR2_X1 U23098 ( .A1(n20428), .A2(n20162), .ZN(n20180) );
  AOI21_X1 U23099 ( .B1(n20225), .B2(n20429), .A(n20180), .ZN(n20163) );
  OAI22_X1 U23100 ( .A1(n20163), .A2(n20509), .B1(n20162), .B2(n20573), .ZN(
        n20181) );
  AOI22_X1 U23101 ( .A1(n20511), .A2(n20181), .B1(n20510), .B2(n20180), .ZN(
        n20167) );
  NOR2_X1 U23102 ( .A1(n20232), .A2(n20509), .ZN(n20228) );
  OAI21_X1 U23103 ( .B1(n20228), .B2(n20432), .A(n20163), .ZN(n20164) );
  OAI211_X1 U23104 ( .C1(n20518), .C2(n20165), .A(n20516), .B(n20164), .ZN(
        n20183) );
  AOI22_X1 U23105 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20519), .ZN(n20166) );
  OAI211_X1 U23106 ( .C1(n20522), .C2(n20186), .A(n20167), .B(n20166), .ZN(
        P1_U3073) );
  AOI22_X1 U23107 ( .A1(n20524), .A2(n20181), .B1(n20523), .B2(n20180), .ZN(
        n20169) );
  INV_X1 U23108 ( .A(n20442), .ZN(n20525) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20525), .ZN(n20168) );
  OAI211_X1 U23110 ( .C1(n20528), .C2(n20186), .A(n20169), .B(n20168), .ZN(
        P1_U3074) );
  AOI22_X1 U23111 ( .A1(n20530), .A2(n20181), .B1(n20529), .B2(n20180), .ZN(
        n20171) );
  AOI22_X1 U23112 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20531), .ZN(n20170) );
  OAI211_X1 U23113 ( .C1(n20534), .C2(n20186), .A(n20171), .B(n20170), .ZN(
        P1_U3075) );
  AOI22_X1 U23114 ( .A1(n20536), .A2(n20181), .B1(n20535), .B2(n20180), .ZN(
        n20173) );
  INV_X1 U23115 ( .A(n20450), .ZN(n20537) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20537), .ZN(n20172) );
  OAI211_X1 U23117 ( .C1(n20540), .C2(n20186), .A(n20173), .B(n20172), .ZN(
        P1_U3076) );
  AOI22_X1 U23118 ( .A1(n20542), .A2(n20180), .B1(n20541), .B2(n20181), .ZN(
        n20175) );
  AOI22_X1 U23119 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20543), .ZN(n20174) );
  OAI211_X1 U23120 ( .C1(n20546), .C2(n20186), .A(n20175), .B(n20174), .ZN(
        P1_U3077) );
  AOI22_X1 U23121 ( .A1(n20548), .A2(n20181), .B1(n20547), .B2(n20180), .ZN(
        n20177) );
  INV_X1 U23122 ( .A(n20458), .ZN(n20549) );
  AOI22_X1 U23123 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20549), .ZN(n20176) );
  OAI211_X1 U23124 ( .C1(n20552), .C2(n20186), .A(n20177), .B(n20176), .ZN(
        P1_U3078) );
  AOI22_X1 U23125 ( .A1(n20554), .A2(n20181), .B1(n20553), .B2(n20180), .ZN(
        n20179) );
  INV_X1 U23126 ( .A(n20462), .ZN(n20555) );
  AOI22_X1 U23127 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20555), .ZN(n20178) );
  OAI211_X1 U23128 ( .C1(n20558), .C2(n20186), .A(n20179), .B(n20178), .ZN(
        P1_U3079) );
  AOI22_X1 U23129 ( .A1(n20562), .A2(n20181), .B1(n20560), .B2(n20180), .ZN(
        n20185) );
  INV_X1 U23130 ( .A(n20470), .ZN(n20563) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20183), .B1(
        n20182), .B2(n20563), .ZN(n20184) );
  OAI211_X1 U23132 ( .C1(n20569), .C2(n20186), .A(n20185), .B(n20184), .ZN(
        P1_U3080) );
  NOR2_X1 U23133 ( .A1(n20507), .A2(n20187), .ZN(n20230) );
  INV_X1 U23134 ( .A(n20230), .ZN(n20226) );
  OR2_X1 U23135 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20226), .ZN(
        n20217) );
  OAI22_X1 U23136 ( .A1(n20243), .A2(n20438), .B1(n20380), .B2(n20217), .ZN(
        n20188) );
  INV_X1 U23137 ( .A(n20188), .ZN(n20198) );
  NAND3_X1 U23138 ( .A1(n20243), .A2(n20218), .A3(n20518), .ZN(n20189) );
  NAND2_X1 U23139 ( .A1(n20189), .A2(n20382), .ZN(n20193) );
  OR2_X1 U23140 ( .A1(n20190), .A2(n12955), .ZN(n20195) );
  AOI22_X1 U23141 ( .A1(n20193), .A2(n20195), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20217), .ZN(n20192) );
  NAND3_X1 U23142 ( .A1(n20480), .A2(n20192), .A3(n20191), .ZN(n20221) );
  INV_X1 U23143 ( .A(n20193), .ZN(n20196) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20221), .B1(
        n20511), .B2(n20220), .ZN(n20197) );
  OAI211_X1 U23145 ( .C1(n20522), .C2(n20218), .A(n20198), .B(n20197), .ZN(
        P1_U3081) );
  OAI22_X1 U23146 ( .A1(n20218), .A2(n20528), .B1(n20394), .B2(n20217), .ZN(
        n20199) );
  INV_X1 U23147 ( .A(n20199), .ZN(n20201) );
  AOI22_X1 U23148 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20221), .B1(
        n20524), .B2(n20220), .ZN(n20200) );
  OAI211_X1 U23149 ( .C1(n20442), .C2(n20243), .A(n20201), .B(n20200), .ZN(
        P1_U3082) );
  OAI22_X1 U23150 ( .A1(n20218), .A2(n20534), .B1(n20398), .B2(n20217), .ZN(
        n20202) );
  INV_X1 U23151 ( .A(n20202), .ZN(n20204) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20221), .B1(
        n20530), .B2(n20220), .ZN(n20203) );
  OAI211_X1 U23153 ( .C1(n20446), .C2(n20243), .A(n20204), .B(n20203), .ZN(
        P1_U3083) );
  OAI22_X1 U23154 ( .A1(n20218), .A2(n20540), .B1(n20402), .B2(n20217), .ZN(
        n20205) );
  INV_X1 U23155 ( .A(n20205), .ZN(n20207) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20221), .B1(
        n20536), .B2(n20220), .ZN(n20206) );
  OAI211_X1 U23157 ( .C1(n20450), .C2(n20243), .A(n20207), .B(n20206), .ZN(
        P1_U3084) );
  OAI22_X1 U23158 ( .A1(n20218), .A2(n20546), .B1(n20406), .B2(n20217), .ZN(
        n20208) );
  INV_X1 U23159 ( .A(n20208), .ZN(n20210) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20221), .B1(
        n20541), .B2(n20220), .ZN(n20209) );
  OAI211_X1 U23161 ( .C1(n20454), .C2(n20243), .A(n20210), .B(n20209), .ZN(
        P1_U3085) );
  OAI22_X1 U23162 ( .A1(n20243), .A2(n20458), .B1(n20410), .B2(n20217), .ZN(
        n20211) );
  INV_X1 U23163 ( .A(n20211), .ZN(n20213) );
  AOI22_X1 U23164 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20221), .B1(
        n20548), .B2(n20220), .ZN(n20212) );
  OAI211_X1 U23165 ( .C1(n20552), .C2(n20218), .A(n20213), .B(n20212), .ZN(
        P1_U3086) );
  OAI22_X1 U23166 ( .A1(n20218), .A2(n20558), .B1(n20414), .B2(n20217), .ZN(
        n20214) );
  INV_X1 U23167 ( .A(n20214), .ZN(n20216) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20221), .B1(
        n20554), .B2(n20220), .ZN(n20215) );
  OAI211_X1 U23169 ( .C1(n20462), .C2(n20243), .A(n20216), .B(n20215), .ZN(
        P1_U3087) );
  OAI22_X1 U23170 ( .A1(n20218), .A2(n20569), .B1(n20419), .B2(n20217), .ZN(
        n20219) );
  INV_X1 U23171 ( .A(n20219), .ZN(n20223) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20221), .B1(
        n20562), .B2(n20220), .ZN(n20222) );
  OAI211_X1 U23173 ( .C1(n20470), .C2(n20243), .A(n20223), .B(n20222), .ZN(
        P1_U3088) );
  INV_X1 U23174 ( .A(n20224), .ZN(n20248) );
  AOI21_X1 U23175 ( .B1(n20225), .B2(n20504), .A(n20248), .ZN(n20227) );
  OAI22_X1 U23176 ( .A1(n20227), .A2(n20509), .B1(n20226), .B2(n20573), .ZN(
        n20249) );
  AOI22_X1 U23177 ( .A1(n20511), .A2(n20249), .B1(n20248), .B2(n20510), .ZN(
        n20234) );
  OAI21_X1 U23178 ( .B1(n20514), .B2(n20228), .A(n20227), .ZN(n20229) );
  OAI211_X1 U23179 ( .C1(n20518), .C2(n20230), .A(n20516), .B(n20229), .ZN(
        n20251) );
  NAND2_X1 U23180 ( .A1(n20232), .A2(n20231), .ZN(n20254) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20251), .B1(
        n20278), .B2(n20519), .ZN(n20233) );
  OAI211_X1 U23182 ( .C1(n20522), .C2(n20243), .A(n20234), .B(n20233), .ZN(
        P1_U3089) );
  AOI22_X1 U23183 ( .A1(n20524), .A2(n20249), .B1(n20248), .B2(n20523), .ZN(
        n20236) );
  INV_X1 U23184 ( .A(n20243), .ZN(n20250) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20251), .B1(
        n20250), .B2(n20439), .ZN(n20235) );
  OAI211_X1 U23186 ( .C1(n20442), .C2(n20254), .A(n20236), .B(n20235), .ZN(
        P1_U3090) );
  AOI22_X1 U23187 ( .A1(n20530), .A2(n20249), .B1(n20248), .B2(n20529), .ZN(
        n20238) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20251), .B1(
        n20278), .B2(n20531), .ZN(n20237) );
  OAI211_X1 U23189 ( .C1(n20534), .C2(n20243), .A(n20238), .B(n20237), .ZN(
        P1_U3091) );
  AOI22_X1 U23190 ( .A1(n20536), .A2(n20249), .B1(n20248), .B2(n20535), .ZN(
        n20240) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20251), .B1(
        n20278), .B2(n20537), .ZN(n20239) );
  OAI211_X1 U23192 ( .C1(n20540), .C2(n20243), .A(n20240), .B(n20239), .ZN(
        P1_U3092) );
  AOI22_X1 U23193 ( .A1(n20542), .A2(n20248), .B1(n20541), .B2(n20249), .ZN(
        n20242) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20251), .B1(
        n20278), .B2(n20543), .ZN(n20241) );
  OAI211_X1 U23195 ( .C1(n20546), .C2(n20243), .A(n20242), .B(n20241), .ZN(
        P1_U3093) );
  AOI22_X1 U23196 ( .A1(n20548), .A2(n20249), .B1(n20248), .B2(n20547), .ZN(
        n20245) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20251), .B1(
        n20250), .B2(n20455), .ZN(n20244) );
  OAI211_X1 U23198 ( .C1(n20458), .C2(n20254), .A(n20245), .B(n20244), .ZN(
        P1_U3094) );
  AOI22_X1 U23199 ( .A1(n20554), .A2(n20249), .B1(n20248), .B2(n20553), .ZN(
        n20247) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20251), .B1(
        n20250), .B2(n20459), .ZN(n20246) );
  OAI211_X1 U23201 ( .C1(n20462), .C2(n20254), .A(n20247), .B(n20246), .ZN(
        P1_U3095) );
  AOI22_X1 U23202 ( .A1(n20562), .A2(n20249), .B1(n20248), .B2(n20560), .ZN(
        n20253) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20251), .B1(
        n20250), .B2(n20465), .ZN(n20252) );
  OAI211_X1 U23204 ( .C1(n20470), .C2(n20254), .A(n20253), .B(n20252), .ZN(
        P1_U3096) );
  AND2_X1 U23205 ( .A1(n20255), .A2(n12770), .ZN(n20349) );
  NAND2_X1 U23206 ( .A1(n20256), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20348) );
  AOI21_X1 U23207 ( .B1(n20349), .B2(n12955), .A(n10078), .ZN(n20260) );
  INV_X1 U23208 ( .A(n20312), .ZN(n20258) );
  NAND2_X1 U23209 ( .A1(n20258), .A2(n20257), .ZN(n20389) );
  OAI22_X1 U23210 ( .A1(n20260), .A2(n20509), .B1(n20318), .B2(n20389), .ZN(
        n20277) );
  AOI22_X1 U23211 ( .A1(n20511), .A2(n20277), .B1(n10078), .B2(n20510), .ZN(
        n20264) );
  INV_X1 U23212 ( .A(n20307), .ZN(n20259) );
  OAI21_X1 U23213 ( .B1(n20259), .B2(n20278), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20261) );
  NAND2_X1 U23214 ( .A1(n20261), .A2(n20260), .ZN(n20262) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20435), .ZN(n20263) );
  OAI211_X1 U23216 ( .C1(n20438), .C2(n20307), .A(n20264), .B(n20263), .ZN(
        P1_U3097) );
  AOI22_X1 U23217 ( .A1(n20524), .A2(n20277), .B1(n10078), .B2(n20523), .ZN(
        n20266) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20439), .ZN(n20265) );
  OAI211_X1 U23219 ( .C1(n20442), .C2(n20307), .A(n20266), .B(n20265), .ZN(
        P1_U3098) );
  AOI22_X1 U23220 ( .A1(n20530), .A2(n20277), .B1(n10078), .B2(n20529), .ZN(
        n20268) );
  AOI22_X1 U23221 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20443), .ZN(n20267) );
  OAI211_X1 U23222 ( .C1(n20446), .C2(n20307), .A(n20268), .B(n20267), .ZN(
        P1_U3099) );
  AOI22_X1 U23223 ( .A1(n20536), .A2(n20277), .B1(n10078), .B2(n20535), .ZN(
        n20270) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20447), .ZN(n20269) );
  OAI211_X1 U23225 ( .C1(n20450), .C2(n20307), .A(n20270), .B(n20269), .ZN(
        P1_U3100) );
  AOI22_X1 U23226 ( .A1(n20542), .A2(n10078), .B1(n20277), .B2(n20541), .ZN(
        n20272) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20451), .ZN(n20271) );
  OAI211_X1 U23228 ( .C1(n20454), .C2(n20307), .A(n20272), .B(n20271), .ZN(
        P1_U3101) );
  AOI22_X1 U23229 ( .A1(n20548), .A2(n20277), .B1(n10078), .B2(n20547), .ZN(
        n20274) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20455), .ZN(n20273) );
  OAI211_X1 U23231 ( .C1(n20458), .C2(n20307), .A(n20274), .B(n20273), .ZN(
        P1_U3102) );
  AOI22_X1 U23232 ( .A1(n20554), .A2(n20277), .B1(n10078), .B2(n20553), .ZN(
        n20276) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20459), .ZN(n20275) );
  OAI211_X1 U23234 ( .C1(n20462), .C2(n20307), .A(n20276), .B(n20275), .ZN(
        P1_U3103) );
  AOI22_X1 U23235 ( .A1(n20562), .A2(n20277), .B1(n10078), .B2(n20560), .ZN(
        n20281) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20465), .ZN(n20280) );
  OAI211_X1 U23237 ( .C1(n20470), .C2(n20307), .A(n20281), .B(n20280), .ZN(
        P1_U3104) );
  NOR2_X1 U23238 ( .A1(n20348), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20286) );
  INV_X1 U23239 ( .A(n20286), .ZN(n20282) );
  NOR2_X1 U23240 ( .A1(n20428), .A2(n20282), .ZN(n20302) );
  AOI21_X1 U23241 ( .B1(n20349), .B2(n20429), .A(n20302), .ZN(n20284) );
  OAI22_X1 U23242 ( .A1(n20284), .A2(n20509), .B1(n20282), .B2(n20573), .ZN(
        n20303) );
  AOI22_X1 U23243 ( .A1(n20511), .A2(n20303), .B1(n20510), .B2(n20302), .ZN(
        n20289) );
  NOR2_X1 U23244 ( .A1(n20283), .A2(n20509), .ZN(n20352) );
  OAI21_X1 U23245 ( .B1(n20352), .B2(n20432), .A(n20284), .ZN(n20285) );
  OAI211_X1 U23246 ( .C1(n20518), .C2(n20286), .A(n20516), .B(n20285), .ZN(
        n20304) );
  AOI22_X1 U23247 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20304), .B1(
        n20310), .B2(n20519), .ZN(n20288) );
  OAI211_X1 U23248 ( .C1(n20522), .C2(n20307), .A(n20289), .B(n20288), .ZN(
        P1_U3105) );
  AOI22_X1 U23249 ( .A1(n20524), .A2(n20303), .B1(n20523), .B2(n20302), .ZN(
        n20291) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20304), .B1(
        n20310), .B2(n20525), .ZN(n20290) );
  OAI211_X1 U23251 ( .C1(n20528), .C2(n20307), .A(n20291), .B(n20290), .ZN(
        P1_U3106) );
  AOI22_X1 U23252 ( .A1(n20530), .A2(n20303), .B1(n20529), .B2(n20302), .ZN(
        n20293) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20304), .B1(
        n20310), .B2(n20531), .ZN(n20292) );
  OAI211_X1 U23254 ( .C1(n20534), .C2(n20307), .A(n20293), .B(n20292), .ZN(
        P1_U3107) );
  AOI22_X1 U23255 ( .A1(n20536), .A2(n20303), .B1(n20535), .B2(n20302), .ZN(
        n20295) );
  AOI22_X1 U23256 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20304), .B1(
        n20310), .B2(n20537), .ZN(n20294) );
  OAI211_X1 U23257 ( .C1(n20540), .C2(n20307), .A(n20295), .B(n20294), .ZN(
        P1_U3108) );
  AOI22_X1 U23258 ( .A1(n20542), .A2(n20302), .B1(n20303), .B2(n20541), .ZN(
        n20297) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20304), .B1(
        n20310), .B2(n20543), .ZN(n20296) );
  OAI211_X1 U23260 ( .C1(n20546), .C2(n20307), .A(n20297), .B(n20296), .ZN(
        P1_U3109) );
  AOI22_X1 U23261 ( .A1(n20548), .A2(n20303), .B1(n20547), .B2(n20302), .ZN(
        n20299) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20304), .B1(
        n20310), .B2(n20549), .ZN(n20298) );
  OAI211_X1 U23263 ( .C1(n20552), .C2(n20307), .A(n20299), .B(n20298), .ZN(
        P1_U3110) );
  AOI22_X1 U23264 ( .A1(n20554), .A2(n20303), .B1(n20553), .B2(n20302), .ZN(
        n20301) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20304), .B1(
        n20310), .B2(n20555), .ZN(n20300) );
  OAI211_X1 U23266 ( .C1(n20558), .C2(n20307), .A(n20301), .B(n20300), .ZN(
        P1_U3111) );
  AOI22_X1 U23267 ( .A1(n20562), .A2(n20303), .B1(n20560), .B2(n20302), .ZN(
        n20306) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20304), .B1(
        n20310), .B2(n20563), .ZN(n20305) );
  OAI211_X1 U23269 ( .C1(n20569), .C2(n20307), .A(n20306), .B(n20305), .ZN(
        P1_U3112) );
  INV_X1 U23270 ( .A(n20474), .ZN(n20308) );
  NOR2_X1 U23271 ( .A1(n20507), .A2(n20348), .ZN(n20354) );
  INV_X1 U23272 ( .A(n20354), .ZN(n20350) );
  NOR2_X1 U23273 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20350), .ZN(
        n20313) );
  INV_X1 U23274 ( .A(n20313), .ZN(n20341) );
  OAI22_X1 U23275 ( .A1(n20342), .A2(n20522), .B1(n20380), .B2(n20341), .ZN(
        n20309) );
  INV_X1 U23276 ( .A(n20309), .ZN(n20322) );
  OAI21_X1 U23277 ( .B1(n20367), .B2(n20310), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20311) );
  NAND2_X1 U23278 ( .A1(n20311), .A2(n20518), .ZN(n20320) );
  AND2_X1 U23279 ( .A1(n20349), .A2(n20471), .ZN(n20317) );
  NAND2_X1 U23280 ( .A1(n20312), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20472) );
  NAND2_X1 U23281 ( .A1(n20472), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20479) );
  OAI21_X1 U23282 ( .B1(n20386), .B2(n20313), .A(n20479), .ZN(n20314) );
  INV_X1 U23283 ( .A(n20314), .ZN(n20316) );
  INV_X1 U23284 ( .A(n20317), .ZN(n20319) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20345), .B1(
        n20511), .B2(n20344), .ZN(n20321) );
  OAI211_X1 U23286 ( .C1(n20438), .C2(n20378), .A(n20322), .B(n20321), .ZN(
        P1_U3113) );
  OAI22_X1 U23287 ( .A1(n20378), .A2(n20442), .B1(n20394), .B2(n20341), .ZN(
        n20323) );
  INV_X1 U23288 ( .A(n20323), .ZN(n20325) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20345), .B1(
        n20524), .B2(n20344), .ZN(n20324) );
  OAI211_X1 U23290 ( .C1(n20528), .C2(n20342), .A(n20325), .B(n20324), .ZN(
        P1_U3114) );
  OAI22_X1 U23291 ( .A1(n20378), .A2(n20446), .B1(n20398), .B2(n20341), .ZN(
        n20326) );
  INV_X1 U23292 ( .A(n20326), .ZN(n20328) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20345), .B1(
        n20530), .B2(n20344), .ZN(n20327) );
  OAI211_X1 U23294 ( .C1(n20534), .C2(n20342), .A(n20328), .B(n20327), .ZN(
        P1_U3115) );
  OAI22_X1 U23295 ( .A1(n20342), .A2(n20540), .B1(n20402), .B2(n20341), .ZN(
        n20329) );
  INV_X1 U23296 ( .A(n20329), .ZN(n20331) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20345), .B1(
        n20536), .B2(n20344), .ZN(n20330) );
  OAI211_X1 U23298 ( .C1(n20450), .C2(n20378), .A(n20331), .B(n20330), .ZN(
        P1_U3116) );
  OAI22_X1 U23299 ( .A1(n20342), .A2(n20546), .B1(n20406), .B2(n20341), .ZN(
        n20332) );
  INV_X1 U23300 ( .A(n20332), .ZN(n20334) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20345), .B1(
        n20541), .B2(n20344), .ZN(n20333) );
  OAI211_X1 U23302 ( .C1(n20454), .C2(n20378), .A(n20334), .B(n20333), .ZN(
        P1_U3117) );
  OAI22_X1 U23303 ( .A1(n20378), .A2(n20458), .B1(n20410), .B2(n20341), .ZN(
        n20335) );
  INV_X1 U23304 ( .A(n20335), .ZN(n20337) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20345), .B1(
        n20548), .B2(n20344), .ZN(n20336) );
  OAI211_X1 U23306 ( .C1(n20552), .C2(n20342), .A(n20337), .B(n20336), .ZN(
        P1_U3118) );
  OAI22_X1 U23307 ( .A1(n20378), .A2(n20462), .B1(n20414), .B2(n20341), .ZN(
        n20338) );
  INV_X1 U23308 ( .A(n20338), .ZN(n20340) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20345), .B1(
        n20554), .B2(n20344), .ZN(n20339) );
  OAI211_X1 U23310 ( .C1(n20558), .C2(n20342), .A(n20340), .B(n20339), .ZN(
        P1_U3119) );
  OAI22_X1 U23311 ( .A1(n20342), .A2(n20569), .B1(n20419), .B2(n20341), .ZN(
        n20343) );
  INV_X1 U23312 ( .A(n20343), .ZN(n20347) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20345), .B1(
        n20562), .B2(n20344), .ZN(n20346) );
  OAI211_X1 U23314 ( .C1(n20470), .C2(n20378), .A(n20347), .B(n20346), .ZN(
        P1_U3120) );
  NOR2_X1 U23315 ( .A1(n20503), .A2(n20348), .ZN(n20372) );
  AOI21_X1 U23316 ( .B1(n20349), .B2(n20504), .A(n20372), .ZN(n20351) );
  OAI22_X1 U23317 ( .A1(n20351), .A2(n20509), .B1(n20350), .B2(n20573), .ZN(
        n20373) );
  AOI22_X1 U23318 ( .A1(n20511), .A2(n20373), .B1(n20510), .B2(n20372), .ZN(
        n20358) );
  OAI21_X1 U23319 ( .B1(n20514), .B2(n20352), .A(n20351), .ZN(n20353) );
  OAI211_X1 U23320 ( .C1(n20518), .C2(n20354), .A(n20516), .B(n20353), .ZN(
        n20375) );
  INV_X1 U23321 ( .A(n20425), .ZN(n20374) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20519), .ZN(n20357) );
  OAI211_X1 U23323 ( .C1(n20522), .C2(n20378), .A(n20358), .B(n20357), .ZN(
        P1_U3121) );
  AOI22_X1 U23324 ( .A1(n20524), .A2(n20373), .B1(n20523), .B2(n20372), .ZN(
        n20360) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20525), .ZN(n20359) );
  OAI211_X1 U23326 ( .C1(n20528), .C2(n20378), .A(n20360), .B(n20359), .ZN(
        P1_U3122) );
  AOI22_X1 U23327 ( .A1(n20530), .A2(n20373), .B1(n20529), .B2(n20372), .ZN(
        n20362) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20375), .B1(
        n20367), .B2(n20443), .ZN(n20361) );
  OAI211_X1 U23329 ( .C1(n20446), .C2(n20425), .A(n20362), .B(n20361), .ZN(
        P1_U3123) );
  AOI22_X1 U23330 ( .A1(n20536), .A2(n20373), .B1(n20535), .B2(n20372), .ZN(
        n20364) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20375), .B1(
        n20367), .B2(n20447), .ZN(n20363) );
  OAI211_X1 U23332 ( .C1(n20450), .C2(n20425), .A(n20364), .B(n20363), .ZN(
        P1_U3124) );
  AOI22_X1 U23333 ( .A1(n20542), .A2(n20372), .B1(n20373), .B2(n20541), .ZN(
        n20366) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20375), .B1(
        n20367), .B2(n20451), .ZN(n20365) );
  OAI211_X1 U23335 ( .C1(n20454), .C2(n20425), .A(n20366), .B(n20365), .ZN(
        P1_U3125) );
  AOI22_X1 U23336 ( .A1(n20548), .A2(n20373), .B1(n20547), .B2(n20372), .ZN(
        n20369) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20375), .B1(
        n20367), .B2(n20455), .ZN(n20368) );
  OAI211_X1 U23338 ( .C1(n20458), .C2(n20425), .A(n20369), .B(n20368), .ZN(
        P1_U3126) );
  AOI22_X1 U23339 ( .A1(n20554), .A2(n20373), .B1(n20553), .B2(n20372), .ZN(
        n20371) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20555), .ZN(n20370) );
  OAI211_X1 U23341 ( .C1(n20558), .C2(n20378), .A(n20371), .B(n20370), .ZN(
        P1_U3127) );
  AOI22_X1 U23342 ( .A1(n20562), .A2(n20373), .B1(n20560), .B2(n20372), .ZN(
        n20377) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20375), .B1(
        n20374), .B2(n20563), .ZN(n20376) );
  OAI211_X1 U23344 ( .C1(n20569), .C2(n20378), .A(n20377), .B(n20376), .ZN(
        P1_U3128) );
  NAND2_X1 U23345 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20506) );
  OR2_X1 U23346 ( .A1(n20379), .A2(n20506), .ZN(n20418) );
  NOR2_X1 U23347 ( .A1(n20380), .A2(n20418), .ZN(n20381) );
  AOI21_X1 U23348 ( .B1(n20466), .B2(n20519), .A(n20381), .ZN(n20393) );
  INV_X1 U23349 ( .A(n20418), .ZN(n20387) );
  NAND2_X1 U23350 ( .A1(n20425), .A2(n20518), .ZN(n20383) );
  OAI21_X1 U23351 ( .B1(n20383), .B2(n20466), .A(n20382), .ZN(n20388) );
  OR2_X1 U23352 ( .A1(n12770), .A2(n20384), .ZN(n20427) );
  OR2_X1 U23353 ( .A1(n20427), .A2(n20471), .ZN(n20390) );
  AOI22_X1 U23354 ( .A1(n20388), .A2(n20390), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20389), .ZN(n20385) );
  OAI211_X1 U23355 ( .C1(n20387), .C2(n20386), .A(n20480), .B(n20385), .ZN(
        n20422) );
  INV_X1 U23356 ( .A(n20388), .ZN(n20391) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20422), .B1(
        n20511), .B2(n20421), .ZN(n20392) );
  OAI211_X1 U23358 ( .C1(n20522), .C2(n20425), .A(n20393), .B(n20392), .ZN(
        P1_U3129) );
  NOR2_X1 U23359 ( .A1(n20394), .A2(n20418), .ZN(n20395) );
  AOI21_X1 U23360 ( .B1(n20466), .B2(n20525), .A(n20395), .ZN(n20397) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20422), .B1(
        n20524), .B2(n20421), .ZN(n20396) );
  OAI211_X1 U23362 ( .C1(n20528), .C2(n20425), .A(n20397), .B(n20396), .ZN(
        P1_U3130) );
  NOR2_X1 U23363 ( .A1(n20398), .A2(n20418), .ZN(n20399) );
  AOI21_X1 U23364 ( .B1(n20466), .B2(n20531), .A(n20399), .ZN(n20401) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20422), .B1(
        n20530), .B2(n20421), .ZN(n20400) );
  OAI211_X1 U23366 ( .C1(n20534), .C2(n20425), .A(n20401), .B(n20400), .ZN(
        P1_U3131) );
  NOR2_X1 U23367 ( .A1(n20402), .A2(n20418), .ZN(n20403) );
  AOI21_X1 U23368 ( .B1(n20466), .B2(n20537), .A(n20403), .ZN(n20405) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20422), .B1(
        n20536), .B2(n20421), .ZN(n20404) );
  OAI211_X1 U23370 ( .C1(n20540), .C2(n20425), .A(n20405), .B(n20404), .ZN(
        P1_U3132) );
  NOR2_X1 U23371 ( .A1(n20406), .A2(n20418), .ZN(n20407) );
  AOI21_X1 U23372 ( .B1(n20466), .B2(n20543), .A(n20407), .ZN(n20409) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20422), .B1(
        n20541), .B2(n20421), .ZN(n20408) );
  OAI211_X1 U23374 ( .C1(n20546), .C2(n20425), .A(n20409), .B(n20408), .ZN(
        P1_U3133) );
  NOR2_X1 U23375 ( .A1(n20410), .A2(n20418), .ZN(n20411) );
  AOI21_X1 U23376 ( .B1(n20466), .B2(n20549), .A(n20411), .ZN(n20413) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20422), .B1(
        n20548), .B2(n20421), .ZN(n20412) );
  OAI211_X1 U23378 ( .C1(n20552), .C2(n20425), .A(n20413), .B(n20412), .ZN(
        P1_U3134) );
  NOR2_X1 U23379 ( .A1(n20414), .A2(n20418), .ZN(n20415) );
  AOI21_X1 U23380 ( .B1(n20466), .B2(n20555), .A(n20415), .ZN(n20417) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20422), .B1(
        n20554), .B2(n20421), .ZN(n20416) );
  OAI211_X1 U23382 ( .C1(n20558), .C2(n20425), .A(n20417), .B(n20416), .ZN(
        P1_U3135) );
  NOR2_X1 U23383 ( .A1(n20419), .A2(n20418), .ZN(n20420) );
  AOI21_X1 U23384 ( .B1(n20466), .B2(n20563), .A(n20420), .ZN(n20424) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20422), .B1(
        n20562), .B2(n20421), .ZN(n20423) );
  OAI211_X1 U23386 ( .C1(n20569), .C2(n20425), .A(n20424), .B(n20423), .ZN(
        P1_U3136) );
  NOR3_X2 U23387 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20428), .A3(
        n20506), .ZN(n20463) );
  AOI21_X1 U23388 ( .B1(n20505), .B2(n20429), .A(n20463), .ZN(n20431) );
  NOR2_X1 U23389 ( .A1(n20506), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20434) );
  INV_X1 U23390 ( .A(n20434), .ZN(n20430) );
  OAI22_X1 U23391 ( .A1(n20431), .A2(n20509), .B1(n20430), .B2(n20573), .ZN(
        n20464) );
  AOI22_X1 U23392 ( .A1(n20511), .A2(n20464), .B1(n20510), .B2(n20463), .ZN(
        n20437) );
  NOR2_X1 U23393 ( .A1(n20475), .A2(n20509), .ZN(n20513) );
  OAI21_X1 U23394 ( .B1(n20513), .B2(n20432), .A(n20431), .ZN(n20433) );
  OAI211_X1 U23395 ( .C1(n20518), .C2(n20434), .A(n20516), .B(n20433), .ZN(
        n20467) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20435), .ZN(n20436) );
  OAI211_X1 U23397 ( .C1(n20438), .C2(n20502), .A(n20437), .B(n20436), .ZN(
        P1_U3137) );
  AOI22_X1 U23398 ( .A1(n20524), .A2(n20464), .B1(n20523), .B2(n20463), .ZN(
        n20441) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20439), .ZN(n20440) );
  OAI211_X1 U23400 ( .C1(n20442), .C2(n20502), .A(n20441), .B(n20440), .ZN(
        P1_U3138) );
  AOI22_X1 U23401 ( .A1(n20530), .A2(n20464), .B1(n20529), .B2(n20463), .ZN(
        n20445) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20443), .ZN(n20444) );
  OAI211_X1 U23403 ( .C1(n20446), .C2(n20502), .A(n20445), .B(n20444), .ZN(
        P1_U3139) );
  AOI22_X1 U23404 ( .A1(n20536), .A2(n20464), .B1(n20535), .B2(n20463), .ZN(
        n20449) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20447), .ZN(n20448) );
  OAI211_X1 U23406 ( .C1(n20450), .C2(n20502), .A(n20449), .B(n20448), .ZN(
        P1_U3140) );
  AOI22_X1 U23407 ( .A1(n20542), .A2(n20463), .B1(n20541), .B2(n20464), .ZN(
        n20453) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20451), .ZN(n20452) );
  OAI211_X1 U23409 ( .C1(n20454), .C2(n20502), .A(n20453), .B(n20452), .ZN(
        P1_U3141) );
  AOI22_X1 U23410 ( .A1(n20548), .A2(n20464), .B1(n20547), .B2(n20463), .ZN(
        n20457) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20455), .ZN(n20456) );
  OAI211_X1 U23412 ( .C1(n20458), .C2(n20502), .A(n20457), .B(n20456), .ZN(
        P1_U3142) );
  AOI22_X1 U23413 ( .A1(n20554), .A2(n20464), .B1(n20553), .B2(n20463), .ZN(
        n20461) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20459), .ZN(n20460) );
  OAI211_X1 U23415 ( .C1(n20462), .C2(n20502), .A(n20461), .B(n20460), .ZN(
        P1_U3143) );
  AOI22_X1 U23416 ( .A1(n20562), .A2(n20464), .B1(n20560), .B2(n20463), .ZN(
        n20469) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20467), .B1(
        n20466), .B2(n20465), .ZN(n20468) );
  OAI211_X1 U23418 ( .C1(n20470), .C2(n20502), .A(n20469), .B(n20468), .ZN(
        P1_U3144) );
  NAND2_X1 U23419 ( .A1(n20505), .A2(n20471), .ZN(n20477) );
  OAI22_X1 U23420 ( .A1(n20477), .A2(n20509), .B1(n20473), .B2(n20472), .ZN(
        n20497) );
  NOR3_X2 U23421 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20507), .A3(
        n20506), .ZN(n20496) );
  AOI22_X1 U23422 ( .A1(n20511), .A2(n20497), .B1(n20510), .B2(n20496), .ZN(
        n20483) );
  INV_X1 U23423 ( .A(n20502), .ZN(n20476) );
  OAI21_X1 U23424 ( .B1(n20498), .B2(n20476), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20478) );
  AOI21_X1 U23425 ( .B1(n20478), .B2(n20477), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20481) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20499), .B1(
        n20498), .B2(n20519), .ZN(n20482) );
  OAI211_X1 U23427 ( .C1(n20522), .C2(n20502), .A(n20483), .B(n20482), .ZN(
        P1_U3145) );
  AOI22_X1 U23428 ( .A1(n20524), .A2(n20497), .B1(n20523), .B2(n20496), .ZN(
        n20485) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20499), .B1(
        n20498), .B2(n20525), .ZN(n20484) );
  OAI211_X1 U23430 ( .C1(n20528), .C2(n20502), .A(n20485), .B(n20484), .ZN(
        P1_U3146) );
  AOI22_X1 U23431 ( .A1(n20530), .A2(n20497), .B1(n20529), .B2(n20496), .ZN(
        n20487) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20499), .B1(
        n20498), .B2(n20531), .ZN(n20486) );
  OAI211_X1 U23433 ( .C1(n20534), .C2(n20502), .A(n20487), .B(n20486), .ZN(
        P1_U3147) );
  AOI22_X1 U23434 ( .A1(n20536), .A2(n20497), .B1(n20535), .B2(n20496), .ZN(
        n20489) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20499), .B1(
        n20498), .B2(n20537), .ZN(n20488) );
  OAI211_X1 U23436 ( .C1(n20540), .C2(n20502), .A(n20489), .B(n20488), .ZN(
        P1_U3148) );
  AOI22_X1 U23437 ( .A1(n20542), .A2(n20496), .B1(n20541), .B2(n20497), .ZN(
        n20491) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20499), .B1(
        n20498), .B2(n20543), .ZN(n20490) );
  OAI211_X1 U23439 ( .C1(n20546), .C2(n20502), .A(n20491), .B(n20490), .ZN(
        P1_U3149) );
  AOI22_X1 U23440 ( .A1(n20548), .A2(n20497), .B1(n20547), .B2(n20496), .ZN(
        n20493) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20499), .B1(
        n20498), .B2(n20549), .ZN(n20492) );
  OAI211_X1 U23442 ( .C1(n20552), .C2(n20502), .A(n20493), .B(n20492), .ZN(
        P1_U3150) );
  AOI22_X1 U23443 ( .A1(n20554), .A2(n20497), .B1(n20553), .B2(n20496), .ZN(
        n20495) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20499), .B1(
        n20498), .B2(n20555), .ZN(n20494) );
  OAI211_X1 U23445 ( .C1(n20558), .C2(n20502), .A(n20495), .B(n20494), .ZN(
        P1_U3151) );
  AOI22_X1 U23446 ( .A1(n20562), .A2(n20497), .B1(n20560), .B2(n20496), .ZN(
        n20501) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20499), .B1(
        n20498), .B2(n20563), .ZN(n20500) );
  OAI211_X1 U23448 ( .C1(n20569), .C2(n20502), .A(n20501), .B(n20500), .ZN(
        P1_U3152) );
  NOR2_X1 U23449 ( .A1(n20503), .A2(n20506), .ZN(n20559) );
  AOI21_X1 U23450 ( .B1(n20505), .B2(n20504), .A(n20559), .ZN(n20512) );
  NOR2_X1 U23451 ( .A1(n20507), .A2(n20506), .ZN(n20517) );
  INV_X1 U23452 ( .A(n20517), .ZN(n20508) );
  OAI22_X1 U23453 ( .A1(n20512), .A2(n20509), .B1(n20508), .B2(n20573), .ZN(
        n20561) );
  AOI22_X1 U23454 ( .A1(n20511), .A2(n20561), .B1(n20510), .B2(n20559), .ZN(
        n20521) );
  OAI21_X1 U23455 ( .B1(n20514), .B2(n20513), .A(n20512), .ZN(n20515) );
  OAI211_X1 U23456 ( .C1(n20518), .C2(n20517), .A(n20516), .B(n20515), .ZN(
        n20565) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20519), .ZN(n20520) );
  OAI211_X1 U23458 ( .C1(n20522), .C2(n20568), .A(n20521), .B(n20520), .ZN(
        P1_U3153) );
  AOI22_X1 U23459 ( .A1(n20524), .A2(n20561), .B1(n20523), .B2(n20559), .ZN(
        n20527) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20525), .ZN(n20526) );
  OAI211_X1 U23461 ( .C1(n20528), .C2(n20568), .A(n20527), .B(n20526), .ZN(
        P1_U3154) );
  AOI22_X1 U23462 ( .A1(n20530), .A2(n20561), .B1(n20529), .B2(n20559), .ZN(
        n20533) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20531), .ZN(n20532) );
  OAI211_X1 U23464 ( .C1(n20534), .C2(n20568), .A(n20533), .B(n20532), .ZN(
        P1_U3155) );
  AOI22_X1 U23465 ( .A1(n20536), .A2(n20561), .B1(n20535), .B2(n20559), .ZN(
        n20539) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20537), .ZN(n20538) );
  OAI211_X1 U23467 ( .C1(n20540), .C2(n20568), .A(n20539), .B(n20538), .ZN(
        P1_U3156) );
  AOI22_X1 U23468 ( .A1(n20542), .A2(n20559), .B1(n20541), .B2(n20561), .ZN(
        n20545) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20543), .ZN(n20544) );
  OAI211_X1 U23470 ( .C1(n20546), .C2(n20568), .A(n20545), .B(n20544), .ZN(
        P1_U3157) );
  AOI22_X1 U23471 ( .A1(n20548), .A2(n20561), .B1(n20547), .B2(n20559), .ZN(
        n20551) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20549), .ZN(n20550) );
  OAI211_X1 U23473 ( .C1(n20552), .C2(n20568), .A(n20551), .B(n20550), .ZN(
        P1_U3158) );
  AOI22_X1 U23474 ( .A1(n20554), .A2(n20561), .B1(n20553), .B2(n20559), .ZN(
        n20557) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20555), .ZN(n20556) );
  OAI211_X1 U23476 ( .C1(n20558), .C2(n20568), .A(n20557), .B(n20556), .ZN(
        P1_U3159) );
  AOI22_X1 U23477 ( .A1(n20562), .A2(n20561), .B1(n20560), .B2(n20559), .ZN(
        n20567) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20563), .ZN(n20566) );
  OAI211_X1 U23479 ( .C1(n20569), .C2(n20568), .A(n20567), .B(n20566), .ZN(
        P1_U3160) );
  NOR2_X1 U23480 ( .A1(n20571), .A2(n20570), .ZN(n20574) );
  OAI21_X1 U23481 ( .B1(n20574), .B2(n20573), .A(n20572), .ZN(P1_U3163) );
  AND2_X1 U23482 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20649), .ZN(
        P1_U3164) );
  AND2_X1 U23483 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20649), .ZN(
        P1_U3165) );
  AND2_X1 U23484 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20649), .ZN(
        P1_U3166) );
  AND2_X1 U23485 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20649), .ZN(
        P1_U3167) );
  AND2_X1 U23486 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20649), .ZN(
        P1_U3168) );
  AND2_X1 U23487 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20649), .ZN(
        P1_U3169) );
  AND2_X1 U23488 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20649), .ZN(
        P1_U3170) );
  AND2_X1 U23489 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20649), .ZN(
        P1_U3171) );
  AND2_X1 U23490 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20649), .ZN(
        P1_U3172) );
  AND2_X1 U23491 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20649), .ZN(
        P1_U3173) );
  AND2_X1 U23492 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20649), .ZN(
        P1_U3174) );
  AND2_X1 U23493 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20649), .ZN(
        P1_U3175) );
  AND2_X1 U23494 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20649), .ZN(
        P1_U3176) );
  AND2_X1 U23495 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20649), .ZN(
        P1_U3177) );
  AND2_X1 U23496 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20649), .ZN(
        P1_U3178) );
  AND2_X1 U23497 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20649), .ZN(
        P1_U3179) );
  AND2_X1 U23498 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20649), .ZN(
        P1_U3180) );
  AND2_X1 U23499 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20649), .ZN(
        P1_U3181) );
  AND2_X1 U23500 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20649), .ZN(
        P1_U3182) );
  AND2_X1 U23501 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20649), .ZN(
        P1_U3183) );
  INV_X1 U23502 ( .A(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20772) );
  NOR2_X1 U23503 ( .A1(n20653), .A2(n20772), .ZN(P1_U3184) );
  AND2_X1 U23504 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20649), .ZN(
        P1_U3185) );
  AND2_X1 U23505 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20649), .ZN(P1_U3186) );
  AND2_X1 U23506 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20649), .ZN(P1_U3187) );
  AND2_X1 U23507 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20649), .ZN(P1_U3188) );
  AND2_X1 U23508 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20649), .ZN(P1_U3189) );
  AND2_X1 U23509 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20649), .ZN(P1_U3190) );
  AND2_X1 U23510 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20649), .ZN(P1_U3191) );
  AND2_X1 U23511 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20649), .ZN(P1_U3192) );
  AND2_X1 U23512 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20649), .ZN(P1_U3193) );
  NAND2_X1 U23513 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20575), .ZN(n20586) );
  INV_X1 U23514 ( .A(n20586), .ZN(n20579) );
  INV_X2 U23515 ( .A(n20675), .ZN(n20663) );
  NAND2_X1 U23516 ( .A1(n20587), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20580) );
  AOI22_X1 U23517 ( .A1(HOLD), .A2(n20577), .B1(n20580), .B2(n20576), .ZN(
        n20578) );
  OAI22_X1 U23518 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20579), .B1(n20663), 
        .B2(n20578), .ZN(P1_U3194) );
  INV_X1 U23519 ( .A(n20580), .ZN(n20583) );
  AOI21_X1 U23520 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20592), .A(n20581), .ZN(n20582) );
  AOI21_X1 U23521 ( .B1(n20584), .B2(n20583), .A(n20582), .ZN(n20591) );
  NAND3_X1 U23522 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20585), .A3(n20587), 
        .ZN(n20589) );
  OAI211_X1 U23523 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20587), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20586), .ZN(n20588) );
  OAI221_X1 U23524 ( .B1(n20591), .B2(n20590), .C1(n20591), .C2(n20589), .A(
        n20588), .ZN(P1_U3196) );
  INV_X1 U23525 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20593) );
  NAND2_X1 U23526 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20663), .ZN(n20642) );
  OAI222_X1 U23527 ( .A1(n20639), .A2(n12715), .B1(n20593), .B2(n20663), .C1(
        n12892), .C2(n20642), .ZN(P1_U3197) );
  INV_X1 U23528 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20594) );
  OAI222_X1 U23529 ( .A1(n20642), .A2(n12715), .B1(n20594), .B2(n20663), .C1(
        n12905), .C2(n20639), .ZN(P1_U3198) );
  OAI222_X1 U23530 ( .A1(n20642), .A2(n12905), .B1(n20595), .B2(n20663), .C1(
        n20597), .C2(n20639), .ZN(P1_U3199) );
  INV_X1 U23531 ( .A(n20639), .ZN(n20630) );
  AOI22_X1 U23532 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20630), .ZN(n20596) );
  OAI21_X1 U23533 ( .B1(n20597), .B2(n20642), .A(n20596), .ZN(P1_U3200) );
  INV_X1 U23534 ( .A(n20642), .ZN(n20631) );
  AOI22_X1 U23535 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20631), .ZN(n20598) );
  OAI21_X1 U23536 ( .B1(n20600), .B2(n20639), .A(n20598), .ZN(P1_U3201) );
  INV_X1 U23537 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20599) );
  OAI222_X1 U23538 ( .A1(n20642), .A2(n20600), .B1(n20599), .B2(n20663), .C1(
        n20757), .C2(n20639), .ZN(P1_U3202) );
  INV_X1 U23539 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20601) );
  OAI222_X1 U23540 ( .A1(n20642), .A2(n20757), .B1(n20601), .B2(n20663), .C1(
        n20603), .C2(n20639), .ZN(P1_U3203) );
  INV_X1 U23541 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20602) );
  OAI222_X1 U23542 ( .A1(n20642), .A2(n20603), .B1(n20602), .B2(n20663), .C1(
        n20605), .C2(n20639), .ZN(P1_U3204) );
  INV_X1 U23543 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20604) );
  INV_X1 U23544 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20606) );
  OAI222_X1 U23545 ( .A1(n20642), .A2(n20605), .B1(n20604), .B2(n20663), .C1(
        n20606), .C2(n20639), .ZN(P1_U3205) );
  INV_X1 U23546 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20607) );
  OAI222_X1 U23547 ( .A1(n20639), .A2(n20609), .B1(n20607), .B2(n20663), .C1(
        n20606), .C2(n20642), .ZN(P1_U3206) );
  AOI22_X1 U23548 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20630), .ZN(n20608) );
  OAI21_X1 U23549 ( .B1(n20609), .B2(n20642), .A(n20608), .ZN(P1_U3207) );
  AOI22_X1 U23550 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20631), .ZN(n20610) );
  OAI21_X1 U23551 ( .B1(n14702), .B2(n20639), .A(n20610), .ZN(P1_U3208) );
  INV_X1 U23552 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20611) );
  OAI222_X1 U23553 ( .A1(n20642), .A2(n14702), .B1(n20611), .B2(n20663), .C1(
        n20612), .C2(n20639), .ZN(P1_U3209) );
  INV_X1 U23554 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20613) );
  OAI222_X1 U23555 ( .A1(n20639), .A2(n14689), .B1(n20613), .B2(n20663), .C1(
        n20612), .C2(n20642), .ZN(P1_U3210) );
  INV_X1 U23556 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20614) );
  OAI222_X1 U23557 ( .A1(n20642), .A2(n14689), .B1(n20614), .B2(n20663), .C1(
        n14817), .C2(n20639), .ZN(P1_U3211) );
  AOI22_X1 U23558 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20630), .ZN(n20615) );
  OAI21_X1 U23559 ( .B1(n14817), .B2(n20642), .A(n20615), .ZN(P1_U3212) );
  INV_X1 U23560 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20618) );
  AOI22_X1 U23561 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20631), .ZN(n20616) );
  OAI21_X1 U23562 ( .B1(n20618), .B2(n20639), .A(n20616), .ZN(P1_U3213) );
  AOI22_X1 U23563 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20630), .ZN(n20617) );
  OAI21_X1 U23564 ( .B1(n20618), .B2(n20642), .A(n20617), .ZN(P1_U3214) );
  AOI22_X1 U23565 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20631), .ZN(n20619) );
  OAI21_X1 U23566 ( .B1(n20621), .B2(n20639), .A(n20619), .ZN(P1_U3215) );
  INV_X1 U23567 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20620) );
  OAI222_X1 U23568 ( .A1(n20642), .A2(n20621), .B1(n20620), .B2(n20663), .C1(
        n20623), .C2(n20639), .ZN(P1_U3216) );
  INV_X1 U23569 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20622) );
  OAI222_X1 U23570 ( .A1(n20642), .A2(n20623), .B1(n20622), .B2(n20663), .C1(
        n20823), .C2(n20639), .ZN(P1_U3217) );
  INV_X1 U23571 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20624) );
  OAI222_X1 U23572 ( .A1(n20642), .A2(n20823), .B1(n20624), .B2(n20663), .C1(
        n20627), .C2(n20639), .ZN(P1_U3218) );
  INV_X1 U23573 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20626) );
  OAI222_X1 U23574 ( .A1(n20642), .A2(n20627), .B1(n20626), .B2(n20663), .C1(
        n20625), .C2(n20639), .ZN(P1_U3219) );
  AOI222_X1 U23575 ( .A1(n20631), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20630), .ZN(n20628) );
  INV_X1 U23576 ( .A(n20628), .ZN(P1_U3220) );
  AOI222_X1 U23577 ( .A1(n20631), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20630), .ZN(n20629) );
  INV_X1 U23578 ( .A(n20629), .ZN(P1_U3221) );
  AOI222_X1 U23579 ( .A1(n20631), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20630), .ZN(n20632) );
  INV_X1 U23580 ( .A(n20632), .ZN(P1_U3222) );
  INV_X1 U23581 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20633) );
  OAI222_X1 U23582 ( .A1(n20642), .A2(n20634), .B1(n20633), .B2(n20663), .C1(
        n20636), .C2(n20639), .ZN(P1_U3223) );
  INV_X1 U23583 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20635) );
  OAI222_X1 U23584 ( .A1(n20642), .A2(n20636), .B1(n20635), .B2(n20663), .C1(
        n20638), .C2(n20639), .ZN(P1_U3224) );
  INV_X1 U23585 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20637) );
  OAI222_X1 U23586 ( .A1(n20642), .A2(n20638), .B1(n20637), .B2(n20663), .C1(
        n20807), .C2(n20639), .ZN(P1_U3225) );
  INV_X1 U23587 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20641) );
  OAI222_X1 U23588 ( .A1(n20642), .A2(n20807), .B1(n20641), .B2(n20663), .C1(
        n20640), .C2(n20639), .ZN(P1_U3226) );
  INV_X1 U23589 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20643) );
  AOI22_X1 U23590 ( .A1(n20663), .A2(n20758), .B1(n20643), .B2(n20675), .ZN(
        P1_U3458) );
  INV_X1 U23591 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20655) );
  INV_X1 U23592 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20644) );
  AOI22_X1 U23593 ( .A1(n20663), .A2(n20655), .B1(n20644), .B2(n20675), .ZN(
        P1_U3459) );
  INV_X1 U23594 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20645) );
  AOI22_X1 U23595 ( .A1(n20663), .A2(n20646), .B1(n20645), .B2(n20675), .ZN(
        P1_U3460) );
  INV_X1 U23596 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20661) );
  INV_X1 U23597 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20647) );
  AOI22_X1 U23598 ( .A1(n20663), .A2(n20661), .B1(n20647), .B2(n20675), .ZN(
        P1_U3461) );
  INV_X1 U23599 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20650) );
  INV_X1 U23600 ( .A(n20651), .ZN(n20648) );
  AOI21_X1 U23601 ( .B1(n20650), .B2(n20649), .A(n20648), .ZN(P1_U3464) );
  OAI21_X1 U23602 ( .B1(n20653), .B2(n20652), .A(n20651), .ZN(P1_U3465) );
  AOI21_X1 U23603 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20654) );
  AOI22_X1 U23604 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20654), .B2(n12892), .ZN(n20656) );
  AOI22_X1 U23605 ( .A1(n20657), .A2(n20656), .B1(n20655), .B2(n20660), .ZN(
        P1_U3481) );
  NOR2_X1 U23606 ( .A1(n20660), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20658) );
  AOI22_X1 U23607 ( .A1(n20661), .A2(n20660), .B1(n20659), .B2(n20658), .ZN(
        P1_U3482) );
  AOI22_X1 U23608 ( .A1(n20663), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20662), 
        .B2(n20675), .ZN(P1_U3483) );
  AOI211_X1 U23609 ( .C1(n20667), .C2(n20666), .A(n20665), .B(n20664), .ZN(
        n20674) );
  OAI211_X1 U23610 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n9590), .A(n20668), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20671) );
  AOI21_X1 U23611 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20671), .A(n20670), 
        .ZN(n20673) );
  NAND2_X1 U23612 ( .A1(n20674), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20672) );
  OAI21_X1 U23613 ( .B1(n20674), .B2(n20673), .A(n20672), .ZN(P1_U3485) );
  INV_X1 U23614 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20738) );
  INV_X1 U23615 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20676) );
  AOI22_X1 U23616 ( .A1(n20663), .A2(n20738), .B1(n20676), .B2(n20675), .ZN(
        P1_U3486) );
  AOI22_X1 U23617 ( .A1(n20679), .A2(keyinput58), .B1(keyinput28), .B2(n20678), 
        .ZN(n20677) );
  OAI221_X1 U23618 ( .B1(n20679), .B2(keyinput58), .C1(n20678), .C2(keyinput28), .A(n20677), .ZN(n20691) );
  INV_X1 U23619 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20681) );
  AOI22_X1 U23620 ( .A1(n20682), .A2(keyinput59), .B1(n20681), .B2(keyinput27), 
        .ZN(n20680) );
  OAI221_X1 U23621 ( .B1(n20682), .B2(keyinput59), .C1(n20681), .C2(keyinput27), .A(n20680), .ZN(n20690) );
  AOI22_X1 U23622 ( .A1(n20685), .A2(keyinput43), .B1(n20684), .B2(keyinput35), 
        .ZN(n20683) );
  OAI221_X1 U23623 ( .B1(n20685), .B2(keyinput43), .C1(n20684), .C2(keyinput35), .A(n20683), .ZN(n20689) );
  AOI22_X1 U23624 ( .A1(n11050), .A2(keyinput16), .B1(keyinput44), .B2(n20687), 
        .ZN(n20686) );
  OAI221_X1 U23625 ( .B1(n11050), .B2(keyinput16), .C1(n20687), .C2(keyinput44), .A(n20686), .ZN(n20688) );
  NOR4_X1 U23626 ( .A1(n20691), .A2(n20690), .A3(n20689), .A4(n20688), .ZN(
        n20736) );
  AOI22_X1 U23627 ( .A1(n20694), .A2(keyinput36), .B1(n20693), .B2(keyinput31), 
        .ZN(n20692) );
  OAI221_X1 U23628 ( .B1(n20694), .B2(keyinput36), .C1(n20693), .C2(keyinput31), .A(n20692), .ZN(n20707) );
  AOI22_X1 U23629 ( .A1(n20697), .A2(keyinput1), .B1(n20696), .B2(keyinput63), 
        .ZN(n20695) );
  OAI221_X1 U23630 ( .B1(n20697), .B2(keyinput1), .C1(n20696), .C2(keyinput63), 
        .A(n20695), .ZN(n20706) );
  AOI22_X1 U23631 ( .A1(n20700), .A2(keyinput23), .B1(n20699), .B2(keyinput38), 
        .ZN(n20698) );
  OAI221_X1 U23632 ( .B1(n20700), .B2(keyinput23), .C1(n20699), .C2(keyinput38), .A(n20698), .ZN(n20705) );
  AOI22_X1 U23633 ( .A1(n20703), .A2(keyinput25), .B1(keyinput52), .B2(n20702), 
        .ZN(n20701) );
  OAI221_X1 U23634 ( .B1(n20703), .B2(keyinput25), .C1(n20702), .C2(keyinput52), .A(n20701), .ZN(n20704) );
  NOR4_X1 U23635 ( .A1(n20707), .A2(n20706), .A3(n20705), .A4(n20704), .ZN(
        n20735) );
  AOI22_X1 U23636 ( .A1(n20709), .A2(keyinput40), .B1(n14959), .B2(keyinput19), 
        .ZN(n20708) );
  OAI221_X1 U23637 ( .B1(n20709), .B2(keyinput40), .C1(n14959), .C2(keyinput19), .A(n20708), .ZN(n20719) );
  AOI22_X1 U23638 ( .A1(n20712), .A2(keyinput15), .B1(n20711), .B2(keyinput61), 
        .ZN(n20710) );
  OAI221_X1 U23639 ( .B1(n20712), .B2(keyinput15), .C1(n20711), .C2(keyinput61), .A(n20710), .ZN(n20718) );
  AOI22_X1 U23640 ( .A1(n14348), .A2(keyinput29), .B1(keyinput7), .B2(n20714), 
        .ZN(n20713) );
  OAI221_X1 U23641 ( .B1(n14348), .B2(keyinput29), .C1(n20714), .C2(keyinput7), 
        .A(n20713), .ZN(n20717) );
  INV_X1 U23642 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20816) );
  AOI22_X1 U23643 ( .A1(n20823), .A2(keyinput51), .B1(n20816), .B2(keyinput34), 
        .ZN(n20715) );
  OAI221_X1 U23644 ( .B1(n20823), .B2(keyinput51), .C1(n20816), .C2(keyinput34), .A(n20715), .ZN(n20716) );
  NOR4_X1 U23645 ( .A1(n20719), .A2(n20718), .A3(n20717), .A4(n20716), .ZN(
        n20734) );
  AOI22_X1 U23646 ( .A1(n20721), .A2(keyinput53), .B1(keyinput32), .B2(n20813), 
        .ZN(n20720) );
  OAI221_X1 U23647 ( .B1(n20721), .B2(keyinput53), .C1(n20813), .C2(keyinput32), .A(n20720), .ZN(n20725) );
  XOR2_X1 U23648 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B(keyinput13), .Z(
        n20724) );
  XNOR2_X1 U23649 ( .A(n20722), .B(keyinput54), .ZN(n20723) );
  OR3_X1 U23650 ( .A1(n20725), .A2(n20724), .A3(n20723), .ZN(n20732) );
  AOI22_X1 U23651 ( .A1(n20727), .A2(keyinput57), .B1(n20814), .B2(keyinput20), 
        .ZN(n20726) );
  OAI221_X1 U23652 ( .B1(n20727), .B2(keyinput57), .C1(n20814), .C2(keyinput20), .A(n20726), .ZN(n20731) );
  AOI22_X1 U23653 ( .A1(n20815), .A2(keyinput21), .B1(keyinput22), .B2(n20729), 
        .ZN(n20728) );
  OAI221_X1 U23654 ( .B1(n20815), .B2(keyinput21), .C1(n20729), .C2(keyinput22), .A(n20728), .ZN(n20730) );
  NOR3_X1 U23655 ( .A1(n20732), .A2(n20731), .A3(n20730), .ZN(n20733) );
  NAND4_X1 U23656 ( .A1(n20736), .A2(n20735), .A3(n20734), .A4(n20733), .ZN(
        n20799) );
  AOI22_X1 U23657 ( .A1(n20739), .A2(keyinput42), .B1(n20738), .B2(keyinput48), 
        .ZN(n20737) );
  OAI221_X1 U23658 ( .B1(n20739), .B2(keyinput42), .C1(n20738), .C2(keyinput48), .A(n20737), .ZN(n20752) );
  AOI22_X1 U23659 ( .A1(n20742), .A2(keyinput12), .B1(n20741), .B2(keyinput62), 
        .ZN(n20740) );
  OAI221_X1 U23660 ( .B1(n20742), .B2(keyinput12), .C1(n20741), .C2(keyinput62), .A(n20740), .ZN(n20751) );
  INV_X1 U23661 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n20745) );
  AOI22_X1 U23662 ( .A1(n20745), .A2(keyinput60), .B1(keyinput14), .B2(n20744), 
        .ZN(n20743) );
  OAI221_X1 U23663 ( .B1(n20745), .B2(keyinput60), .C1(n20744), .C2(keyinput14), .A(n20743), .ZN(n20750) );
  INV_X1 U23664 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n20747) );
  AOI22_X1 U23665 ( .A1(n20748), .A2(keyinput41), .B1(n20747), .B2(keyinput30), 
        .ZN(n20746) );
  OAI221_X1 U23666 ( .B1(n20748), .B2(keyinput41), .C1(n20747), .C2(keyinput30), .A(n20746), .ZN(n20749) );
  NOR4_X1 U23667 ( .A1(n20752), .A2(n20751), .A3(n20750), .A4(n20749), .ZN(
        n20797) );
  INV_X1 U23668 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n20755) );
  AOI22_X1 U23669 ( .A1(n20755), .A2(keyinput3), .B1(keyinput24), .B2(n20754), 
        .ZN(n20753) );
  OAI221_X1 U23670 ( .B1(n20755), .B2(keyinput3), .C1(n20754), .C2(keyinput24), 
        .A(n20753), .ZN(n20768) );
  AOI22_X1 U23671 ( .A1(n20758), .A2(keyinput47), .B1(n20757), .B2(keyinput26), 
        .ZN(n20756) );
  OAI221_X1 U23672 ( .B1(n20758), .B2(keyinput47), .C1(n20757), .C2(keyinput26), .A(n20756), .ZN(n20767) );
  AOI22_X1 U23673 ( .A1(n20761), .A2(keyinput18), .B1(keyinput4), .B2(n20760), 
        .ZN(n20759) );
  OAI221_X1 U23674 ( .B1(n20761), .B2(keyinput18), .C1(n20760), .C2(keyinput4), 
        .A(n20759), .ZN(n20766) );
  INV_X1 U23675 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n20763) );
  AOI22_X1 U23676 ( .A1(n20764), .A2(keyinput56), .B1(keyinput49), .B2(n20763), 
        .ZN(n20762) );
  OAI221_X1 U23677 ( .B1(n20764), .B2(keyinput56), .C1(n20763), .C2(keyinput49), .A(n20762), .ZN(n20765) );
  NOR4_X1 U23678 ( .A1(n20768), .A2(n20767), .A3(n20766), .A4(n20765), .ZN(
        n20796) );
  AOI22_X1 U23679 ( .A1(n14010), .A2(keyinput46), .B1(keyinput11), .B2(n20819), 
        .ZN(n20769) );
  OAI221_X1 U23680 ( .B1(n14010), .B2(keyinput46), .C1(n20819), .C2(keyinput11), .A(n20769), .ZN(n20778) );
  INV_X1 U23681 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n20771) );
  AOI22_X1 U23682 ( .A1(n20772), .A2(keyinput6), .B1(n20771), .B2(keyinput37), 
        .ZN(n20770) );
  OAI221_X1 U23683 ( .B1(n20772), .B2(keyinput6), .C1(n20771), .C2(keyinput37), 
        .A(n20770), .ZN(n20777) );
  AOI22_X1 U23684 ( .A1(n20808), .A2(keyinput33), .B1(keyinput50), .B2(n20807), 
        .ZN(n20773) );
  OAI221_X1 U23685 ( .B1(n20808), .B2(keyinput33), .C1(n20807), .C2(keyinput50), .A(n20773), .ZN(n20776) );
  AOI22_X1 U23686 ( .A1(n20809), .A2(keyinput17), .B1(n20810), .B2(keyinput8), 
        .ZN(n20774) );
  OAI221_X1 U23687 ( .B1(n20809), .B2(keyinput17), .C1(n20810), .C2(keyinput8), 
        .A(n20774), .ZN(n20775) );
  NOR4_X1 U23688 ( .A1(n20778), .A2(n20777), .A3(n20776), .A4(n20775), .ZN(
        n20795) );
  AOI22_X1 U23689 ( .A1(n20780), .A2(keyinput39), .B1(n20820), .B2(keyinput45), 
        .ZN(n20779) );
  OAI221_X1 U23690 ( .B1(n20780), .B2(keyinput39), .C1(n20820), .C2(keyinput45), .A(n20779), .ZN(n20793) );
  AOI22_X1 U23691 ( .A1(n20783), .A2(keyinput0), .B1(keyinput10), .B2(n20782), 
        .ZN(n20781) );
  OAI221_X1 U23692 ( .B1(n20783), .B2(keyinput0), .C1(n20782), .C2(keyinput10), 
        .A(n20781), .ZN(n20792) );
  AOI22_X1 U23693 ( .A1(n20786), .A2(keyinput5), .B1(keyinput55), .B2(n20785), 
        .ZN(n20784) );
  OAI221_X1 U23694 ( .B1(n20786), .B2(keyinput5), .C1(n20785), .C2(keyinput55), 
        .A(n20784), .ZN(n20791) );
  INV_X1 U23695 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20789) );
  AOI22_X1 U23696 ( .A1(n20789), .A2(keyinput9), .B1(n20788), .B2(keyinput2), 
        .ZN(n20787) );
  OAI221_X1 U23697 ( .B1(n20789), .B2(keyinput9), .C1(n20788), .C2(keyinput2), 
        .A(n20787), .ZN(n20790) );
  NOR4_X1 U23698 ( .A1(n20793), .A2(n20792), .A3(n20791), .A4(n20790), .ZN(
        n20794) );
  NAND4_X1 U23699 ( .A1(n20797), .A2(n20796), .A3(n20795), .A4(n20794), .ZN(
        n20798) );
  NOR2_X1 U23700 ( .A1(n20799), .A2(n20798), .ZN(n20839) );
  AOI22_X1 U23701 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20800), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17234), .ZN(n20801) );
  OAI21_X1 U23702 ( .B1(n20802), .B2(n17244), .A(n20801), .ZN(n20837) );
  NOR4_X1 U23703 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(P1_DATAO_REG_30__SCAN_IN), 
        .A3(P1_DATAO_REG_21__SCAN_IN), .A4(P1_DATAO_REG_11__SCAN_IN), .ZN(
        n20806) );
  NOR4_X1 U23704 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(P2_UWORD_REG_13__SCAN_IN), 
        .A4(P3_LWORD_REG_7__SCAN_IN), .ZN(n20805) );
  NOR4_X1 U23705 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_0__SCAN_IN), .A4(BUF2_REG_2__SCAN_IN), .ZN(n20804) );
  NOR4_X1 U23706 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_12__2__SCAN_IN), .A3(P1_EAX_REG_12__SCAN_IN), .A4(
        P2_DATAO_REG_28__SCAN_IN), .ZN(n20803) );
  NAND4_X1 U23707 ( .A1(n20806), .A2(n20805), .A3(n20804), .A4(n20803), .ZN(
        n20835) );
  NAND4_X1 U23708 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(DATAI_8_), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20834) );
  NOR4_X1 U23709 ( .A1(n20810), .A2(n20809), .A3(n20808), .A4(n20807), .ZN(
        n20811) );
  NAND3_X1 U23710 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20811), .A3(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20812) );
  NOR4_X1 U23711 ( .A1(n20814), .A2(n20813), .A3(n20812), .A4(n20712), .ZN(
        n20818) );
  NOR3_X1 U23712 ( .A1(n20816), .A2(n20815), .A3(n14959), .ZN(n20817) );
  NAND2_X1 U23713 ( .A1(n20818), .A2(n20817), .ZN(n20833) );
  NOR4_X1 U23714 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .A3(P3_M_IO_N_REG_SCAN_IN), .A4(
        P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20831) );
  NOR4_X1 U23715 ( .A1(P1_EAX_REG_3__SCAN_IN), .A2(P1_DATAO_REG_10__SCAN_IN), 
        .A3(P3_ADDRESS_REG_28__SCAN_IN), .A4(P1_BYTEENABLE_REG_3__SCAN_IN), 
        .ZN(n20830) );
  NAND4_X1 U23716 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_2__3__SCAN_IN), .A3(n20820), .A4(n20819), .ZN(n20821)
         );
  NOR4_X1 U23717 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_0__5__SCAN_IN), .A3(n20822), .A4(n20821), .ZN(n20829)
         );
  NAND4_X1 U23718 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_3__2__SCAN_IN), .A3(n14010), .A4(n20823), .ZN(n20827)
         );
  NAND4_X1 U23719 ( .A1(DATAI_11_), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .A3(P3_EBX_REG_3__SCAN_IN), .A4(P3_ADDRESS_REG_11__SCAN_IN), .ZN(
        n20826) );
  NAND4_X1 U23720 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_REIP_REG_7__SCAN_IN), .A3(DATAI_13_), .A4(P3_DATAO_REG_26__SCAN_IN), 
        .ZN(n20825) );
  NAND4_X1 U23721 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_REIP_REG_0__SCAN_IN), .A3(P1_MEMORYFETCH_REG_SCAN_IN), .A4(
        P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20824) );
  NOR4_X1 U23722 ( .A1(n20827), .A2(n20826), .A3(n20825), .A4(n20824), .ZN(
        n20828) );
  NAND4_X1 U23723 ( .A1(n20831), .A2(n20830), .A3(n20829), .A4(n20828), .ZN(
        n20832) );
  NOR4_X1 U23724 ( .A1(n20835), .A2(n20834), .A3(n20833), .A4(n20832), .ZN(
        n20836) );
  XNOR2_X1 U23725 ( .A(n20837), .B(n20836), .ZN(n20838) );
  XNOR2_X1 U23726 ( .A(n20839), .B(n20838), .ZN(P3_U2783) );
  NAND2_X1 U11084 ( .A1(n11778), .A2(n11777), .ZN(n12261) );
  CLKBUF_X1 U11041 ( .A(n13731), .Z(n13889) );
  CLKBUF_X1 U11042 ( .A(n11581), .Z(n13879) );
  CLKBUF_X1 U11043 ( .A(n11602), .Z(n13888) );
  NOR2_X1 U11049 ( .A1(n11666), .A2(n11679), .ZN(n11707) );
  CLKBUF_X1 U11074 ( .A(n10268), .Z(n13993) );
  CLKBUF_X1 U11076 ( .A(n10416), .Z(n13042) );
  INV_X1 U11083 ( .A(n19972), .ZN(n12926) );
  CLKBUF_X1 U11085 ( .A(n12025), .Z(n12114) );
  CLKBUF_X1 U11117 ( .A(n20669), .Z(n9590) );
  CLKBUF_X1 U11129 ( .A(n10756), .Z(n9566) );
  CLKBUF_X1 U11136 ( .A(n10417), .Z(n19123) );
  NAND2_X1 U11195 ( .A1(n12261), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11786) );
  CLKBUF_X3 U11369 ( .A(n10226), .Z(n19683) );
  CLKBUF_X1 U11406 ( .A(n17524), .Z(n9600) );
  CLKBUF_X1 U11678 ( .A(n16206), .Z(n9570) );
  CLKBUF_X1 U12213 ( .A(n17623), .Z(n9597) );
  CLKBUF_X1 U12286 ( .A(n16300), .Z(n16298) );
endmodule

