

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862;

  INV_X1 U2387 ( .A(n4492), .ZN(n4232) );
  CLKBUF_X2 U2388 ( .A(n3584), .Z(n2152) );
  INV_X1 U2389 ( .A(n2879), .ZN(n3594) );
  CLKBUF_X2 U2390 ( .A(n3597), .Z(n2154) );
  INV_X2 U2391 ( .A(n2153), .ZN(n2872) );
  CLKBUF_X2 U2392 ( .A(n2424), .Z(n3779) );
  NAND2_X1 U2393 ( .A1(n2865), .A2(n2983), .ZN(n2873) );
  INV_X1 U2394 ( .A(n2873), .ZN(n3584) );
  INV_X1 U2395 ( .A(n3585), .ZN(n2884) );
  CLKBUF_X3 U2396 ( .A(n2873), .Z(n3562) );
  AOI211_X1 U2399 ( .C1(n2195), .C2(n3951), .A(n2940), .B(n2939), .ZN(n2959)
         );
  INV_X1 U2400 ( .A(n2417), .ZN(n2145) );
  AND2_X1 U2401 ( .A1(n4355), .A2(n2387), .ZN(n2417) );
  NAND2_X2 U2402 ( .A1(n3650), .A2(n3580), .ZN(n3710) );
  INV_X2 U2403 ( .A(IR_REG_11__SCAN_IN), .ZN(n2518) );
  NAND2_X2 U2404 ( .A1(n3524), .A2(n3703), .ZN(n3656) );
  AOI22_X1 U2405 ( .A1(n3949), .A2(n3584), .B1(n2155), .B2(n2971), .ZN(n2883)
         );
  INV_X4 U2406 ( .A(n2145), .ZN(n2146) );
  AND2_X1 U2407 ( .A1(n2386), .A2(n2387), .ZN(n2416) );
  CLKBUF_X1 U2408 ( .A(n2873), .Z(n2149) );
  INV_X1 U2409 ( .A(n2879), .ZN(n2150) );
  NAND2_X4 U2410 ( .A1(n2155), .A2(n2871), .ZN(n2879) );
  BUF_X2 U2411 ( .A(n2726), .Z(n2151) );
  XNOR2_X1 U2412 ( .A(n2680), .B(IR_REG_21__SCAN_IN), .ZN(n2726) );
  NAND2_X1 U2413 ( .A1(n3080), .A2(n3079), .ZN(n3081) );
  NAND4_X1 U2414 ( .A1(n2442), .A2(n2441), .A3(n2440), .A4(n2439), .ZN(n3088)
         );
  AND3_X1 U2415 ( .A1(n2423), .A2(n2422), .A3(n2421), .ZN(n3009) );
  INV_X1 U2416 ( .A(IR_REG_16__SCAN_IN), .ZN(n4650) );
  CLKBUF_X2 U2417 ( .A(IR_REG_0__SCAN_IN), .Z(n4652) );
  INV_X2 U2418 ( .A(IR_REG_0__SCAN_IN), .ZN(n2195) );
  NAND2_X1 U2419 ( .A1(n3577), .A2(n3576), .ZN(n3711) );
  NAND2_X1 U2420 ( .A1(n3669), .A2(n3722), .ZN(n3721) );
  NOR2_X1 U2421 ( .A1(n4441), .A2(REG1_REG_16__SCAN_IN), .ZN(n4442) );
  NOR2_X1 U2422 ( .A1(n3689), .A2(n3508), .ZN(n3515) );
  NAND2_X1 U2423 ( .A1(n4386), .A2(n3161), .ZN(n4397) );
  NOR2_X2 U2424 ( .A1(n2926), .A2(n2927), .ZN(n2989) );
  AOI21_X1 U2425 ( .B1(n3157), .B2(REG1_REG_8__SCAN_IN), .A(n2270), .ZN(n3158)
         );
  NAND2_X1 U2426 ( .A1(n2283), .A2(n2192), .ZN(n2285) );
  NOR2_X1 U2427 ( .A1(n2271), .A2(n3174), .ZN(n2270) );
  XNOR2_X1 U2428 ( .A(n2271), .B(n2246), .ZN(n3157) );
  NAND2_X1 U2429 ( .A1(n2272), .A2(n2194), .ZN(n2271) );
  NAND2_X1 U2430 ( .A1(n2912), .A2(n2911), .ZN(n2272) );
  NOR2_X1 U2431 ( .A1(n2841), .A2(n2273), .ZN(n2912) );
  AND2_X2 U2432 ( .A1(n2969), .A2(n4114), .ZN(n4492) );
  NAND2_X2 U2433 ( .A1(n3814), .A2(n2716), .ZN(n4196) );
  AND2_X1 U2434 ( .A1(n2278), .A2(n2277), .ZN(n2276) );
  NAND4_X1 U2435 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .ZN(n2992)
         );
  NAND2_X1 U2436 ( .A1(n2953), .A2(n2281), .ZN(n2280) );
  AND4_X1 U2437 ( .A1(n2403), .A2(n2404), .A3(n2405), .A4(n2402), .ZN(n2973)
         );
  NAND4_X1 U2438 ( .A1(n2410), .A2(n2409), .A3(n2408), .A4(n2407), .ZN(n3949)
         );
  OR2_X1 U2439 ( .A1(n2726), .A2(n4360), .ZN(n4510) );
  NAND2_X1 U2440 ( .A1(n2413), .A2(n2412), .ZN(n2971) );
  NAND3_X1 U2441 ( .A1(n4358), .A2(n4359), .A3(n2772), .ZN(n2983) );
  NAND2_X1 U2442 ( .A1(n4366), .A2(REG1_REG_5__SCAN_IN), .ZN(n2277) );
  AND2_X1 U2443 ( .A1(n2585), .A2(n2584), .ZN(n2589) );
  AND2_X1 U2444 ( .A1(n2258), .A2(n2375), .ZN(n2731) );
  AND2_X1 U2445 ( .A1(n2544), .A2(n2372), .ZN(n2375) );
  AND2_X1 U2446 ( .A1(n2359), .A2(n2395), .ZN(n2358) );
  AND2_X1 U2447 ( .A1(n2320), .A2(n2374), .ZN(n2472) );
  AND2_X1 U2448 ( .A1(n2540), .A2(n2369), .ZN(n2544) );
  AND2_X1 U2449 ( .A1(n2360), .A2(n2171), .ZN(n2359) );
  NOR2_X1 U2450 ( .A1(n2368), .A2(IR_REG_9__SCAN_IN), .ZN(n2540) );
  AND2_X1 U2451 ( .A1(n2373), .A2(n2321), .ZN(n2320) );
  NAND3_X1 U2452 ( .A1(n2195), .A2(n2196), .A3(n2247), .ZN(n2431) );
  AND2_X1 U2453 ( .A1(n2376), .A2(n2361), .ZN(n2360) );
  AND2_X1 U2454 ( .A1(n2539), .A2(n4657), .ZN(n2369) );
  AND2_X1 U2455 ( .A1(n2471), .A2(n2261), .ZN(n2260) );
  NOR2_X1 U2456 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2373)
         );
  INV_X1 U2457 ( .A(IR_REG_14__SCAN_IN), .ZN(n4651) );
  INV_X1 U2458 ( .A(IR_REG_18__SCAN_IN), .ZN(n4577) );
  INV_X1 U2459 ( .A(IR_REG_20__SCAN_IN), .ZN(n2676) );
  NOR2_X1 U2460 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n4576)
         );
  NOR2_X1 U2461 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2376)
         );
  INV_X1 U2462 ( .A(IR_REG_15__SCAN_IN), .ZN(n2583) );
  NOR2_X1 U2463 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2539)
         );
  NAND2_X2 U2464 ( .A1(n2684), .A2(n2151), .ZN(n2868) );
  NAND2_X2 U2465 ( .A1(n3542), .A2(n3541), .ZN(n3669) );
  NAND2_X1 U2466 ( .A1(n2674), .A2(n2610), .ZN(n4010) );
  NAND2_X1 U2467 ( .A1(n2674), .A2(IR_REG_31__SCAN_IN), .ZN(n2675) );
  INV_X4 U2468 ( .A(n2406), .ZN(n2721) );
  NAND2_X2 U2470 ( .A1(n2868), .A2(n2983), .ZN(n3597) );
  NAND2_X2 U2471 ( .A1(n3711), .A2(n3582), .ZN(n3680) );
  AOI21_X2 U2472 ( .B1(n3294), .B2(n2166), .A(n2310), .ZN(n3435) );
  OAI21_X2 U2473 ( .B1(n2306), .B2(n2305), .A(n2174), .ZN(n3632) );
  AOI21_X2 U2474 ( .B1(n3213), .B2(n3214), .A(n3202), .ZN(n3248) );
  INV_X1 U2475 ( .A(n3597), .ZN(n2155) );
  XNOR2_X2 U2476 ( .A(n2675), .B(n2676), .ZN(n2684) );
  INV_X1 U2477 ( .A(n3055), .ZN(n2289) );
  NAND2_X1 U2478 ( .A1(n4396), .A2(n3162), .ZN(n3163) );
  INV_X1 U2479 ( .A(n2353), .ZN(n2349) );
  OR2_X1 U2480 ( .A1(n2693), .A2(n2200), .ZN(n2197) );
  AND3_X1 U2481 ( .A1(n2583), .A2(n4651), .A3(n4650), .ZN(n2584) );
  NAND2_X1 U2482 ( .A1(n2394), .A2(n2393), .ZN(n2397) );
  INV_X1 U2483 ( .A(n3290), .ZN(n3321) );
  NAND2_X1 U2484 ( .A1(n4397), .A2(n4398), .ZN(n4396) );
  AOI22_X1 U2485 ( .A1(n4044), .A2(n2659), .B1(n3599), .B2(n3940), .ZN(n4026)
         );
  NAND2_X1 U2486 ( .A1(n4155), .A2(n2627), .ZN(n2347) );
  NOR2_X1 U2487 ( .A1(n2363), .A2(n2173), .ZN(n2342) );
  NAND2_X1 U2488 ( .A1(n4045), .A2(n4245), .ZN(n4030) );
  AND2_X1 U2489 ( .A1(n4111), .A2(n2268), .ZN(n4045) );
  AND2_X1 U2490 ( .A1(n2163), .A2(n4249), .ZN(n2268) );
  AND2_X1 U2491 ( .A1(n2472), .A2(n2259), .ZN(n2257) );
  AND2_X1 U2492 ( .A1(n2360), .A2(n2260), .ZN(n2259) );
  INV_X1 U2493 ( .A(n3801), .ZN(n2212) );
  AND2_X1 U2494 ( .A1(n4191), .A2(n2701), .ZN(n3863) );
  INV_X1 U2495 ( .A(n3835), .ZN(n2200) );
  INV_X1 U2496 ( .A(n3317), .ZN(n2315) );
  AND2_X1 U2497 ( .A1(n3890), .A2(n4091), .ZN(n3871) );
  INV_X1 U2498 ( .A(n2245), .ZN(n2238) );
  AND2_X1 U2499 ( .A1(n2644), .A2(REG3_REG_25__SCAN_IN), .ZN(n2649) );
  NAND2_X1 U2500 ( .A1(n2205), .A2(n4043), .ZN(n2204) );
  INV_X1 U2501 ( .A(n2207), .ZN(n2205) );
  AND2_X1 U2502 ( .A1(n4064), .A2(n3599), .ZN(n3802) );
  AND2_X1 U2503 ( .A1(n3875), .A2(n2212), .ZN(n2209) );
  OR2_X1 U2504 ( .A1(n3878), .A2(n3802), .ZN(n3923) );
  NAND2_X1 U2505 ( .A1(n2329), .A2(n2328), .ZN(n2327) );
  INV_X1 U2506 ( .A(n2330), .ZN(n2328) );
  NAND2_X1 U2507 ( .A1(n4095), .A2(n4078), .ZN(n2335) );
  NAND2_X1 U2508 ( .A1(n4126), .A2(n4262), .ZN(n2336) );
  AND2_X1 U2509 ( .A1(n3862), .A2(n3787), .ZN(n2218) );
  INV_X1 U2510 ( .A(n4295), .ZN(n2757) );
  OAI21_X1 U2511 ( .B1(n2576), .B2(n2340), .A(n2592), .ZN(n2339) );
  NOR2_X1 U2512 ( .A1(n2509), .A2(n2354), .ZN(n2353) );
  INV_X1 U2513 ( .A(n2500), .ZN(n2354) );
  INV_X1 U2514 ( .A(n2199), .ZN(n2198) );
  OAI21_X1 U2515 ( .B1(n3834), .B2(n2200), .A(n3833), .ZN(n2199) );
  OR2_X1 U2516 ( .A1(n3101), .A2(n2692), .ZN(n2693) );
  NAND2_X1 U2517 ( .A1(n2437), .A2(n2436), .ZN(n3018) );
  NAND2_X1 U2518 ( .A1(n3455), .A2(n3461), .ZN(n2265) );
  INV_X1 U2519 ( .A(IR_REG_28__SCAN_IN), .ZN(n2395) );
  INV_X1 U2520 ( .A(IR_REG_22__SCAN_IN), .ZN(n2261) );
  INV_X1 U2521 ( .A(IR_REG_6__SCAN_IN), .ZN(n2471) );
  INV_X1 U2522 ( .A(IR_REG_17__SCAN_IN), .ZN(n2588) );
  OR2_X1 U2523 ( .A1(n2561), .A2(IR_REG_14__SCAN_IN), .ZN(n2562) );
  INV_X1 U2524 ( .A(IR_REG_1__SCAN_IN), .ZN(n2196) );
  NAND2_X1 U2525 ( .A1(n3282), .A2(n3281), .ZN(n3283) );
  NOR2_X1 U2526 ( .A1(n2304), .A2(n2303), .ZN(n2302) );
  INV_X1 U2527 ( .A(n2181), .ZN(n2304) );
  NAND2_X1 U2528 ( .A1(n2181), .A2(n2300), .ZN(n2299) );
  NAND2_X1 U2529 ( .A1(n2301), .A2(n3751), .ZN(n2300) );
  INV_X1 U2530 ( .A(n3682), .ZN(n2301) );
  OAI21_X1 U2531 ( .B1(n2424), .B2(n2793), .A(n2401), .ZN(n3034) );
  NAND2_X1 U2532 ( .A1(n2424), .A2(DATAI_1_), .ZN(n2401) );
  INV_X1 U2533 ( .A(n2314), .ZN(n2313) );
  OAI21_X1 U2534 ( .B1(n3293), .B2(n2315), .A(n3374), .ZN(n2314) );
  INV_X1 U2535 ( .A(n2317), .ZN(n2316) );
  OAI21_X1 U2536 ( .B1(n3293), .B2(n2318), .A(n3373), .ZN(n2317) );
  NAND2_X1 U2537 ( .A1(n2313), .A2(n2315), .ZN(n2311) );
  NAND2_X1 U2538 ( .A1(n2290), .A2(n2289), .ZN(n2288) );
  NAND2_X1 U2539 ( .A1(n2877), .A2(REG1_REG_0__SCAN_IN), .ZN(n2878) );
  INV_X1 U2540 ( .A(n3734), .ZN(n3563) );
  NAND2_X1 U2541 ( .A1(n2621), .A2(REG3_REG_21__SCAN_IN), .ZN(n2630) );
  INV_X1 U2542 ( .A(n4487), .ZN(n2929) );
  OR2_X1 U2543 ( .A1(n2579), .A2(n2578), .ZN(n2594) );
  NAND2_X1 U2544 ( .A1(n2226), .A2(n2231), .ZN(n2224) );
  NAND2_X1 U2545 ( .A1(n2246), .A2(REG2_REG_8__SCAN_IN), .ZN(n2245) );
  NOR2_X1 U2546 ( .A1(n2243), .A2(n2241), .ZN(n2240) );
  INV_X1 U2547 ( .A(n4376), .ZN(n2241) );
  NAND2_X1 U2548 ( .A1(n4407), .A2(n3164), .ZN(n3167) );
  NAND2_X1 U2549 ( .A1(n3167), .A2(n3166), .ZN(n3970) );
  NOR2_X1 U2550 ( .A1(n4427), .A2(n2223), .ZN(n3988) );
  AND2_X1 U2551 ( .A1(n3986), .A2(REG2_REG_15__SCAN_IN), .ZN(n2223) );
  NAND2_X1 U2552 ( .A1(n4432), .A2(n3974), .ZN(n3975) );
  NAND2_X1 U2553 ( .A1(n4000), .A2(n2254), .ZN(n2253) );
  OR2_X1 U2554 ( .A1(n4363), .A2(REG2_REG_17__SCAN_IN), .ZN(n2254) );
  AND2_X1 U2555 ( .A1(n2649), .A2(REG3_REG_26__SCAN_IN), .ZN(n2661) );
  AOI21_X1 U2556 ( .B1(n4054), .B2(n2653), .A(n2334), .ZN(n4044) );
  NOR2_X1 U2557 ( .A1(n4061), .A2(n4038), .ZN(n2334) );
  NOR2_X1 U2558 ( .A1(n2332), .A2(n2331), .ZN(n2330) );
  INV_X1 U2559 ( .A(n2336), .ZN(n2332) );
  INV_X1 U2560 ( .A(n2636), .ZN(n2331) );
  NAND2_X1 U2561 ( .A1(n2620), .A2(n3899), .ZN(n4155) );
  NAND2_X1 U2562 ( .A1(n3450), .A2(n3448), .ZN(n2219) );
  NAND2_X1 U2563 ( .A1(n2156), .A2(n2576), .ZN(n3449) );
  NOR2_X1 U2564 ( .A1(n2176), .A2(n2345), .ZN(n2344) );
  INV_X1 U2565 ( .A(n2530), .ZN(n2345) );
  AND2_X1 U2566 ( .A1(n2355), .A2(n2356), .ZN(n2351) );
  OR2_X1 U2567 ( .A1(n3321), .A2(n3346), .ZN(n2356) );
  NAND2_X1 U2568 ( .A1(n2501), .A2(n2353), .ZN(n2352) );
  NAND2_X1 U2569 ( .A1(n2695), .A2(n3847), .ZN(n3263) );
  INV_X1 U2570 ( .A(n3252), .ZN(n3257) );
  AND2_X1 U2571 ( .A1(n2895), .A2(n2860), .ZN(n4217) );
  NAND2_X1 U2572 ( .A1(n2972), .A2(n2971), .ZN(n3030) );
  INV_X1 U2573 ( .A(n4220), .ZN(n4476) );
  INV_X1 U2574 ( .A(n3034), .ZN(n3040) );
  NAND2_X1 U2575 ( .A1(n4111), .A2(n2163), .ZN(n4065) );
  NOR2_X1 U2576 ( .A1(n4143), .A2(n4112), .ZN(n4111) );
  NAND2_X1 U2577 ( .A1(n3339), .A2(n3441), .ZN(n3412) );
  XNOR2_X1 U2578 ( .A(n2380), .B(n2379), .ZN(n2386) );
  INV_X1 U2579 ( .A(IR_REG_30__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U2580 ( .A1(n2776), .A2(n2383), .ZN(n2387) );
  NAND2_X1 U2581 ( .A1(n2382), .A2(n2381), .ZN(n2383) );
  NOR2_X1 U2582 ( .A1(n2371), .A2(n2370), .ZN(n2372) );
  AND2_X1 U2583 ( .A1(n2498), .A2(n2517), .ZN(n3173) );
  NAND2_X1 U2584 ( .A1(n2196), .A2(n2195), .ZN(n2399) );
  NOR2_X1 U2585 ( .A1(n2175), .A2(n2307), .ZN(n2305) );
  INV_X1 U2586 ( .A(n4152), .ZN(n3674) );
  AOI21_X1 U2587 ( .B1(n2297), .B2(n2299), .A(n2296), .ZN(n2295) );
  INV_X1 U2588 ( .A(n3625), .ZN(n2296) );
  INV_X1 U2589 ( .A(n2302), .ZN(n2297) );
  INV_X1 U2590 ( .A(n2299), .ZN(n2298) );
  INV_X1 U2591 ( .A(n2992), .ZN(n4480) );
  AND2_X1 U2592 ( .A1(n2894), .A2(n4114), .ZN(n3772) );
  XNOR2_X1 U2593 ( .A(n2836), .B(n4365), .ZN(n2838) );
  XNOR2_X1 U2594 ( .A(n3975), .B(n3987), .ZN(n4441) );
  NAND2_X1 U2595 ( .A1(n2252), .A2(n4410), .ZN(n2251) );
  NAND2_X1 U2596 ( .A1(n2253), .A2(n4448), .ZN(n2252) );
  AOI21_X1 U2597 ( .B1(n4450), .B2(ADDR_REG_18__SCAN_IN), .A(n4449), .ZN(n2250) );
  NOR2_X1 U2598 ( .A1(n2253), .A2(n4448), .ZN(n4447) );
  NOR2_X1 U2599 ( .A1(n4004), .A2(n4005), .ZN(n4453) );
  NAND2_X1 U2600 ( .A1(n4453), .A2(n4454), .ZN(n4451) );
  AND2_X1 U2601 ( .A1(n3953), .A2(n3950), .ZN(n4452) );
  OAI21_X1 U2602 ( .B1(n2758), .B2(n3795), .A(n4239), .ZN(n3619) );
  OR2_X1 U2603 ( .A1(n3619), .A2(n4300), .ZN(n2765) );
  OR2_X1 U2604 ( .A1(n3619), .A2(n4352), .ZN(n2760) );
  AND2_X1 U2605 ( .A1(n4244), .A2(n2221), .ZN(n4313) );
  AOI21_X1 U2606 ( .B1(n4246), .B2(n4542), .A(n2222), .ZN(n2221) );
  NOR2_X1 U2607 ( .A1(n4294), .A2(n4245), .ZN(n2222) );
  INV_X1 U2608 ( .A(n3279), .ZN(n3282) );
  AND2_X1 U2609 ( .A1(n2713), .A2(n4055), .ZN(n3880) );
  INV_X1 U2610 ( .A(n2228), .ZN(n2226) );
  NAND2_X1 U2611 ( .A1(n2208), .A2(n2212), .ZN(n2207) );
  INV_X1 U2612 ( .A(n3880), .ZN(n2208) );
  NAND2_X1 U2613 ( .A1(n3263), .A2(n3849), .ZN(n3302) );
  AND2_X1 U2614 ( .A1(n3826), .A2(n3829), .ZN(n3905) );
  AND2_X1 U2615 ( .A1(n3823), .A2(n3820), .ZN(n4473) );
  OAI21_X1 U2616 ( .B1(n2686), .B2(n3030), .A(n3819), .ZN(n4472) );
  NAND2_X1 U2617 ( .A1(n2973), .A2(n3034), .ZN(n3819) );
  INV_X1 U2618 ( .A(IR_REG_26__SCAN_IN), .ZN(n4669) );
  NOR2_X1 U2619 ( .A1(n4078), .A2(n3575), .ZN(n2269) );
  AND2_X1 U2620 ( .A1(n3017), .A2(n3020), .ZN(n3016) );
  AND2_X1 U2621 ( .A1(n2258), .A2(n2170), .ZN(n2719) );
  INV_X1 U2622 ( .A(n3492), .ZN(n2309) );
  AND2_X1 U2623 ( .A1(n3436), .A2(n2308), .ZN(n2307) );
  INV_X1 U2624 ( .A(n3491), .ZN(n2308) );
  OR3_X1 U2625 ( .A1(n2630), .A2(n4636), .A3(n3735), .ZN(n2637) );
  INV_X1 U2626 ( .A(n3292), .ZN(n3293) );
  INV_X1 U2627 ( .A(n3949), .ZN(n2972) );
  AND2_X1 U2628 ( .A1(n3779), .A2(DATAI_21_), .ZN(n3555) );
  AND2_X1 U2629 ( .A1(n3579), .A2(n3578), .ZN(n3580) );
  NAND2_X1 U2630 ( .A1(n3721), .A2(n2159), .ZN(n2282) );
  NAND2_X1 U2631 ( .A1(n3081), .A2(n2289), .ZN(n2286) );
  NAND2_X1 U2632 ( .A1(n2285), .A2(n3081), .ZN(n2284) );
  NOR2_X1 U2633 ( .A1(n2547), .A2(n3639), .ZN(n2555) );
  OR2_X1 U2634 ( .A1(n2661), .A2(n2650), .ZN(n3753) );
  AND2_X1 U2635 ( .A1(n2447), .A2(n2446), .ZN(n3083) );
  NAND2_X1 U2636 ( .A1(n2941), .A2(n2236), .ZN(n2235) );
  NAND2_X1 U2637 ( .A1(n4369), .A2(REG2_REG_2__SCAN_IN), .ZN(n2236) );
  AOI21_X1 U2638 ( .B1(n2801), .B2(REG2_REG_3__SCAN_IN), .A(n2234), .ZN(n2802)
         );
  AND2_X1 U2639 ( .A1(n2235), .A2(n4368), .ZN(n2234) );
  AOI21_X1 U2640 ( .B1(n2233), .B2(n2229), .A(n2829), .ZN(n2228) );
  NAND2_X1 U2641 ( .A1(n2280), .A2(n2279), .ZN(n2278) );
  INV_X1 U2642 ( .A(n2826), .ZN(n2279) );
  AOI21_X1 U2643 ( .B1(n2238), .B2(n2240), .A(n2182), .ZN(n2237) );
  INV_X1 U2644 ( .A(n2240), .ZN(n2239) );
  XNOR2_X1 U2645 ( .A(n3163), .B(n4503), .ZN(n4408) );
  INV_X1 U2646 ( .A(IR_REG_10__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U2647 ( .A1(n3970), .A2(n3971), .ZN(n3972) );
  OAI21_X1 U2648 ( .B1(n3982), .B2(n3981), .A(n3980), .ZN(n3983) );
  OR2_X1 U2649 ( .A1(n4030), .A2(n3800), .ZN(n4239) );
  AND2_X1 U2650 ( .A1(n2209), .A2(n4043), .ZN(n2206) );
  NAND2_X1 U2651 ( .A1(n2204), .A2(n2203), .ZN(n2202) );
  INV_X1 U2652 ( .A(n3802), .ZN(n2203) );
  NAND2_X1 U2653 ( .A1(n2201), .A2(n2207), .ZN(n4037) );
  NAND2_X1 U2654 ( .A1(n2712), .A2(n2209), .ZN(n2201) );
  INV_X1 U2655 ( .A(n3923), .ZN(n4043) );
  OAI22_X1 U2656 ( .A1(n4110), .A2(n2325), .B1(n2324), .B2(n2168), .ZN(n4054)
         );
  INV_X1 U2657 ( .A(n2335), .ZN(n2324) );
  NAND2_X1 U2658 ( .A1(n2329), .A2(n2335), .ZN(n2325) );
  NAND2_X1 U2659 ( .A1(n2712), .A2(n3875), .ZN(n4056) );
  NAND2_X1 U2660 ( .A1(n2712), .A2(n3889), .ZN(n4076) );
  NAND2_X1 U2661 ( .A1(n2705), .A2(n3789), .ZN(n4151) );
  OAI21_X1 U2662 ( .B1(n3450), .B2(n2216), .A(n2213), .ZN(n2705) );
  AND2_X1 U2663 ( .A1(n3867), .A2(n2214), .ZN(n2213) );
  NAND2_X1 U2664 ( .A1(n2215), .A2(n2576), .ZN(n2214) );
  AND2_X1 U2665 ( .A1(n2613), .A2(n2385), .ZN(n2621) );
  NAND2_X1 U2666 ( .A1(n2219), .A2(n2215), .ZN(n4165) );
  AND2_X1 U2667 ( .A1(n2219), .A2(n2218), .ZN(n4190) );
  OR3_X1 U2668 ( .A1(n3511), .A2(n2265), .A3(n2757), .ZN(n2264) );
  OAI22_X1 U2669 ( .A1(n2156), .A2(n2337), .B1(n2338), .B2(n2591), .ZN(n4212)
         );
  NAND2_X1 U2670 ( .A1(n2341), .A2(n2577), .ZN(n2337) );
  INV_X1 U2671 ( .A(n2339), .ZN(n2338) );
  NAND2_X1 U2672 ( .A1(n4212), .A2(n4214), .ZN(n4211) );
  AND2_X1 U2673 ( .A1(n2582), .A2(n2581), .ZN(n4221) );
  AND2_X1 U2674 ( .A1(n2555), .A2(REG3_REG_15__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U2675 ( .A1(n2567), .A2(REG3_REG_16__SCAN_IN), .ZN(n2579) );
  OAI21_X1 U2676 ( .B1(n3302), .B2(n3852), .A(n3854), .ZN(n3785) );
  NAND2_X1 U2677 ( .A1(n2531), .A2(n2530), .ZN(n3402) );
  INV_X1 U2678 ( .A(n3944), .ZN(n3338) );
  OAI21_X1 U2679 ( .B1(n2501), .B2(n2350), .A(n2348), .ZN(n3308) );
  AOI21_X1 U2680 ( .B1(n2351), .B2(n2349), .A(n2179), .ZN(n2348) );
  INV_X1 U2681 ( .A(n2351), .ZN(n2350) );
  INV_X1 U2682 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U2683 ( .A1(n2197), .A2(n2180), .ZN(n2694) );
  OR2_X1 U2684 ( .A1(n2502), .A2(n4635), .ZN(n2511) );
  NAND2_X1 U2685 ( .A1(n2197), .A2(n2198), .ZN(n3140) );
  OAI21_X1 U2686 ( .B1(n4537), .B2(n2172), .A(n2322), .ZN(n3144) );
  INV_X1 U2687 ( .A(n2323), .ZN(n2322) );
  OAI21_X1 U2688 ( .B1(n2479), .B2(n2172), .A(n2488), .ZN(n2323) );
  INV_X1 U2689 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2489) );
  OR2_X1 U2690 ( .A1(n2490), .A2(n2489), .ZN(n2502) );
  NAND2_X1 U2691 ( .A1(n2693), .A2(n3834), .ZN(n3236) );
  AND2_X1 U2692 ( .A1(n2483), .A2(n2482), .ZN(n3256) );
  NAND2_X1 U2693 ( .A1(n2456), .A2(REG3_REG_6__SCAN_IN), .ZN(n2465) );
  INV_X1 U2694 ( .A(n3050), .ZN(n3020) );
  AND2_X1 U2695 ( .A1(n3033), .A2(n2415), .ZN(n2364) );
  INV_X1 U2696 ( .A(n4473), .ZN(n2425) );
  NAND2_X1 U2697 ( .A1(n2364), .A2(n2425), .ZN(n4470) );
  NAND2_X1 U2698 ( .A1(n3816), .A2(n3819), .ZN(n2686) );
  INV_X1 U2699 ( .A(n4217), .ZN(n4479) );
  INV_X1 U2700 ( .A(IR_REG_13__SCAN_IN), .ZN(n4657) );
  NOR2_X1 U2701 ( .A1(n4239), .A2(n4240), .ZN(n4238) );
  INV_X1 U2702 ( .A(n4034), .ZN(n4245) );
  NAND2_X1 U2703 ( .A1(n4111), .A2(n2269), .ZN(n4083) );
  NAND2_X1 U2704 ( .A1(n4111), .A2(n4262), .ZN(n4102) );
  INV_X1 U2705 ( .A(n4123), .ZN(n4112) );
  AND2_X1 U2706 ( .A1(n3779), .A2(DATAI_22_), .ZN(n4144) );
  NOR3_X1 U2707 ( .A1(n4225), .A2(n4198), .A3(n4180), .ZN(n4179) );
  OR2_X1 U2708 ( .A1(n4224), .A2(n4216), .ZN(n4225) );
  NOR3_X1 U2709 ( .A1(n3412), .A2(n3511), .A3(n3638), .ZN(n3456) );
  INV_X1 U2710 ( .A(n3439), .ZN(n3441) );
  AND2_X1 U2711 ( .A1(n3231), .A2(n2185), .ZN(n3339) );
  NAND2_X1 U2712 ( .A1(n3231), .A2(n2157), .ZN(n3270) );
  NAND2_X1 U2713 ( .A1(n3231), .A2(n3257), .ZN(n3225) );
  NOR2_X1 U2714 ( .A1(n3106), .A2(n3197), .ZN(n3234) );
  AND2_X1 U2715 ( .A1(n3234), .A2(n3233), .ZN(n3231) );
  OR2_X1 U2716 ( .A1(n3096), .A2(n3133), .ZN(n3106) );
  NOR2_X1 U2717 ( .A1(n4484), .A2(n3012), .ZN(n3017) );
  OR2_X1 U2718 ( .A1(n4486), .A2(n4487), .ZN(n4484) );
  MUX2_X1 U2719 ( .A(n4369), .B(DATAI_2_), .S(n2424), .Z(n4487) );
  XNOR2_X1 U2720 ( .A(n2735), .B(n2361), .ZN(n2741) );
  XNOR2_X1 U2721 ( .A(n2733), .B(n2732), .ZN(n2755) );
  NAND2_X1 U2722 ( .A1(n2607), .A2(n4577), .ZN(n2679) );
  AND2_X1 U2723 ( .A1(n2573), .A2(n2564), .ZN(n3986) );
  AND2_X1 U2724 ( .A1(n2520), .A2(n2527), .ZN(n3172) );
  INV_X1 U2725 ( .A(IR_REG_3__SCAN_IN), .ZN(n2432) );
  MUX2_X1 U2726 ( .A(IR_REG_31__SCAN_IN), .B(n2398), .S(IR_REG_1__SCAN_IN), 
        .Z(n2400) );
  OR2_X1 U2727 ( .A1(n4028), .A2(n2384), .ZN(n2669) );
  NAND2_X1 U2728 ( .A1(n2294), .A2(n2299), .ZN(n3626) );
  NAND2_X1 U2729 ( .A1(n3294), .A2(n3293), .ZN(n3318) );
  AND2_X1 U2730 ( .A1(n2292), .A2(n3606), .ZN(n2291) );
  INV_X1 U2731 ( .A(n3555), .ZN(n4277) );
  NAND2_X1 U2732 ( .A1(n2312), .A2(n2311), .ZN(n2310) );
  NAND2_X1 U2733 ( .A1(n2316), .A2(n2318), .ZN(n2312) );
  AND2_X1 U2734 ( .A1(n2642), .A2(n2641), .ZN(n4126) );
  INV_X1 U2735 ( .A(n3943), .ZN(n3696) );
  INV_X1 U2736 ( .A(n3947), .ZN(n3130) );
  INV_X1 U2737 ( .A(n2285), .ZN(n2287) );
  NAND2_X1 U2738 ( .A1(n2288), .A2(n2192), .ZN(n3056) );
  NAND2_X1 U2739 ( .A1(n2411), .A2(n4652), .ZN(n2413) );
  INV_X1 U2740 ( .A(n3772), .ZN(n3755) );
  NAND2_X1 U2741 ( .A1(n2282), .A2(n3668), .ZN(n3733) );
  AND2_X1 U2742 ( .A1(n2658), .A2(n2657), .ZN(n4064) );
  INV_X1 U2743 ( .A(n3758), .ZN(n3774) );
  OAI211_X1 U2744 ( .C1(n3684), .C2(n2384), .A(n2647), .B(n2646), .ZN(n4095)
         );
  INV_X1 U2745 ( .A(n3083), .ZN(n3132) );
  INV_X1 U2746 ( .A(n3009), .ZN(n3035) );
  CLKBUF_X1 U2747 ( .A(U4043), .Z(n2937) );
  OR2_X1 U2748 ( .A1(n2983), .A2(n4495), .ZN(n3948) );
  NAND2_X1 U2749 ( .A1(n2942), .A2(n2943), .ZN(n2941) );
  XNOR2_X1 U2750 ( .A(n2235), .B(n2796), .ZN(n2801) );
  AOI21_X1 U2751 ( .B1(n2952), .B2(REG2_REG_4__SCAN_IN), .A(n2230), .ZN(n2830)
         );
  NAND2_X1 U2752 ( .A1(n2374), .A2(n2373), .ZN(n2448) );
  NOR2_X1 U2753 ( .A1(n2276), .A2(n2274), .ZN(n2273) );
  INV_X1 U2754 ( .A(n4365), .ZN(n2274) );
  AOI22_X1 U2755 ( .A1(n2838), .A2(REG2_REG_6__SCAN_IN), .B1(n4365), .B2(n2837), .ZN(n2840) );
  XNOR2_X1 U2756 ( .A(n3175), .B(n3174), .ZN(n3177) );
  NAND2_X1 U2757 ( .A1(n2242), .A2(n2240), .ZN(n4375) );
  NAND2_X1 U2758 ( .A1(n3175), .A2(n2245), .ZN(n2242) );
  XNOR2_X1 U2759 ( .A(n3972), .B(n4426), .ZN(n4423) );
  NOR2_X1 U2760 ( .A1(n4429), .A2(n4428), .ZN(n4427) );
  XNOR2_X1 U2761 ( .A(n3988), .B(n3987), .ZN(n4438) );
  NAND2_X1 U2762 ( .A1(n4438), .A2(n4780), .ZN(n4437) );
  NOR2_X1 U2763 ( .A1(n4442), .A2(n3976), .ZN(n3979) );
  XNOR2_X1 U2764 ( .A(n2275), .B(n4007), .ZN(n4012) );
  NAND2_X1 U2765 ( .A1(n4451), .A2(n2193), .ZN(n2275) );
  XNOR2_X1 U2766 ( .A(n4026), .B(n4021), .ZN(n4246) );
  NAND2_X1 U2767 ( .A1(n2326), .A2(n2329), .ZN(n4074) );
  NAND2_X1 U2768 ( .A1(n4110), .A2(n2330), .ZN(n2326) );
  AND2_X1 U2769 ( .A1(n2333), .A2(n2165), .ZN(n4101) );
  NAND2_X1 U2770 ( .A1(n4110), .A2(n2636), .ZN(n2333) );
  NAND2_X1 U2771 ( .A1(n2347), .A2(n2628), .ZN(n4132) );
  NOR2_X1 U2772 ( .A1(n2217), .A2(n3858), .ZN(n3471) );
  INV_X1 U2773 ( .A(n2219), .ZN(n2217) );
  NAND2_X1 U2774 ( .A1(n3449), .A2(n2577), .ZN(n3473) );
  AND2_X1 U2775 ( .A1(n2343), .A2(n2346), .ZN(n3420) );
  NAND2_X1 U2776 ( .A1(n2352), .A2(n2351), .ZN(n3269) );
  NAND2_X1 U2777 ( .A1(n2352), .A2(n2356), .ZN(n3267) );
  NAND2_X1 U2778 ( .A1(n2501), .A2(n2500), .ZN(n3224) );
  NAND2_X1 U2779 ( .A1(n4537), .A2(n2479), .ZN(n3235) );
  INV_X1 U2780 ( .A(n4235), .ZN(n4156) );
  INV_X1 U2781 ( .A(n4207), .ZN(n4488) );
  INV_X1 U2782 ( .A(n4483), .ZN(n4114) );
  OAI21_X1 U2783 ( .B1(n4047), .B2(n4249), .A(n4046), .ZN(n4318) );
  NAND2_X1 U2784 ( .A1(n2779), .A2(n2963), .ZN(n4493) );
  NAND2_X1 U2785 ( .A1(n2167), .A2(n2258), .ZN(n2776) );
  INV_X1 U2786 ( .A(n2895), .ZN(n4357) );
  XNOR2_X1 U2787 ( .A(n2738), .B(IR_REG_26__SCAN_IN), .ZN(n2772) );
  INV_X1 U2788 ( .A(n2741), .ZN(n4358) );
  INV_X1 U2789 ( .A(n2755), .ZN(n4359) );
  XNOR2_X1 U2790 ( .A(n2682), .B(IR_REG_22__SCAN_IN), .ZN(n4360) );
  INV_X1 U2791 ( .A(n4010), .ZN(n4362) );
  INV_X1 U2792 ( .A(n2249), .ZN(n4456) );
  OAI21_X1 U2793 ( .B1(n4447), .B2(n2251), .A(n2250), .ZN(n2249) );
  AND2_X1 U2794 ( .A1(n2765), .A2(n2362), .ZN(n2766) );
  OAI21_X1 U2795 ( .B1(n4313), .B2(n4557), .A(n2160), .ZN(U3546) );
  OR2_X1 U2796 ( .A1(n4314), .A2(n4300), .ZN(n2220) );
  AND2_X1 U2797 ( .A1(n2760), .A2(n2759), .ZN(n2761) );
  OAI21_X1 U2798 ( .B1(n4313), .B2(n4544), .A(n2161), .ZN(U3514) );
  OR2_X1 U2799 ( .A1(n4314), .A2(n4352), .ZN(n2357) );
  AND2_X1 U2800 ( .A1(n2566), .A2(n2565), .ZN(n2156) );
  XNOR2_X1 U2801 ( .A(n2248), .B(n2247), .ZN(n4369) );
  INV_X1 U2802 ( .A(n2147), .ZN(n2820) );
  AND2_X1 U2803 ( .A1(n3257), .A2(n3346), .ZN(n2157) );
  INV_X1 U2804 ( .A(n3174), .ZN(n2246) );
  OR2_X1 U2805 ( .A1(n4225), .A2(n2255), .ZN(n2158) );
  AND2_X1 U2806 ( .A1(n2189), .A2(n3724), .ZN(n2159) );
  AND2_X1 U2807 ( .A1(n2220), .A2(n2190), .ZN(n2160) );
  AND2_X1 U2808 ( .A1(n2357), .A2(n2191), .ZN(n2161) );
  NAND2_X1 U2809 ( .A1(n2169), .A2(n2336), .ZN(n2329) );
  AND2_X1 U2810 ( .A1(n2157), .A2(n3357), .ZN(n2162) );
  AND2_X1 U2811 ( .A1(n2269), .A2(n4066), .ZN(n2163) );
  AND2_X1 U2812 ( .A1(n2242), .A2(n2244), .ZN(n2164) );
  INV_X4 U2813 ( .A(n2384), .ZN(n2420) );
  NAND2_X1 U2814 ( .A1(n2400), .A2(n2399), .ZN(n2793) );
  NAND2_X1 U2815 ( .A1(n4137), .A2(n4112), .ZN(n2165) );
  AND2_X1 U2816 ( .A1(n2443), .A2(n2434), .ZN(n4368) );
  NAND2_X1 U2817 ( .A1(n2262), .A2(n2375), .ZN(n2681) );
  OR2_X1 U2818 ( .A1(n2316), .A2(n2313), .ZN(n2166) );
  AND3_X1 U2819 ( .A1(n2358), .A2(n2375), .A3(n2378), .ZN(n2167) );
  AND2_X1 U2820 ( .A1(n2327), .A2(n2648), .ZN(n2168) );
  NAND2_X1 U2821 ( .A1(n2643), .A2(n2165), .ZN(n2169) );
  NAND2_X1 U2822 ( .A1(n2608), .A2(n2677), .ZN(n2674) );
  AND2_X1 U2823 ( .A1(n2358), .A2(n2375), .ZN(n2170) );
  INV_X1 U2824 ( .A(n2233), .ZN(n2230) );
  NAND2_X1 U2825 ( .A1(n2803), .A2(n4367), .ZN(n2233) );
  AND2_X1 U2826 ( .A1(n4669), .A2(n2377), .ZN(n2171) );
  INV_X1 U2827 ( .A(IR_REG_2__SCAN_IN), .ZN(n2247) );
  INV_X1 U2828 ( .A(IR_REG_25__SCAN_IN), .ZN(n2361) );
  OR2_X1 U2829 ( .A1(n3887), .A2(n2211), .ZN(n2210) );
  AND2_X1 U2830 ( .A1(n3256), .A2(n3233), .ZN(n2172) );
  AND2_X1 U2831 ( .A1(n2545), .A2(n2544), .ZN(n2585) );
  AND2_X1 U2832 ( .A1(n2472), .A2(n2471), .ZN(n2545) );
  AND2_X1 U2833 ( .A1(n2472), .A2(n2471), .ZN(n2262) );
  NAND2_X1 U2834 ( .A1(n3318), .A2(n3317), .ZN(n3375) );
  INV_X1 U2835 ( .A(IR_REG_5__SCAN_IN), .ZN(n2321) );
  OAI211_X1 U2836 ( .C1(n3753), .C2(n2384), .A(n2652), .B(n2651), .ZN(n4038)
         );
  INV_X1 U2837 ( .A(IR_REG_31__SCAN_IN), .ZN(n2730) );
  INV_X1 U2838 ( .A(n3889), .ZN(n2211) );
  NOR2_X1 U2839 ( .A1(n3803), .A2(n3798), .ZN(n4027) );
  AND2_X1 U2840 ( .A1(n3943), .A2(n3511), .ZN(n2173) );
  INV_X1 U2841 ( .A(n3271), .ZN(n3357) );
  INV_X1 U2842 ( .A(n3681), .ZN(n2303) );
  OR2_X1 U2843 ( .A1(n3491), .A2(n3492), .ZN(n2174) );
  NOR3_X1 U2844 ( .A1(n4225), .A2(n2255), .A3(n4144), .ZN(n2256) );
  AND2_X1 U2845 ( .A1(n3436), .A2(n2309), .ZN(n2175) );
  OR2_X1 U2846 ( .A1(n3401), .A2(n2554), .ZN(n2176) );
  INV_X1 U2847 ( .A(n2577), .ZN(n2340) );
  NAND2_X1 U2848 ( .A1(n3251), .A2(n3257), .ZN(n2177) );
  AND2_X1 U2849 ( .A1(n3537), .A2(n3536), .ZN(n2178) );
  AND2_X1 U2850 ( .A1(n3387), .A2(n3357), .ZN(n2179) );
  AND2_X1 U2851 ( .A1(n2198), .A2(n2177), .ZN(n2180) );
  INV_X1 U2852 ( .A(n3379), .ZN(n3388) );
  NAND2_X1 U2853 ( .A1(n3596), .A2(n3595), .ZN(n2181) );
  NAND2_X1 U2854 ( .A1(n4366), .A2(REG2_REG_5__SCAN_IN), .ZN(n2231) );
  AND2_X1 U2855 ( .A1(n3173), .A2(REG2_REG_9__SCAN_IN), .ZN(n2182) );
  INV_X1 U2856 ( .A(n2591), .ZN(n2341) );
  INV_X1 U2857 ( .A(n2216), .ZN(n2215) );
  NAND2_X1 U2858 ( .A1(n3863), .A2(n2218), .ZN(n2216) );
  AND2_X1 U2859 ( .A1(n4119), .A2(n2708), .ZN(n4135) );
  INV_X1 U2860 ( .A(n4135), .ZN(n2629) );
  AND2_X1 U2861 ( .A1(n3563), .A2(n3668), .ZN(n2183) );
  AND2_X1 U2862 ( .A1(n2629), .A2(n2628), .ZN(n2184) );
  AND2_X1 U2863 ( .A1(n2162), .A2(n3388), .ZN(n2185) );
  INV_X1 U2864 ( .A(IR_REG_27__SCAN_IN), .ZN(n2377) );
  AND2_X1 U2865 ( .A1(n3231), .A2(n2162), .ZN(n2186) );
  OR2_X1 U2866 ( .A1(n4225), .A2(n4198), .ZN(n2187) );
  INV_X1 U2867 ( .A(n3908), .ZN(n2355) );
  INV_X1 U2868 ( .A(n2263), .ZN(n4301) );
  NOR3_X1 U2869 ( .A1(n3412), .A2(n3511), .A3(n2265), .ZN(n2263) );
  AND2_X1 U2870 ( .A1(n2691), .A2(n3834), .ZN(n3906) );
  INV_X1 U2871 ( .A(n3906), .ZN(n2477) );
  NOR2_X1 U2872 ( .A1(n3412), .A2(n3638), .ZN(n2267) );
  AND2_X1 U2873 ( .A1(n2288), .A2(n2287), .ZN(n2188) );
  NOR2_X1 U2874 ( .A1(n3412), .A2(n2264), .ZN(n2266) );
  NAND2_X1 U2875 ( .A1(n3557), .A2(n3558), .ZN(n2189) );
  INV_X1 U2876 ( .A(n4180), .ZN(n3727) );
  INV_X1 U2877 ( .A(n2363), .ZN(n2346) );
  INV_X1 U2878 ( .A(n4559), .ZN(n4557) );
  NAND2_X1 U2879 ( .A1(n2970), .A2(n2684), .ZN(n2871) );
  AND2_X1 U2880 ( .A1(n3953), .A2(n2788), .ZN(n4410) );
  OR2_X1 U2881 ( .A1(n4559), .A2(n4247), .ZN(n2190) );
  OR2_X1 U2882 ( .A1(n4545), .A2(n4735), .ZN(n2191) );
  OR2_X1 U2883 ( .A1(n3053), .A2(n3052), .ZN(n2192) );
  INV_X1 U2884 ( .A(n3575), .ZN(n4262) );
  AND2_X1 U2885 ( .A1(n3779), .A2(DATAI_24_), .ZN(n3575) );
  INV_X1 U2886 ( .A(n2244), .ZN(n2243) );
  NAND2_X1 U2887 ( .A1(n3174), .A2(n3176), .ZN(n2244) );
  INV_X1 U2888 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2229) );
  OR2_X1 U2889 ( .A1(n4497), .A2(n4006), .ZN(n2193) );
  NAND2_X1 U2890 ( .A1(n2845), .A2(n4555), .ZN(n2194) );
  AND2_X1 U2891 ( .A1(n2399), .A2(IR_REG_31__SCAN_IN), .ZN(n2248) );
  AOI21_X1 U2892 ( .B1(n2712), .B2(n2206), .A(n2202), .ZN(n4022) );
  NAND2_X1 U2893 ( .A1(n2225), .A2(n2224), .ZN(n2836) );
  NAND3_X1 U2894 ( .A1(n2227), .A2(n2231), .A3(n2233), .ZN(n2225) );
  OAI21_X1 U2895 ( .B1(n2952), .B2(n2230), .A(n2228), .ZN(n2232) );
  INV_X1 U2896 ( .A(n2952), .ZN(n2227) );
  INV_X1 U2897 ( .A(n2232), .ZN(n2828) );
  OAI21_X1 U2898 ( .B1(n3175), .B2(n2239), .A(n2237), .ZN(n3178) );
  NAND3_X1 U2899 ( .A1(n4203), .A2(n3727), .A3(n4277), .ZN(n2255) );
  INV_X1 U2900 ( .A(n2256), .ZN(n4143) );
  AND2_X1 U2901 ( .A1(n2472), .A2(n2260), .ZN(n2258) );
  NAND2_X1 U2902 ( .A1(n2257), .A2(n2375), .ZN(n2737) );
  INV_X1 U2903 ( .A(n2266), .ZN(n4224) );
  INV_X1 U2904 ( .A(n2267), .ZN(n3427) );
  INV_X1 U2905 ( .A(n2280), .ZN(n2827) );
  INV_X1 U2906 ( .A(n2278), .ZN(n2825) );
  NAND2_X1 U2907 ( .A1(n2808), .A2(n4367), .ZN(n2281) );
  NAND2_X1 U2908 ( .A1(IR_REG_31__SCAN_IN), .A2(n4652), .ZN(n2398) );
  NAND2_X1 U2909 ( .A1(n2431), .A2(IR_REG_31__SCAN_IN), .ZN(n2433) );
  NAND2_X1 U2910 ( .A1(n2497), .A2(IR_REG_31__SCAN_IN), .ZN(n2496) );
  NAND2_X1 U2911 ( .A1(n2561), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U2912 ( .A1(n2734), .A2(IR_REG_31__SCAN_IN), .ZN(n2735) );
  OAI21_X1 U2913 ( .B1(n2517), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2519) );
  NAND2_X1 U2914 ( .A1(n2776), .A2(IR_REG_31__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U2915 ( .A1(n2737), .A2(IR_REG_31__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U2916 ( .A1(n2679), .A2(IR_REG_31__SCAN_IN), .ZN(n2608) );
  OAI21_X1 U2917 ( .B1(n2737), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2392) );
  OAI21_X1 U2918 ( .B1(n2679), .B2(n2678), .A(IR_REG_31__SCAN_IN), .ZN(n2680)
         );
  NAND2_X1 U2919 ( .A1(n2282), .A2(n2183), .ZN(n3647) );
  NAND2_X1 U2920 ( .A1(n3721), .A2(n3724), .ZN(n3673) );
  INV_X1 U2921 ( .A(n3057), .ZN(n2283) );
  OAI21_X2 U2922 ( .B1(n3054), .B2(n2286), .A(n2284), .ZN(n3128) );
  INV_X1 U2923 ( .A(n3054), .ZN(n2290) );
  OAI21_X2 U2924 ( .B1(n3128), .B2(n3127), .A(n3126), .ZN(n3191) );
  NAND2_X1 U2925 ( .A1(n3680), .A2(n2302), .ZN(n2294) );
  AOI21_X1 U2926 ( .B1(n3680), .B2(n3681), .A(n3682), .ZN(n3750) );
  OAI21_X1 U2927 ( .B1(n3680), .B2(n2298), .A(n2295), .ZN(n3615) );
  NAND2_X1 U2928 ( .A1(n2293), .A2(n2291), .ZN(n3614) );
  NAND2_X1 U2929 ( .A1(n2295), .A2(n2298), .ZN(n2292) );
  NAND2_X1 U2930 ( .A1(n3680), .A2(n2295), .ZN(n2293) );
  INV_X1 U2931 ( .A(n3437), .ZN(n2306) );
  NAND2_X1 U2932 ( .A1(n3437), .A2(n3436), .ZN(n3490) );
  OAI21_X2 U2933 ( .B1(n3632), .B2(n3635), .A(n3633), .ZN(n3510) );
  NAND2_X1 U2934 ( .A1(n3317), .A2(n2319), .ZN(n2318) );
  INV_X1 U2935 ( .A(n3374), .ZN(n2319) );
  INV_X1 U2936 ( .A(n3144), .ZN(n2499) );
  NAND2_X1 U2937 ( .A1(n2343), .A2(n2342), .ZN(n2566) );
  NAND2_X1 U2938 ( .A1(n2531), .A2(n2344), .ZN(n2343) );
  NAND2_X1 U2939 ( .A1(n2347), .A2(n2184), .ZN(n4134) );
  NAND2_X1 U2940 ( .A1(n2731), .A2(n2376), .ZN(n2734) );
  AND2_X1 U2941 ( .A1(n2731), .A2(n2359), .ZN(n2717) );
  NAND2_X1 U2942 ( .A1(n3191), .A2(n3189), .ZN(n3192) );
  NAND2_X1 U2943 ( .A1(n2883), .A2(n2884), .ZN(n2885) );
  NAND2_X1 U2944 ( .A1(n2386), .A2(n4356), .ZN(n2406) );
  AOI21_X2 U2945 ( .B1(n2991), .B2(n2990), .A(n2989), .ZN(n3054) );
  OR2_X1 U2946 ( .A1(n4559), .A2(n2672), .ZN(n2362) );
  AND2_X1 U2947 ( .A1(n3534), .A2(n3533), .ZN(n3741) );
  INV_X1 U2948 ( .A(n3742), .ZN(n3535) );
  NAND2_X1 U2949 ( .A1(n3647), .A2(n3570), .ZN(n3650) );
  NOR2_X1 U2950 ( .A1(n2554), .A2(n3404), .ZN(n2363) );
  NAND2_X1 U2951 ( .A1(n3251), .A2(n3252), .ZN(n2365) );
  AND2_X1 U2952 ( .A1(n3861), .A2(n3787), .ZN(n3448) );
  INV_X1 U2953 ( .A(n3448), .ZN(n2576) );
  NAND2_X1 U2954 ( .A1(n2883), .A2(n2878), .ZN(n2904) );
  INV_X1 U2955 ( .A(n2971), .ZN(n2880) );
  NAND2_X1 U2956 ( .A1(n3535), .A2(n3657), .ZN(n3536) );
  INV_X1 U2957 ( .A(IR_REG_12__SCAN_IN), .ZN(n2366) );
  INV_X1 U2958 ( .A(n3692), .ZN(n3508) );
  INV_X1 U2959 ( .A(n3280), .ZN(n3281) );
  OR2_X1 U2960 ( .A1(n2392), .A2(n2377), .ZN(n2394) );
  NAND2_X1 U2961 ( .A1(n2921), .A2(n2923), .ZN(n2924) );
  AND2_X1 U2962 ( .A1(n4164), .A2(n2704), .ZN(n3867) );
  NAND2_X1 U2963 ( .A1(n3009), .A2(n4487), .ZN(n3820) );
  INV_X1 U2964 ( .A(IR_REG_19__SCAN_IN), .ZN(n2677) );
  INV_X1 U2965 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2464) );
  NOR2_X1 U2966 ( .A1(n2637), .A2(n3715), .ZN(n2644) );
  OAI22_X1 U2967 ( .A1(n2880), .A2(n2873), .B1(n2195), .B2(n2983), .ZN(n2881)
         );
  INV_X1 U2968 ( .A(n3689), .ZN(n3764) );
  AND2_X1 U2969 ( .A1(n3939), .A2(n4245), .ZN(n3798) );
  AND2_X1 U2970 ( .A1(n4040), .A2(n4034), .ZN(n3803) );
  AND2_X1 U2971 ( .A1(n3301), .A2(n3849), .ZN(n3908) );
  AND2_X1 U2972 ( .A1(n3779), .A2(DATAI_20_), .ZN(n4180) );
  INV_X1 U2973 ( .A(n3693), .ZN(n3455) );
  NAND2_X1 U2974 ( .A1(IR_REG_31__SCAN_IN), .A2(n2378), .ZN(n2381) );
  NOR2_X1 U2975 ( .A1(n2465), .A2(n2464), .ZN(n2480) );
  AND2_X1 U2976 ( .A1(n3608), .A2(n3767), .ZN(n3605) );
  INV_X1 U2977 ( .A(n3305), .ZN(n3387) );
  AND3_X1 U2978 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U2979 ( .A1(n2424), .A2(DATAI_0_), .ZN(n2412) );
  OR2_X1 U2980 ( .A1(n2533), .A2(n2532), .ZN(n2547) );
  NOR2_X1 U2981 ( .A1(n2511), .A2(n2510), .ZN(n2521) );
  NOR2_X1 U2982 ( .A1(n2594), .A2(n2593), .ZN(n2613) );
  INV_X1 U2983 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4635) );
  INV_X1 U2984 ( .A(n4294), .ZN(n4475) );
  INV_X1 U2985 ( .A(n4144), .ZN(n4140) );
  INV_X1 U2986 ( .A(n3497), .ZN(n3770) );
  INV_X1 U2987 ( .A(n3251), .ZN(n3296) );
  AND2_X1 U2988 ( .A1(n2151), .A2(n4360), .ZN(n2860) );
  AND2_X1 U2989 ( .A1(n3779), .A2(DATAI_27_), .ZN(n3599) );
  OR2_X1 U2990 ( .A1(n2684), .A2(n4510), .ZN(n4294) );
  AND2_X1 U2991 ( .A1(n2739), .A2(n2772), .ZN(n2778) );
  OR2_X1 U2992 ( .A1(n2497), .A2(IR_REG_9__SCAN_IN), .ZN(n2517) );
  AND2_X1 U2993 ( .A1(n3607), .A2(n3605), .ZN(n3606) );
  XOR2_X1 U2994 ( .A(n3279), .B(n3280), .Z(n3277) );
  INV_X1 U2995 ( .A(n3769), .ZN(n3754) );
  AND3_X1 U2996 ( .A1(n2967), .A2(n2858), .A3(n2857), .ZN(n2898) );
  AND2_X1 U2997 ( .A1(n2669), .A2(n2668), .ZN(n4040) );
  INV_X1 U2998 ( .A(n4221), .ZN(n3744) );
  NAND4_X1 U2999 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n3290)
         );
  OR2_X1 U3000 ( .A1(n2546), .A2(n2585), .ZN(n3170) );
  AND2_X1 U3001 ( .A1(n2790), .A2(n2789), .ZN(n3953) );
  AND2_X1 U3002 ( .A1(n3779), .A2(DATAI_28_), .ZN(n4034) );
  AOI21_X1 U3003 ( .B1(n2778), .B2(n4668), .A(n2782), .ZN(n2858) );
  AND2_X1 U3004 ( .A1(n4174), .A2(n4523), .ZN(n4533) );
  INV_X1 U3005 ( .A(n2871), .ZN(n4516) );
  INV_X1 U3006 ( .A(n4533), .ZN(n4542) );
  AND3_X1 U3007 ( .A1(n2754), .A2(n2753), .A3(n2856), .ZN(n2763) );
  AND2_X1 U3008 ( .A1(n2983), .A2(n2781), .ZN(n2963) );
  AND2_X1 U3009 ( .A1(n2791), .A2(n2790), .ZN(n4450) );
  NAND2_X1 U3010 ( .A1(n2898), .A2(n2890), .ZN(n3762) );
  INV_X1 U3011 ( .A(n3747), .ZN(n3778) );
  INV_X1 U3012 ( .A(n4126), .ZN(n4079) );
  NAND4_X1 U3013 ( .A1(n2572), .A2(n2571), .A3(n2570), .A4(n2569), .ZN(n3942)
         );
  NAND4_X1 U3014 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n3944)
         );
  INV_X1 U3015 ( .A(n4410), .ZN(n4446) );
  NAND2_X1 U3016 ( .A1(n4232), .A2(n3075), .ZN(n4235) );
  NAND2_X1 U3017 ( .A1(n4559), .A2(n4516), .ZN(n4300) );
  NAND2_X1 U3018 ( .A1(n4545), .A2(n4516), .ZN(n4352) );
  INV_X1 U3019 ( .A(n4545), .ZN(n4544) );
  INV_X1 U3020 ( .A(n4493), .ZN(n4494) );
  INV_X1 U3021 ( .A(n2387), .ZN(n4356) );
  AND2_X1 U3022 ( .A1(n2476), .A2(n2484), .ZN(n4364) );
  INV_X1 U3023 ( .A(n3948), .ZN(U4043) );
  NAND2_X1 U3024 ( .A1(n2762), .A2(n2761), .ZN(U3515) );
  NAND3_X1 U3025 ( .A1(n2518), .A2(n2367), .A3(n2366), .ZN(n2368) );
  NAND4_X1 U3026 ( .A1(n4577), .A2(n2583), .A3(n4650), .A4(n2676), .ZN(n2371)
         );
  NAND3_X1 U3027 ( .A1(n4576), .A2(n2677), .A3(n4651), .ZN(n2370) );
  INV_X1 U3028 ( .A(n2431), .ZN(n2374) );
  INV_X1 U3029 ( .A(IR_REG_29__SCAN_IN), .ZN(n2378) );
  OAI21_X1 U3030 ( .B1(n2719), .B2(n2730), .A(IR_REG_29__SCAN_IN), .ZN(n2382)
         );
  NAND2_X1 U3031 ( .A1(n2148), .A2(REG0_REG_22__SCAN_IN), .ZN(n2391) );
  INV_X1 U3032 ( .A(n2386), .ZN(n4355) );
  NAND2_X1 U3033 ( .A1(n4355), .A2(n4356), .ZN(n2384) );
  NAND2_X1 U3034 ( .A1(n2480), .A2(REG3_REG_8__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U3035 ( .A1(n2521), .A2(REG3_REG_12__SCAN_IN), .ZN(n2533) );
  INV_X1 U3036 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2532) );
  INV_X1 U3037 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3639) );
  INV_X1 U3038 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2578) );
  INV_X1 U3039 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2593) );
  AND2_X1 U3040 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2385) );
  XNOR2_X1 U3041 ( .A(n2630), .B(REG3_REG_22__SCAN_IN), .ZN(n4145) );
  NAND2_X1 U3042 ( .A1(n2420), .A2(n4145), .ZN(n2390) );
  NAND2_X1 U3043 ( .A1(n2721), .A2(REG1_REG_22__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U3044 ( .A1(n2146), .A2(REG2_REG_22__SCAN_IN), .ZN(n2388) );
  NAND4_X1 U3045 ( .A1(n2391), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n4152)
         );
  NAND2_X1 U3046 ( .A1(n2392), .A2(n2395), .ZN(n2393) );
  NAND2_X1 U3047 ( .A1(n2395), .A2(IR_REG_27__SCAN_IN), .ZN(n2396) );
  NAND2_X2 U3048 ( .A1(n2397), .A2(n2396), .ZN(n2424) );
  NAND2_X1 U3049 ( .A1(n2420), .A2(REG3_REG_1__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U3050 ( .A1(n2417), .A2(REG2_REG_1__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3051 ( .A1(n2416), .A2(REG0_REG_1__SCAN_IN), .ZN(n2402) );
  NAND2_X1 U3052 ( .A1(n2721), .A2(REG1_REG_1__SCAN_IN), .ZN(n2404) );
  INV_X1 U3053 ( .A(n2793), .ZN(n4370) );
  NAND4_X1 U3054 ( .A1(n2405), .A2(n2404), .A3(n2403), .A4(n2402), .ZN(n2875)
         );
  NAND2_X1 U3055 ( .A1(n2875), .A2(n3040), .ZN(n3816) );
  NAND2_X1 U3056 ( .A1(n2721), .A2(REG1_REG_0__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3057 ( .A1(n2420), .A2(REG3_REG_0__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U3058 ( .A1(n2146), .A2(REG2_REG_0__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U3059 ( .A1(n2147), .A2(REG0_REG_0__SCAN_IN), .ZN(n2407) );
  INV_X1 U3060 ( .A(n2424), .ZN(n2411) );
  AND2_X1 U3061 ( .A1(n3949), .A2(n2971), .ZN(n3031) );
  NAND2_X1 U3062 ( .A1(n2686), .A2(n3031), .ZN(n3033) );
  INV_X1 U3063 ( .A(n2973), .ZN(n2414) );
  NAND2_X1 U3064 ( .A1(n2414), .A2(n3034), .ZN(n2415) );
  NAND2_X1 U3065 ( .A1(n2147), .A2(REG0_REG_2__SCAN_IN), .ZN(n2419) );
  NAND2_X1 U3066 ( .A1(n2146), .A2(REG2_REG_2__SCAN_IN), .ZN(n2418) );
  AND2_X1 U3067 ( .A1(n2419), .A2(n2418), .ZN(n2423) );
  NAND2_X1 U3068 ( .A1(n2721), .A2(REG1_REG_2__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3069 ( .A1(n2420), .A2(REG3_REG_2__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U3070 ( .A1(n3035), .A2(n2929), .ZN(n3823) );
  NAND2_X1 U3071 ( .A1(n3009), .A2(n2929), .ZN(n2426) );
  NAND2_X1 U3072 ( .A1(n4470), .A2(n2426), .ZN(n3003) );
  NAND2_X1 U3073 ( .A1(n2148), .A2(REG0_REG_3__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3074 ( .A1(n2420), .A2(n4638), .ZN(n2429) );
  NAND2_X1 U3075 ( .A1(n2721), .A2(REG1_REG_3__SCAN_IN), .ZN(n2428) );
  NAND2_X1 U3076 ( .A1(n2146), .A2(REG2_REG_3__SCAN_IN), .ZN(n2427) );
  NAND2_X1 U3077 ( .A1(n2433), .A2(n2432), .ZN(n2443) );
  OR2_X1 U3078 ( .A1(n2433), .A2(n2432), .ZN(n2434) );
  MUX2_X1 U3079 ( .A(n4368), .B(DATAI_3_), .S(n3779), .Z(n3012) );
  NAND2_X1 U3080 ( .A1(n2992), .A2(n3012), .ZN(n2435) );
  NAND2_X1 U3081 ( .A1(n3003), .A2(n2435), .ZN(n2437) );
  INV_X1 U3082 ( .A(n3012), .ZN(n2998) );
  NAND2_X1 U3083 ( .A1(n4480), .A2(n2998), .ZN(n2436) );
  NAND2_X1 U3084 ( .A1(n2148), .A2(REG0_REG_4__SCAN_IN), .ZN(n2442) );
  INV_X1 U3085 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2438) );
  XNOR2_X1 U3086 ( .A(n2438), .B(REG3_REG_3__SCAN_IN), .ZN(n3060) );
  NAND2_X1 U3087 ( .A1(n2420), .A2(n3060), .ZN(n2441) );
  NAND2_X1 U3088 ( .A1(n2146), .A2(REG2_REG_4__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U3089 ( .A1(n2721), .A2(REG1_REG_4__SCAN_IN), .ZN(n2439) );
  INV_X1 U3090 ( .A(n3088), .ZN(n2997) );
  NAND2_X1 U3091 ( .A1(n2443), .A2(IR_REG_31__SCAN_IN), .ZN(n2444) );
  XNOR2_X1 U3092 ( .A(n2444), .B(IR_REG_4__SCAN_IN), .ZN(n4367) );
  MUX2_X1 U3093 ( .A(n4367), .B(DATAI_4_), .S(n3779), .Z(n3050) );
  NAND2_X1 U3094 ( .A1(n2997), .A2(n3050), .ZN(n3826) );
  NAND2_X1 U3095 ( .A1(n3088), .A2(n3020), .ZN(n3829) );
  AOI22_X1 U3096 ( .A1(n2147), .A2(REG0_REG_5__SCAN_IN), .B1(n2721), .B2(
        REG1_REG_5__SCAN_IN), .ZN(n2447) );
  AOI21_X1 U3097 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2445) );
  NOR2_X1 U3098 ( .A1(n2445), .A2(n2456), .ZN(n3068) );
  AOI22_X1 U3099 ( .A1(n2420), .A2(n3068), .B1(n2146), .B2(REG2_REG_5__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3100 ( .A1(n2448), .A2(IR_REG_31__SCAN_IN), .ZN(n2449) );
  XNOR2_X1 U3101 ( .A(n2449), .B(n2321), .ZN(n2832) );
  INV_X1 U3102 ( .A(DATAI_5_), .ZN(n2450) );
  MUX2_X1 U3103 ( .A(n2832), .B(n2450), .S(n3779), .Z(n3117) );
  AND2_X1 U3104 ( .A1(n3083), .A2(n3117), .ZN(n2453) );
  OR2_X1 U3105 ( .A1(n3905), .A2(n2453), .ZN(n2455) );
  NAND2_X1 U3106 ( .A1(n3088), .A2(n3050), .ZN(n3071) );
  INV_X1 U3107 ( .A(n3117), .ZN(n3067) );
  NAND2_X1 U3108 ( .A1(n3132), .A2(n3067), .ZN(n2451) );
  AND2_X1 U3109 ( .A1(n3071), .A2(n2451), .ZN(n2452) );
  OR2_X1 U3110 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  OAI21_X1 U3111 ( .B1(n3018), .B2(n2455), .A(n2454), .ZN(n3094) );
  NAND2_X1 U3112 ( .A1(n2147), .A2(REG0_REG_6__SCAN_IN), .ZN(n2461) );
  OAI21_X1 U3113 ( .B1(n2456), .B2(REG3_REG_6__SCAN_IN), .A(n2465), .ZN(n2457)
         );
  INV_X1 U3114 ( .A(n2457), .ZN(n3137) );
  NAND2_X1 U3115 ( .A1(n2420), .A2(n3137), .ZN(n2460) );
  NAND2_X1 U3116 ( .A1(n2146), .A2(REG2_REG_6__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U3117 ( .A1(n2721), .A2(REG1_REG_6__SCAN_IN), .ZN(n2458) );
  NAND4_X1 U3118 ( .A1(n2461), .A2(n2460), .A3(n2459), .A4(n2458), .ZN(n3947)
         );
  OR2_X1 U3119 ( .A1(n2472), .A2(n2730), .ZN(n2462) );
  XNOR2_X1 U3120 ( .A(n2462), .B(IR_REG_6__SCAN_IN), .ZN(n4365) );
  MUX2_X1 U3121 ( .A(n4365), .B(DATAI_6_), .S(n3779), .Z(n3133) );
  AND2_X1 U3122 ( .A1(n3947), .A2(n3133), .ZN(n2463) );
  OAI22_X1 U3123 ( .A1(n3094), .A2(n2463), .B1(n3133), .B2(n3947), .ZN(n3110)
         );
  INV_X1 U3124 ( .A(n3110), .ZN(n2478) );
  NAND2_X1 U3125 ( .A1(n2148), .A2(REG0_REG_7__SCAN_IN), .ZN(n2470) );
  AND2_X1 U3126 ( .A1(n2465), .A2(n2464), .ZN(n2466) );
  NOR2_X1 U3127 ( .A1(n2480), .A2(n2466), .ZN(n3218) );
  NAND2_X1 U3128 ( .A1(n2420), .A2(n3218), .ZN(n2469) );
  NAND2_X1 U3129 ( .A1(n2146), .A2(REG2_REG_7__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U3130 ( .A1(n2721), .A2(REG1_REG_7__SCAN_IN), .ZN(n2467) );
  NAND4_X1 U3131 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), .ZN(n3946)
         );
  INV_X1 U3132 ( .A(n3946), .ZN(n3209) );
  NOR2_X1 U3133 ( .A1(n2262), .A2(n2730), .ZN(n2473) );
  NAND2_X1 U3134 ( .A1(n2473), .A2(IR_REG_7__SCAN_IN), .ZN(n2476) );
  INV_X1 U3135 ( .A(n2473), .ZN(n2475) );
  INV_X1 U3136 ( .A(IR_REG_7__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3137 ( .A1(n2475), .A2(n2474), .ZN(n2484) );
  MUX2_X1 U3138 ( .A(n4364), .B(DATAI_7_), .S(n3779), .Z(n3197) );
  NAND2_X1 U3139 ( .A1(n3209), .A2(n3197), .ZN(n2691) );
  INV_X1 U3140 ( .A(n3197), .ZN(n3215) );
  NAND2_X1 U3141 ( .A1(n3946), .A2(n3215), .ZN(n3834) );
  NAND2_X1 U3142 ( .A1(n2478), .A2(n2477), .ZN(n4537) );
  NAND2_X1 U3143 ( .A1(n3946), .A2(n3197), .ZN(n2479) );
  AOI22_X1 U3144 ( .A1(n2147), .A2(REG0_REG_8__SCAN_IN), .B1(n2721), .B2(
        REG1_REG_8__SCAN_IN), .ZN(n2483) );
  OR2_X1 U3145 ( .A1(n2480), .A2(REG3_REG_8__SCAN_IN), .ZN(n2481) );
  AND2_X1 U3146 ( .A1(n2490), .A2(n2481), .ZN(n4458) );
  AOI22_X1 U3147 ( .A1(n2420), .A2(n4458), .B1(n2146), .B2(REG2_REG_8__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U31480 ( .A1(n2484), .A2(IR_REG_31__SCAN_IN), .ZN(n2486) );
  INV_X1 U31490 ( .A(IR_REG_8__SCAN_IN), .ZN(n2485) );
  XNOR2_X1 U3150 ( .A(n2486), .B(n2485), .ZN(n3174) );
  INV_X1 U3151 ( .A(DATAI_8_), .ZN(n2487) );
  MUX2_X1 U3152 ( .A(n3174), .B(n2487), .S(n3779), .Z(n3233) );
  INV_X1 U3153 ( .A(n3256), .ZN(n3945) );
  INV_X1 U3154 ( .A(n3233), .ZN(n3238) );
  NAND2_X1 U3155 ( .A1(n3945), .A2(n3238), .ZN(n2488) );
  NAND2_X1 U3156 ( .A1(n2148), .A2(REG0_REG_9__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3157 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  AND2_X1 U3158 ( .A1(n2502), .A2(n2491), .ZN(n3259) );
  NAND2_X1 U3159 ( .A1(n2420), .A2(n3259), .ZN(n2494) );
  NAND2_X1 U3160 ( .A1(n2146), .A2(REG2_REG_9__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3161 ( .A1(n2721), .A2(REG1_REG_9__SCAN_IN), .ZN(n2492) );
  NAND4_X1 U3162 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n3251)
         );
  NAND2_X1 U3163 ( .A1(n2262), .A2(n2539), .ZN(n2497) );
  MUX2_X1 U3164 ( .A(IR_REG_31__SCAN_IN), .B(n2496), .S(IR_REG_9__SCAN_IN), 
        .Z(n2498) );
  MUX2_X1 U3165 ( .A(n3173), .B(DATAI_9_), .S(n3779), .Z(n3252) );
  NAND2_X1 U3166 ( .A1(n2499), .A2(n2365), .ZN(n2501) );
  NAND2_X1 U3167 ( .A1(n3296), .A2(n3257), .ZN(n2500) );
  NAND2_X1 U3168 ( .A1(n2148), .A2(REG0_REG_10__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3169 ( .A1(n2502), .A2(n4635), .ZN(n2503) );
  AND2_X1 U3170 ( .A1(n2511), .A2(n2503), .ZN(n3276) );
  NAND2_X1 U3171 ( .A1(n2420), .A2(n3276), .ZN(n2506) );
  NAND2_X1 U3172 ( .A1(n2721), .A2(REG1_REG_10__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U3173 ( .A1(n2146), .A2(REG2_REG_10__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U3174 ( .A1(n2517), .A2(IR_REG_31__SCAN_IN), .ZN(n2508) );
  XNOR2_X1 U3175 ( .A(n2508), .B(IR_REG_10__SCAN_IN), .ZN(n4506) );
  MUX2_X1 U3176 ( .A(n4506), .B(DATAI_10_), .S(n3779), .Z(n3288) );
  NOR2_X1 U3177 ( .A1(n3290), .A2(n3288), .ZN(n2509) );
  INV_X1 U3178 ( .A(n3288), .ZN(n3346) );
  NAND2_X1 U3179 ( .A1(n2147), .A2(REG0_REG_11__SCAN_IN), .ZN(n2516) );
  AND2_X1 U3180 ( .A1(n2511), .A2(n2510), .ZN(n2512) );
  NOR2_X1 U3181 ( .A1(n2521), .A2(n2512), .ZN(n3323) );
  NAND2_X1 U3182 ( .A1(n2420), .A2(n3323), .ZN(n2515) );
  NAND2_X1 U3183 ( .A1(n2721), .A2(REG1_REG_11__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U3184 ( .A1(n2146), .A2(REG2_REG_11__SCAN_IN), .ZN(n2513) );
  NAND4_X1 U3185 ( .A1(n2516), .A2(n2515), .A3(n2514), .A4(n2513), .ZN(n3305)
         );
  OR2_X1 U3186 ( .A1(n2519), .A2(n2518), .ZN(n2520) );
  NAND2_X1 U3187 ( .A1(n2519), .A2(n2518), .ZN(n2527) );
  MUX2_X1 U3188 ( .A(n3172), .B(DATAI_11_), .S(n3779), .Z(n3271) );
  NAND2_X1 U3189 ( .A1(n3387), .A2(n3271), .ZN(n3301) );
  NAND2_X1 U3190 ( .A1(n3305), .A2(n3357), .ZN(n3849) );
  NAND2_X1 U3191 ( .A1(n2147), .A2(REG0_REG_12__SCAN_IN), .ZN(n2526) );
  OR2_X1 U3192 ( .A1(n2521), .A2(REG3_REG_12__SCAN_IN), .ZN(n2522) );
  AND2_X1 U3193 ( .A1(n2522), .A2(n2533), .ZN(n3390) );
  NAND2_X1 U3194 ( .A1(n2420), .A2(n3390), .ZN(n2525) );
  NAND2_X1 U3195 ( .A1(n2146), .A2(REG2_REG_12__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U3196 ( .A1(n2721), .A2(REG1_REG_12__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U3197 ( .A1(n2527), .A2(IR_REG_31__SCAN_IN), .ZN(n2528) );
  XNOR2_X1 U3198 ( .A(n2528), .B(IR_REG_12__SCAN_IN), .ZN(n3181) );
  MUX2_X1 U3199 ( .A(n3181), .B(DATAI_12_), .S(n3779), .Z(n3379) );
  NAND2_X1 U3200 ( .A1(n3944), .A2(n3379), .ZN(n2529) );
  NAND2_X1 U3201 ( .A1(n3308), .A2(n2529), .ZN(n2531) );
  NAND2_X1 U3202 ( .A1(n3338), .A2(n3388), .ZN(n2530) );
  NAND2_X1 U3203 ( .A1(n2148), .A2(REG0_REG_13__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U3204 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  AND2_X1 U3205 ( .A1(n2547), .A2(n2534), .ZN(n3444) );
  NAND2_X1 U3206 ( .A1(n2420), .A2(n3444), .ZN(n2537) );
  NAND2_X1 U3207 ( .A1(n2721), .A2(REG1_REG_13__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U3208 ( .A1(n2146), .A2(REG2_REG_13__SCAN_IN), .ZN(n2535) );
  NAND4_X1 U3209 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), .ZN(n3637)
         );
  AND2_X1 U32100 ( .A1(n2262), .A2(n2539), .ZN(n2541) );
  AND2_X1 U32110 ( .A1(n2541), .A2(n2540), .ZN(n2542) );
  NOR2_X1 U32120 ( .A1(n2542), .A2(n2730), .ZN(n2543) );
  MUX2_X1 U32130 ( .A(n2730), .B(n2543), .S(IR_REG_13__SCAN_IN), .Z(n2546) );
  INV_X1 U32140 ( .A(n3170), .ZN(n2769) );
  MUX2_X1 U32150 ( .A(n2769), .B(DATAI_13_), .S(n3779), .Z(n3439) );
  NOR2_X1 U32160 ( .A1(n3637), .A2(n3439), .ZN(n3401) );
  NAND2_X1 U32170 ( .A1(n2148), .A2(REG0_REG_14__SCAN_IN), .ZN(n2552) );
  AND2_X1 U32180 ( .A1(n2547), .A2(n3639), .ZN(n2548) );
  NOR2_X1 U32190 ( .A1(n2555), .A2(n2548), .ZN(n3644) );
  NAND2_X1 U32200 ( .A1(n2420), .A2(n3644), .ZN(n2551) );
  NAND2_X1 U32210 ( .A1(n2721), .A2(REG1_REG_14__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32220 ( .A1(n2146), .A2(REG2_REG_14__SCAN_IN), .ZN(n2549) );
  NAND4_X1 U32230 ( .A1(n2552), .A2(n2551), .A3(n2550), .A4(n2549), .ZN(n3497)
         );
  INV_X1 U32240 ( .A(n2585), .ZN(n2561) );
  XNOR2_X1 U32250 ( .A(n2553), .B(IR_REG_14__SCAN_IN), .ZN(n4501) );
  MUX2_X1 U32260 ( .A(n4501), .B(DATAI_14_), .S(n3779), .Z(n3638) );
  INV_X1 U32270 ( .A(n3638), .ZN(n3461) );
  AND2_X1 U32280 ( .A1(n3770), .A2(n3461), .ZN(n2554) );
  NAND2_X1 U32290 ( .A1(n3770), .A2(n3638), .ZN(n3781) );
  NAND2_X1 U32300 ( .A1(n3497), .A2(n3461), .ZN(n3782) );
  NAND2_X1 U32310 ( .A1(n3781), .A2(n3782), .ZN(n3916) );
  NAND2_X1 U32320 ( .A1(n3637), .A2(n3439), .ZN(n3403) );
  AND2_X1 U32330 ( .A1(n3916), .A2(n3403), .ZN(n3404) );
  NAND2_X1 U32340 ( .A1(n2147), .A2(REG0_REG_15__SCAN_IN), .ZN(n2560) );
  NOR2_X1 U32350 ( .A1(n2555), .A2(REG3_REG_15__SCAN_IN), .ZN(n2556) );
  OR2_X1 U32360 ( .A1(n2567), .A2(n2556), .ZN(n3777) );
  INV_X1 U32370 ( .A(n3777), .ZN(n3429) );
  NAND2_X1 U32380 ( .A1(n2420), .A2(n3429), .ZN(n2559) );
  NAND2_X1 U32390 ( .A1(n2146), .A2(REG2_REG_15__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U32400 ( .A1(n2721), .A2(REG1_REG_15__SCAN_IN), .ZN(n2557) );
  NAND4_X1 U32410 ( .A1(n2560), .A2(n2559), .A3(n2558), .A4(n2557), .ZN(n3943)
         );
  NAND2_X1 U32420 ( .A1(n2562), .A2(IR_REG_31__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32430 ( .A1(n2563), .A2(n2583), .ZN(n2573) );
  OR2_X1 U32440 ( .A1(n2563), .A2(n2583), .ZN(n2564) );
  MUX2_X1 U32450 ( .A(n3986), .B(DATAI_15_), .S(n2424), .Z(n3511) );
  INV_X1 U32460 ( .A(n3511), .ZN(n3771) );
  NAND2_X1 U32470 ( .A1(n3696), .A2(n3771), .ZN(n2565) );
  NAND2_X1 U32480 ( .A1(n2148), .A2(REG0_REG_16__SCAN_IN), .ZN(n2572) );
  OR2_X1 U32490 ( .A1(n2567), .A2(REG3_REG_16__SCAN_IN), .ZN(n2568) );
  AND2_X1 U32500 ( .A1(n2579), .A2(n2568), .ZN(n3698) );
  NAND2_X1 U32510 ( .A1(n2420), .A2(n3698), .ZN(n2571) );
  NAND2_X1 U32520 ( .A1(n2146), .A2(REG2_REG_16__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U32530 ( .A1(n2721), .A2(REG1_REG_16__SCAN_IN), .ZN(n2569) );
  INV_X1 U32540 ( .A(n3942), .ZN(n2575) );
  NAND2_X1 U32550 ( .A1(n2573), .A2(IR_REG_31__SCAN_IN), .ZN(n2574) );
  XNOR2_X1 U32560 ( .A(n2574), .B(IR_REG_16__SCAN_IN), .ZN(n3987) );
  MUX2_X1 U32570 ( .A(n3987), .B(DATAI_16_), .S(n2424), .Z(n3693) );
  NAND2_X1 U32580 ( .A1(n2575), .A2(n3693), .ZN(n3861) );
  NAND2_X1 U32590 ( .A1(n3942), .A2(n3455), .ZN(n3787) );
  NAND2_X1 U32600 ( .A1(n3942), .A2(n3693), .ZN(n2577) );
  AOI22_X1 U32610 ( .A1(n2148), .A2(REG0_REG_17__SCAN_IN), .B1(n2721), .B2(
        REG1_REG_17__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U32620 ( .A1(n2579), .A2(n2578), .ZN(n2580) );
  AND2_X1 U32630 ( .A1(n2594), .A2(n2580), .ZN(n3706) );
  AOI22_X1 U32640 ( .A1(n2420), .A2(n3706), .B1(n2146), .B2(
        REG2_REG_17__SCAN_IN), .ZN(n2581) );
  NOR2_X1 U32650 ( .A1(n2589), .A2(n2730), .ZN(n2586) );
  MUX2_X1 U32660 ( .A(n2730), .B(n2586), .S(IR_REG_17__SCAN_IN), .Z(n2587) );
  INV_X1 U32670 ( .A(n2587), .ZN(n2590) );
  NAND2_X1 U32680 ( .A1(n2589), .A2(n2588), .ZN(n2606) );
  NAND2_X1 U32690 ( .A1(n2590), .A2(n2606), .ZN(n3993) );
  INV_X1 U32700 ( .A(DATAI_17_), .ZN(n4616) );
  MUX2_X1 U32710 ( .A(n3993), .B(n4616), .S(n2424), .Z(n4295) );
  NAND2_X1 U32720 ( .A1(n4221), .A2(n4295), .ZN(n2592) );
  AND2_X1 U32730 ( .A1(n3744), .A2(n2757), .ZN(n2591) );
  NAND2_X1 U32740 ( .A1(n2148), .A2(REG0_REG_18__SCAN_IN), .ZN(n2599) );
  AND2_X1 U32750 ( .A1(n2594), .A2(n2593), .ZN(n2595) );
  NOR2_X1 U32760 ( .A1(n2613), .A2(n2595), .ZN(n4228) );
  NAND2_X1 U32770 ( .A1(n2420), .A2(n4228), .ZN(n2598) );
  NAND2_X1 U32780 ( .A1(n2721), .A2(REG1_REG_18__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U32790 ( .A1(n2146), .A2(REG2_REG_18__SCAN_IN), .ZN(n2596) );
  NAND4_X1 U32800 ( .A1(n2599), .A2(n2598), .A3(n2597), .A4(n2596), .ZN(n3941)
         );
  INV_X1 U32810 ( .A(n3941), .ZN(n4202) );
  NAND2_X1 U32820 ( .A1(n2606), .A2(IR_REG_31__SCAN_IN), .ZN(n2600) );
  XNOR2_X1 U32830 ( .A(n2600), .B(IR_REG_18__SCAN_IN), .ZN(n4003) );
  MUX2_X1 U32840 ( .A(n4003), .B(DATAI_18_), .S(n3779), .Z(n4216) );
  NAND2_X1 U32850 ( .A1(n4202), .A2(n4216), .ZN(n4193) );
  INV_X1 U32860 ( .A(n4216), .ZN(n4226) );
  NAND2_X1 U32870 ( .A1(n3941), .A2(n4226), .ZN(n4191) );
  NAND2_X1 U32880 ( .A1(n4193), .A2(n4191), .ZN(n4214) );
  NAND2_X1 U32890 ( .A1(n4202), .A2(n4226), .ZN(n4186) );
  NAND2_X1 U32900 ( .A1(n2147), .A2(REG0_REG_19__SCAN_IN), .ZN(n2605) );
  INV_X1 U32910 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2601) );
  XNOR2_X1 U32920 ( .A(n2613), .B(n2601), .ZN(n4205) );
  NAND2_X1 U32930 ( .A1(n2420), .A2(n4205), .ZN(n2604) );
  NAND2_X1 U32940 ( .A1(n2146), .A2(REG2_REG_19__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U32950 ( .A1(n2721), .A2(REG1_REG_19__SCAN_IN), .ZN(n2602) );
  NAND4_X1 U32960 ( .A1(n2605), .A2(n2604), .A3(n2603), .A4(n2602), .ZN(n4218)
         );
  INV_X1 U32970 ( .A(n4218), .ZN(n4169) );
  INV_X1 U32980 ( .A(n2606), .ZN(n2607) );
  INV_X1 U32990 ( .A(n2608), .ZN(n2609) );
  NAND2_X1 U33000 ( .A1(n2609), .A2(IR_REG_19__SCAN_IN), .ZN(n2610) );
  MUX2_X1 U33010 ( .A(n4362), .B(DATAI_19_), .S(n2424), .Z(n4198) );
  INV_X1 U33020 ( .A(n4198), .ZN(n4203) );
  NAND2_X1 U33030 ( .A1(n4169), .A2(n4203), .ZN(n2611) );
  AND2_X1 U33040 ( .A1(n4186), .A2(n2611), .ZN(n2612) );
  NAND2_X1 U33050 ( .A1(n4211), .A2(n2612), .ZN(n4171) );
  NAND2_X1 U33060 ( .A1(n4218), .A2(n4198), .ZN(n4170) );
  NAND2_X1 U33070 ( .A1(n2148), .A2(REG0_REG_20__SCAN_IN), .ZN(n2618) );
  AOI21_X1 U33080 ( .B1(n2613), .B2(REG3_REG_19__SCAN_IN), .A(
        REG3_REG_20__SCAN_IN), .ZN(n2614) );
  NOR2_X1 U33090 ( .A1(n2621), .A2(n2614), .ZN(n4178) );
  NAND2_X1 U33100 ( .A1(n2420), .A2(n4178), .ZN(n2617) );
  NAND2_X1 U33110 ( .A1(n2721), .A2(REG1_REG_20__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U33120 ( .A1(n2146), .A2(REG2_REG_20__SCAN_IN), .ZN(n2615) );
  NAND4_X1 U33130 ( .A1(n2618), .A2(n2617), .A3(n2616), .A4(n2615), .ZN(n4199)
         );
  NAND2_X1 U33140 ( .A1(n4199), .A2(n4180), .ZN(n3898) );
  AND2_X1 U33150 ( .A1(n4170), .A2(n3898), .ZN(n2619) );
  NAND2_X1 U33160 ( .A1(n4171), .A2(n2619), .ZN(n2620) );
  INV_X1 U33170 ( .A(n4199), .ZN(n3675) );
  NAND2_X1 U33180 ( .A1(n3675), .A2(n3727), .ZN(n3899) );
  NAND2_X1 U33190 ( .A1(n2147), .A2(REG0_REG_21__SCAN_IN), .ZN(n2626) );
  OR2_X1 U33200 ( .A1(n2621), .A2(REG3_REG_21__SCAN_IN), .ZN(n2622) );
  AND2_X1 U33210 ( .A1(n2630), .A2(n2622), .ZN(n4157) );
  NAND2_X1 U33220 ( .A1(n2420), .A2(n4157), .ZN(n2625) );
  NAND2_X1 U33230 ( .A1(n2146), .A2(REG2_REG_21__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U33240 ( .A1(n2721), .A2(REG1_REG_21__SCAN_IN), .ZN(n2623) );
  NAND4_X1 U33250 ( .A1(n2626), .A2(n2625), .A3(n2624), .A4(n2623), .ZN(n4167)
         );
  NAND2_X1 U33260 ( .A1(n4167), .A2(n3555), .ZN(n2627) );
  INV_X1 U33270 ( .A(n4167), .ZN(n3736) );
  NAND2_X1 U33280 ( .A1(n3736), .A2(n4277), .ZN(n2628) );
  NAND2_X1 U33290 ( .A1(n3674), .A2(n4144), .ZN(n4119) );
  NAND2_X1 U33300 ( .A1(n4152), .A2(n4140), .ZN(n2708) );
  OAI21_X1 U33310 ( .B1(n3674), .B2(n4140), .A(n4134), .ZN(n4110) );
  NAND2_X1 U33320 ( .A1(n2147), .A2(REG0_REG_23__SCAN_IN), .ZN(n2635) );
  INV_X1 U33330 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3735) );
  INV_X1 U33340 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4636) );
  OAI21_X1 U33350 ( .B1(n2630), .B2(n3735), .A(n4636), .ZN(n2631) );
  AND2_X1 U33360 ( .A1(n2631), .A2(n2637), .ZN(n4113) );
  NAND2_X1 U33370 ( .A1(n2420), .A2(n4113), .ZN(n2634) );
  NAND2_X1 U33380 ( .A1(n2721), .A2(REG1_REG_23__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U33390 ( .A1(n2146), .A2(REG2_REG_23__SCAN_IN), .ZN(n2632) );
  NAND4_X1 U33400 ( .A1(n2635), .A2(n2634), .A3(n2633), .A4(n2632), .ZN(n4137)
         );
  INV_X1 U33410 ( .A(n4137), .ZN(n4097) );
  NAND2_X1 U33420 ( .A1(n2424), .A2(DATAI_23_), .ZN(n4123) );
  NAND2_X1 U33430 ( .A1(n4097), .A2(n4123), .ZN(n2636) );
  INV_X1 U33440 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3715) );
  AND2_X1 U33450 ( .A1(n2637), .A2(n3715), .ZN(n2638) );
  OR2_X1 U33460 ( .A1(n2638), .A2(n2644), .ZN(n3714) );
  NAND2_X1 U33470 ( .A1(n2721), .A2(REG1_REG_24__SCAN_IN), .ZN(n2639) );
  OAI21_X1 U33480 ( .B1(n3714), .B2(n2384), .A(n2639), .ZN(n2640) );
  INV_X1 U33490 ( .A(n2640), .ZN(n2642) );
  AOI22_X1 U33500 ( .A1(n2147), .A2(REG0_REG_24__SCAN_IN), .B1(n2146), .B2(
        REG2_REG_24__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U33510 ( .A1(n4079), .A2(n3575), .ZN(n2643) );
  NOR2_X1 U33520 ( .A1(n2644), .A2(REG3_REG_25__SCAN_IN), .ZN(n2645) );
  OR2_X1 U3353 ( .A1(n2649), .A2(n2645), .ZN(n3684) );
  AOI22_X1 U33540 ( .A1(n2148), .A2(REG0_REG_25__SCAN_IN), .B1(n2721), .B2(
        REG1_REG_25__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U3355 ( .A1(n2146), .A2(REG2_REG_25__SCAN_IN), .ZN(n2646) );
  INV_X1 U3356 ( .A(n4095), .ZN(n3716) );
  NAND2_X1 U3357 ( .A1(n2424), .A2(DATAI_25_), .ZN(n4084) );
  NAND2_X1 U3358 ( .A1(n3716), .A2(n4084), .ZN(n2648) );
  INV_X1 U3359 ( .A(n4084), .ZN(n4078) );
  NOR2_X1 U3360 ( .A1(n2649), .A2(REG3_REG_26__SCAN_IN), .ZN(n2650) );
  AOI22_X1 U3361 ( .A1(n2148), .A2(REG0_REG_26__SCAN_IN), .B1(n2721), .B2(
        REG1_REG_26__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U3362 ( .A1(n2146), .A2(REG2_REG_26__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U3363 ( .A1(n2424), .A2(DATAI_26_), .ZN(n4066) );
  INV_X1 U3364 ( .A(n4066), .ZN(n4061) );
  NAND2_X1 U3365 ( .A1(n4038), .A2(n4061), .ZN(n2653) );
  INV_X1 U3366 ( .A(n4038), .ZN(n4082) );
  INV_X1 U3367 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3627) );
  XNOR2_X1 U3368 ( .A(n2661), .B(n3627), .ZN(n4048) );
  NAND2_X1 U3369 ( .A1(n4048), .A2(n2420), .ZN(n2658) );
  INV_X1 U3370 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4316) );
  NAND2_X1 U3371 ( .A1(n2146), .A2(REG2_REG_27__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3372 ( .A1(n2721), .A2(REG1_REG_27__SCAN_IN), .ZN(n2654) );
  OAI211_X1 U3373 ( .C1(n2820), .C2(n4316), .A(n2655), .B(n2654), .ZN(n2656)
         );
  INV_X1 U3374 ( .A(n2656), .ZN(n2657) );
  INV_X1 U3375 ( .A(n3599), .ZN(n4249) );
  NAND2_X1 U3376 ( .A1(n4064), .A2(n4249), .ZN(n2659) );
  INV_X1 U3377 ( .A(n4064), .ZN(n3940) );
  AND2_X1 U3378 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2660) );
  NAND2_X1 U3379 ( .A1(n2661), .A2(n2660), .ZN(n3618) );
  INV_X1 U3380 ( .A(n2661), .ZN(n2663) );
  INV_X1 U3381 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2662) );
  OAI21_X1 U3382 ( .B1(n2663), .B2(n3627), .A(n2662), .ZN(n2664) );
  NAND2_X1 U3383 ( .A1(n3618), .A2(n2664), .ZN(n4028) );
  INV_X1 U3384 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U3385 ( .A1(n2146), .A2(REG2_REG_28__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3386 ( .A1(n2721), .A2(REG1_REG_28__SCAN_IN), .ZN(n2665) );
  OAI211_X1 U3387 ( .C1(n2820), .C2(n4735), .A(n2666), .B(n2665), .ZN(n2667)
         );
  INV_X1 U3388 ( .A(n2667), .ZN(n2668) );
  INV_X1 U3389 ( .A(n4040), .ZN(n3939) );
  OAI22_X1 U3390 ( .A1(n4026), .A2(n4027), .B1(n4040), .B2(n4245), .ZN(n2673)
         );
  INV_X1 U3391 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2672) );
  OR2_X1 U3392 ( .A1(n3618), .A2(n2384), .ZN(n2671) );
  AOI22_X1 U3393 ( .A1(n2146), .A2(REG2_REG_29__SCAN_IN), .B1(n2147), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n2670) );
  OAI211_X1 U3394 ( .C1(n2672), .C2(n2406), .A(n2671), .B(n2670), .ZN(n3797)
         );
  NAND2_X1 U3395 ( .A1(n2424), .A2(DATAI_29_), .ZN(n3795) );
  XNOR2_X1 U3396 ( .A(n3797), .B(n3795), .ZN(n3903) );
  XNOR2_X1 U3397 ( .A(n2673), .B(n3903), .ZN(n3624) );
  NAND2_X1 U3398 ( .A1(n2677), .A2(n2676), .ZN(n2678) );
  NAND2_X1 U3399 ( .A1(n2681), .A2(IR_REG_31__SCAN_IN), .ZN(n2682) );
  XNOR2_X1 U3400 ( .A(n2868), .B(n4360), .ZN(n2683) );
  NAND2_X1 U3401 ( .A1(n2683), .A2(n4010), .ZN(n4174) );
  NOR2_X1 U3402 ( .A1(n4010), .A2(n4360), .ZN(n2685) );
  NAND2_X1 U3403 ( .A1(n2684), .A2(n2685), .ZN(n4523) );
  NAND2_X1 U3404 ( .A1(n4472), .A2(n4473), .ZN(n4471) );
  NAND2_X1 U3405 ( .A1(n4471), .A2(n3820), .ZN(n3005) );
  NAND2_X1 U3406 ( .A1(n4480), .A2(n3012), .ZN(n3825) );
  NAND2_X1 U3407 ( .A1(n2992), .A2(n2998), .ZN(n3822) );
  AND2_X1 U3408 ( .A1(n3825), .A2(n3822), .ZN(n3004) );
  NAND2_X1 U3409 ( .A1(n3005), .A2(n3004), .ZN(n2687) );
  NAND2_X1 U3410 ( .A1(n2687), .A2(n3825), .ZN(n3022) );
  INV_X1 U3411 ( .A(n3826), .ZN(n2688) );
  OR2_X1 U3412 ( .A1(n3022), .A2(n2688), .ZN(n2689) );
  NAND2_X1 U3413 ( .A1(n2689), .A2(n3829), .ZN(n3063) );
  AND2_X1 U3414 ( .A1(n3132), .A2(n3117), .ZN(n3062) );
  NAND2_X1 U3415 ( .A1(n3083), .A2(n3067), .ZN(n3839) );
  OAI21_X1 U3416 ( .B1(n3063), .B2(n3062), .A(n3839), .ZN(n3092) );
  INV_X1 U3417 ( .A(n3133), .ZN(n3150) );
  NAND2_X1 U3418 ( .A1(n3947), .A2(n3150), .ZN(n3840) );
  NAND2_X1 U3419 ( .A1(n3092), .A2(n3840), .ZN(n2690) );
  NAND2_X1 U3420 ( .A1(n3130), .A2(n3133), .ZN(n3831) );
  NAND2_X1 U3421 ( .A1(n2690), .A2(n3831), .ZN(n3101) );
  INV_X1 U3422 ( .A(n2691), .ZN(n2692) );
  NAND2_X1 U3423 ( .A1(n3256), .A2(n3238), .ZN(n3835) );
  NAND2_X1 U3424 ( .A1(n3945), .A2(n3233), .ZN(n3833) );
  NAND2_X1 U3425 ( .A1(n3296), .A2(n3252), .ZN(n3836) );
  NAND2_X1 U3426 ( .A1(n2694), .A2(n3836), .ZN(n3222) );
  NAND2_X1 U3427 ( .A1(n3290), .A2(n3346), .ZN(n3848) );
  NAND2_X1 U3428 ( .A1(n3222), .A2(n3848), .ZN(n2695) );
  NAND2_X1 U3429 ( .A1(n3321), .A2(n3288), .ZN(n3847) );
  NAND2_X1 U3430 ( .A1(n3944), .A2(n3388), .ZN(n3331) );
  NAND2_X1 U3431 ( .A1(n3637), .A2(n3441), .ZN(n3327) );
  NAND2_X1 U3432 ( .A1(n3331), .A2(n3327), .ZN(n3852) );
  NAND2_X1 U3433 ( .A1(n3338), .A2(n3379), .ZN(n3330) );
  NAND2_X1 U3434 ( .A1(n3301), .A2(n3330), .ZN(n2697) );
  INV_X1 U3435 ( .A(n3852), .ZN(n2696) );
  NOR2_X1 U3436 ( .A1(n3637), .A2(n3441), .ZN(n3328) );
  AOI21_X1 U3437 ( .B1(n2697), .B2(n2696), .A(n3328), .ZN(n3854) );
  INV_X1 U3438 ( .A(n3916), .ZN(n3408) );
  NAND2_X1 U3439 ( .A1(n3785), .A2(n3408), .ZN(n3421) );
  NAND2_X1 U3440 ( .A1(n3696), .A2(n3511), .ZN(n3784) );
  NAND2_X1 U3441 ( .A1(n3943), .A2(n3771), .ZN(n3783) );
  NAND2_X1 U3442 ( .A1(n3784), .A2(n3783), .ZN(n3422) );
  INV_X1 U3443 ( .A(n3781), .ZN(n2698) );
  NOR2_X1 U3444 ( .A1(n3422), .A2(n2698), .ZN(n2699) );
  NAND2_X1 U3445 ( .A1(n3421), .A2(n2699), .ZN(n2700) );
  NAND2_X1 U3446 ( .A1(n2700), .A2(n3783), .ZN(n3450) );
  INV_X1 U3447 ( .A(n3787), .ZN(n3858) );
  NAND2_X1 U3448 ( .A1(n3744), .A2(n4295), .ZN(n3862) );
  NAND2_X1 U3449 ( .A1(n4218), .A2(n4203), .ZN(n2701) );
  NAND2_X1 U3450 ( .A1(n4221), .A2(n2757), .ZN(n4188) );
  NAND2_X1 U3451 ( .A1(n4193), .A2(n4188), .ZN(n2703) );
  NOR2_X1 U3452 ( .A1(n4218), .A2(n4203), .ZN(n2702) );
  AOI21_X1 U3453 ( .B1(n2703), .B2(n3863), .A(n2702), .ZN(n4164) );
  NAND2_X1 U3454 ( .A1(n3675), .A2(n4180), .ZN(n2704) );
  NAND2_X1 U3455 ( .A1(n4199), .A2(n3727), .ZN(n3789) );
  NAND2_X1 U3456 ( .A1(n3736), .A2(n3555), .ZN(n4117) );
  NAND2_X1 U3457 ( .A1(n4119), .A2(n4117), .ZN(n3869) );
  INV_X1 U34580 ( .A(n3869), .ZN(n2706) );
  NAND2_X1 U34590 ( .A1(n4151), .A2(n2706), .ZN(n2711) );
  NAND2_X1 U3460 ( .A1(n4137), .A2(n4123), .ZN(n2707) );
  NAND2_X1 U3461 ( .A1(n2708), .A2(n2707), .ZN(n3872) );
  INV_X1 U3462 ( .A(n3872), .ZN(n2710) );
  AND2_X1 U3463 ( .A1(n4167), .A2(n4277), .ZN(n4116) );
  NAND2_X1 U3464 ( .A1(n4119), .A2(n4116), .ZN(n2709) );
  AND2_X1 U3465 ( .A1(n2710), .A2(n2709), .ZN(n3791) );
  NAND2_X1 U3466 ( .A1(n2711), .A2(n3791), .ZN(n4092) );
  NAND2_X1 U34670 ( .A1(n4126), .A2(n3575), .ZN(n3890) );
  NAND2_X1 U3468 ( .A1(n4097), .A2(n4112), .ZN(n4091) );
  NAND2_X1 U34690 ( .A1(n4092), .A2(n3871), .ZN(n2712) );
  NAND2_X1 U3470 ( .A1(n4079), .A2(n4262), .ZN(n3889) );
  AND2_X1 U34710 ( .A1(n4095), .A2(n4084), .ZN(n3887) );
  OR2_X1 U3472 ( .A1(n4038), .A2(n4066), .ZN(n2713) );
  OR2_X1 U34730 ( .A1(n4095), .A2(n4084), .ZN(n4055) );
  AND2_X1 U3474 ( .A1(n4038), .A2(n4066), .ZN(n3801) );
  NOR2_X1 U34750 ( .A1(n4064), .A2(n3599), .ZN(n3878) );
  INV_X1 U3476 ( .A(n3803), .ZN(n2714) );
  OAI21_X1 U34770 ( .B1(n4022), .B2(n3798), .A(n2714), .ZN(n2715) );
  XOR2_X1 U3478 ( .A(n3903), .B(n2715), .Z(n2729) );
  INV_X1 U34790 ( .A(n2684), .ZN(n4361) );
  NAND2_X1 U3480 ( .A1(n4361), .A2(n2151), .ZN(n3814) );
  NAND2_X1 U34810 ( .A1(n4362), .A2(n4360), .ZN(n2716) );
  NOR2_X1 U3482 ( .A1(n2717), .A2(n2730), .ZN(n2718) );
  MUX2_X1 U34830 ( .A(n2730), .B(n2718), .S(IR_REG_28__SCAN_IN), .Z(n2720) );
  OR2_X1 U3484 ( .A1(n2720), .A2(n2719), .ZN(n2895) );
  NAND2_X1 U34850 ( .A1(n4357), .A2(n2860), .ZN(n4220) );
  NOR2_X1 U3486 ( .A1(n4040), .A2(n4220), .ZN(n2728) );
  INV_X1 U34870 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U3488 ( .A1(n2146), .A2(REG2_REG_30__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U34890 ( .A1(n2721), .A2(REG1_REG_30__SCAN_IN), .ZN(n2722) );
  OAI211_X1 U3490 ( .C1(n2820), .C2(n2724), .A(n2723), .B(n2722), .ZN(n3780)
         );
  INV_X1 U34910 ( .A(n3780), .ZN(n3794) );
  XNOR2_X1 U3492 ( .A(n2392), .B(IR_REG_27__SCAN_IN), .ZN(n2935) );
  NAND2_X1 U34930 ( .A1(n2935), .A2(B_REG_SCAN_IN), .ZN(n2725) );
  NAND2_X1 U3494 ( .A1(n4217), .A2(n2725), .ZN(n4015) );
  OAI22_X1 U34950 ( .A1(n3794), .A2(n4015), .B1(n3795), .B2(n4294), .ZN(n2727)
         );
  AOI211_X1 U3496 ( .C1(n2729), .C2(n4196), .A(n2728), .B(n2727), .ZN(n3617)
         );
  OAI21_X1 U34970 ( .B1(n3624), .B2(n4533), .A(n3617), .ZN(n2764) );
  OR2_X1 U3498 ( .A1(n2731), .A2(n2730), .ZN(n2744) );
  INV_X1 U34990 ( .A(IR_REG_23__SCAN_IN), .ZN(n2743) );
  NAND2_X1 U3500 ( .A1(n2744), .A2(n2743), .ZN(n2742) );
  NAND2_X1 U35010 ( .A1(n2742), .A2(IR_REG_31__SCAN_IN), .ZN(n2733) );
  INV_X1 U3502 ( .A(IR_REG_24__SCAN_IN), .ZN(n2732) );
  NAND2_X1 U35030 ( .A1(n2755), .A2(n2741), .ZN(n2736) );
  MUX2_X1 U3504 ( .A(n2755), .B(n2736), .S(B_REG_SCAN_IN), .Z(n2739) );
  INV_X1 U35050 ( .A(D_REG_1__SCAN_IN), .ZN(n2740) );
  NAND2_X1 U35060 ( .A1(n2778), .A2(n2740), .ZN(n2857) );
  INV_X1 U35070 ( .A(n2772), .ZN(n2756) );
  NAND2_X1 U35080 ( .A1(n2756), .A2(n2741), .ZN(n2855) );
  NAND2_X1 U35090 ( .A1(n2857), .A2(n2855), .ZN(n2754) );
  OAI21_X1 U35100 ( .B1(n2744), .B2(n2743), .A(n2742), .ZN(n2982) );
  NAND2_X1 U35110 ( .A1(n2982), .A2(STATE_REG_SCAN_IN), .ZN(n4495) );
  INV_X1 U35120 ( .A(n4495), .ZN(n2781) );
  OR2_X1 U35130 ( .A1(n4523), .A2(n2151), .ZN(n2892) );
  NAND2_X1 U35140 ( .A1(n2684), .A2(n4010), .ZN(n2859) );
  NAND2_X1 U35150 ( .A1(n2859), .A2(n2860), .ZN(n2966) );
  AND3_X1 U35160 ( .A1(n2963), .A2(n2892), .A3(n2966), .ZN(n2753) );
  NOR4_X1 U35170 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2748) );
  NOR4_X1 U35180 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2747) );
  NOR4_X1 U35190 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2746) );
  NOR4_X1 U35200 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2745) );
  NAND4_X1 U35210 ( .A1(n2748), .A2(n2747), .A3(n2746), .A4(n2745), .ZN(n2752)
         );
  INV_X1 U35220 ( .A(D_REG_8__SCAN_IN), .ZN(n4839) );
  INV_X1 U35230 ( .A(D_REG_3__SCAN_IN), .ZN(n4679) );
  INV_X1 U35240 ( .A(D_REG_5__SCAN_IN), .ZN(n4680) );
  INV_X1 U35250 ( .A(D_REG_22__SCAN_IN), .ZN(n4699) );
  NAND4_X1 U35260 ( .A1(n4839), .A2(n4679), .A3(n4680), .A4(n4699), .ZN(n2749)
         );
  NOR3_X1 U35270 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(n2749), 
        .ZN(n4587) );
  NOR4_X1 U35280 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n4574) );
  NOR4_X1 U35290 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2750) );
  NAND3_X1 U35300 ( .A1(n4587), .A2(n4574), .A3(n2750), .ZN(n2751) );
  OAI21_X1 U35310 ( .B1(n2752), .B2(n2751), .A(n2778), .ZN(n2856) );
  INV_X1 U35320 ( .A(D_REG_0__SCAN_IN), .ZN(n4668) );
  AND2_X1 U35330 ( .A1(n2756), .A2(n2755), .ZN(n2782) );
  INV_X1 U35340 ( .A(n2858), .ZN(n2968) );
  AND2_X2 U35350 ( .A1(n2763), .A2(n2968), .ZN(n4545) );
  NAND2_X1 U35360 ( .A1(n2764), .A2(n4545), .ZN(n2762) );
  NAND2_X1 U35370 ( .A1(n3040), .A2(n2880), .ZN(n4486) );
  NAND2_X1 U35380 ( .A1(n3016), .A2(n3117), .ZN(n3096) );
  INV_X1 U35390 ( .A(n4030), .ZN(n2758) );
  INV_X1 U35400 ( .A(n3795), .ZN(n3800) );
  INV_X1 U35410 ( .A(n4510), .ZN(n2970) );
  NAND2_X1 U35420 ( .A1(n4544), .A2(REG0_REG_29__SCAN_IN), .ZN(n2759) );
  AND2_X2 U35430 ( .A1(n2763), .A2(n2858), .ZN(n4559) );
  NAND2_X1 U35440 ( .A1(n2764), .A2(n4559), .ZN(n2767) );
  NAND2_X1 U35450 ( .A1(n2767), .A2(n2766), .ZN(U3547) );
  INV_X2 U35460 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  MUX2_X1 U35470 ( .A(n3174), .B(n2487), .S(U3149), .Z(n2768) );
  INV_X1 U35480 ( .A(n2768), .ZN(U3344) );
  INV_X1 U35490 ( .A(DATAI_13_), .ZN(n2771) );
  NAND2_X1 U35500 ( .A1(n2769), .A2(STATE_REG_SCAN_IN), .ZN(n2770) );
  OAI21_X1 U35510 ( .B1(STATE_REG_SCAN_IN), .B2(n2771), .A(n2770), .ZN(U3339)
         );
  INV_X1 U35520 ( .A(DATAI_26_), .ZN(n4610) );
  NAND2_X1 U35530 ( .A1(n2772), .A2(STATE_REG_SCAN_IN), .ZN(n2773) );
  OAI21_X1 U35540 ( .B1(STATE_REG_SCAN_IN), .B2(n4610), .A(n2773), .ZN(U3326)
         );
  INV_X1 U35550 ( .A(DATAI_27_), .ZN(n2775) );
  NAND2_X1 U35560 ( .A1(n2935), .A2(STATE_REG_SCAN_IN), .ZN(n2774) );
  OAI21_X1 U35570 ( .B1(STATE_REG_SCAN_IN), .B2(n2775), .A(n2774), .ZN(U3325)
         );
  INV_X1 U35580 ( .A(DATAI_31_), .ZN(n4608) );
  OR4_X1 U35590 ( .A1(n2776), .A2(IR_REG_30__SCAN_IN), .A3(n2730), .A4(U3149), 
        .ZN(n2777) );
  OAI21_X1 U35600 ( .B1(STATE_REG_SCAN_IN), .B2(n4608), .A(n2777), .ZN(U3321)
         );
  INV_X1 U35610 ( .A(n2778), .ZN(n2779) );
  INV_X1 U35620 ( .A(n2855), .ZN(n2780) );
  AOI22_X1 U35630 ( .A1(n4493), .A2(n2740), .B1(n2780), .B2(n2781), .ZN(U3459)
         );
  AOI22_X1 U35640 ( .A1(n4493), .A2(n4668), .B1(n2782), .B2(n2781), .ZN(U3458)
         );
  XNOR2_X1 U35650 ( .A(n2793), .B(REG2_REG_1__SCAN_IN), .ZN(n3964) );
  AND2_X1 U35660 ( .A1(n4652), .A2(REG2_REG_0__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U35670 ( .A1(n3964), .A2(n2783), .ZN(n3963) );
  NAND2_X1 U35680 ( .A1(n4370), .A2(REG2_REG_1__SCAN_IN), .ZN(n2784) );
  NAND2_X1 U35690 ( .A1(n3963), .A2(n2784), .ZN(n2942) );
  INV_X1 U35700 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2785) );
  MUX2_X1 U35710 ( .A(REG2_REG_2__SCAN_IN), .B(n2785), .S(n4369), .Z(n2943) );
  XNOR2_X1 U35720 ( .A(n2801), .B(REG2_REG_3__SCAN_IN), .ZN(n2800) );
  OR2_X1 U35730 ( .A1(n2982), .A2(U3149), .ZN(n3937) );
  INV_X1 U35740 ( .A(n3937), .ZN(n2786) );
  OR2_X1 U35750 ( .A1(n2963), .A2(n2786), .ZN(n2790) );
  NAND2_X1 U35760 ( .A1(n2860), .A2(n2982), .ZN(n2787) );
  AND2_X1 U35770 ( .A1(n3779), .A2(n2787), .ZN(n2789) );
  NAND2_X1 U35780 ( .A1(n4357), .A2(n2935), .ZN(n3934) );
  INV_X1 U35790 ( .A(n3934), .ZN(n2788) );
  INV_X1 U35800 ( .A(n2789), .ZN(n2791) );
  INV_X1 U35810 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4638) );
  NOR2_X1 U3582 ( .A1(STATE_REG_SCAN_IN), .A2(n4638), .ZN(n3000) );
  NAND2_X1 U3583 ( .A1(n3953), .A2(n2895), .ZN(n4457) );
  INV_X1 U3584 ( .A(n4368), .ZN(n2796) );
  NOR2_X1 U3585 ( .A1(n4457), .A2(n2796), .ZN(n2792) );
  AOI211_X1 U3586 ( .C1(n4450), .C2(ADDR_REG_3__SCAN_IN), .A(n3000), .B(n2792), 
        .ZN(n2799) );
  XNOR2_X1 U3587 ( .A(n2793), .B(REG1_REG_1__SCAN_IN), .ZN(n3961) );
  AND2_X1 U3588 ( .A1(n4652), .A2(REG1_REG_0__SCAN_IN), .ZN(n3960) );
  NAND2_X1 U3589 ( .A1(n3961), .A2(n3960), .ZN(n3959) );
  NAND2_X1 U3590 ( .A1(n4370), .A2(REG1_REG_1__SCAN_IN), .ZN(n2794) );
  NAND2_X1 U3591 ( .A1(n3959), .A2(n2794), .ZN(n2945) );
  INV_X1 U3592 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4552) );
  MUX2_X1 U3593 ( .A(REG1_REG_2__SCAN_IN), .B(n4552), .S(n4369), .Z(n2946) );
  NAND2_X1 U3594 ( .A1(n2945), .A2(n2946), .ZN(n2944) );
  NAND2_X1 U3595 ( .A1(n4369), .A2(REG1_REG_2__SCAN_IN), .ZN(n2795) );
  NAND2_X1 U3596 ( .A1(n2944), .A2(n2795), .ZN(n2805) );
  XNOR2_X1 U3597 ( .A(n2805), .B(n2796), .ZN(n2797) );
  INV_X1 U3598 ( .A(n2935), .ZN(n3950) );
  NAND2_X1 U3599 ( .A1(n2797), .A2(REG1_REG_3__SCAN_IN), .ZN(n2807) );
  OAI211_X1 U3600 ( .C1(REG1_REG_3__SCAN_IN), .C2(n2797), .A(n4452), .B(n2807), 
        .ZN(n2798) );
  OAI211_X1 U3601 ( .C1(n2800), .C2(n4446), .A(n2799), .B(n2798), .ZN(U3243)
         );
  INV_X1 U3602 ( .A(n2832), .ZN(n4366) );
  XNOR2_X1 U3603 ( .A(n2802), .B(n4367), .ZN(n2952) );
  INV_X1 U3604 ( .A(n2802), .ZN(n2803) );
  INV_X1 U3605 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4762) );
  MUX2_X1 U3606 ( .A(REG2_REG_5__SCAN_IN), .B(n4762), .S(n2832), .Z(n2829) );
  XNOR2_X1 U3607 ( .A(n2838), .B(REG2_REG_6__SCAN_IN), .ZN(n2814) );
  INV_X1 U3608 ( .A(n4457), .ZN(n3958) );
  INV_X1 U3609 ( .A(n4450), .ZN(n4378) );
  INV_X1 U3610 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n2804) );
  NAND2_X1 U3611 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3134) );
  OAI21_X1 U3612 ( .B1(n4378), .B2(n2804), .A(n3134), .ZN(n2812) );
  INV_X1 U3613 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2810) );
  NAND2_X1 U3614 ( .A1(n2805), .A2(n4368), .ZN(n2806) );
  NAND2_X1 U3615 ( .A1(n2807), .A2(n2806), .ZN(n2808) );
  INV_X1 U3616 ( .A(n4367), .ZN(n2958) );
  XNOR2_X1 U3617 ( .A(n2808), .B(n2958), .ZN(n2954) );
  NAND2_X1 U3618 ( .A1(n2954), .A2(REG1_REG_4__SCAN_IN), .ZN(n2953) );
  XNOR2_X1 U3619 ( .A(n4366), .B(REG1_REG_5__SCAN_IN), .ZN(n2826) );
  XOR2_X1 U3620 ( .A(n4365), .B(n2276), .Z(n2809) );
  INV_X1 U3621 ( .A(n4452), .ZN(n3998) );
  NOR2_X1 U3622 ( .A1(n2809), .A2(n2810), .ZN(n2841) );
  AOI211_X1 U3623 ( .C1(n2810), .C2(n2809), .A(n3998), .B(n2841), .ZN(n2811)
         );
  AOI211_X1 U3624 ( .C1(n3958), .C2(n4365), .A(n2812), .B(n2811), .ZN(n2813)
         );
  OAI21_X1 U3625 ( .B1(n2814), .B2(n4446), .A(n2813), .ZN(U3246) );
  NOR2_X1 U3626 ( .A1(n4450), .A2(n2937), .ZN(U3148) );
  INV_X1 U3627 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4814) );
  NAND2_X1 U3628 ( .A1(n3088), .A2(U4043), .ZN(n2815) );
  OAI21_X1 U3629 ( .B1(n2937), .B2(n4814), .A(n2815), .ZN(U3554) );
  INV_X1 U3630 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U3631 ( .A1(n3744), .A2(U4043), .ZN(n2816) );
  OAI21_X1 U3632 ( .B1(n2937), .B2(n4826), .A(n2816), .ZN(U3567) );
  INV_X1 U3633 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4827) );
  NAND2_X1 U3634 ( .A1(n3497), .A2(U4043), .ZN(n2817) );
  OAI21_X1 U3635 ( .B1(n2937), .B2(n4827), .A(n2817), .ZN(U3564) );
  INV_X1 U3636 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4843) );
  INV_X1 U3637 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4306) );
  NAND2_X1 U3638 ( .A1(n2146), .A2(REG2_REG_31__SCAN_IN), .ZN(n2819) );
  NAND2_X1 U3639 ( .A1(n2721), .A2(REG1_REG_31__SCAN_IN), .ZN(n2818) );
  OAI211_X1 U3640 ( .C1(n2820), .C2(n4306), .A(n2819), .B(n2818), .ZN(n4017)
         );
  NAND2_X1 U3641 ( .A1(n4017), .A2(U4043), .ZN(n2821) );
  OAI21_X1 U3642 ( .B1(n2937), .B2(n4843), .A(n2821), .ZN(U3581) );
  INV_X1 U3643 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U3644 ( .A1(n3780), .A2(U4043), .ZN(n2822) );
  OAI21_X1 U3645 ( .B1(n2937), .B2(n4842), .A(n2822), .ZN(U3580) );
  INV_X1 U3646 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U3647 ( .A1(n3132), .A2(U4043), .ZN(n2823) );
  OAI21_X1 U3648 ( .B1(n2937), .B2(n4813), .A(n2823), .ZN(U3555) );
  INV_X1 U3649 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4811) );
  NAND2_X1 U3650 ( .A1(n2992), .A2(U4043), .ZN(n2824) );
  OAI21_X1 U3651 ( .B1(n2937), .B2(n4811), .A(n2824), .ZN(U3553) );
  AOI211_X1 U3652 ( .C1(n2827), .C2(n2826), .A(n2825), .B(n3998), .ZN(n2835)
         );
  AOI211_X1 U3653 ( .C1(n2830), .C2(n2829), .A(n2828), .B(n4446), .ZN(n2834)
         );
  AND2_X1 U3654 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3087) );
  AOI21_X1 U3655 ( .B1(n4450), .B2(ADDR_REG_5__SCAN_IN), .A(n3087), .ZN(n2831)
         );
  OAI21_X1 U3656 ( .B1(n2832), .B2(n4457), .A(n2831), .ZN(n2833) );
  OR3_X1 U3657 ( .A1(n2835), .A2(n2834), .A3(n2833), .ZN(U3245) );
  INV_X1 U3658 ( .A(n2836), .ZN(n2837) );
  INV_X1 U3659 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4760) );
  MUX2_X1 U3660 ( .A(n4760), .B(REG2_REG_7__SCAN_IN), .S(n4364), .Z(n2839) );
  NOR2_X1 U3661 ( .A1(n2840), .A2(n2839), .ZN(n2913) );
  AOI211_X1 U3662 ( .C1(n2840), .C2(n2839), .A(n4446), .B(n2913), .ZN(n2848)
         );
  INV_X1 U3663 ( .A(n4364), .ZN(n2845) );
  INV_X1 U3664 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4555) );
  NAND2_X1 U3665 ( .A1(n4364), .A2(REG1_REG_7__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U3666 ( .A1(n2194), .A2(n2911), .ZN(n2843) );
  OAI21_X1 U3667 ( .B1(n2912), .B2(n2843), .A(n4452), .ZN(n2842) );
  AOI21_X1 U3668 ( .B1(n2912), .B2(n2843), .A(n2842), .ZN(n2847) );
  AND2_X1 U3669 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3217) );
  AOI21_X1 U3670 ( .B1(n4450), .B2(ADDR_REG_7__SCAN_IN), .A(n3217), .ZN(n2844)
         );
  OAI21_X1 U3671 ( .B1(n2845), .B2(n4457), .A(n2844), .ZN(n2846) );
  OR3_X1 U3672 ( .A1(n2848), .A2(n2847), .A3(n2846), .ZN(U3247) );
  INV_X1 U3673 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4823) );
  NAND2_X1 U3674 ( .A1(n3637), .A2(n2937), .ZN(n2849) );
  OAI21_X1 U3675 ( .B1(n2937), .B2(n4823), .A(n2849), .ZN(U3563) );
  INV_X1 U3676 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4816) );
  NAND2_X1 U3677 ( .A1(n3290), .A2(n2937), .ZN(n2850) );
  OAI21_X1 U3678 ( .B1(n2937), .B2(n4816), .A(n2850), .ZN(U3560) );
  INV_X1 U3679 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4817) );
  NAND2_X1 U3680 ( .A1(n3251), .A2(n2937), .ZN(n2851) );
  OAI21_X1 U3681 ( .B1(n2937), .B2(n4817), .A(n2851), .ZN(U3559) );
  INV_X1 U3682 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4829) );
  NAND2_X1 U3683 ( .A1(n4167), .A2(n2937), .ZN(n2852) );
  OAI21_X1 U3684 ( .B1(n2937), .B2(n4829), .A(n2852), .ZN(U3571) );
  INV_X1 U3685 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U3686 ( .A1(n3305), .A2(n2937), .ZN(n2853) );
  OAI21_X1 U3687 ( .B1(n2937), .B2(n4824), .A(n2853), .ZN(U3561) );
  INV_X1 U3688 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U3689 ( .A1(n3035), .A2(n2937), .ZN(n2854) );
  OAI21_X1 U3690 ( .B1(n2937), .B2(n4810), .A(n2854), .ZN(U3552) );
  AND2_X1 U3691 ( .A1(n2856), .A2(n2855), .ZN(n2967) );
  INV_X1 U3692 ( .A(n2898), .ZN(n2867) );
  NAND2_X1 U3693 ( .A1(n2970), .A2(n2859), .ZN(n2862) );
  INV_X1 U3694 ( .A(n2860), .ZN(n2861) );
  NAND2_X1 U3695 ( .A1(n2862), .A2(n2861), .ZN(n2888) );
  NAND2_X1 U3696 ( .A1(n2888), .A2(n4294), .ZN(n2864) );
  INV_X1 U3697 ( .A(n2966), .ZN(n2863) );
  AOI21_X1 U3698 ( .B1(n2867), .B2(n2864), .A(n2863), .ZN(n2984) );
  INV_X1 U3699 ( .A(n2868), .ZN(n2865) );
  NAND2_X1 U3700 ( .A1(n4010), .A2(n4360), .ZN(n2869) );
  OR3_X1 U3701 ( .A1(n3562), .A2(n4495), .A3(n2869), .ZN(n3933) );
  INV_X1 U3702 ( .A(n3933), .ZN(n2866) );
  NAND2_X1 U3703 ( .A1(n2867), .A2(n2866), .ZN(n2985) );
  NAND3_X1 U3704 ( .A1(n2984), .A2(n2963), .A3(n2985), .ZN(n2931) );
  INV_X1 U3705 ( .A(n2931), .ZN(n2903) );
  INV_X1 U3706 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2902) );
  OAI22_X1 U3707 ( .A1(n2973), .A2(n2873), .B1(n2154), .B2(n3040), .ZN(n2870)
         );
  NAND2_X4 U3708 ( .A1(n2868), .A2(n2869), .ZN(n3585) );
  XNOR2_X1 U3709 ( .A(n2870), .B(n3585), .ZN(n2921) );
  AND2_X1 U3710 ( .A1(n3034), .A2(n3584), .ZN(n2874) );
  AOI21_X2 U3711 ( .B1(n2875), .B2(n2150), .A(n2874), .ZN(n2922) );
  XNOR2_X1 U3712 ( .A(n2921), .B(n2922), .ZN(n2886) );
  INV_X1 U3713 ( .A(n2983), .ZN(n2877) );
  INV_X1 U3714 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2876) );
  INV_X1 U3715 ( .A(n2881), .ZN(n2882) );
  OAI21_X1 U3716 ( .B1(n2972), .B2(n2879), .A(n2882), .ZN(n2906) );
  NAND2_X1 U3717 ( .A1(n2904), .A2(n2906), .ZN(n2905) );
  NAND2_X1 U3718 ( .A1(n2905), .A2(n2885), .ZN(n2887) );
  NAND2_X1 U3719 ( .A1(n2887), .A2(n2886), .ZN(n2925) );
  INV_X1 U3720 ( .A(n2888), .ZN(n2889) );
  AND2_X1 U3721 ( .A1(n2889), .A2(n2963), .ZN(n2890) );
  INV_X1 U3722 ( .A(n3762), .ZN(n3767) );
  OAI211_X1 U3723 ( .C1(n2886), .C2(n2887), .A(n2925), .B(n3767), .ZN(n2901)
         );
  AND2_X1 U3724 ( .A1(n4475), .A2(n2963), .ZN(n2891) );
  NAND2_X1 U3725 ( .A1(n2898), .A2(n2891), .ZN(n2894) );
  INV_X1 U3726 ( .A(n2892), .ZN(n2893) );
  AND2_X2 U3727 ( .A1(n2893), .A2(n2963), .ZN(n4483) );
  NOR2_X1 U3728 ( .A1(n3933), .A2(n2895), .ZN(n2896) );
  NAND2_X1 U3729 ( .A1(n2898), .A2(n2896), .ZN(n3769) );
  NOR2_X1 U3730 ( .A1(n3933), .A2(n4357), .ZN(n2897) );
  NAND2_X1 U3731 ( .A1(n2898), .A2(n2897), .ZN(n3758) );
  OAI22_X1 U3732 ( .A1(n2972), .A2(n3769), .B1(n3009), .B2(n3758), .ZN(n2899)
         );
  AOI21_X1 U3733 ( .B1(n3034), .B2(n3755), .A(n2899), .ZN(n2900) );
  OAI211_X1 U3734 ( .C1(n2903), .C2(n2902), .A(n2901), .B(n2900), .ZN(U3219)
         );
  OAI21_X1 U3735 ( .B1(n2906), .B2(n2904), .A(n2905), .ZN(n2938) );
  AOI22_X1 U3736 ( .A1(n3755), .A2(n2971), .B1(n3774), .B2(n2414), .ZN(n2908)
         );
  NAND2_X1 U3737 ( .A1(n2931), .A2(REG3_REG_0__SCAN_IN), .ZN(n2907) );
  OAI211_X1 U3738 ( .C1(n2938), .C2(n3762), .A(n2908), .B(n2907), .ZN(U3229)
         );
  INV_X1 U3739 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4833) );
  NAND2_X1 U3740 ( .A1(n3797), .A2(U4043), .ZN(n2909) );
  OAI21_X1 U3741 ( .B1(U4043), .B2(n4833), .A(n2909), .ZN(U3579) );
  INV_X1 U3742 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U3743 ( .A1(n4095), .A2(U4043), .ZN(n2910) );
  OAI21_X1 U3744 ( .B1(n2937), .B2(n4830), .A(n2910), .ZN(U3575) );
  XNOR2_X1 U3745 ( .A(n3157), .B(REG1_REG_8__SCAN_IN), .ZN(n2919) );
  AOI21_X1 U3746 ( .B1(n4364), .B2(REG2_REG_7__SCAN_IN), .A(n2913), .ZN(n3175)
         );
  XNOR2_X1 U3747 ( .A(REG2_REG_8__SCAN_IN), .B(n3177), .ZN(n2914) );
  NAND2_X1 U3748 ( .A1(n4410), .A2(n2914), .ZN(n2915) );
  NAND2_X1 U3749 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3207) );
  NAND2_X1 U3750 ( .A1(n2915), .A2(n3207), .ZN(n2917) );
  NOR2_X1 U3751 ( .A1(n4457), .A2(n3174), .ZN(n2916) );
  AOI211_X1 U3752 ( .C1(n4450), .C2(ADDR_REG_8__SCAN_IN), .A(n2917), .B(n2916), 
        .ZN(n2918) );
  OAI21_X1 U3753 ( .B1(n2919), .B2(n3998), .A(n2918), .ZN(U3248) );
  OAI22_X1 U3754 ( .A1(n3009), .A2(n2149), .B1(n2929), .B2(n2154), .ZN(n2920)
         );
  XNOR2_X1 U3755 ( .A(n2920), .B(n3585), .ZN(n2988) );
  OAI22_X1 U3756 ( .A1(n3009), .A2(n2879), .B1(n2929), .B2(n3562), .ZN(n2987)
         );
  XNOR2_X1 U3757 ( .A(n2988), .B(n2987), .ZN(n2927) );
  INV_X1 U3758 ( .A(n2922), .ZN(n2923) );
  NAND2_X1 U3759 ( .A1(n2925), .A2(n2924), .ZN(n2926) );
  AOI21_X1 U3760 ( .B1(n2927), .B2(n2926), .A(n2989), .ZN(n2933) );
  AOI22_X1 U3761 ( .A1(n3774), .A2(n2992), .B1(n3754), .B2(n2414), .ZN(n2928)
         );
  OAI21_X1 U3762 ( .B1(n3772), .B2(n2929), .A(n2928), .ZN(n2930) );
  AOI21_X1 U3763 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2931), .A(n2930), .ZN(n2932)
         );
  OAI21_X1 U3764 ( .B1(n2933), .B2(n3762), .A(n2932), .ZN(U3234) );
  INV_X1 U3765 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U3766 ( .A1(n4038), .A2(U4043), .ZN(n2934) );
  OAI21_X1 U3767 ( .B1(n2937), .B2(n4832), .A(n2934), .ZN(U3576) );
  INV_X1 U3768 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2976) );
  NAND2_X1 U3769 ( .A1(n2935), .A2(n2976), .ZN(n2936) );
  NAND2_X1 U3770 ( .A1(n4357), .A2(n2936), .ZN(n3951) );
  NAND2_X1 U3771 ( .A1(n4652), .A2(REG2_REG_0__SCAN_IN), .ZN(n3962) );
  OAI21_X1 U3772 ( .B1(n3934), .B2(n3962), .A(n2937), .ZN(n2940) );
  AND3_X1 U3773 ( .A1(n2938), .A2(n4357), .A3(n3950), .ZN(n2939) );
  OAI211_X1 U3774 ( .C1(n2943), .C2(n2942), .A(n4410), .B(n2941), .ZN(n2950)
         );
  NAND2_X1 U3775 ( .A1(n3958), .A2(n4369), .ZN(n2949) );
  OAI211_X1 U3776 ( .C1(n2946), .C2(n2945), .A(n4452), .B(n2944), .ZN(n2948)
         );
  AOI22_X1 U3777 ( .A1(n4450), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2947) );
  NAND4_X1 U3778 ( .A1(n2950), .A2(n2949), .A3(n2948), .A4(n2947), .ZN(n2951)
         );
  OR2_X1 U3779 ( .A1(n2959), .A2(n2951), .ZN(U3242) );
  XOR2_X1 U3780 ( .A(REG2_REG_4__SCAN_IN), .B(n2952), .Z(n2961) );
  OAI211_X1 U3781 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2954), .A(n4452), .B(n2953), 
        .ZN(n2957) );
  NAND2_X1 U3782 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3045) );
  INV_X1 U3783 ( .A(n3045), .ZN(n2955) );
  AOI21_X1 U3784 ( .B1(n4450), .B2(ADDR_REG_4__SCAN_IN), .A(n2955), .ZN(n2956)
         );
  OAI211_X1 U3785 ( .C1(n4457), .C2(n2958), .A(n2957), .B(n2956), .ZN(n2960)
         );
  AOI211_X1 U3786 ( .C1(n4410), .C2(n2961), .A(n2960), .B(n2959), .ZN(n2962)
         );
  INV_X1 U3787 ( .A(n2962), .ZN(U3244) );
  NAND2_X1 U3788 ( .A1(n2963), .A2(D_REG_1__SCAN_IN), .ZN(n2964) );
  NAND2_X1 U3789 ( .A1(n4493), .A2(n2964), .ZN(n2965) );
  NAND4_X1 U3790 ( .A1(n2968), .A2(n2967), .A3(n2966), .A4(n2965), .ZN(n2969)
         );
  INV_X2 U3791 ( .A(n4232), .ZN(n4371) );
  NOR2_X1 U3792 ( .A1(n4371), .A2(n4362), .ZN(n4227) );
  NOR2_X1 U3793 ( .A1(n4371), .A2(n4294), .ZN(n4033) );
  AOI21_X1 U3794 ( .B1(n4227), .B2(n2970), .A(n4033), .ZN(n2981) );
  NOR2_X1 U3795 ( .A1(n2972), .A2(n2971), .ZN(n3815) );
  INV_X1 U3796 ( .A(n3030), .ZN(n3818) );
  NOR2_X1 U3797 ( .A1(n3815), .A2(n3818), .ZN(n4511) );
  INV_X1 U3798 ( .A(n4174), .ZN(n4482) );
  NOR2_X1 U3799 ( .A1(n4482), .A2(n4196), .ZN(n2974) );
  OAI22_X1 U3800 ( .A1(n4511), .A2(n2974), .B1(n2973), .B2(n4479), .ZN(n4513)
         );
  INV_X1 U3801 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2975) );
  OAI22_X1 U3802 ( .A1(n4232), .A2(n2976), .B1(n2975), .B2(n4114), .ZN(n2979)
         );
  OR2_X1 U3803 ( .A1(n2868), .A2(n4010), .ZN(n3074) );
  INV_X1 U3804 ( .A(n3074), .ZN(n2977) );
  NAND2_X1 U3805 ( .A1(n4232), .A2(n2977), .ZN(n4183) );
  NOR2_X1 U3806 ( .A1(n4511), .A2(n4183), .ZN(n2978) );
  AOI211_X1 U3807 ( .C1(n4232), .C2(n4513), .A(n2979), .B(n2978), .ZN(n2980)
         );
  OAI21_X1 U3808 ( .B1(n2981), .B2(n2880), .A(n2980), .ZN(U3290) );
  AND3_X1 U3809 ( .A1(n2984), .A2(n2983), .A3(n2982), .ZN(n2986) );
  OAI21_X2 U3810 ( .B1(n2986), .B2(U3149), .A(n2985), .ZN(n3747) );
  INV_X1 U3811 ( .A(n2987), .ZN(n2991) );
  INV_X1 U3812 ( .A(n2988), .ZN(n2990) );
  NAND2_X1 U3813 ( .A1(n2992), .A2(n3584), .ZN(n2994) );
  NAND2_X1 U3814 ( .A1(n3012), .A2(n2872), .ZN(n2993) );
  NAND2_X1 U3815 ( .A1(n2994), .A2(n2993), .ZN(n2995) );
  XNOR2_X1 U3816 ( .A(n2995), .B(n3585), .ZN(n3053) );
  OAI22_X1 U3817 ( .A1(n4480), .A2(n2879), .B1(n2998), .B2(n3562), .ZN(n3052)
         );
  XNOR2_X1 U3818 ( .A(n3053), .B(n3052), .ZN(n3055) );
  XNOR2_X1 U3819 ( .A(n3054), .B(n3055), .ZN(n2996) );
  NAND2_X1 U3820 ( .A1(n2996), .A2(n3767), .ZN(n3002) );
  OAI22_X1 U3821 ( .A1(n3772), .A2(n2998), .B1(n2997), .B2(n3758), .ZN(n2999)
         );
  AOI211_X1 U3822 ( .C1(n3754), .C2(n3035), .A(n3000), .B(n2999), .ZN(n3001)
         );
  OAI211_X1 U3823 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3778), .A(n3002), .B(n3001), 
        .ZN(U3215) );
  INV_X1 U3824 ( .A(n4523), .ZN(n4530) );
  INV_X1 U3825 ( .A(n3004), .ZN(n3914) );
  XNOR2_X1 U3826 ( .A(n3003), .B(n3914), .ZN(n4466) );
  XNOR2_X1 U3827 ( .A(n3005), .B(n3004), .ZN(n3006) );
  NAND2_X1 U3828 ( .A1(n3006), .A2(n4196), .ZN(n3008) );
  AOI22_X1 U3829 ( .A1(n3088), .A2(n4217), .B1(n4475), .B2(n3012), .ZN(n3007)
         );
  OAI211_X1 U3830 ( .C1(n3009), .C2(n4220), .A(n3008), .B(n3007), .ZN(n3010)
         );
  AOI21_X1 U3831 ( .B1(n4482), .B2(n4466), .A(n3010), .ZN(n4469) );
  INV_X1 U3832 ( .A(n4469), .ZN(n3011) );
  AOI21_X1 U3833 ( .B1(n4530), .B2(n4466), .A(n3011), .ZN(n3015) );
  AOI21_X1 U3834 ( .B1(n3012), .B2(n4484), .A(n3017), .ZN(n4465) );
  INV_X1 U3835 ( .A(n4300), .ZN(n4549) );
  AOI22_X1 U3836 ( .A1(n4465), .A2(n4549), .B1(REG1_REG_3__SCAN_IN), .B2(n4557), .ZN(n3013) );
  OAI21_X1 U3837 ( .B1(n3015), .B2(n4557), .A(n3013), .ZN(U3521) );
  INV_X1 U3838 ( .A(n4352), .ZN(n4525) );
  AOI22_X1 U3839 ( .A1(n4465), .A2(n4525), .B1(REG0_REG_3__SCAN_IN), .B2(n4544), .ZN(n3014) );
  OAI21_X1 U3840 ( .B1(n3015), .B2(n4544), .A(n3014), .ZN(U3473) );
  INV_X1 U3841 ( .A(n3016), .ZN(n3066) );
  OAI211_X1 U3842 ( .C1(n3017), .C2(n3020), .A(n3066), .B(n4516), .ZN(n4527)
         );
  NOR2_X1 U3843 ( .A1(n4527), .A2(n4362), .ZN(n3026) );
  OR2_X1 U3844 ( .A1(n3018), .A2(n3905), .ZN(n3072) );
  NAND2_X1 U3845 ( .A1(n3018), .A2(n3905), .ZN(n3019) );
  NAND2_X1 U3846 ( .A1(n3072), .A2(n3019), .ZN(n3027) );
  OAI22_X1 U3847 ( .A1(n4480), .A2(n4220), .B1(n3020), .B2(n4294), .ZN(n3021)
         );
  AOI21_X1 U3848 ( .B1(n4217), .B2(n3132), .A(n3021), .ZN(n3025) );
  XNOR2_X1 U3849 ( .A(n3022), .B(n3905), .ZN(n3023) );
  NAND2_X1 U3850 ( .A1(n3023), .A2(n4196), .ZN(n3024) );
  OAI211_X1 U3851 ( .C1(n3027), .C2(n4174), .A(n3025), .B(n3024), .ZN(n4528)
         );
  AOI211_X1 U3852 ( .C1(n4483), .C2(n3060), .A(n3026), .B(n4528), .ZN(n3029)
         );
  INV_X1 U3853 ( .A(n3027), .ZN(n4531) );
  INV_X1 U3854 ( .A(n4183), .ZN(n4489) );
  AOI22_X1 U3855 ( .A1(n4531), .A2(n4489), .B1(REG2_REG_4__SCAN_IN), .B2(n4371), .ZN(n3028) );
  OAI21_X1 U3856 ( .B1(n3029), .B2(n4371), .A(n3028), .ZN(U3286) );
  XNOR2_X1 U3857 ( .A(n2686), .B(n3030), .ZN(n3039) );
  OR2_X1 U3858 ( .A1(n2686), .A2(n3031), .ZN(n3032) );
  NAND2_X1 U3859 ( .A1(n3033), .A2(n3032), .ZN(n4518) );
  AOI22_X1 U3860 ( .A1(n3035), .A2(n4217), .B1(n4475), .B2(n3034), .ZN(n3037)
         );
  NAND2_X1 U3861 ( .A1(n3949), .A2(n4476), .ZN(n3036) );
  OAI211_X1 U3862 ( .C1(n4518), .C2(n4174), .A(n3037), .B(n3036), .ZN(n3038)
         );
  AOI21_X1 U3863 ( .B1(n4196), .B2(n3039), .A(n3038), .ZN(n4515) );
  NAND2_X1 U3864 ( .A1(n4227), .A2(n4516), .ZN(n4207) );
  OAI21_X1 U3865 ( .B1(n2880), .B2(n3040), .A(n4486), .ZN(n4517) );
  INV_X1 U3866 ( .A(n4517), .ZN(n3043) );
  AOI22_X1 U3867 ( .A1(n4492), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4483), .ZN(n3041) );
  OAI21_X1 U3868 ( .B1(n4518), .B2(n4183), .A(n3041), .ZN(n3042) );
  AOI21_X1 U3869 ( .B1(n4488), .B2(n3043), .A(n3042), .ZN(n3044) );
  OAI21_X1 U3870 ( .B1(n4515), .B2(n4371), .A(n3044), .ZN(U3289) );
  INV_X1 U3871 ( .A(n3778), .ZN(n3760) );
  AOI22_X1 U3872 ( .A1(n3755), .A2(n3050), .B1(n3132), .B2(n3774), .ZN(n3046)
         );
  OAI211_X1 U3873 ( .C1(n4480), .C2(n3769), .A(n3046), .B(n3045), .ZN(n3059)
         );
  NAND2_X1 U3874 ( .A1(n3088), .A2(n3584), .ZN(n3048) );
  NAND2_X1 U3875 ( .A1(n3050), .A2(n2872), .ZN(n3047) );
  NAND2_X1 U3876 ( .A1(n3048), .A2(n3047), .ZN(n3049) );
  XNOR2_X1 U3877 ( .A(n3049), .B(n3585), .ZN(n3080) );
  AND2_X1 U3878 ( .A1(n3050), .A2(n3584), .ZN(n3051) );
  AOI21_X1 U3879 ( .B1(n3088), .B2(n3594), .A(n3051), .ZN(n3078) );
  XOR2_X1 U3880 ( .A(n3080), .B(n3078), .Z(n3057) );
  AOI211_X1 U3881 ( .C1(n3057), .C2(n3056), .A(n3762), .B(n2188), .ZN(n3058)
         );
  AOI211_X1 U3882 ( .C1(n3060), .C2(n3760), .A(n3059), .B(n3058), .ZN(n3061)
         );
  INV_X1 U3883 ( .A(n3061), .ZN(U3227) );
  INV_X1 U3884 ( .A(n3062), .ZN(n3828) );
  NAND2_X1 U3885 ( .A1(n3828), .A2(n3839), .ZN(n3910) );
  XNOR2_X1 U3886 ( .A(n3063), .B(n3910), .ZN(n3064) );
  AOI222_X1 U3887 ( .A1(n4196), .A2(n3064), .B1(n3947), .B2(n4217), .C1(n3088), 
        .C2(n4476), .ZN(n3116) );
  INV_X1 U3888 ( .A(n3096), .ZN(n3065) );
  AOI21_X1 U3889 ( .B1(n3067), .B2(n3066), .A(n3065), .ZN(n3121) );
  INV_X1 U3890 ( .A(n4033), .ZN(n4159) );
  NOR2_X1 U3891 ( .A1(n4159), .A2(n3117), .ZN(n3070) );
  INV_X1 U3892 ( .A(n3068), .ZN(n3091) );
  OAI22_X1 U3893 ( .A1(n4232), .A2(n4762), .B1(n3091), .B2(n4114), .ZN(n3069)
         );
  AOI211_X1 U3894 ( .C1(n3121), .C2(n4488), .A(n3070), .B(n3069), .ZN(n3077)
         );
  NAND2_X1 U3895 ( .A1(n3072), .A2(n3071), .ZN(n3073) );
  XOR2_X1 U3896 ( .A(n3910), .B(n3073), .Z(n3119) );
  NAND2_X1 U3897 ( .A1(n4174), .A2(n3074), .ZN(n3075) );
  NAND2_X1 U3898 ( .A1(n3119), .A2(n4156), .ZN(n3076) );
  OAI211_X1 U3899 ( .C1(n3116), .C2(n4371), .A(n3077), .B(n3076), .ZN(U3285)
         );
  INV_X1 U3900 ( .A(n3078), .ZN(n3079) );
  OAI22_X1 U3901 ( .A1(n3083), .A2(n3562), .B1(n2153), .B2(n3117), .ZN(n3082)
         );
  XNOR2_X1 U3902 ( .A(n3082), .B(n3585), .ZN(n3124) );
  OAI22_X1 U3903 ( .A1(n3083), .A2(n2879), .B1(n3562), .B2(n3117), .ZN(n3125)
         );
  XNOR2_X1 U3904 ( .A(n3124), .B(n3125), .ZN(n3127) );
  AOI21_X1 U3905 ( .B1(n3128), .B2(n3127), .A(n3762), .ZN(n3085) );
  OR2_X1 U3906 ( .A1(n3128), .A2(n3127), .ZN(n3084) );
  NAND2_X1 U3907 ( .A1(n3085), .A2(n3084), .ZN(n3090) );
  OAI22_X1 U3908 ( .A1(n3772), .A2(n3117), .B1(n3130), .B2(n3758), .ZN(n3086)
         );
  AOI211_X1 U3909 ( .C1(n3754), .C2(n3088), .A(n3087), .B(n3086), .ZN(n3089)
         );
  OAI211_X1 U3910 ( .C1(n3778), .C2(n3091), .A(n3090), .B(n3089), .ZN(U3224)
         );
  NAND2_X1 U3911 ( .A1(n3831), .A2(n3840), .ZN(n3915) );
  XOR2_X1 U3912 ( .A(n3915), .B(n3092), .Z(n3093) );
  AOI222_X1 U3913 ( .A1(n4196), .A2(n3093), .B1(n3946), .B2(n4217), .C1(n3132), 
        .C2(n4476), .ZN(n3149) );
  XOR2_X1 U3914 ( .A(n3915), .B(n3094), .Z(n3152) );
  INV_X1 U3915 ( .A(n3106), .ZN(n3095) );
  AOI21_X1 U3916 ( .B1(n3133), .B2(n3096), .A(n3095), .ZN(n3154) );
  NAND2_X1 U3917 ( .A1(n3154), .A2(n4488), .ZN(n3098) );
  AOI22_X1 U3918 ( .A1(n4492), .A2(REG2_REG_6__SCAN_IN), .B1(n3137), .B2(n4483), .ZN(n3097) );
  OAI211_X1 U3919 ( .C1(n4159), .C2(n3150), .A(n3098), .B(n3097), .ZN(n3099)
         );
  AOI21_X1 U3920 ( .B1(n3152), .B2(n4156), .A(n3099), .ZN(n3100) );
  OAI21_X1 U3921 ( .B1(n3149), .B2(n4371), .A(n3100), .ZN(U3284) );
  XNOR2_X1 U3922 ( .A(n3101), .B(n3906), .ZN(n3102) );
  NAND2_X1 U3923 ( .A1(n3102), .A2(n4196), .ZN(n3105) );
  OAI22_X1 U3924 ( .A1(n3256), .A2(n4479), .B1(n3215), .B2(n4294), .ZN(n3103)
         );
  INV_X1 U3925 ( .A(n3103), .ZN(n3104) );
  OAI211_X1 U3926 ( .C1(n3130), .C2(n4220), .A(n3105), .B(n3104), .ZN(n4535)
         );
  INV_X1 U3927 ( .A(n4535), .ZN(n3115) );
  NAND2_X1 U3928 ( .A1(n3106), .A2(n3197), .ZN(n3107) );
  NAND2_X1 U3929 ( .A1(n3107), .A2(n4516), .ZN(n3108) );
  NOR2_X1 U3930 ( .A1(n3234), .A2(n3108), .ZN(n4536) );
  INV_X1 U3931 ( .A(n3218), .ZN(n3109) );
  OAI22_X1 U3932 ( .A1(n4232), .A2(n4760), .B1(n3109), .B2(n4114), .ZN(n3113)
         );
  INV_X1 U3933 ( .A(n4537), .ZN(n3111) );
  AND2_X1 U3934 ( .A1(n3110), .A2(n3906), .ZN(n4534) );
  NOR3_X1 U3935 ( .A1(n3111), .A2(n4534), .A3(n4235), .ZN(n3112) );
  AOI211_X1 U3936 ( .C1(n4227), .C2(n4536), .A(n3113), .B(n3112), .ZN(n3114)
         );
  OAI21_X1 U3937 ( .B1(n4371), .B2(n3115), .A(n3114), .ZN(U3283) );
  OAI21_X1 U3938 ( .B1(n3117), .B2(n4294), .A(n3116), .ZN(n3118) );
  AOI21_X1 U3939 ( .B1(n3119), .B2(n4542), .A(n3118), .ZN(n3123) );
  AOI22_X1 U3940 ( .A1(n3121), .A2(n4549), .B1(REG1_REG_5__SCAN_IN), .B2(n4557), .ZN(n3120) );
  OAI21_X1 U3941 ( .B1(n3123), .B2(n4557), .A(n3120), .ZN(U3523) );
  AOI22_X1 U3942 ( .A1(n3121), .A2(n4525), .B1(REG0_REG_5__SCAN_IN), .B2(n4544), .ZN(n3122) );
  OAI21_X1 U3943 ( .B1(n3123), .B2(n4544), .A(n3122), .ZN(U3477) );
  NAND2_X1 U3944 ( .A1(n3124), .A2(n3125), .ZN(n3126) );
  OAI22_X1 U3945 ( .A1(n3130), .A2(n3562), .B1(n2154), .B2(n3150), .ZN(n3129)
         );
  XNOR2_X1 U3946 ( .A(n3129), .B(n3585), .ZN(n3188) );
  OAI22_X1 U3947 ( .A1(n3130), .A2(n2879), .B1(n3562), .B2(n3150), .ZN(n3189)
         );
  INV_X1 U3948 ( .A(n3189), .ZN(n3190) );
  XNOR2_X1 U3949 ( .A(n3188), .B(n3190), .ZN(n3131) );
  XNOR2_X1 U3950 ( .A(n3191), .B(n3131), .ZN(n3139) );
  AOI22_X1 U3951 ( .A1(n3755), .A2(n3133), .B1(n3132), .B2(n3754), .ZN(n3135)
         );
  OAI211_X1 U3952 ( .C1(n3209), .C2(n3758), .A(n3135), .B(n3134), .ZN(n3136)
         );
  AOI21_X1 U3953 ( .B1(n3137), .B2(n3760), .A(n3136), .ZN(n3138) );
  OAI21_X1 U3954 ( .B1(n3139), .B2(n3762), .A(n3138), .ZN(U3236) );
  NAND2_X1 U3955 ( .A1(n2177), .A2(n3836), .ZN(n3891) );
  XNOR2_X1 U3956 ( .A(n3140), .B(n3891), .ZN(n3143) );
  AOI22_X1 U3957 ( .A1(n3290), .A2(n4217), .B1(n4475), .B2(n3252), .ZN(n3141)
         );
  OAI21_X1 U3958 ( .B1(n3256), .B2(n4220), .A(n3141), .ZN(n3142) );
  AOI21_X1 U3959 ( .B1(n3143), .B2(n4196), .A(n3142), .ZN(n4539) );
  XOR2_X1 U3960 ( .A(n3891), .B(n3144), .Z(n4543) );
  OR2_X1 U3961 ( .A1(n3231), .A2(n3257), .ZN(n3145) );
  NAND2_X1 U3962 ( .A1(n3225), .A2(n3145), .ZN(n4540) );
  AOI22_X1 U3963 ( .A1(n4492), .A2(REG2_REG_9__SCAN_IN), .B1(n3259), .B2(n4483), .ZN(n3146) );
  OAI21_X1 U3964 ( .B1(n4540), .B2(n4207), .A(n3146), .ZN(n3147) );
  AOI21_X1 U3965 ( .B1(n4543), .B2(n4156), .A(n3147), .ZN(n3148) );
  OAI21_X1 U3966 ( .B1(n4492), .B2(n4539), .A(n3148), .ZN(U3281) );
  OAI21_X1 U3967 ( .B1(n3150), .B2(n4294), .A(n3149), .ZN(n3151) );
  AOI21_X1 U3968 ( .B1(n3152), .B2(n4542), .A(n3151), .ZN(n3156) );
  AOI22_X1 U3969 ( .A1(n3154), .A2(n4525), .B1(n4544), .B2(REG0_REG_6__SCAN_IN), .ZN(n3153) );
  OAI21_X1 U3970 ( .B1(n3156), .B2(n4544), .A(n3153), .ZN(U3479) );
  AOI22_X1 U3971 ( .A1(n3154), .A2(n4549), .B1(n4557), .B2(REG1_REG_6__SCAN_IN), .ZN(n3155) );
  OAI21_X1 U3972 ( .B1(n3156), .B2(n4557), .A(n3155), .ZN(U3524) );
  NAND2_X1 U3973 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3172), .ZN(n3162) );
  INV_X1 U3974 ( .A(n3172), .ZN(n4505) );
  INV_X1 U3975 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4747) );
  AOI22_X1 U3976 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3172), .B1(n4505), .B2(
        n4747), .ZN(n4398) );
  NAND2_X1 U3977 ( .A1(n3173), .A2(REG1_REG_9__SCAN_IN), .ZN(n3159) );
  INV_X1 U3978 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4744) );
  INV_X1 U3979 ( .A(n3173), .ZN(n4509) );
  AOI22_X1 U3980 ( .A1(n3173), .A2(REG1_REG_9__SCAN_IN), .B1(n4744), .B2(n4509), .ZN(n4383) );
  INV_X1 U3981 ( .A(n3158), .ZN(n4382) );
  NAND2_X1 U3982 ( .A1(n4383), .A2(n4382), .ZN(n4381) );
  NAND2_X1 U3983 ( .A1(n3159), .A2(n4381), .ZN(n3160) );
  NAND2_X1 U3984 ( .A1(n4506), .A2(n3160), .ZN(n3161) );
  INV_X1 U3985 ( .A(n4506), .ZN(n4392) );
  XNOR2_X1 U3986 ( .A(n3160), .B(n4392), .ZN(n4387) );
  NAND2_X1 U3987 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4387), .ZN(n4386) );
  NAND2_X1 U3988 ( .A1(n3181), .A2(n3163), .ZN(n3164) );
  INV_X1 U3989 ( .A(n3181), .ZN(n4503) );
  NAND2_X1 U3990 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4408), .ZN(n4407) );
  INV_X1 U3991 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3165) );
  NOR2_X1 U3992 ( .A1(n3170), .A2(n3165), .ZN(n3969) );
  AOI21_X1 U3993 ( .B1(n3165), .B2(n3170), .A(n3969), .ZN(n3166) );
  OAI211_X1 U3994 ( .C1(n3167), .C2(n3166), .A(n4452), .B(n3970), .ZN(n3169)
         );
  AND2_X1 U3995 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3443) );
  AOI21_X1 U3996 ( .B1(n4450), .B2(ADDR_REG_13__SCAN_IN), .A(n3443), .ZN(n3168) );
  OAI211_X1 U3997 ( .C1(n4457), .C2(n3170), .A(n3169), .B(n3168), .ZN(n3187)
         );
  INV_X1 U3998 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4777) );
  NOR2_X1 U3999 ( .A1(n3170), .A2(n4777), .ZN(n3981) );
  NAND2_X1 U4000 ( .A1(n3170), .A2(n4777), .ZN(n3980) );
  INV_X1 U4001 ( .A(n3980), .ZN(n3171) );
  NOR2_X1 U4002 ( .A1(n3981), .A2(n3171), .ZN(n3185) );
  NAND2_X1 U4003 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3172), .ZN(n3180) );
  INV_X1 U4004 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4776) );
  AOI22_X1 U4005 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3172), .B1(n4505), .B2(
        n4776), .ZN(n4401) );
  INV_X1 U4006 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4773) );
  AOI22_X1 U4007 ( .A1(n3173), .A2(REG2_REG_9__SCAN_IN), .B1(n4773), .B2(n4509), .ZN(n4376) );
  INV_X1 U4008 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4009 ( .A1(n4506), .A2(n3178), .ZN(n3179) );
  XNOR2_X1 U4010 ( .A(n3178), .B(n4392), .ZN(n4389) );
  NAND2_X1 U4011 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4389), .ZN(n4388) );
  NAND2_X1 U4012 ( .A1(n3179), .A2(n4388), .ZN(n4400) );
  NAND2_X1 U4013 ( .A1(n4401), .A2(n4400), .ZN(n4399) );
  NAND2_X1 U4014 ( .A1(n3180), .A2(n4399), .ZN(n3182) );
  NAND2_X1 U4015 ( .A1(n3181), .A2(n3182), .ZN(n3183) );
  XNOR2_X1 U4016 ( .A(n3182), .B(n4503), .ZN(n4411) );
  NAND2_X1 U4017 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4411), .ZN(n4409) );
  NAND2_X1 U4018 ( .A1(n3183), .A2(n4409), .ZN(n3982) );
  OAI21_X1 U4019 ( .B1(n3185), .B2(n3982), .A(n4410), .ZN(n3184) );
  AOI21_X1 U4020 ( .B1(n3185), .B2(n3982), .A(n3184), .ZN(n3186) );
  OR2_X1 U4021 ( .A1(n3187), .A2(n3186), .ZN(U3253) );
  OAI21_X1 U4022 ( .B1(n3191), .B2(n3189), .A(n3188), .ZN(n3193) );
  NAND2_X1 U4023 ( .A1(n3193), .A2(n3192), .ZN(n3213) );
  NAND2_X1 U4024 ( .A1(n3946), .A2(n2152), .ZN(n3195) );
  NAND2_X1 U4025 ( .A1(n3197), .A2(n2872), .ZN(n3194) );
  NAND2_X1 U4026 ( .A1(n3195), .A2(n3194), .ZN(n3196) );
  XNOR2_X1 U4027 ( .A(n3196), .B(n3585), .ZN(n3199) );
  AND2_X1 U4028 ( .A1(n3197), .A2(n2152), .ZN(n3198) );
  AOI21_X1 U4029 ( .B1(n3946), .B2(n3594), .A(n3198), .ZN(n3200) );
  XNOR2_X1 U4030 ( .A(n3199), .B(n3200), .ZN(n3214) );
  INV_X1 U4031 ( .A(n3199), .ZN(n3201) );
  NOR2_X1 U4032 ( .A1(n3201), .A2(n3200), .ZN(n3202) );
  OAI22_X1 U4033 ( .A1(n3256), .A2(n3562), .B1(n2153), .B2(n3233), .ZN(n3203)
         );
  XNOR2_X1 U4034 ( .A(n3203), .B(n3585), .ZN(n3205) );
  OAI22_X1 U4035 ( .A1(n3256), .A2(n2879), .B1(n3562), .B2(n3233), .ZN(n3204)
         );
  OR2_X1 U4036 ( .A1(n3205), .A2(n3204), .ZN(n3249) );
  NAND2_X1 U4037 ( .A1(n3205), .A2(n3204), .ZN(n3247) );
  NAND2_X1 U4038 ( .A1(n3249), .A2(n3247), .ZN(n3206) );
  XNOR2_X1 U4039 ( .A(n3248), .B(n3206), .ZN(n3212) );
  AOI22_X1 U4040 ( .A1(n3755), .A2(n3238), .B1(n3774), .B2(n3251), .ZN(n3208)
         );
  OAI211_X1 U4041 ( .C1(n3209), .C2(n3769), .A(n3208), .B(n3207), .ZN(n3210)
         );
  AOI21_X1 U4042 ( .B1(n4458), .B2(n3760), .A(n3210), .ZN(n3211) );
  OAI21_X1 U40430 ( .B1(n3212), .B2(n3762), .A(n3211), .ZN(U3218) );
  XNOR2_X1 U4044 ( .A(n3213), .B(n3214), .ZN(n3221) );
  OAI22_X1 U4045 ( .A1(n3772), .A2(n3215), .B1(n3256), .B2(n3758), .ZN(n3216)
         );
  AOI211_X1 U4046 ( .C1(n3754), .C2(n3947), .A(n3217), .B(n3216), .ZN(n3220)
         );
  NAND2_X1 U4047 ( .A1(n3747), .A2(n3218), .ZN(n3219) );
  OAI211_X1 U4048 ( .C1(n3221), .C2(n3762), .A(n3220), .B(n3219), .ZN(U3210)
         );
  NAND2_X1 U4049 ( .A1(n3847), .A2(n3848), .ZN(n3913) );
  XOR2_X1 U4050 ( .A(n3222), .B(n3913), .Z(n3223) );
  AOI222_X1 U4051 ( .A1(n4196), .A2(n3223), .B1(n3305), .B2(n4217), .C1(n3251), 
        .C2(n4476), .ZN(n3345) );
  XNOR2_X1 U4052 ( .A(n3224), .B(n3913), .ZN(n3348) );
  INV_X1 U4053 ( .A(n3225), .ZN(n3226) );
  OAI21_X1 U4054 ( .B1(n3226), .B2(n3346), .A(n3270), .ZN(n3353) );
  AOI22_X1 U4055 ( .A1(n4492), .A2(REG2_REG_10__SCAN_IN), .B1(n3276), .B2(
        n4483), .ZN(n3228) );
  NAND2_X1 U4056 ( .A1(n4033), .A2(n3288), .ZN(n3227) );
  OAI211_X1 U4057 ( .C1(n3353), .C2(n4207), .A(n3228), .B(n3227), .ZN(n3229)
         );
  AOI21_X1 U4058 ( .B1(n3348), .B2(n4156), .A(n3229), .ZN(n3230) );
  OAI21_X1 U4059 ( .B1(n3345), .B2(n4371), .A(n3230), .ZN(U3280) );
  INV_X1 U4060 ( .A(n3231), .ZN(n3232) );
  OAI21_X1 U4061 ( .B1(n3234), .B2(n3233), .A(n3232), .ZN(n4459) );
  INV_X1 U4062 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U4063 ( .A1(n3835), .A2(n3833), .ZN(n3909) );
  XOR2_X1 U4064 ( .A(n3909), .B(n3235), .Z(n4461) );
  XNOR2_X1 U4065 ( .A(n3236), .B(n3909), .ZN(n3237) );
  NAND2_X1 U4066 ( .A1(n3237), .A2(n4196), .ZN(n3240) );
  AOI22_X1 U4067 ( .A1(n3946), .A2(n4476), .B1(n4475), .B2(n3238), .ZN(n3239)
         );
  OAI211_X1 U4068 ( .C1(n3296), .C2(n4479), .A(n3240), .B(n3239), .ZN(n3241)
         );
  AOI21_X1 U4069 ( .B1(n4461), .B2(n4482), .A(n3241), .ZN(n4464) );
  INV_X1 U4070 ( .A(n4464), .ZN(n3242) );
  AOI21_X1 U4071 ( .B1(n4530), .B2(n4461), .A(n3242), .ZN(n3244) );
  MUX2_X1 U4072 ( .A(n4720), .B(n3244), .S(n4545), .Z(n3243) );
  OAI21_X1 U4073 ( .B1(n4459), .B2(n4352), .A(n3243), .ZN(U3483) );
  INV_X1 U4074 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3245) );
  MUX2_X1 U4075 ( .A(n3245), .B(n3244), .S(n4559), .Z(n3246) );
  OAI21_X1 U4076 ( .B1(n4459), .B2(n4300), .A(n3246), .ZN(U3526) );
  NAND2_X1 U4077 ( .A1(n3248), .A2(n3247), .ZN(n3250) );
  NAND2_X1 U4078 ( .A1(n3250), .A2(n3249), .ZN(n3278) );
  NAND2_X1 U4079 ( .A1(n3251), .A2(n2152), .ZN(n3254) );
  NAND2_X1 U4080 ( .A1(n3252), .A2(n2872), .ZN(n3253) );
  NAND2_X1 U4081 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  XNOR2_X1 U4082 ( .A(n3255), .B(n3585), .ZN(n3279) );
  OAI22_X1 U4083 ( .A1(n3296), .A2(n2879), .B1(n3257), .B2(n3562), .ZN(n3280)
         );
  XOR2_X1 U4084 ( .A(n3278), .B(n3277), .Z(n3262) );
  AND2_X1 U4085 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4380) );
  OAI22_X1 U4086 ( .A1(n3772), .A2(n3257), .B1(n3256), .B2(n3769), .ZN(n3258)
         );
  AOI211_X1 U4087 ( .C1(n3774), .C2(n3290), .A(n4380), .B(n3258), .ZN(n3261)
         );
  NAND2_X1 U4088 ( .A1(n3747), .A2(n3259), .ZN(n3260) );
  OAI211_X1 U4089 ( .C1(n3262), .C2(n3762), .A(n3261), .B(n3260), .ZN(U3228)
         );
  XNOR2_X1 U4090 ( .A(n3263), .B(n3908), .ZN(n3264) );
  NAND2_X1 U4091 ( .A1(n3264), .A2(n4196), .ZN(n3266) );
  AOI22_X1 U4092 ( .A1(n4217), .A2(n3944), .B1(n3290), .B2(n4476), .ZN(n3265)
         );
  AND2_X1 U4093 ( .A1(n3266), .A2(n3265), .ZN(n3355) );
  NAND2_X1 U4094 ( .A1(n3267), .A2(n3908), .ZN(n3268) );
  NAND2_X1 U4095 ( .A1(n3269), .A2(n3268), .ZN(n3354) );
  AOI21_X1 U4096 ( .B1(n3271), .B2(n3270), .A(n2186), .ZN(n3362) );
  NAND2_X1 U4097 ( .A1(n3362), .A2(n4488), .ZN(n3273) );
  AOI22_X1 U4098 ( .A1(n4492), .A2(REG2_REG_11__SCAN_IN), .B1(n3323), .B2(
        n4483), .ZN(n3272) );
  OAI211_X1 U4099 ( .C1(n4159), .C2(n3357), .A(n3273), .B(n3272), .ZN(n3274)
         );
  AOI21_X1 U4100 ( .B1(n3354), .B2(n4156), .A(n3274), .ZN(n3275) );
  OAI21_X1 U4101 ( .B1(n4371), .B2(n3355), .A(n3275), .ZN(U3279) );
  INV_X1 U4102 ( .A(n3276), .ZN(n3300) );
  NAND2_X1 U4103 ( .A1(n3278), .A2(n3277), .ZN(n3284) );
  NAND2_X1 U4104 ( .A1(n3284), .A2(n3283), .ZN(n3291) );
  NAND2_X1 U4105 ( .A1(n3290), .A2(n2152), .ZN(n3286) );
  NAND2_X1 U4106 ( .A1(n3288), .A2(n2872), .ZN(n3285) );
  NAND2_X1 U4107 ( .A1(n3286), .A2(n3285), .ZN(n3287) );
  XNOR2_X1 U4108 ( .A(n3287), .B(n3585), .ZN(n3316) );
  AND2_X1 U4109 ( .A1(n3288), .A2(n2152), .ZN(n3289) );
  AOI21_X1 U4110 ( .B1(n3290), .B2(n3594), .A(n3289), .ZN(n3314) );
  XOR2_X1 U4111 ( .A(n3316), .B(n3314), .Z(n3292) );
  AOI21_X1 U4112 ( .B1(n3291), .B2(n3292), .A(n3762), .ZN(n3295) );
  INV_X1 U4113 ( .A(n3291), .ZN(n3294) );
  NAND2_X1 U4114 ( .A1(n3295), .A2(n3318), .ZN(n3299) );
  NOR2_X1 U4115 ( .A1(STATE_REG_SCAN_IN), .A2(n4635), .ZN(n4394) );
  OAI22_X1 U4116 ( .A1(n3772), .A2(n3346), .B1(n3296), .B2(n3769), .ZN(n3297)
         );
  AOI211_X1 U4117 ( .C1(n3774), .C2(n3305), .A(n4394), .B(n3297), .ZN(n3298)
         );
  OAI211_X1 U4118 ( .C1(n3778), .C2(n3300), .A(n3299), .B(n3298), .ZN(U3214)
         );
  NAND2_X1 U4119 ( .A1(n3302), .A2(n3301), .ZN(n3333) );
  NAND2_X1 U4120 ( .A1(n3330), .A2(n3331), .ZN(n3892) );
  INV_X1 U4121 ( .A(n3892), .ZN(n3303) );
  XNOR2_X1 U4122 ( .A(n3333), .B(n3303), .ZN(n3304) );
  NAND2_X1 U4123 ( .A1(n3304), .A2(n4196), .ZN(n3307) );
  AOI22_X1 U4124 ( .A1(n4476), .A2(n3305), .B1(n3637), .B2(n4217), .ZN(n3306)
         );
  AND2_X1 U4125 ( .A1(n3307), .A2(n3306), .ZN(n3365) );
  XNOR2_X1 U4126 ( .A(n3308), .B(n3892), .ZN(n3364) );
  NOR2_X1 U4127 ( .A1(n2186), .A2(n3388), .ZN(n3309) );
  OR2_X1 U4128 ( .A1(n3339), .A2(n3309), .ZN(n3372) );
  AOI22_X1 U4129 ( .A1(n4492), .A2(REG2_REG_12__SCAN_IN), .B1(n3390), .B2(
        n4483), .ZN(n3311) );
  NAND2_X1 U4130 ( .A1(n4033), .A2(n3379), .ZN(n3310) );
  OAI211_X1 U4131 ( .C1(n3372), .C2(n4207), .A(n3311), .B(n3310), .ZN(n3312)
         );
  AOI21_X1 U4132 ( .B1(n3364), .B2(n4156), .A(n3312), .ZN(n3313) );
  OAI21_X1 U4133 ( .B1(n4371), .B2(n3365), .A(n3313), .ZN(U3278) );
  INV_X1 U4134 ( .A(n3314), .ZN(n3315) );
  NAND2_X1 U4135 ( .A1(n3316), .A2(n3315), .ZN(n3317) );
  OAI22_X1 U4136 ( .A1(n3387), .A2(n2879), .B1(n3562), .B2(n3357), .ZN(n3374)
         );
  OAI22_X1 U4137 ( .A1(n3387), .A2(n3562), .B1(n2154), .B2(n3357), .ZN(n3319)
         );
  XNOR2_X1 U4138 ( .A(n3319), .B(n3585), .ZN(n3373) );
  XOR2_X1 U4139 ( .A(n3374), .B(n3373), .Z(n3320) );
  XNOR2_X1 U4140 ( .A(n3375), .B(n3320), .ZN(n3326) );
  AND2_X1 U4141 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4405) );
  OAI22_X1 U4142 ( .A1(n3772), .A2(n3357), .B1(n3321), .B2(n3769), .ZN(n3322)
         );
  AOI211_X1 U4143 ( .C1(n3774), .C2(n3944), .A(n4405), .B(n3322), .ZN(n3325)
         );
  NAND2_X1 U4144 ( .A1(n3747), .A2(n3323), .ZN(n3324) );
  OAI211_X1 U4145 ( .C1(n3326), .C2(n3762), .A(n3325), .B(n3324), .ZN(U3233)
         );
  INV_X1 U4146 ( .A(n3327), .ZN(n3329) );
  OR2_X1 U4147 ( .A1(n3329), .A2(n3328), .ZN(n3897) );
  XNOR2_X1 U4148 ( .A(n3402), .B(n3897), .ZN(n3395) );
  INV_X1 U4149 ( .A(n3395), .ZN(n3344) );
  INV_X1 U4150 ( .A(n3330), .ZN(n3332) );
  OAI21_X1 U4151 ( .B1(n3333), .B2(n3332), .A(n3331), .ZN(n3334) );
  XNOR2_X1 U4152 ( .A(n3334), .B(n3897), .ZN(n3335) );
  NAND2_X1 U4153 ( .A1(n3335), .A2(n4196), .ZN(n3337) );
  AOI22_X1 U4154 ( .A1(n3497), .A2(n4217), .B1(n4475), .B2(n3439), .ZN(n3336)
         );
  OAI211_X1 U4155 ( .C1(n3338), .C2(n4220), .A(n3337), .B(n3336), .ZN(n3394)
         );
  OR2_X1 U4156 ( .A1(n3339), .A2(n3441), .ZN(n3340) );
  NAND2_X1 U4157 ( .A1(n3412), .A2(n3340), .ZN(n3400) );
  AOI22_X1 U4158 ( .A1(n4492), .A2(REG2_REG_13__SCAN_IN), .B1(n3444), .B2(
        n4483), .ZN(n3341) );
  OAI21_X1 U4159 ( .B1(n3400), .B2(n4207), .A(n3341), .ZN(n3342) );
  AOI21_X1 U4160 ( .B1(n3394), .B2(n4232), .A(n3342), .ZN(n3343) );
  OAI21_X1 U4161 ( .B1(n3344), .B2(n4235), .A(n3343), .ZN(U3277) );
  INV_X1 U4162 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4731) );
  OAI21_X1 U4163 ( .B1(n3346), .B2(n4294), .A(n3345), .ZN(n3347) );
  AOI21_X1 U4164 ( .B1(n4542), .B2(n3348), .A(n3347), .ZN(n3350) );
  MUX2_X1 U4165 ( .A(n4731), .B(n3350), .S(n4545), .Z(n3349) );
  OAI21_X1 U4166 ( .B1(n3353), .B2(n4352), .A(n3349), .ZN(U3487) );
  INV_X1 U4167 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3351) );
  MUX2_X1 U4168 ( .A(n3351), .B(n3350), .S(n4559), .Z(n3352) );
  OAI21_X1 U4169 ( .B1(n3353), .B2(n4300), .A(n3352), .ZN(U3528) );
  NAND2_X1 U4170 ( .A1(n3354), .A2(n4542), .ZN(n3356) );
  OAI211_X1 U4171 ( .C1(n4294), .C2(n3357), .A(n3356), .B(n3355), .ZN(n3360)
         );
  MUX2_X1 U4172 ( .A(REG0_REG_11__SCAN_IN), .B(n3360), .S(n4545), .Z(n3358) );
  AOI21_X1 U4173 ( .B1(n3362), .B2(n4525), .A(n3358), .ZN(n3359) );
  INV_X1 U4174 ( .A(n3359), .ZN(U3489) );
  MUX2_X1 U4175 ( .A(REG1_REG_11__SCAN_IN), .B(n3360), .S(n4559), .Z(n3361) );
  AOI21_X1 U4176 ( .B1(n4549), .B2(n3362), .A(n3361), .ZN(n3363) );
  INV_X1 U4177 ( .A(n3363), .ZN(U3529) );
  NAND2_X1 U4178 ( .A1(n3364), .A2(n4542), .ZN(n3366) );
  OAI211_X1 U4179 ( .C1(n4294), .C2(n3388), .A(n3366), .B(n3365), .ZN(n3369)
         );
  MUX2_X1 U4180 ( .A(REG1_REG_12__SCAN_IN), .B(n3369), .S(n4559), .Z(n3367) );
  INV_X1 U4181 ( .A(n3367), .ZN(n3368) );
  OAI21_X1 U4182 ( .B1(n4300), .B2(n3372), .A(n3368), .ZN(U3530) );
  MUX2_X1 U4183 ( .A(REG0_REG_12__SCAN_IN), .B(n3369), .S(n4545), .Z(n3370) );
  INV_X1 U4184 ( .A(n3370), .ZN(n3371) );
  OAI21_X1 U4185 ( .B1(n3372), .B2(n4352), .A(n3371), .ZN(U3491) );
  NAND2_X1 U4186 ( .A1(n3944), .A2(n2152), .ZN(n3377) );
  NAND2_X1 U4187 ( .A1(n3379), .A2(n2872), .ZN(n3376) );
  NAND2_X1 U4188 ( .A1(n3377), .A2(n3376), .ZN(n3378) );
  XNOR2_X1 U4189 ( .A(n3378), .B(n3585), .ZN(n3382) );
  NAND2_X1 U4190 ( .A1(n3944), .A2(n3594), .ZN(n3381) );
  NAND2_X1 U4191 ( .A1(n3379), .A2(n2152), .ZN(n3380) );
  NAND2_X1 U4192 ( .A1(n3381), .A2(n3380), .ZN(n3383) );
  NAND2_X1 U4193 ( .A1(n3382), .A2(n3383), .ZN(n3434) );
  INV_X1 U4194 ( .A(n3382), .ZN(n3385) );
  INV_X1 U4195 ( .A(n3383), .ZN(n3384) );
  NAND2_X1 U4196 ( .A1(n3385), .A2(n3384), .ZN(n3436) );
  NAND2_X1 U4197 ( .A1(n3434), .A2(n3436), .ZN(n3386) );
  XNOR2_X1 U4198 ( .A(n3435), .B(n3386), .ZN(n3393) );
  INV_X1 U4199 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4640) );
  NOR2_X1 U4200 ( .A1(STATE_REG_SCAN_IN), .A2(n4640), .ZN(n4415) );
  OAI22_X1 U4201 ( .A1(n3772), .A2(n3388), .B1(n3387), .B2(n3769), .ZN(n3389)
         );
  AOI211_X1 U4202 ( .C1(n3774), .C2(n3637), .A(n4415), .B(n3389), .ZN(n3392)
         );
  NAND2_X1 U4203 ( .A1(n3747), .A2(n3390), .ZN(n3391) );
  OAI211_X1 U4204 ( .C1(n3393), .C2(n3762), .A(n3392), .B(n3391), .ZN(U3221)
         );
  INV_X1 U4205 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3396) );
  AOI21_X1 U4206 ( .B1(n4542), .B2(n3395), .A(n3394), .ZN(n3398) );
  MUX2_X1 U4207 ( .A(n3396), .B(n3398), .S(n4545), .Z(n3397) );
  OAI21_X1 U4208 ( .B1(n3400), .B2(n4352), .A(n3397), .ZN(U3493) );
  MUX2_X1 U4209 ( .A(n3165), .B(n3398), .S(n4559), .Z(n3399) );
  OAI21_X1 U4210 ( .B1(n4300), .B2(n3400), .A(n3399), .ZN(U3531) );
  OR2_X1 U4211 ( .A1(n3402), .A2(n3401), .ZN(n3405) );
  AND2_X1 U4212 ( .A1(n3405), .A2(n3403), .ZN(n3407) );
  NAND2_X1 U4213 ( .A1(n3405), .A2(n3404), .ZN(n3406) );
  OAI21_X1 U4214 ( .B1(n3407), .B2(n3916), .A(n3406), .ZN(n3464) );
  INV_X1 U4215 ( .A(n3464), .ZN(n3419) );
  AOI22_X1 U4216 ( .A1(n4217), .A2(n3943), .B1(n3637), .B2(n4476), .ZN(n3411)
         );
  OAI21_X1 U4217 ( .B1(n3408), .B2(n3785), .A(n3421), .ZN(n3409) );
  NAND2_X1 U4218 ( .A1(n3409), .A2(n4196), .ZN(n3410) );
  OAI211_X1 U4219 ( .C1(n3419), .C2(n4174), .A(n3411), .B(n3410), .ZN(n3462)
         );
  NAND2_X1 U4220 ( .A1(n3462), .A2(n4232), .ZN(n3418) );
  INV_X1 U4221 ( .A(n3412), .ZN(n3413) );
  OAI21_X1 U4222 ( .B1(n3413), .B2(n3461), .A(n3427), .ZN(n3470) );
  INV_X1 U4223 ( .A(n3470), .ZN(n3416) );
  AOI22_X1 U4224 ( .A1(n4492), .A2(REG2_REG_14__SCAN_IN), .B1(n3644), .B2(
        n4483), .ZN(n3414) );
  OAI21_X1 U4225 ( .B1(n4159), .B2(n3461), .A(n3414), .ZN(n3415) );
  AOI21_X1 U4226 ( .B1(n3416), .B2(n4488), .A(n3415), .ZN(n3417) );
  OAI211_X1 U4227 ( .C1(n3419), .C2(n4183), .A(n3418), .B(n3417), .ZN(U3276)
         );
  XNOR2_X1 U4228 ( .A(n3420), .B(n3422), .ZN(n3480) );
  INV_X1 U4229 ( .A(n3480), .ZN(n3433) );
  NAND2_X1 U4230 ( .A1(n3421), .A2(n3781), .ZN(n3423) );
  INV_X1 U4231 ( .A(n3422), .ZN(n3921) );
  XNOR2_X1 U4232 ( .A(n3423), .B(n3921), .ZN(n3424) );
  NAND2_X1 U4233 ( .A1(n3424), .A2(n4196), .ZN(n3426) );
  AOI22_X1 U4234 ( .A1(n3942), .A2(n4217), .B1(n4475), .B2(n3511), .ZN(n3425)
         );
  OAI211_X1 U4235 ( .C1(n3770), .C2(n4220), .A(n3426), .B(n3425), .ZN(n3479)
         );
  INV_X1 U4236 ( .A(n3456), .ZN(n3428) );
  OAI21_X1 U4237 ( .B1(n2267), .B2(n3771), .A(n3428), .ZN(n3485) );
  AOI22_X1 U4238 ( .A1(n4371), .A2(REG2_REG_15__SCAN_IN), .B1(n3429), .B2(
        n4483), .ZN(n3430) );
  OAI21_X1 U4239 ( .B1(n3485), .B2(n4207), .A(n3430), .ZN(n3431) );
  AOI21_X1 U4240 ( .B1(n3479), .B2(n4232), .A(n3431), .ZN(n3432) );
  OAI21_X1 U4241 ( .B1(n3433), .B2(n4235), .A(n3432), .ZN(U3275) );
  NAND2_X1 U4242 ( .A1(n3435), .A2(n3434), .ZN(n3437) );
  AOI22_X1 U4243 ( .A1(n3637), .A2(n2152), .B1(n2872), .B2(n3439), .ZN(n3438)
         );
  XNOR2_X1 U4244 ( .A(n3438), .B(n3585), .ZN(n3491) );
  AOI22_X1 U4245 ( .A1(n3637), .A2(n3594), .B1(n2152), .B2(n3439), .ZN(n3492)
         );
  XNOR2_X1 U4246 ( .A(n3491), .B(n3492), .ZN(n3440) );
  XNOR2_X1 U4247 ( .A(n3490), .B(n3440), .ZN(n3447) );
  OAI22_X1 U4248 ( .A1(n3772), .A2(n3441), .B1(n3770), .B2(n3758), .ZN(n3442)
         );
  AOI211_X1 U4249 ( .C1(n3754), .C2(n3944), .A(n3443), .B(n3442), .ZN(n3446)
         );
  NAND2_X1 U4250 ( .A1(n3747), .A2(n3444), .ZN(n3445) );
  OAI211_X1 U4251 ( .C1(n3447), .C2(n3762), .A(n3446), .B(n3445), .ZN(U3231)
         );
  OAI21_X1 U4252 ( .B1(n2156), .B2(n2576), .A(n3449), .ZN(n4305) );
  XNOR2_X1 U4253 ( .A(n3450), .B(n2576), .ZN(n3454) );
  NAND2_X1 U4254 ( .A1(n3693), .A2(n4475), .ZN(n3452) );
  NAND2_X1 U4255 ( .A1(n3943), .A2(n4476), .ZN(n3451) );
  OAI211_X1 U4256 ( .C1(n4221), .C2(n4479), .A(n3452), .B(n3451), .ZN(n3453)
         );
  AOI21_X1 U4257 ( .B1(n3454), .B2(n4196), .A(n3453), .ZN(n4304) );
  AOI22_X1 U4258 ( .A1(n4492), .A2(REG2_REG_16__SCAN_IN), .B1(n3698), .B2(
        n4483), .ZN(n3458) );
  OR2_X1 U4259 ( .A1(n3456), .A2(n3455), .ZN(n4302) );
  NAND3_X1 U4260 ( .A1(n4301), .A2(n4302), .A3(n4488), .ZN(n3457) );
  OAI211_X1 U4261 ( .C1(n4304), .C2(n4371), .A(n3458), .B(n3457), .ZN(n3459)
         );
  INV_X1 U4262 ( .A(n3459), .ZN(n3460) );
  OAI21_X1 U4263 ( .B1(n4305), .B2(n4235), .A(n3460), .ZN(U3274) );
  INV_X1 U4264 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3465) );
  NOR2_X1 U4265 ( .A1(n3461), .A2(n4294), .ZN(n3463) );
  AOI211_X1 U4266 ( .C1(n4530), .C2(n3464), .A(n3463), .B(n3462), .ZN(n3467)
         );
  MUX2_X1 U4267 ( .A(n3465), .B(n3467), .S(n4545), .Z(n3466) );
  OAI21_X1 U4268 ( .B1(n3470), .B2(n4352), .A(n3466), .ZN(U3495) );
  INV_X1 U4269 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3468) );
  MUX2_X1 U4270 ( .A(n3468), .B(n3467), .S(n4559), .Z(n3469) );
  OAI21_X1 U4271 ( .B1(n4300), .B2(n3470), .A(n3469), .ZN(U3532) );
  NAND2_X1 U4272 ( .A1(n4188), .A2(n3862), .ZN(n3912) );
  XOR2_X1 U4273 ( .A(n3912), .B(n3471), .Z(n3472) );
  AOI222_X1 U4274 ( .A1(n4196), .A2(n3472), .B1(n3941), .B2(n4217), .C1(n3942), 
        .C2(n4476), .ZN(n4293) );
  XOR2_X1 U4275 ( .A(n3912), .B(n3473), .Z(n4297) );
  NAND2_X1 U4276 ( .A1(n4297), .A2(n4156), .ZN(n3478) );
  OAI21_X1 U4277 ( .B1(n2263), .B2(n4295), .A(n4224), .ZN(n4353) );
  INV_X1 U4278 ( .A(n4353), .ZN(n3476) );
  AOI22_X1 U4279 ( .A1(n4492), .A2(REG2_REG_17__SCAN_IN), .B1(n3706), .B2(
        n4483), .ZN(n3474) );
  OAI21_X1 U4280 ( .B1(n4159), .B2(n4295), .A(n3474), .ZN(n3475) );
  AOI21_X1 U4281 ( .B1(n3476), .B2(n4488), .A(n3475), .ZN(n3477) );
  OAI211_X1 U4282 ( .C1(n4371), .C2(n4293), .A(n3478), .B(n3477), .ZN(U3273)
         );
  AOI21_X1 U4283 ( .B1(n3480), .B2(n4542), .A(n3479), .ZN(n3483) );
  MUX2_X1 U4284 ( .A(n3483), .B(n4748), .S(n4557), .Z(n3481) );
  OAI21_X1 U4285 ( .B1(n4300), .B2(n3485), .A(n3481), .ZN(U3533) );
  INV_X1 U4286 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3482) );
  MUX2_X1 U4287 ( .A(n3483), .B(n3482), .S(n4544), .Z(n3484) );
  OAI21_X1 U4288 ( .B1(n3485), .B2(n4352), .A(n3484), .ZN(U3497) );
  OAI22_X1 U4289 ( .A1(n4040), .A2(n3562), .B1(n4245), .B2(n2154), .ZN(n3486)
         );
  XNOR2_X1 U4290 ( .A(n3486), .B(n2884), .ZN(n3488) );
  OAI22_X1 U4291 ( .A1(n4040), .A2(n2879), .B1(n4245), .B2(n3562), .ZN(n3487)
         );
  XNOR2_X1 U4292 ( .A(n3488), .B(n3487), .ZN(n3607) );
  INV_X1 U4293 ( .A(n3607), .ZN(n3489) );
  NAND2_X1 U4294 ( .A1(n3489), .A2(n3767), .ZN(n3616) );
  NAND2_X1 U4295 ( .A1(n3497), .A2(n2152), .ZN(n3494) );
  NAND2_X1 U4296 ( .A1(n3638), .A2(n2872), .ZN(n3493) );
  NAND2_X1 U4297 ( .A1(n3494), .A2(n3493), .ZN(n3495) );
  XNOR2_X1 U4298 ( .A(n3495), .B(n2884), .ZN(n3499) );
  AND2_X1 U4299 ( .A1(n3638), .A2(n2152), .ZN(n3496) );
  AOI21_X1 U4300 ( .B1(n3497), .B2(n3594), .A(n3496), .ZN(n3498) );
  NOR2_X1 U4301 ( .A1(n3499), .A2(n3498), .ZN(n3635) );
  NAND2_X1 U4302 ( .A1(n3499), .A2(n3498), .ZN(n3633) );
  OAI22_X1 U4303 ( .A1(n3696), .A2(n3562), .B1(n2153), .B2(n3771), .ZN(n3500)
         );
  XOR2_X1 U4304 ( .A(n3585), .B(n3500), .Z(n3509) );
  NOR2_X1 U4305 ( .A1(n3510), .A2(n3509), .ZN(n3689) );
  NAND2_X1 U4306 ( .A1(n3942), .A2(n2152), .ZN(n3502) );
  NAND2_X1 U4307 ( .A1(n3693), .A2(n2872), .ZN(n3501) );
  NAND2_X1 U4308 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  XNOR2_X1 U4309 ( .A(n3503), .B(n3585), .ZN(n3507) );
  NAND2_X1 U4310 ( .A1(n3942), .A2(n3594), .ZN(n3505) );
  NAND2_X1 U4311 ( .A1(n3693), .A2(n2152), .ZN(n3504) );
  NAND2_X1 U4312 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  NOR2_X1 U4313 ( .A1(n3507), .A2(n3506), .ZN(n3516) );
  AOI21_X1 U4314 ( .B1(n3507), .B2(n3506), .A(n3516), .ZN(n3692) );
  NAND2_X1 U4315 ( .A1(n3510), .A2(n3509), .ZN(n3690) );
  NAND2_X1 U4316 ( .A1(n3943), .A2(n3594), .ZN(n3513) );
  NAND2_X1 U4317 ( .A1(n3511), .A2(n2152), .ZN(n3512) );
  NAND2_X1 U4318 ( .A1(n3513), .A2(n3512), .ZN(n3765) );
  NAND2_X1 U4319 ( .A1(n3690), .A2(n3765), .ZN(n3514) );
  NAND2_X1 U4320 ( .A1(n3515), .A2(n3514), .ZN(n3518) );
  INV_X1 U4321 ( .A(n3516), .ZN(n3517) );
  NAND2_X1 U4322 ( .A1(n3518), .A2(n3517), .ZN(n3701) );
  OAI22_X1 U4323 ( .A1(n4221), .A2(n3562), .B1(n2154), .B2(n4295), .ZN(n3519)
         );
  XNOR2_X1 U4324 ( .A(n3519), .B(n3585), .ZN(n3520) );
  OAI22_X1 U4325 ( .A1(n4221), .A2(n2879), .B1(n3562), .B2(n4295), .ZN(n3521)
         );
  NAND2_X1 U4326 ( .A1(n3520), .A2(n3521), .ZN(n3702) );
  NAND2_X1 U4327 ( .A1(n3701), .A2(n3702), .ZN(n3524) );
  INV_X1 U4328 ( .A(n3520), .ZN(n3523) );
  INV_X1 U4329 ( .A(n3521), .ZN(n3522) );
  NAND2_X1 U4330 ( .A1(n3523), .A2(n3522), .ZN(n3703) );
  NAND2_X1 U4331 ( .A1(n4218), .A2(n2152), .ZN(n3526) );
  NAND2_X1 U4332 ( .A1(n4198), .A2(n2872), .ZN(n3525) );
  NAND2_X1 U4333 ( .A1(n3526), .A2(n3525), .ZN(n3527) );
  XNOR2_X1 U4334 ( .A(n3527), .B(n3585), .ZN(n3539) );
  NAND2_X1 U4335 ( .A1(n4218), .A2(n3594), .ZN(n3529) );
  NAND2_X1 U4336 ( .A1(n4198), .A2(n2152), .ZN(n3528) );
  NAND2_X1 U4337 ( .A1(n3529), .A2(n3528), .ZN(n3538) );
  NAND2_X1 U4338 ( .A1(n3539), .A2(n3538), .ZN(n3537) );
  NAND2_X1 U4339 ( .A1(n3941), .A2(n2152), .ZN(n3531) );
  NAND2_X1 U4340 ( .A1(n4216), .A2(n2872), .ZN(n3530) );
  NAND2_X1 U4341 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  XNOR2_X1 U4342 ( .A(n3532), .B(n2884), .ZN(n3742) );
  NAND2_X1 U4343 ( .A1(n3941), .A2(n3594), .ZN(n3534) );
  NAND2_X1 U4344 ( .A1(n4216), .A2(n2152), .ZN(n3533) );
  NAND2_X1 U4345 ( .A1(n3656), .A2(n2178), .ZN(n3542) );
  INV_X1 U4346 ( .A(n3537), .ZN(n3660) );
  INV_X1 U4347 ( .A(n3741), .ZN(n3657) );
  NOR3_X1 U4348 ( .A1(n3660), .A2(n3657), .A3(n3535), .ZN(n3540) );
  NOR2_X1 U4349 ( .A1(n3539), .A2(n3538), .ZN(n3661) );
  NOR2_X1 U4350 ( .A1(n3540), .A2(n3661), .ZN(n3541) );
  NAND2_X1 U4351 ( .A1(n4199), .A2(n2152), .ZN(n3544) );
  NAND2_X1 U4352 ( .A1(n4180), .A2(n2872), .ZN(n3543) );
  NAND2_X1 U4353 ( .A1(n3544), .A2(n3543), .ZN(n3545) );
  XNOR2_X1 U4354 ( .A(n3545), .B(n3585), .ZN(n3548) );
  NAND2_X1 U4355 ( .A1(n4199), .A2(n3594), .ZN(n3547) );
  NAND2_X1 U4356 ( .A1(n4180), .A2(n2152), .ZN(n3546) );
  NAND2_X1 U4357 ( .A1(n3547), .A2(n3546), .ZN(n3549) );
  NAND2_X1 U4358 ( .A1(n3548), .A2(n3549), .ZN(n3722) );
  INV_X1 U4359 ( .A(n3548), .ZN(n3551) );
  INV_X1 U4360 ( .A(n3549), .ZN(n3550) );
  NAND2_X1 U4361 ( .A1(n3551), .A2(n3550), .ZN(n3724) );
  NAND2_X1 U4362 ( .A1(n4167), .A2(n2152), .ZN(n3553) );
  NAND2_X1 U4363 ( .A1(n3555), .A2(n2872), .ZN(n3552) );
  NAND2_X1 U4364 ( .A1(n3553), .A2(n3552), .ZN(n3554) );
  XNOR2_X1 U4365 ( .A(n3554), .B(n2884), .ZN(n3557) );
  AND2_X1 U4366 ( .A1(n3555), .A2(n2152), .ZN(n3556) );
  AOI21_X1 U4367 ( .B1(n4167), .B2(n3594), .A(n3556), .ZN(n3558) );
  INV_X1 U4368 ( .A(n3557), .ZN(n3560) );
  INV_X1 U4369 ( .A(n3558), .ZN(n3559) );
  NAND2_X1 U4370 ( .A1(n3560), .A2(n3559), .ZN(n3668) );
  OAI22_X1 U4371 ( .A1(n3674), .A2(n3562), .B1(n4140), .B2(n2153), .ZN(n3561)
         );
  XNOR2_X1 U4372 ( .A(n3561), .B(n3585), .ZN(n3565) );
  OAI22_X1 U4373 ( .A1(n3674), .A2(n2879), .B1(n4140), .B2(n3562), .ZN(n3564)
         );
  XNOR2_X1 U4374 ( .A(n3565), .B(n3564), .ZN(n3734) );
  NOR2_X1 U4375 ( .A1(n3565), .A2(n3564), .ZN(n3649) );
  NAND2_X1 U4376 ( .A1(n4137), .A2(n2152), .ZN(n3567) );
  OR2_X1 U4377 ( .A1(n4123), .A2(n2153), .ZN(n3566) );
  NAND2_X1 U4378 ( .A1(n3567), .A2(n3566), .ZN(n3568) );
  XNOR2_X1 U4379 ( .A(n3568), .B(n2884), .ZN(n3571) );
  NOR2_X1 U4380 ( .A1(n4123), .A2(n3562), .ZN(n3569) );
  AOI21_X1 U4381 ( .B1(n4137), .B2(n3594), .A(n3569), .ZN(n3572) );
  XNOR2_X1 U4382 ( .A(n3571), .B(n3572), .ZN(n3648) );
  NOR2_X1 U4383 ( .A1(n3649), .A2(n3648), .ZN(n3570) );
  INV_X1 U4384 ( .A(n3571), .ZN(n3574) );
  INV_X1 U4385 ( .A(n3572), .ZN(n3573) );
  NAND2_X1 U4386 ( .A1(n3574), .A2(n3573), .ZN(n3579) );
  NAND2_X1 U4387 ( .A1(n3650), .A2(n3579), .ZN(n3577) );
  AOI22_X1 U4388 ( .A1(n4079), .A2(n3594), .B1(n2152), .B2(n3575), .ZN(n3578)
         );
  INV_X1 U4389 ( .A(n3578), .ZN(n3576) );
  OAI22_X1 U4390 ( .A1(n4126), .A2(n3562), .B1(n2153), .B2(n4262), .ZN(n3581)
         );
  XNOR2_X1 U4391 ( .A(n3581), .B(n3585), .ZN(n3713) );
  NAND2_X1 U4392 ( .A1(n3710), .A2(n3713), .ZN(n3582) );
  NOR2_X1 U4393 ( .A1(n4084), .A2(n2154), .ZN(n3583) );
  AOI21_X1 U4394 ( .B1(n4095), .B2(n2152), .A(n3583), .ZN(n3586) );
  XNOR2_X1 U4395 ( .A(n3586), .B(n3585), .ZN(n3589) );
  NOR2_X1 U4396 ( .A1(n4084), .A2(n3562), .ZN(n3587) );
  AOI21_X1 U4397 ( .B1(n4095), .B2(n3594), .A(n3587), .ZN(n3588) );
  NAND2_X1 U4398 ( .A1(n3589), .A2(n3588), .ZN(n3681) );
  NOR2_X1 U4399 ( .A1(n3589), .A2(n3588), .ZN(n3682) );
  NAND2_X1 U4400 ( .A1(n4038), .A2(n2152), .ZN(n3591) );
  OR2_X1 U4401 ( .A1(n4066), .A2(n2154), .ZN(n3590) );
  NAND2_X1 U4402 ( .A1(n3591), .A2(n3590), .ZN(n3592) );
  XNOR2_X1 U4403 ( .A(n3592), .B(n2884), .ZN(n3596) );
  NOR2_X1 U4404 ( .A1(n4066), .A2(n3562), .ZN(n3593) );
  AOI21_X1 U4405 ( .B1(n4038), .B2(n3594), .A(n3593), .ZN(n3595) );
  OR2_X1 U4406 ( .A1(n3596), .A2(n3595), .ZN(n3751) );
  OAI22_X1 U4407 ( .A1(n4064), .A2(n3562), .B1(n2153), .B2(n4249), .ZN(n3598)
         );
  XNOR2_X1 U4408 ( .A(n3598), .B(n2884), .ZN(n3602) );
  OR2_X1 U4409 ( .A1(n4064), .A2(n2879), .ZN(n3601) );
  NAND2_X1 U4410 ( .A1(n3599), .A2(n2152), .ZN(n3600) );
  NAND2_X1 U4411 ( .A1(n3601), .A2(n3600), .ZN(n3603) );
  XNOR2_X1 U4412 ( .A(n3602), .B(n3603), .ZN(n3625) );
  INV_X1 U4413 ( .A(n3602), .ZN(n3604) );
  NAND2_X1 U4414 ( .A1(n3604), .A2(n3603), .ZN(n3608) );
  NOR3_X1 U4415 ( .A1(n3608), .A2(n3607), .A3(n3762), .ZN(n3612) );
  AOI22_X1 U4416 ( .A1(n3940), .A2(n3754), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3610) );
  AOI22_X1 U4417 ( .A1(n3755), .A2(n4034), .B1(n3797), .B2(n3774), .ZN(n3609)
         );
  OAI211_X1 U4418 ( .C1(n3778), .C2(n4028), .A(n3610), .B(n3609), .ZN(n3611)
         );
  NOR2_X1 U4419 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  OAI211_X1 U4420 ( .C1(n3616), .C2(n3615), .A(n3614), .B(n3613), .ZN(U3217)
         );
  INV_X1 U4421 ( .A(n3617), .ZN(n3621) );
  OAI22_X1 U4422 ( .A1(n3619), .A2(n4207), .B1(n3618), .B2(n4114), .ZN(n3620)
         );
  OAI21_X1 U4423 ( .B1(n3621), .B2(n3620), .A(n4232), .ZN(n3623) );
  NAND2_X1 U4424 ( .A1(n4371), .A2(REG2_REG_29__SCAN_IN), .ZN(n3622) );
  OAI211_X1 U4425 ( .C1(n3624), .C2(n4235), .A(n3623), .B(n3622), .ZN(U3354)
         );
  XNOR2_X1 U4426 ( .A(n3626), .B(n3625), .ZN(n3631) );
  OAI22_X1 U4427 ( .A1(n4040), .A2(n3758), .B1(STATE_REG_SCAN_IN), .B2(n3627), 
        .ZN(n3629) );
  OAI22_X1 U4428 ( .A1(n4082), .A2(n3769), .B1(n3772), .B2(n4249), .ZN(n3628)
         );
  AOI211_X1 U4429 ( .C1(n4048), .C2(n3747), .A(n3629), .B(n3628), .ZN(n3630)
         );
  OAI21_X1 U4430 ( .B1(n3631), .B2(n3762), .A(n3630), .ZN(U3211) );
  INV_X1 U4431 ( .A(n3633), .ZN(n3634) );
  NOR2_X1 U4432 ( .A1(n3635), .A2(n3634), .ZN(n3636) );
  XNOR2_X1 U4433 ( .A(n3632), .B(n3636), .ZN(n3646) );
  INV_X1 U4434 ( .A(n3637), .ZN(n3642) );
  AOI22_X1 U4435 ( .A1(n3755), .A2(n3638), .B1(n3774), .B2(n3943), .ZN(n3641)
         );
  NOR2_X1 U4436 ( .A1(n3639), .A2(STATE_REG_SCAN_IN), .ZN(n4421) );
  INV_X1 U4437 ( .A(n4421), .ZN(n3640) );
  OAI211_X1 U4438 ( .C1(n3642), .C2(n3769), .A(n3641), .B(n3640), .ZN(n3643)
         );
  AOI21_X1 U4439 ( .B1(n3644), .B2(n3747), .A(n3643), .ZN(n3645) );
  OAI21_X1 U4440 ( .B1(n3646), .B2(n3762), .A(n3645), .ZN(U3212) );
  INV_X1 U4441 ( .A(n3647), .ZN(n3732) );
  OAI21_X1 U4442 ( .B1(n3732), .B2(n3649), .A(n3648), .ZN(n3651) );
  NAND3_X1 U4443 ( .A1(n3651), .A2(n3767), .A3(n3650), .ZN(n3655) );
  OAI22_X1 U4444 ( .A1(n4126), .A2(n3758), .B1(STATE_REG_SCAN_IN), .B2(n4636), 
        .ZN(n3653) );
  OAI22_X1 U4445 ( .A1(n3772), .A2(n4123), .B1(n3674), .B2(n3769), .ZN(n3652)
         );
  AOI211_X1 U4446 ( .C1(n3747), .C2(n4113), .A(n3653), .B(n3652), .ZN(n3654)
         );
  NAND2_X1 U4447 ( .A1(n3655), .A2(n3654), .ZN(U3213) );
  INV_X1 U4448 ( .A(n3656), .ZN(n3658) );
  OAI21_X1 U4449 ( .B1(n3658), .B2(n3657), .A(n3535), .ZN(n3659) );
  OAI21_X1 U4450 ( .B1(n3741), .B2(n3656), .A(n3659), .ZN(n3663) );
  NOR2_X1 U4451 ( .A1(n3661), .A2(n3660), .ZN(n3662) );
  XNOR2_X1 U4452 ( .A(n3663), .B(n3662), .ZN(n3667) );
  AOI22_X1 U4453 ( .A1(n3755), .A2(n4198), .B1(n3754), .B2(n3941), .ZN(n3664)
         );
  NAND2_X1 U4454 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4009) );
  OAI211_X1 U4455 ( .C1(n3675), .C2(n3758), .A(n3664), .B(n4009), .ZN(n3665)
         );
  AOI21_X1 U4456 ( .B1(n4205), .B2(n3747), .A(n3665), .ZN(n3666) );
  OAI21_X1 U4457 ( .B1(n3667), .B2(n3762), .A(n3666), .ZN(U3216) );
  NAND2_X1 U4458 ( .A1(n2189), .A2(n3668), .ZN(n3672) );
  INV_X1 U4459 ( .A(n3724), .ZN(n3670) );
  OAI211_X1 U4460 ( .C1(n3669), .C2(n3670), .A(n3722), .B(n3672), .ZN(n3671)
         );
  OAI211_X1 U4461 ( .C1(n3673), .C2(n3672), .A(n3767), .B(n3671), .ZN(n3679)
         );
  INV_X1 U4462 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4641) );
  OAI22_X1 U4463 ( .A1(n3674), .A2(n3758), .B1(STATE_REG_SCAN_IN), .B2(n4641), 
        .ZN(n3677) );
  OAI22_X1 U4464 ( .A1(n3772), .A2(n4277), .B1(n3675), .B2(n3769), .ZN(n3676)
         );
  AOI211_X1 U4465 ( .C1(n3747), .C2(n4157), .A(n3677), .B(n3676), .ZN(n3678)
         );
  NAND2_X1 U4466 ( .A1(n3679), .A2(n3678), .ZN(U3220) );
  NOR2_X1 U4467 ( .A1(n3682), .A2(n2303), .ZN(n3683) );
  XNOR2_X1 U4468 ( .A(n3680), .B(n3683), .ZN(n3688) );
  INV_X1 U4469 ( .A(n3684), .ZN(n4086) );
  OAI22_X1 U4470 ( .A1(n3772), .A2(n4084), .B1(n4126), .B2(n3769), .ZN(n3686)
         );
  OAI22_X1 U4471 ( .A1(n4082), .A2(n3758), .B1(STATE_REG_SCAN_IN), .B2(n4644), 
        .ZN(n3685) );
  AOI211_X1 U4472 ( .C1(n4086), .C2(n3760), .A(n3686), .B(n3685), .ZN(n3687)
         );
  OAI21_X1 U4473 ( .B1(n3688), .B2(n3762), .A(n3687), .ZN(U3222) );
  OAI21_X1 U4474 ( .B1(n3689), .B2(n3765), .A(n3690), .ZN(n3691) );
  XOR2_X1 U4475 ( .A(n3692), .B(n3691), .Z(n3700) );
  AOI22_X1 U4476 ( .A1(n3755), .A2(n3693), .B1(n3744), .B2(n3774), .ZN(n3695)
         );
  INV_X1 U4477 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4643) );
  NOR2_X1 U4478 ( .A1(n4643), .A2(STATE_REG_SCAN_IN), .ZN(n4440) );
  INV_X1 U4479 ( .A(n4440), .ZN(n3694) );
  OAI211_X1 U4480 ( .C1(n3696), .C2(n3769), .A(n3695), .B(n3694), .ZN(n3697)
         );
  AOI21_X1 U4481 ( .B1(n3698), .B2(n3747), .A(n3697), .ZN(n3699) );
  OAI21_X1 U4482 ( .B1(n3700), .B2(n3762), .A(n3699), .ZN(U3223) );
  NAND2_X1 U4483 ( .A1(n3703), .A2(n3702), .ZN(n3704) );
  XNOR2_X1 U4484 ( .A(n3701), .B(n3704), .ZN(n3709) );
  AND2_X1 U4485 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3995) );
  OAI22_X1 U4486 ( .A1(n3772), .A2(n4295), .B1(n4202), .B2(n3758), .ZN(n3705)
         );
  AOI211_X1 U4487 ( .C1(n3754), .C2(n3942), .A(n3995), .B(n3705), .ZN(n3708)
         );
  NAND2_X1 U4488 ( .A1(n3747), .A2(n3706), .ZN(n3707) );
  OAI211_X1 U4489 ( .C1(n3709), .C2(n3762), .A(n3708), .B(n3707), .ZN(U3225)
         );
  NAND2_X1 U4490 ( .A1(n3711), .A2(n3710), .ZN(n3712) );
  XOR2_X1 U4491 ( .A(n3713), .B(n3712), .Z(n3720) );
  INV_X1 U4492 ( .A(n3714), .ZN(n4103) );
  OAI22_X1 U4493 ( .A1(n3772), .A2(n4262), .B1(n4097), .B2(n3769), .ZN(n3718)
         );
  OAI22_X1 U4494 ( .A1(n3716), .A2(n3758), .B1(STATE_REG_SCAN_IN), .B2(n3715), 
        .ZN(n3717) );
  AOI211_X1 U4495 ( .C1(n3747), .C2(n4103), .A(n3718), .B(n3717), .ZN(n3719)
         );
  OAI21_X1 U4496 ( .B1(n3720), .B2(n3762), .A(n3719), .ZN(U3226) );
  INV_X1 U4497 ( .A(n3721), .ZN(n3725) );
  AOI21_X1 U4498 ( .B1(n3722), .B2(n3724), .A(n3669), .ZN(n3723) );
  AOI21_X1 U4499 ( .B1(n3725), .B2(n3724), .A(n3723), .ZN(n3731) );
  INV_X1 U4500 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3726) );
  OAI22_X1 U4501 ( .A1(n3736), .A2(n3758), .B1(STATE_REG_SCAN_IN), .B2(n3726), 
        .ZN(n3729) );
  OAI22_X1 U4502 ( .A1(n3772), .A2(n3727), .B1(n4169), .B2(n3769), .ZN(n3728)
         );
  AOI211_X1 U4503 ( .C1(n3747), .C2(n4178), .A(n3729), .B(n3728), .ZN(n3730)
         );
  OAI21_X1 U4504 ( .B1(n3731), .B2(n3762), .A(n3730), .ZN(U3230) );
  AOI21_X1 U4505 ( .B1(n3734), .B2(n3733), .A(n3732), .ZN(n3740) );
  OAI22_X1 U4506 ( .A1(n4097), .A2(n3758), .B1(STATE_REG_SCAN_IN), .B2(n3735), 
        .ZN(n3738) );
  OAI22_X1 U4507 ( .A1(n3772), .A2(n4140), .B1(n3736), .B2(n3769), .ZN(n3737)
         );
  AOI211_X1 U4508 ( .C1(n3747), .C2(n4145), .A(n3738), .B(n3737), .ZN(n3739)
         );
  OAI21_X1 U4509 ( .B1(n3740), .B2(n3762), .A(n3739), .ZN(U3232) );
  XNOR2_X1 U4510 ( .A(n3742), .B(n3741), .ZN(n3743) );
  XNOR2_X1 U4511 ( .A(n3656), .B(n3743), .ZN(n3749) );
  AOI22_X1 U4512 ( .A1(n3755), .A2(n4216), .B1(n3744), .B2(n3754), .ZN(n3745)
         );
  NAND2_X1 U4513 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4445) );
  OAI211_X1 U4514 ( .C1(n4169), .C2(n3758), .A(n3745), .B(n4445), .ZN(n3746)
         );
  AOI21_X1 U4515 ( .B1(n4228), .B2(n3747), .A(n3746), .ZN(n3748) );
  OAI21_X1 U4516 ( .B1(n3749), .B2(n3762), .A(n3748), .ZN(U3235) );
  NAND2_X1 U4517 ( .A1(n2181), .A2(n3751), .ZN(n3752) );
  XNOR2_X1 U4518 ( .A(n3750), .B(n3752), .ZN(n3763) );
  INV_X1 U4519 ( .A(n3753), .ZN(n4068) );
  AOI22_X1 U4520 ( .A1(n3755), .A2(n4061), .B1(n3754), .B2(n4095), .ZN(n3757)
         );
  NAND2_X1 U4521 ( .A1(U3149), .A2(REG3_REG_26__SCAN_IN), .ZN(n3756) );
  OAI211_X1 U4522 ( .C1(n4064), .C2(n3758), .A(n3757), .B(n3756), .ZN(n3759)
         );
  AOI21_X1 U4523 ( .B1(n4068), .B2(n3760), .A(n3759), .ZN(n3761) );
  OAI21_X1 U4524 ( .B1(n3763), .B2(n3762), .A(n3761), .ZN(U3237) );
  NAND2_X1 U4525 ( .A1(n3764), .A2(n3690), .ZN(n3766) );
  XNOR2_X1 U4526 ( .A(n3766), .B(n3765), .ZN(n3768) );
  NAND2_X1 U4527 ( .A1(n3768), .A2(n3767), .ZN(n3776) );
  INV_X1 U4528 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4844) );
  NOR2_X1 U4529 ( .A1(STATE_REG_SCAN_IN), .A2(n4844), .ZN(n4431) );
  OAI22_X1 U4530 ( .A1(n3772), .A2(n3771), .B1(n3770), .B2(n3769), .ZN(n3773)
         );
  AOI211_X1 U4531 ( .C1(n3774), .C2(n3942), .A(n4431), .B(n3773), .ZN(n3775)
         );
  OAI211_X1 U4532 ( .C1(n3778), .C2(n3777), .A(n3776), .B(n3775), .ZN(U3238)
         );
  NAND2_X1 U4533 ( .A1(n2424), .A2(DATAI_31_), .ZN(n4018) );
  AND2_X1 U4534 ( .A1(n3779), .A2(DATAI_30_), .ZN(n4240) );
  INV_X1 U4535 ( .A(n4240), .ZN(n3808) );
  NAND2_X1 U4536 ( .A1(n3780), .A2(n3808), .ZN(n3883) );
  NOR2_X1 U4537 ( .A1(n3887), .A2(n2211), .ZN(n3875) );
  NAND2_X1 U4538 ( .A1(n3781), .A2(n3784), .ZN(n3856) );
  NAND2_X1 U4539 ( .A1(n3783), .A2(n3782), .ZN(n3838) );
  NAND2_X1 U4540 ( .A1(n3838), .A2(n3784), .ZN(n3855) );
  OAI21_X1 U4541 ( .B1(n3785), .B2(n3856), .A(n3855), .ZN(n3786) );
  NAND2_X1 U4542 ( .A1(n3786), .A2(n3861), .ZN(n3788) );
  NAND4_X1 U4543 ( .A1(n3788), .A2(n3863), .A3(n3787), .A4(n3862), .ZN(n3790)
         );
  INV_X1 U4544 ( .A(n3789), .ZN(n3866) );
  AOI21_X1 U4545 ( .B1(n3790), .B2(n3867), .A(n3866), .ZN(n3792) );
  OAI21_X1 U4546 ( .B1(n3792), .B2(n3869), .A(n3791), .ZN(n3793) );
  OAI221_X1 U4547 ( .B1(n2210), .B2(n3871), .C1(n2210), .C2(n3793), .A(n3880), 
        .ZN(n3796) );
  NAND2_X1 U4548 ( .A1(n4017), .A2(n4018), .ZN(n3893) );
  NAND2_X1 U4549 ( .A1(n3794), .A2(n4240), .ZN(n3894) );
  OAI211_X1 U4550 ( .C1(n3797), .C2(n3795), .A(n3893), .B(n3894), .ZN(n3804)
         );
  NOR4_X1 U4551 ( .A1(n3796), .A2(n3803), .A3(n3802), .A4(n3804), .ZN(n3810)
         );
  INV_X1 U4552 ( .A(n3797), .ZN(n4023) );
  INV_X1 U4553 ( .A(n3798), .ZN(n3799) );
  OAI21_X1 U4554 ( .B1(n4023), .B2(n3800), .A(n3799), .ZN(n3806) );
  NOR2_X1 U4555 ( .A1(n3806), .A2(n3801), .ZN(n3876) );
  NOR2_X1 U4556 ( .A1(n3803), .A2(n3802), .ZN(n3807) );
  INV_X1 U4557 ( .A(n3804), .ZN(n3805) );
  OAI21_X1 U4558 ( .B1(n3807), .B2(n3806), .A(n3805), .ZN(n3881) );
  AOI21_X1 U4559 ( .B1(n4043), .B2(n3876), .A(n3881), .ZN(n3809) );
  OAI22_X1 U4560 ( .A1(n3810), .A2(n3809), .B1(n4017), .B2(n3808), .ZN(n3813)
         );
  INV_X1 U4561 ( .A(n4017), .ZN(n3812) );
  INV_X1 U4562 ( .A(n4018), .ZN(n3811) );
  NAND2_X1 U4563 ( .A1(n3812), .A2(n3811), .ZN(n3884) );
  OAI211_X1 U4564 ( .C1(n4018), .C2(n3883), .A(n3813), .B(n3884), .ZN(n3931)
         );
  INV_X1 U4565 ( .A(n3814), .ZN(n3930) );
  INV_X1 U4566 ( .A(n3815), .ZN(n3817) );
  OAI211_X1 U4567 ( .C1(n3818), .C2(n2151), .A(n3817), .B(n3816), .ZN(n3821)
         );
  NAND3_X1 U4568 ( .A1(n3821), .A2(n3820), .A3(n3819), .ZN(n3824) );
  NAND3_X1 U4569 ( .A1(n3824), .A2(n3823), .A3(n3822), .ZN(n3827) );
  NAND3_X1 U4570 ( .A1(n3827), .A2(n3826), .A3(n3825), .ZN(n3830) );
  NAND4_X1 U4571 ( .A1(n3830), .A2(n3829), .A3(n3828), .A4(n3840), .ZN(n3832)
         );
  AND3_X1 U4572 ( .A1(n3832), .A2(n3906), .A3(n3831), .ZN(n3837) );
  NAND2_X1 U4573 ( .A1(n3834), .A2(n3833), .ZN(n3842) );
  OAI211_X1 U4574 ( .C1(n3837), .C2(n3842), .A(n3836), .B(n3835), .ZN(n3846)
         );
  INV_X1 U4575 ( .A(n3838), .ZN(n3845) );
  INV_X1 U4576 ( .A(n3839), .ZN(n3841) );
  NAND2_X1 U4577 ( .A1(n3841), .A2(n3840), .ZN(n3843) );
  OAI21_X1 U4578 ( .B1(n3843), .B2(n3842), .A(n3847), .ZN(n3844) );
  AOI22_X1 U4579 ( .A1(n3846), .A2(n3845), .B1(n3855), .B2(n3844), .ZN(n3853)
         );
  INV_X1 U4580 ( .A(n3847), .ZN(n3850) );
  OAI211_X1 U4581 ( .C1(n3850), .C2(n2177), .A(n3849), .B(n3848), .ZN(n3851)
         );
  OR3_X1 U4582 ( .A1(n3853), .A2(n3852), .A3(n3851), .ZN(n3860) );
  INV_X1 U4583 ( .A(n3854), .ZN(n3857) );
  OAI21_X1 U4584 ( .B1(n3857), .B2(n3856), .A(n3855), .ZN(n3859) );
  AOI21_X1 U4585 ( .B1(n3860), .B2(n3859), .A(n3858), .ZN(n3865) );
  INV_X1 U4586 ( .A(n3861), .ZN(n3864) );
  OAI211_X1 U4587 ( .C1(n3865), .C2(n3864), .A(n3863), .B(n3862), .ZN(n3868)
         );
  AOI211_X1 U4588 ( .C1(n3868), .C2(n3867), .A(n3866), .B(n4116), .ZN(n3870)
         );
  NOR2_X1 U4589 ( .A1(n3870), .A2(n3869), .ZN(n3873) );
  OAI21_X1 U4590 ( .B1(n3873), .B2(n3872), .A(n3871), .ZN(n3874) );
  NAND2_X1 U4591 ( .A1(n3875), .A2(n3874), .ZN(n3879) );
  INV_X1 U4592 ( .A(n3876), .ZN(n3877) );
  AOI211_X1 U4593 ( .C1(n3880), .C2(n3879), .A(n3878), .B(n3877), .ZN(n3882)
         );
  OR2_X1 U4594 ( .A1(n3882), .A2(n3881), .ZN(n3886) );
  NAND2_X1 U4595 ( .A1(n3884), .A2(n3883), .ZN(n3896) );
  NAND2_X1 U4596 ( .A1(n3896), .A2(n3893), .ZN(n3885) );
  NAND2_X1 U4597 ( .A1(n3886), .A2(n3885), .ZN(n3928) );
  INV_X1 U4598 ( .A(n4055), .ZN(n3888) );
  NOR2_X1 U4599 ( .A1(n3888), .A2(n3887), .ZN(n4073) );
  INV_X1 U4600 ( .A(n4073), .ZN(n4075) );
  NAND2_X1 U4601 ( .A1(n3890), .A2(n3889), .ZN(n4100) );
  NOR4_X1 U4602 ( .A1(n4075), .A2(n4100), .A3(n3892), .A4(n3891), .ZN(n3902)
         );
  NAND2_X1 U4603 ( .A1(n3894), .A2(n3893), .ZN(n3895) );
  NOR2_X1 U4604 ( .A1(n3896), .A2(n3895), .ZN(n3901) );
  INV_X1 U4605 ( .A(n3897), .ZN(n3900) );
  NAND2_X1 U4606 ( .A1(n3899), .A2(n3898), .ZN(n4172) );
  NAND4_X1 U4607 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n4172), .ZN(n3904)
         );
  XNOR2_X1 U4608 ( .A(n4038), .B(n4066), .ZN(n4057) );
  XNOR2_X1 U4609 ( .A(n4218), .B(n4203), .ZN(n4195) );
  NOR4_X1 U4610 ( .A1(n3904), .A2(n3903), .A3(n4057), .A4(n4195), .ZN(n3926)
         );
  INV_X1 U4611 ( .A(n3905), .ZN(n3907) );
  NOR4_X1 U4612 ( .A1(n3907), .A2(n2425), .A3(n2477), .A4(n2686), .ZN(n3920)
         );
  NOR4_X1 U4613 ( .A1(n2355), .A2(n3910), .A3(n4214), .A4(n3909), .ZN(n3919)
         );
  INV_X1 U4614 ( .A(n4116), .ZN(n3911) );
  NAND2_X1 U4615 ( .A1(n3911), .A2(n4117), .ZN(n4154) );
  NOR4_X1 U4616 ( .A1(n3914), .A2(n4154), .A3(n3913), .A4(n3912), .ZN(n3918)
         );
  NOR4_X1 U4617 ( .A1(n2629), .A2(n2576), .A3(n3916), .A4(n3915), .ZN(n3917)
         );
  NAND4_X1 U4618 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3924)
         );
  XNOR2_X1 U4619 ( .A(n4137), .B(n4123), .ZN(n4109) );
  INV_X1 U4620 ( .A(n4109), .ZN(n4121) );
  NAND4_X1 U4621 ( .A1(n4027), .A2(n3921), .A3(n4121), .A4(n4511), .ZN(n3922)
         );
  NOR3_X1 U4622 ( .A1(n3924), .A2(n3923), .A3(n3922), .ZN(n3925) );
  AOI21_X1 U4623 ( .B1(n3926), .B2(n3925), .A(n2151), .ZN(n3927) );
  MUX2_X1 U4624 ( .A(n3928), .B(n3927), .S(n4361), .Z(n3929) );
  AOI21_X1 U4625 ( .B1(n3931), .B2(n3930), .A(n3929), .ZN(n3932) );
  XNOR2_X1 U4626 ( .A(n3932), .B(n4362), .ZN(n3938) );
  NOR2_X1 U4627 ( .A1(n3934), .A2(n3933), .ZN(n3936) );
  OAI21_X1 U4628 ( .B1(n3937), .B2(n4360), .A(B_REG_SCAN_IN), .ZN(n3935) );
  OAI22_X1 U4629 ( .A1(n3938), .A2(n3937), .B1(n3936), .B2(n3935), .ZN(U3239)
         );
  MUX2_X1 U4630 ( .A(DATAO_REG_28__SCAN_IN), .B(n3939), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4631 ( .A(DATAO_REG_27__SCAN_IN), .B(n3940), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4632 ( .A(DATAO_REG_24__SCAN_IN), .B(n4079), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4633 ( .A(n4137), .B(DATAO_REG_23__SCAN_IN), .S(n3948), .Z(U3573)
         );
  MUX2_X1 U4634 ( .A(n4152), .B(DATAO_REG_22__SCAN_IN), .S(n3948), .Z(U3572)
         );
  MUX2_X1 U4635 ( .A(n4199), .B(DATAO_REG_20__SCAN_IN), .S(n3948), .Z(U3570)
         );
  MUX2_X1 U4636 ( .A(n4218), .B(DATAO_REG_19__SCAN_IN), .S(n3948), .Z(U3569)
         );
  MUX2_X1 U4637 ( .A(n3941), .B(DATAO_REG_18__SCAN_IN), .S(n3948), .Z(U3568)
         );
  MUX2_X1 U4638 ( .A(n3942), .B(DATAO_REG_16__SCAN_IN), .S(n3948), .Z(U3566)
         );
  MUX2_X1 U4639 ( .A(n3943), .B(DATAO_REG_15__SCAN_IN), .S(n3948), .Z(U3565)
         );
  MUX2_X1 U4640 ( .A(n3944), .B(DATAO_REG_12__SCAN_IN), .S(n3948), .Z(U3562)
         );
  MUX2_X1 U4641 ( .A(DATAO_REG_8__SCAN_IN), .B(n3945), .S(U4043), .Z(U3558) );
  MUX2_X1 U4642 ( .A(n3946), .B(DATAO_REG_7__SCAN_IN), .S(n3948), .Z(U3557) );
  MUX2_X1 U4643 ( .A(n3947), .B(DATAO_REG_6__SCAN_IN), .S(n3948), .Z(U3556) );
  MUX2_X1 U4644 ( .A(n2414), .B(DATAO_REG_1__SCAN_IN), .S(n3948), .Z(U3551) );
  MUX2_X1 U4645 ( .A(n3949), .B(DATAO_REG_0__SCAN_IN), .S(n3948), .Z(U3550) );
  AOI21_X1 U4646 ( .B1(n2876), .B2(n3950), .A(n3951), .ZN(n3952) );
  MUX2_X1 U4647 ( .A(n3952), .B(n3951), .S(n4652), .Z(n3954) );
  NAND2_X1 U4648 ( .A1(n3954), .A2(n3953), .ZN(n3957) );
  AOI22_X1 U4649 ( .A1(n4450), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3956) );
  NAND3_X1 U4650 ( .A1(n4452), .A2(n4652), .A3(n2876), .ZN(n3955) );
  NAND3_X1 U4651 ( .A1(n3957), .A2(n3956), .A3(n3955), .ZN(U3240) );
  NAND2_X1 U4652 ( .A1(n3958), .A2(n4370), .ZN(n3968) );
  OAI211_X1 U4653 ( .C1(n3961), .C2(n3960), .A(n4452), .B(n3959), .ZN(n3967)
         );
  OAI211_X1 U4654 ( .C1(n3964), .C2(n2783), .A(n4410), .B(n3963), .ZN(n3966)
         );
  AOI22_X1 U4655 ( .A1(n4450), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3965) );
  NAND4_X1 U4656 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(U3241)
         );
  NAND2_X1 U4657 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3986), .ZN(n3974) );
  INV_X1 U4658 ( .A(n3986), .ZN(n4500) );
  INV_X1 U4659 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4748) );
  AOI22_X1 U4660 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3986), .B1(n4500), .B2(
        n4748), .ZN(n4434) );
  INV_X1 U4661 ( .A(n3969), .ZN(n3971) );
  NAND2_X1 U4662 ( .A1(n4501), .A2(n3972), .ZN(n3973) );
  INV_X1 U4663 ( .A(n4501), .ZN(n4426) );
  NAND2_X1 U4664 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4423), .ZN(n4422) );
  NAND2_X1 U4665 ( .A1(n3973), .A2(n4422), .ZN(n4433) );
  NAND2_X1 U4666 ( .A1(n4434), .A2(n4433), .ZN(n4432) );
  NOR2_X1 U4667 ( .A1(n3987), .A2(n3975), .ZN(n3976) );
  INV_X1 U4668 ( .A(n3987), .ZN(n4499) );
  INV_X1 U4669 ( .A(n3993), .ZN(n4363) );
  NOR2_X1 U4670 ( .A1(n4363), .A2(REG1_REG_17__SCAN_IN), .ZN(n4005) );
  INV_X1 U4671 ( .A(n4005), .ZN(n3977) );
  OAI21_X1 U4672 ( .B1(n4298), .B2(n3993), .A(n3977), .ZN(n3978) );
  NOR2_X1 U4673 ( .A1(n3979), .A2(n3978), .ZN(n4004) );
  AOI21_X1 U4674 ( .B1(n3979), .B2(n3978), .A(n4004), .ZN(n3999) );
  XNOR2_X1 U4675 ( .A(n3993), .B(REG2_REG_17__SCAN_IN), .ZN(n3991) );
  NOR2_X1 U4676 ( .A1(n4426), .A2(n3983), .ZN(n3984) );
  INV_X1 U4677 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4419) );
  XOR2_X1 U4678 ( .A(n4501), .B(n3983), .Z(n4418) );
  NOR2_X1 U4679 ( .A1(n4419), .A2(n4418), .ZN(n4417) );
  NOR2_X1 U4680 ( .A1(n3984), .A2(n4417), .ZN(n4429) );
  NAND2_X1 U4681 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3986), .ZN(n3985) );
  OAI21_X1 U4682 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3986), .A(n3985), .ZN(n4428) );
  NAND2_X1 U4683 ( .A1(n3988), .A2(n4499), .ZN(n3989) );
  INV_X1 U4684 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4780) );
  NAND2_X1 U4685 ( .A1(n3989), .A2(n4437), .ZN(n3990) );
  NAND2_X1 U4686 ( .A1(n3990), .A2(n3991), .ZN(n4000) );
  AOI221_X1 U4687 ( .B1(n3991), .B2(n4000), .C1(n3990), .C2(n4000), .A(n4446), 
        .ZN(n3992) );
  INV_X1 U4688 ( .A(n3992), .ZN(n3997) );
  NOR2_X1 U4689 ( .A1(n4457), .A2(n3993), .ZN(n3994) );
  AOI211_X1 U4690 ( .C1(n4450), .C2(ADDR_REG_17__SCAN_IN), .A(n3995), .B(n3994), .ZN(n3996) );
  OAI211_X1 U4691 ( .C1(n3999), .C2(n3998), .A(n3997), .B(n3996), .ZN(U3257)
         );
  INV_X1 U4692 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4794) );
  MUX2_X1 U4693 ( .A(n4794), .B(REG2_REG_19__SCAN_IN), .S(n4010), .Z(n4002) );
  INV_X1 U4694 ( .A(n4003), .ZN(n4497) );
  INV_X1 U4695 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4782) );
  AOI22_X1 U4696 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4497), .B1(n4003), .B2(
        n4782), .ZN(n4448) );
  AOI21_X1 U4697 ( .B1(n4003), .B2(REG2_REG_18__SCAN_IN), .A(n4447), .ZN(n4001) );
  XOR2_X1 U4698 ( .A(n4002), .B(n4001), .Z(n4014) );
  INV_X1 U4699 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4700 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4003), .B1(n4497), .B2(
        n4006), .ZN(n4454) );
  INV_X1 U4701 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4751) );
  MUX2_X1 U4702 ( .A(REG1_REG_19__SCAN_IN), .B(n4751), .S(n4010), .Z(n4007) );
  NAND2_X1 U4703 ( .A1(n4450), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4008) );
  OAI211_X1 U4704 ( .C1(n4457), .C2(n4010), .A(n4009), .B(n4008), .ZN(n4011)
         );
  AOI21_X1 U4705 ( .B1(n4012), .B2(n4452), .A(n4011), .ZN(n4013) );
  OAI21_X1 U4706 ( .B1(n4014), .B2(n4446), .A(n4013), .ZN(U3259) );
  XNOR2_X1 U4707 ( .A(n4238), .B(n4018), .ZN(n4310) );
  INV_X1 U4708 ( .A(n4015), .ZN(n4016) );
  NAND2_X1 U4709 ( .A1(n4017), .A2(n4016), .ZN(n4242) );
  OAI21_X1 U4710 ( .B1(n4018), .B2(n4294), .A(n4242), .ZN(n4308) );
  NAND2_X1 U4711 ( .A1(n4232), .A2(n4308), .ZN(n4020) );
  NAND2_X1 U4712 ( .A1(n4371), .A2(REG2_REG_31__SCAN_IN), .ZN(n4019) );
  OAI211_X1 U4713 ( .C1(n4310), .C2(n4207), .A(n4020), .B(n4019), .ZN(U3260)
         );
  INV_X1 U4714 ( .A(n4027), .ZN(n4021) );
  XNOR2_X1 U4715 ( .A(n4022), .B(n4021), .ZN(n4025) );
  OAI22_X1 U4716 ( .A1(n4064), .A2(n4220), .B1(n4023), .B2(n4479), .ZN(n4024)
         );
  AOI21_X1 U4717 ( .B1(n4025), .B2(n4196), .A(n4024), .ZN(n4244) );
  NAND2_X1 U4718 ( .A1(n4246), .A2(n4156), .ZN(n4036) );
  INV_X1 U4719 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4029) );
  OAI22_X1 U4720 ( .A1(n4232), .A2(n4029), .B1(n4028), .B2(n4114), .ZN(n4032)
         );
  OAI21_X1 U4721 ( .B1(n4045), .B2(n4245), .A(n4030), .ZN(n4314) );
  NOR2_X1 U4722 ( .A1(n4314), .A2(n4207), .ZN(n4031) );
  AOI211_X1 U4723 ( .C1(n4034), .C2(n4033), .A(n4032), .B(n4031), .ZN(n4035)
         );
  OAI211_X1 U4724 ( .C1(n4244), .C2(n4371), .A(n4036), .B(n4035), .ZN(U3262)
         );
  XNOR2_X1 U4725 ( .A(n4037), .B(n4043), .ZN(n4042) );
  NAND2_X1 U4726 ( .A1(n4038), .A2(n4476), .ZN(n4039) );
  OAI21_X1 U4727 ( .B1(n4040), .B2(n4479), .A(n4039), .ZN(n4041) );
  AOI21_X1 U4728 ( .B1(n4042), .B2(n4196), .A(n4041), .ZN(n4248) );
  XNOR2_X1 U4729 ( .A(n4044), .B(n4043), .ZN(n4251) );
  NAND2_X1 U4730 ( .A1(n4251), .A2(n4156), .ZN(n4053) );
  INV_X1 U4731 ( .A(n4065), .ZN(n4047) );
  INV_X1 U4732 ( .A(n4045), .ZN(n4046) );
  INV_X1 U4733 ( .A(n4318), .ZN(n4051) );
  AOI22_X1 U4734 ( .A1(n4048), .A2(n4483), .B1(n4492), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4049) );
  OAI21_X1 U4735 ( .B1(n4159), .B2(n4249), .A(n4049), .ZN(n4050) );
  AOI21_X1 U4736 ( .B1(n4051), .B2(n4488), .A(n4050), .ZN(n4052) );
  OAI211_X1 U4737 ( .C1(n4248), .C2(n4371), .A(n4053), .B(n4052), .ZN(U3263)
         );
  XNOR2_X1 U4738 ( .A(n4054), .B(n4057), .ZN(n4255) );
  INV_X1 U4739 ( .A(n4255), .ZN(n4072) );
  NAND2_X1 U4740 ( .A1(n4056), .A2(n4055), .ZN(n4059) );
  INV_X1 U4741 ( .A(n4057), .ZN(n4058) );
  XNOR2_X1 U4742 ( .A(n4059), .B(n4058), .ZN(n4060) );
  NAND2_X1 U4743 ( .A1(n4060), .A2(n4196), .ZN(n4063) );
  AOI22_X1 U4744 ( .A1(n4095), .A2(n4476), .B1(n4061), .B2(n4475), .ZN(n4062)
         );
  OAI211_X1 U4745 ( .C1(n4064), .C2(n4479), .A(n4063), .B(n4062), .ZN(n4254)
         );
  INV_X1 U4746 ( .A(n4083), .ZN(n4067) );
  OAI21_X1 U4747 ( .B1(n4067), .B2(n4066), .A(n4065), .ZN(n4322) );
  AOI22_X1 U4748 ( .A1(n4068), .A2(n4483), .B1(n4492), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n4069) );
  OAI21_X1 U4749 ( .B1(n4322), .B2(n4207), .A(n4069), .ZN(n4070) );
  AOI21_X1 U4750 ( .B1(n4254), .B2(n4232), .A(n4070), .ZN(n4071) );
  OAI21_X1 U4751 ( .B1(n4072), .B2(n4235), .A(n4071), .ZN(U3264) );
  XNOR2_X1 U4752 ( .A(n4074), .B(n4073), .ZN(n4258) );
  INV_X1 U4753 ( .A(n4258), .ZN(n4090) );
  XNOR2_X1 U4754 ( .A(n4076), .B(n4075), .ZN(n4077) );
  NAND2_X1 U4755 ( .A1(n4077), .A2(n4196), .ZN(n4081) );
  AOI22_X1 U4756 ( .A1(n4079), .A2(n4476), .B1(n4078), .B2(n4475), .ZN(n4080)
         );
  OAI211_X1 U4757 ( .C1(n4082), .C2(n4479), .A(n4081), .B(n4080), .ZN(n4257)
         );
  INV_X1 U4758 ( .A(n4102), .ZN(n4085) );
  OAI21_X1 U4759 ( .B1(n4085), .B2(n4084), .A(n4083), .ZN(n4326) );
  AOI22_X1 U4760 ( .A1(n4492), .A2(REG2_REG_25__SCAN_IN), .B1(n4086), .B2(
        n4483), .ZN(n4087) );
  OAI21_X1 U4761 ( .B1(n4326), .B2(n4207), .A(n4087), .ZN(n4088) );
  AOI21_X1 U4762 ( .B1(n4257), .B2(n4232), .A(n4088), .ZN(n4089) );
  OAI21_X1 U4763 ( .B1(n4090), .B2(n4235), .A(n4089), .ZN(U3265) );
  NAND2_X1 U4764 ( .A1(n4092), .A2(n4091), .ZN(n4094) );
  INV_X1 U4765 ( .A(n4100), .ZN(n4093) );
  XNOR2_X1 U4766 ( .A(n4094), .B(n4093), .ZN(n4099) );
  NAND2_X1 U4767 ( .A1(n4095), .A2(n4217), .ZN(n4096) );
  OAI21_X1 U4768 ( .B1(n4097), .B2(n4220), .A(n4096), .ZN(n4098) );
  AOI21_X1 U4769 ( .B1(n4099), .B2(n4196), .A(n4098), .ZN(n4261) );
  XNOR2_X1 U4770 ( .A(n4101), .B(n4100), .ZN(n4264) );
  NAND2_X1 U4771 ( .A1(n4264), .A2(n4156), .ZN(n4108) );
  OAI21_X1 U4772 ( .B1(n4111), .B2(n4262), .A(n4102), .ZN(n4330) );
  INV_X1 U4773 ( .A(n4330), .ZN(n4106) );
  AOI22_X1 U4774 ( .A1(n4492), .A2(REG2_REG_24__SCAN_IN), .B1(n4103), .B2(
        n4483), .ZN(n4104) );
  OAI21_X1 U4775 ( .B1(n4159), .B2(n4262), .A(n4104), .ZN(n4105) );
  AOI21_X1 U4776 ( .B1(n4106), .B2(n4488), .A(n4105), .ZN(n4107) );
  OAI211_X1 U4777 ( .C1(n4492), .C2(n4261), .A(n4108), .B(n4107), .ZN(U3266)
         );
  XNOR2_X1 U4778 ( .A(n4110), .B(n4109), .ZN(n4268) );
  AOI21_X1 U4779 ( .B1(n4112), .B2(n4143), .A(n4111), .ZN(n4333) );
  INV_X1 U4780 ( .A(n4113), .ZN(n4115) );
  OAI22_X1 U4781 ( .A1(n4232), .A2(n4796), .B1(n4115), .B2(n4114), .ZN(n4130)
         );
  OR2_X1 U4782 ( .A1(n4151), .A2(n4116), .ZN(n4118) );
  NAND2_X1 U4783 ( .A1(n4118), .A2(n4117), .ZN(n4136) );
  NAND2_X1 U4784 ( .A1(n4136), .A2(n4135), .ZN(n4120) );
  NAND2_X1 U4785 ( .A1(n4120), .A2(n4119), .ZN(n4122) );
  XNOR2_X1 U4786 ( .A(n4122), .B(n4121), .ZN(n4128) );
  OR2_X1 U4787 ( .A1(n4294), .A2(n4123), .ZN(n4125) );
  NAND2_X1 U4788 ( .A1(n4152), .A2(n4476), .ZN(n4124) );
  OAI211_X1 U4789 ( .C1(n4126), .C2(n4479), .A(n4125), .B(n4124), .ZN(n4127)
         );
  AOI21_X1 U4790 ( .B1(n4128), .B2(n4196), .A(n4127), .ZN(n4267) );
  NOR2_X1 U4791 ( .A1(n4267), .A2(n4371), .ZN(n4129) );
  AOI211_X1 U4792 ( .C1(n4333), .C2(n4488), .A(n4130), .B(n4129), .ZN(n4131)
         );
  OAI21_X1 U4793 ( .B1(n4268), .B2(n4235), .A(n4131), .ZN(U3267) );
  NAND2_X1 U4794 ( .A1(n4132), .A2(n4135), .ZN(n4133) );
  NAND2_X1 U4795 ( .A1(n4134), .A2(n4133), .ZN(n4271) );
  XNOR2_X1 U4796 ( .A(n4136), .B(n4135), .ZN(n4142) );
  NAND2_X1 U4797 ( .A1(n4167), .A2(n4476), .ZN(n4139) );
  NAND2_X1 U4798 ( .A1(n4137), .A2(n4217), .ZN(n4138) );
  OAI211_X1 U4799 ( .C1(n4294), .C2(n4140), .A(n4139), .B(n4138), .ZN(n4141)
         );
  AOI21_X1 U4800 ( .B1(n4142), .B2(n4196), .A(n4141), .ZN(n4272) );
  INV_X1 U4801 ( .A(n4272), .ZN(n4149) );
  AOI21_X1 U4802 ( .B1(n4144), .B2(n2158), .A(n2256), .ZN(n4337) );
  INV_X1 U4803 ( .A(n4337), .ZN(n4147) );
  AOI22_X1 U4804 ( .A1(n4371), .A2(REG2_REG_22__SCAN_IN), .B1(n4145), .B2(
        n4483), .ZN(n4146) );
  OAI21_X1 U4805 ( .B1(n4147), .B2(n4207), .A(n4146), .ZN(n4148) );
  AOI21_X1 U4806 ( .B1(n4149), .B2(n4232), .A(n4148), .ZN(n4150) );
  OAI21_X1 U4807 ( .B1(n4271), .B2(n4235), .A(n4150), .ZN(U3268) );
  XNOR2_X1 U4808 ( .A(n4151), .B(n4154), .ZN(n4153) );
  AOI222_X1 U4809 ( .A1(n4196), .A2(n4153), .B1(n4152), .B2(n4217), .C1(n4199), 
        .C2(n4476), .ZN(n4276) );
  XNOR2_X1 U4810 ( .A(n4155), .B(n4154), .ZN(n4279) );
  NAND2_X1 U4811 ( .A1(n4279), .A2(n4156), .ZN(n4163) );
  OAI21_X1 U4812 ( .B1(n4179), .B2(n4277), .A(n2158), .ZN(n4342) );
  INV_X1 U4813 ( .A(n4342), .ZN(n4161) );
  AOI22_X1 U4814 ( .A1(n4371), .A2(REG2_REG_21__SCAN_IN), .B1(n4157), .B2(
        n4483), .ZN(n4158) );
  OAI21_X1 U4815 ( .B1(n4159), .B2(n4277), .A(n4158), .ZN(n4160) );
  AOI21_X1 U4816 ( .B1(n4161), .B2(n4488), .A(n4160), .ZN(n4162) );
  OAI211_X1 U4817 ( .C1(n4371), .C2(n4276), .A(n4163), .B(n4162), .ZN(U3269)
         );
  NAND2_X1 U4818 ( .A1(n4165), .A2(n4164), .ZN(n4166) );
  XNOR2_X1 U4819 ( .A(n4166), .B(n4172), .ZN(n4177) );
  AOI22_X1 U4820 ( .A1(n4167), .A2(n4217), .B1(n4180), .B2(n4475), .ZN(n4168)
         );
  OAI21_X1 U4821 ( .B1(n4169), .B2(n4220), .A(n4168), .ZN(n4176) );
  AND2_X1 U4822 ( .A1(n4171), .A2(n4170), .ZN(n4173) );
  XNOR2_X1 U4823 ( .A(n4173), .B(n4172), .ZN(n4286) );
  NOR2_X1 U4824 ( .A1(n4286), .A2(n4174), .ZN(n4175) );
  AOI211_X1 U4825 ( .C1(n4196), .C2(n4177), .A(n4176), .B(n4175), .ZN(n4285)
         );
  AOI22_X1 U4826 ( .A1(n4371), .A2(REG2_REG_20__SCAN_IN), .B1(n4178), .B2(
        n4483), .ZN(n4182) );
  INV_X1 U4827 ( .A(n4179), .ZN(n4283) );
  NAND2_X1 U4828 ( .A1(n2187), .A2(n4180), .ZN(n4282) );
  NAND3_X1 U4829 ( .A1(n4283), .A2(n4488), .A3(n4282), .ZN(n4181) );
  OAI211_X1 U4830 ( .C1(n4286), .C2(n4183), .A(n4182), .B(n4181), .ZN(n4184)
         );
  INV_X1 U4831 ( .A(n4184), .ZN(n4185) );
  OAI21_X1 U4832 ( .B1(n4285), .B2(n4371), .A(n4185), .ZN(U3270) );
  NAND2_X1 U4833 ( .A1(n4211), .A2(n4186), .ZN(n4187) );
  XNOR2_X1 U4834 ( .A(n4187), .B(n4195), .ZN(n4288) );
  INV_X1 U4835 ( .A(n4288), .ZN(n4210) );
  INV_X1 U4836 ( .A(n4188), .ZN(n4189) );
  NOR2_X1 U4837 ( .A1(n4190), .A2(n4189), .ZN(n4215) );
  INV_X1 U4838 ( .A(n4191), .ZN(n4192) );
  AOI21_X1 U4839 ( .B1(n4215), .B2(n4193), .A(n4192), .ZN(n4194) );
  XOR2_X1 U4840 ( .A(n4195), .B(n4194), .Z(n4197) );
  NAND2_X1 U4841 ( .A1(n4197), .A2(n4196), .ZN(n4201) );
  AOI22_X1 U4842 ( .A1(n4199), .A2(n4217), .B1(n4475), .B2(n4198), .ZN(n4200)
         );
  OAI211_X1 U4843 ( .C1(n4202), .C2(n4220), .A(n4201), .B(n4200), .ZN(n4287)
         );
  INV_X1 U4844 ( .A(n4225), .ZN(n4204) );
  OAI21_X1 U4845 ( .B1(n4204), .B2(n4203), .A(n2187), .ZN(n4347) );
  AOI22_X1 U4846 ( .A1(n4371), .A2(REG2_REG_19__SCAN_IN), .B1(n4205), .B2(
        n4483), .ZN(n4206) );
  OAI21_X1 U4847 ( .B1(n4347), .B2(n4207), .A(n4206), .ZN(n4208) );
  AOI21_X1 U4848 ( .B1(n4287), .B2(n4232), .A(n4208), .ZN(n4209) );
  OAI21_X1 U4849 ( .B1(n4210), .B2(n4235), .A(n4209), .ZN(U3271) );
  OAI21_X1 U4850 ( .B1(n4212), .B2(n4214), .A(n4211), .ZN(n4213) );
  INV_X1 U4851 ( .A(n4213), .ZN(n4292) );
  XNOR2_X1 U4852 ( .A(n4215), .B(n4214), .ZN(n4223) );
  AOI22_X1 U4853 ( .A1(n4218), .A2(n4217), .B1(n4216), .B2(n4475), .ZN(n4219)
         );
  OAI21_X1 U4854 ( .B1(n4221), .B2(n4220), .A(n4219), .ZN(n4222) );
  AOI21_X1 U4855 ( .B1(n4223), .B2(n4196), .A(n4222), .ZN(n4291) );
  INV_X1 U4856 ( .A(n4291), .ZN(n4233) );
  OAI211_X1 U4857 ( .C1(n2266), .C2(n4226), .A(n4516), .B(n4225), .ZN(n4290)
         );
  INV_X1 U4858 ( .A(n4227), .ZN(n4230) );
  AOI22_X1 U4859 ( .A1(n4492), .A2(REG2_REG_18__SCAN_IN), .B1(n4228), .B2(
        n4483), .ZN(n4229) );
  OAI21_X1 U4860 ( .B1(n4290), .B2(n4230), .A(n4229), .ZN(n4231) );
  AOI21_X1 U4861 ( .B1(n4233), .B2(n4232), .A(n4231), .ZN(n4234) );
  OAI21_X1 U4862 ( .B1(n4292), .B2(n4235), .A(n4234), .ZN(U3272) );
  NAND2_X1 U4863 ( .A1(n4308), .A2(n4559), .ZN(n4237) );
  NAND2_X1 U4864 ( .A1(n4557), .A2(REG1_REG_31__SCAN_IN), .ZN(n4236) );
  OAI211_X1 U4865 ( .C1(n4310), .C2(n4300), .A(n4237), .B(n4236), .ZN(U3549)
         );
  AOI21_X1 U4866 ( .B1(n4240), .B2(n4239), .A(n4238), .ZN(n4372) );
  INV_X1 U4867 ( .A(n4372), .ZN(n4312) );
  NAND2_X1 U4868 ( .A1(n4240), .A2(n4475), .ZN(n4241) );
  AND2_X1 U4869 ( .A1(n4242), .A2(n4241), .ZN(n4374) );
  INV_X1 U4870 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4765) );
  MUX2_X1 U4871 ( .A(n4374), .B(n4765), .S(n4557), .Z(n4243) );
  OAI21_X1 U4872 ( .B1(n4312), .B2(n4300), .A(n4243), .ZN(U3548) );
  INV_X1 U4873 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4247) );
  INV_X1 U4874 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4252) );
  OAI21_X1 U4875 ( .B1(n4249), .B2(n4294), .A(n4248), .ZN(n4250) );
  AOI21_X1 U4876 ( .B1(n4251), .B2(n4542), .A(n4250), .ZN(n4315) );
  MUX2_X1 U4877 ( .A(n4252), .B(n4315), .S(n4559), .Z(n4253) );
  OAI21_X1 U4878 ( .B1(n4300), .B2(n4318), .A(n4253), .ZN(U3545) );
  INV_X1 U4879 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4753) );
  AOI21_X1 U4880 ( .B1(n4255), .B2(n4542), .A(n4254), .ZN(n4319) );
  MUX2_X1 U4881 ( .A(n4753), .B(n4319), .S(n4559), .Z(n4256) );
  OAI21_X1 U4882 ( .B1(n4300), .B2(n4322), .A(n4256), .ZN(U3544) );
  INV_X1 U4883 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4259) );
  AOI21_X1 U4884 ( .B1(n4258), .B2(n4542), .A(n4257), .ZN(n4323) );
  MUX2_X1 U4885 ( .A(n4259), .B(n4323), .S(n4559), .Z(n4260) );
  OAI21_X1 U4886 ( .B1(n4300), .B2(n4326), .A(n4260), .ZN(U3543) );
  INV_X1 U4887 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4265) );
  OAI21_X1 U4888 ( .B1(n4262), .B2(n4294), .A(n4261), .ZN(n4263) );
  AOI21_X1 U4889 ( .B1(n4264), .B2(n4542), .A(n4263), .ZN(n4327) );
  MUX2_X1 U4890 ( .A(n4265), .B(n4327), .S(n4559), .Z(n4266) );
  OAI21_X1 U4891 ( .B1(n4300), .B2(n4330), .A(n4266), .ZN(U3542) );
  OAI21_X1 U4892 ( .B1(n4268), .B2(n4533), .A(n4267), .ZN(n4331) );
  MUX2_X1 U4893 ( .A(REG1_REG_23__SCAN_IN), .B(n4331), .S(n4559), .Z(n4269) );
  AOI21_X1 U4894 ( .B1(n4549), .B2(n4333), .A(n4269), .ZN(n4270) );
  INV_X1 U4895 ( .A(n4270), .ZN(U3541) );
  OR2_X1 U4896 ( .A1(n4271), .A2(n4533), .ZN(n4273) );
  NAND2_X1 U4897 ( .A1(n4273), .A2(n4272), .ZN(n4335) );
  MUX2_X1 U4898 ( .A(n4335), .B(REG1_REG_22__SCAN_IN), .S(n4557), .Z(n4274) );
  AOI21_X1 U4899 ( .B1(n4549), .B2(n4337), .A(n4274), .ZN(n4275) );
  INV_X1 U4900 ( .A(n4275), .ZN(U3540) );
  INV_X1 U4901 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4280) );
  OAI21_X1 U4902 ( .B1(n4277), .B2(n4294), .A(n4276), .ZN(n4278) );
  AOI21_X1 U4903 ( .B1(n4279), .B2(n4542), .A(n4278), .ZN(n4339) );
  MUX2_X1 U4904 ( .A(n4280), .B(n4339), .S(n4559), .Z(n4281) );
  OAI21_X1 U4905 ( .B1(n4300), .B2(n4342), .A(n4281), .ZN(U3539) );
  NAND3_X1 U4906 ( .A1(n4283), .A2(n4516), .A3(n4282), .ZN(n4284) );
  OAI211_X1 U4907 ( .C1(n4286), .C2(n4523), .A(n4285), .B(n4284), .ZN(n4343)
         );
  MUX2_X1 U4908 ( .A(REG1_REG_20__SCAN_IN), .B(n4343), .S(n4559), .Z(U3538) );
  AOI21_X1 U4909 ( .B1(n4288), .B2(n4542), .A(n4287), .ZN(n4344) );
  MUX2_X1 U4910 ( .A(n4751), .B(n4344), .S(n4559), .Z(n4289) );
  OAI21_X1 U4911 ( .B1(n4300), .B2(n4347), .A(n4289), .ZN(U3537) );
  OAI211_X1 U4912 ( .C1(n4292), .C2(n4533), .A(n4291), .B(n4290), .ZN(n4348)
         );
  MUX2_X1 U4913 ( .A(REG1_REG_18__SCAN_IN), .B(n4348), .S(n4559), .Z(U3536) );
  OAI21_X1 U4914 ( .B1(n4295), .B2(n4294), .A(n4293), .ZN(n4296) );
  AOI21_X1 U4915 ( .B1(n4297), .B2(n4542), .A(n4296), .ZN(n4350) );
  INV_X1 U4916 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4298) );
  MUX2_X1 U4917 ( .A(n4350), .B(n4298), .S(n4557), .Z(n4299) );
  OAI21_X1 U4918 ( .B1(n4300), .B2(n4353), .A(n4299), .ZN(U3535) );
  NAND3_X1 U4919 ( .A1(n4302), .A2(n4301), .A3(n4516), .ZN(n4303) );
  OAI211_X1 U4920 ( .C1(n4305), .C2(n4533), .A(n4304), .B(n4303), .ZN(n4354)
         );
  MUX2_X1 U4921 ( .A(REG1_REG_16__SCAN_IN), .B(n4354), .S(n4559), .Z(U3534) );
  NOR2_X1 U4922 ( .A1(n4545), .A2(n4306), .ZN(n4307) );
  AOI21_X1 U4923 ( .B1(n4545), .B2(n4308), .A(n4307), .ZN(n4309) );
  OAI21_X1 U4924 ( .B1(n4310), .B2(n4352), .A(n4309), .ZN(U3517) );
  MUX2_X1 U4925 ( .A(n4374), .B(n2724), .S(n4544), .Z(n4311) );
  OAI21_X1 U4926 ( .B1(n4312), .B2(n4352), .A(n4311), .ZN(U3516) );
  MUX2_X1 U4927 ( .A(n4316), .B(n4315), .S(n4545), .Z(n4317) );
  OAI21_X1 U4928 ( .B1(n4318), .B2(n4352), .A(n4317), .ZN(U3513) );
  INV_X1 U4929 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4320) );
  MUX2_X1 U4930 ( .A(n4320), .B(n4319), .S(n4545), .Z(n4321) );
  OAI21_X1 U4931 ( .B1(n4322), .B2(n4352), .A(n4321), .ZN(U3512) );
  INV_X1 U4932 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4324) );
  MUX2_X1 U4933 ( .A(n4324), .B(n4323), .S(n4545), .Z(n4325) );
  OAI21_X1 U4934 ( .B1(n4326), .B2(n4352), .A(n4325), .ZN(U3511) );
  INV_X1 U4935 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4328) );
  MUX2_X1 U4936 ( .A(n4328), .B(n4327), .S(n4545), .Z(n4329) );
  OAI21_X1 U4937 ( .B1(n4330), .B2(n4352), .A(n4329), .ZN(U3510) );
  MUX2_X1 U4938 ( .A(REG0_REG_23__SCAN_IN), .B(n4331), .S(n4545), .Z(n4332) );
  AOI21_X1 U4939 ( .B1(n4333), .B2(n4525), .A(n4332), .ZN(n4334) );
  INV_X1 U4940 ( .A(n4334), .ZN(U3509) );
  MUX2_X1 U4941 ( .A(n4335), .B(REG0_REG_22__SCAN_IN), .S(n4544), .Z(n4336) );
  AOI21_X1 U4942 ( .B1(n4337), .B2(n4525), .A(n4336), .ZN(n4338) );
  INV_X1 U4943 ( .A(n4338), .ZN(U3508) );
  INV_X1 U4944 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4340) );
  MUX2_X1 U4945 ( .A(n4340), .B(n4339), .S(n4545), .Z(n4341) );
  OAI21_X1 U4946 ( .B1(n4342), .B2(n4352), .A(n4341), .ZN(U3507) );
  MUX2_X1 U4947 ( .A(REG0_REG_20__SCAN_IN), .B(n4343), .S(n4545), .Z(U3506) );
  INV_X1 U4948 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4345) );
  MUX2_X1 U4949 ( .A(n4345), .B(n4344), .S(n4545), .Z(n4346) );
  OAI21_X1 U4950 ( .B1(n4347), .B2(n4352), .A(n4346), .ZN(U3505) );
  MUX2_X1 U4951 ( .A(REG0_REG_18__SCAN_IN), .B(n4348), .S(n4545), .Z(U3503) );
  INV_X1 U4952 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4349) );
  MUX2_X1 U4953 ( .A(n4350), .B(n4349), .S(n4544), .Z(n4351) );
  OAI21_X1 U4954 ( .B1(n4353), .B2(n4352), .A(n4351), .ZN(U3501) );
  MUX2_X1 U4955 ( .A(REG0_REG_16__SCAN_IN), .B(n4354), .S(n4545), .Z(U3499) );
  MUX2_X1 U4956 ( .A(DATAI_30_), .B(n4355), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4957 ( .A(n4356), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U4958 ( .A(n4357), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U4959 ( .A(DATAI_25_), .B(n4358), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4960 ( .A(n4359), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4961 ( .A(n4360), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4962 ( .A(n2151), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4963 ( .A(DATAI_20_), .B(n4361), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4964 ( .A(n4362), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4965 ( .A(DATAI_17_), .B(n4363), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U4966 ( .A(n4364), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4967 ( .A(n4365), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4968 ( .A(n4366), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4969 ( .A(DATAI_4_), .B(n4367), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4970 ( .A(n4368), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4971 ( .A(n4369), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4972 ( .A(n4370), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U4973 ( .A(DATAI_0_), .B(n4652), .S(STATE_REG_SCAN_IN), .Z(U3352) );
  AOI22_X1 U4974 ( .A1(n4372), .A2(n4488), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4371), .ZN(n4373) );
  OAI21_X1 U4975 ( .B1(n4492), .B2(n4374), .A(n4373), .ZN(U3261) );
  INV_X1 U4976 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4801) );
  OAI211_X1 U4977 ( .C1(n4376), .C2(n2164), .A(n4410), .B(n4375), .ZN(n4377)
         );
  OAI21_X1 U4978 ( .B1(n4801), .B2(n4378), .A(n4377), .ZN(n4379) );
  NOR2_X1 U4979 ( .A1(n4380), .A2(n4379), .ZN(n4385) );
  OAI211_X1 U4980 ( .C1(n4383), .C2(n4382), .A(n4452), .B(n4381), .ZN(n4384)
         );
  OAI211_X1 U4981 ( .C1(n4457), .C2(n4509), .A(n4385), .B(n4384), .ZN(U3249)
         );
  OAI211_X1 U4982 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4387), .A(n4452), .B(n4386), .ZN(n4391) );
  OAI211_X1 U4983 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4389), .A(n4410), .B(n4388), .ZN(n4390) );
  OAI211_X1 U4984 ( .C1(n4457), .C2(n4392), .A(n4391), .B(n4390), .ZN(n4393)
         );
  AOI211_X1 U4985 ( .C1(n4450), .C2(ADDR_REG_10__SCAN_IN), .A(n4394), .B(n4393), .ZN(n4395) );
  INV_X1 U4986 ( .A(n4395), .ZN(U3250) );
  OAI211_X1 U4987 ( .C1(n4398), .C2(n4397), .A(n4452), .B(n4396), .ZN(n4403)
         );
  OAI211_X1 U4988 ( .C1(n4401), .C2(n4400), .A(n4410), .B(n4399), .ZN(n4402)
         );
  OAI211_X1 U4989 ( .C1(n4457), .C2(n4505), .A(n4403), .B(n4402), .ZN(n4404)
         );
  AOI211_X1 U4990 ( .C1(n4450), .C2(ADDR_REG_11__SCAN_IN), .A(n4405), .B(n4404), .ZN(n4406) );
  INV_X1 U4991 ( .A(n4406), .ZN(U3251) );
  OAI211_X1 U4992 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4408), .A(n4452), .B(n4407), .ZN(n4413) );
  OAI211_X1 U4993 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4411), .A(n4410), .B(n4409), .ZN(n4412) );
  OAI211_X1 U4994 ( .C1(n4457), .C2(n4503), .A(n4413), .B(n4412), .ZN(n4414)
         );
  AOI211_X1 U4995 ( .C1(n4450), .C2(ADDR_REG_12__SCAN_IN), .A(n4415), .B(n4414), .ZN(n4416) );
  INV_X1 U4996 ( .A(n4416), .ZN(U3252) );
  AOI211_X1 U4997 ( .C1(n4419), .C2(n4418), .A(n4417), .B(n4446), .ZN(n4420)
         );
  AOI211_X1 U4998 ( .C1(n4450), .C2(ADDR_REG_14__SCAN_IN), .A(n4421), .B(n4420), .ZN(n4425) );
  OAI211_X1 U4999 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4423), .A(n4452), .B(n4422), .ZN(n4424) );
  OAI211_X1 U5000 ( .C1(n4457), .C2(n4426), .A(n4425), .B(n4424), .ZN(U3254)
         );
  AOI211_X1 U5001 ( .C1(n4429), .C2(n4428), .A(n4427), .B(n4446), .ZN(n4430)
         );
  AOI211_X1 U5002 ( .C1(n4450), .C2(ADDR_REG_15__SCAN_IN), .A(n4431), .B(n4430), .ZN(n4436) );
  OAI211_X1 U5003 ( .C1(n4434), .C2(n4433), .A(n4452), .B(n4432), .ZN(n4435)
         );
  OAI211_X1 U5004 ( .C1(n4457), .C2(n4500), .A(n4436), .B(n4435), .ZN(U3255)
         );
  AOI221_X1 U5005 ( .B1(n4438), .B2(n4437), .C1(n4780), .C2(n4437), .A(n4446), 
        .ZN(n4439) );
  AOI211_X1 U5006 ( .C1(n4450), .C2(ADDR_REG_16__SCAN_IN), .A(n4440), .B(n4439), .ZN(n4444) );
  OAI221_X1 U5007 ( .B1(n4442), .B2(REG1_REG_16__SCAN_IN), .C1(n4442), .C2(
        n4441), .A(n4452), .ZN(n4443) );
  OAI211_X1 U5008 ( .C1(n4457), .C2(n4499), .A(n4444), .B(n4443), .ZN(U3256)
         );
  INV_X1 U5009 ( .A(n4445), .ZN(n4449) );
  OAI211_X1 U5010 ( .C1(n4454), .C2(n4453), .A(n4452), .B(n4451), .ZN(n4455)
         );
  OAI211_X1 U5011 ( .C1(n4457), .C2(n4497), .A(n4456), .B(n4455), .ZN(U3258)
         );
  AOI22_X1 U5012 ( .A1(n4492), .A2(REG2_REG_8__SCAN_IN), .B1(n4458), .B2(n4483), .ZN(n4463) );
  INV_X1 U5013 ( .A(n4459), .ZN(n4460) );
  AOI22_X1 U5014 ( .A1(n4461), .A2(n4489), .B1(n4488), .B2(n4460), .ZN(n4462)
         );
  OAI211_X1 U5015 ( .C1(n4371), .C2(n4464), .A(n4463), .B(n4462), .ZN(U3282)
         );
  AOI22_X1 U5016 ( .A1(n4492), .A2(REG2_REG_3__SCAN_IN), .B1(n4483), .B2(n4638), .ZN(n4468) );
  AOI22_X1 U5017 ( .A1(n4466), .A2(n4489), .B1(n4488), .B2(n4465), .ZN(n4467)
         );
  OAI211_X1 U5018 ( .C1(n4492), .C2(n4469), .A(n4468), .B(n4467), .ZN(U3287)
         );
  OAI21_X1 U5019 ( .B1(n2364), .B2(n2425), .A(n4470), .ZN(n4521) );
  OAI21_X1 U5020 ( .B1(n4473), .B2(n4472), .A(n4471), .ZN(n4474) );
  NAND2_X1 U5021 ( .A1(n4474), .A2(n4196), .ZN(n4478) );
  AOI22_X1 U5022 ( .A1(n2414), .A2(n4476), .B1(n4487), .B2(n4475), .ZN(n4477)
         );
  OAI211_X1 U5023 ( .C1(n4480), .C2(n4479), .A(n4478), .B(n4477), .ZN(n4481)
         );
  AOI21_X1 U5024 ( .B1(n4482), .B2(n4521), .A(n4481), .ZN(n4522) );
  AOI22_X1 U5025 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4483), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4492), .ZN(n4491) );
  INV_X1 U5026 ( .A(n4484), .ZN(n4485) );
  AOI21_X1 U5027 ( .B1(n4487), .B2(n4486), .A(n4485), .ZN(n4548) );
  AOI22_X1 U5028 ( .A1(n4521), .A2(n4489), .B1(n4488), .B2(n4548), .ZN(n4490)
         );
  OAI211_X1 U5029 ( .C1(n4492), .C2(n4522), .A(n4491), .B(n4490), .ZN(U3288)
         );
  AND2_X1 U5030 ( .A1(D_REG_31__SCAN_IN), .A2(n4493), .ZN(U3291) );
  AND2_X1 U5031 ( .A1(D_REG_30__SCAN_IN), .A2(n4493), .ZN(U3292) );
  INV_X1 U5032 ( .A(D_REG_29__SCAN_IN), .ZN(n4711) );
  NOR2_X1 U5033 ( .A1(n4494), .A2(n4711), .ZN(U3293) );
  INV_X1 U5034 ( .A(D_REG_28__SCAN_IN), .ZN(n4704) );
  NOR2_X1 U5035 ( .A1(n4494), .A2(n4704), .ZN(U3294) );
  INV_X1 U5036 ( .A(D_REG_27__SCAN_IN), .ZN(n4705) );
  NOR2_X1 U5037 ( .A1(n4494), .A2(n4705), .ZN(U3295) );
  AND2_X1 U5038 ( .A1(D_REG_26__SCAN_IN), .A2(n4493), .ZN(U3296) );
  INV_X1 U5039 ( .A(D_REG_25__SCAN_IN), .ZN(n4702) );
  NOR2_X1 U5040 ( .A1(n4494), .A2(n4702), .ZN(U3297) );
  INV_X1 U5041 ( .A(D_REG_24__SCAN_IN), .ZN(n4701) );
  NOR2_X1 U5042 ( .A1(n4494), .A2(n4701), .ZN(U3298) );
  INV_X1 U5043 ( .A(D_REG_23__SCAN_IN), .ZN(n4698) );
  NOR2_X1 U5044 ( .A1(n4494), .A2(n4698), .ZN(U3299) );
  NOR2_X1 U5045 ( .A1(n4494), .A2(n4699), .ZN(U3300) );
  INV_X1 U5046 ( .A(D_REG_21__SCAN_IN), .ZN(n4695) );
  NOR2_X1 U5047 ( .A1(n4494), .A2(n4695), .ZN(U3301) );
  AND2_X1 U5048 ( .A1(D_REG_20__SCAN_IN), .A2(n4493), .ZN(U3302) );
  INV_X1 U5049 ( .A(D_REG_19__SCAN_IN), .ZN(n4696) );
  NOR2_X1 U5050 ( .A1(n4494), .A2(n4696), .ZN(U3303) );
  AND2_X1 U5051 ( .A1(D_REG_18__SCAN_IN), .A2(n4493), .ZN(U3304) );
  AND2_X1 U5052 ( .A1(D_REG_17__SCAN_IN), .A2(n4493), .ZN(U3305) );
  AND2_X1 U5053 ( .A1(D_REG_16__SCAN_IN), .A2(n4493), .ZN(U3306) );
  INV_X1 U5054 ( .A(D_REG_15__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5055 ( .A1(n4494), .A2(n4689), .ZN(U3307) );
  INV_X1 U5056 ( .A(D_REG_14__SCAN_IN), .ZN(n4688) );
  NOR2_X1 U5057 ( .A1(n4494), .A2(n4688), .ZN(U3308) );
  INV_X1 U5058 ( .A(D_REG_13__SCAN_IN), .ZN(n4685) );
  NOR2_X1 U5059 ( .A1(n4494), .A2(n4685), .ZN(U3309) );
  INV_X1 U5060 ( .A(D_REG_12__SCAN_IN), .ZN(n4686) );
  NOR2_X1 U5061 ( .A1(n4494), .A2(n4686), .ZN(U3310) );
  INV_X1 U5062 ( .A(D_REG_11__SCAN_IN), .ZN(n4683) );
  NOR2_X1 U5063 ( .A1(n4494), .A2(n4683), .ZN(U3311) );
  AND2_X1 U5064 ( .A1(D_REG_10__SCAN_IN), .A2(n4493), .ZN(U3312) );
  INV_X1 U5065 ( .A(D_REG_9__SCAN_IN), .ZN(n4840) );
  NOR2_X1 U5066 ( .A1(n4494), .A2(n4840), .ZN(U3313) );
  NOR2_X1 U5067 ( .A1(n4494), .A2(n4839), .ZN(U3314) );
  AND2_X1 U5068 ( .A1(D_REG_7__SCAN_IN), .A2(n4493), .ZN(U3315) );
  INV_X1 U5069 ( .A(D_REG_6__SCAN_IN), .ZN(n4682) );
  NOR2_X1 U5070 ( .A1(n4494), .A2(n4682), .ZN(U3316) );
  NOR2_X1 U5071 ( .A1(n4494), .A2(n4680), .ZN(U3317) );
  AND2_X1 U5072 ( .A1(D_REG_4__SCAN_IN), .A2(n4493), .ZN(U3318) );
  NOR2_X1 U5073 ( .A1(n4494), .A2(n4679), .ZN(U3319) );
  INV_X1 U5074 ( .A(D_REG_2__SCAN_IN), .ZN(n4667) );
  NOR2_X1 U5075 ( .A1(n4494), .A2(n4667), .ZN(U3320) );
  OAI21_X1 U5076 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4495), .ZN(
        n4496) );
  INV_X1 U5077 ( .A(n4496), .ZN(U3329) );
  INV_X1 U5078 ( .A(DATAI_18_), .ZN(n4613) );
  AOI22_X1 U5079 ( .A1(STATE_REG_SCAN_IN), .A2(n4497), .B1(n4613), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5080 ( .A(DATAI_16_), .ZN(n4498) );
  AOI22_X1 U5081 ( .A1(STATE_REG_SCAN_IN), .A2(n4499), .B1(n4498), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5082 ( .A(DATAI_15_), .ZN(n4617) );
  AOI22_X1 U5083 ( .A1(STATE_REG_SCAN_IN), .A2(n4500), .B1(n4617), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5084 ( .A1(U3149), .A2(n4501), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4502) );
  INV_X1 U5085 ( .A(n4502), .ZN(U3338) );
  INV_X1 U5086 ( .A(DATAI_12_), .ZN(n4623) );
  AOI22_X1 U5087 ( .A1(STATE_REG_SCAN_IN), .A2(n4503), .B1(n4623), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5088 ( .A(DATAI_11_), .ZN(n4504) );
  AOI22_X1 U5089 ( .A1(STATE_REG_SCAN_IN), .A2(n4505), .B1(n4504), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U5090 ( .A1(U3149), .A2(n4506), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4507) );
  INV_X1 U5091 ( .A(n4507), .ZN(U3342) );
  INV_X1 U5092 ( .A(DATAI_9_), .ZN(n4508) );
  AOI22_X1 U5093 ( .A1(STATE_REG_SCAN_IN), .A2(n4509), .B1(n4508), .B2(U3149), 
        .ZN(U3343) );
  OAI22_X1 U5094 ( .A1(n4511), .A2(n4523), .B1(n2880), .B2(n4510), .ZN(n4512)
         );
  NOR2_X1 U5095 ( .A1(n4513), .A2(n4512), .ZN(n4546) );
  INV_X1 U5096 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4514) );
  AOI22_X1 U5097 ( .A1(n4545), .A2(n4546), .B1(n4514), .B2(n4544), .ZN(U3467)
         );
  INV_X1 U5098 ( .A(n4515), .ZN(n4520) );
  OAI22_X1 U5099 ( .A1(n4518), .A2(n4523), .B1(n2871), .B2(n4517), .ZN(n4519)
         );
  NOR2_X1 U5100 ( .A1(n4520), .A2(n4519), .ZN(n4547) );
  INV_X1 U5101 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4712) );
  AOI22_X1 U5102 ( .A1(n4545), .A2(n4547), .B1(n4712), .B2(n4544), .ZN(U3469)
         );
  INV_X1 U5103 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4714) );
  INV_X1 U5104 ( .A(n4521), .ZN(n4524) );
  OAI21_X1 U5105 ( .B1(n4524), .B2(n4523), .A(n4522), .ZN(n4550) );
  AOI22_X1 U5106 ( .A1(n4550), .A2(n4545), .B1(n4525), .B2(n4548), .ZN(n4526)
         );
  OAI21_X1 U5107 ( .B1(n4545), .B2(n4714), .A(n4526), .ZN(U3471) );
  INV_X1 U5108 ( .A(n4527), .ZN(n4529) );
  AOI211_X1 U5109 ( .C1(n4531), .C2(n4530), .A(n4529), .B(n4528), .ZN(n4554)
         );
  INV_X1 U5110 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4532) );
  AOI22_X1 U5111 ( .A1(n4545), .A2(n4554), .B1(n4532), .B2(n4544), .ZN(U3475)
         );
  NOR2_X1 U5112 ( .A1(n4534), .A2(n4533), .ZN(n4538) );
  AOI211_X1 U5113 ( .C1(n4538), .C2(n4537), .A(n4536), .B(n4535), .ZN(n4556)
         );
  INV_X1 U5114 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4717) );
  AOI22_X1 U5115 ( .A1(n4545), .A2(n4556), .B1(n4717), .B2(n4544), .ZN(U3481)
         );
  OAI21_X1 U5116 ( .B1(n2871), .B2(n4540), .A(n4539), .ZN(n4541) );
  AOI21_X1 U5117 ( .B1(n4543), .B2(n4542), .A(n4541), .ZN(n4558) );
  INV_X1 U5118 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4721) );
  AOI22_X1 U5119 ( .A1(n4545), .A2(n4558), .B1(n4721), .B2(n4544), .ZN(U3485)
         );
  AOI22_X1 U5120 ( .A1(n4559), .A2(n4546), .B1(n2876), .B2(n4557), .ZN(U3518)
         );
  INV_X1 U5121 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4738) );
  AOI22_X1 U5122 ( .A1(n4559), .A2(n4547), .B1(n4738), .B2(n4557), .ZN(U3519)
         );
  AOI22_X1 U5123 ( .A1(n4550), .A2(n4559), .B1(n4549), .B2(n4548), .ZN(n4551)
         );
  OAI21_X1 U5124 ( .B1(n4559), .B2(n4552), .A(n4551), .ZN(U3520) );
  INV_X1 U5125 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4553) );
  AOI22_X1 U5126 ( .A1(n4559), .A2(n4554), .B1(n4553), .B2(n4557), .ZN(U3522)
         );
  AOI22_X1 U5127 ( .A1(n4559), .A2(n4556), .B1(n4555), .B2(n4557), .ZN(U3525)
         );
  AOI22_X1 U5128 ( .A1(n4559), .A2(n4558), .B1(n4744), .B2(n4557), .ZN(n4605)
         );
  NAND4_X1 U5129 ( .A1(REG1_REG_22__SCAN_IN), .A2(REG0_REG_20__SCAN_IN), .A3(
        REG1_REG_16__SCAN_IN), .A4(REG1_REG_30__SCAN_IN), .ZN(n4603) );
  NAND4_X1 U5130 ( .A1(REG3_REG_23__SCAN_IN), .A2(DATAI_26_), .A3(
        REG0_REG_31__SCAN_IN), .A4(ADDR_REG_18__SCAN_IN), .ZN(n4602) );
  NAND4_X1 U5131 ( .A1(DATAI_17_), .A2(DATAI_12_), .A3(DATAO_REG_2__SCAN_IN), 
        .A4(DATAO_REG_25__SCAN_IN), .ZN(n4560) );
  NOR3_X1 U5132 ( .A1(REG2_REG_27__SCAN_IN), .A2(n4844), .A3(n4560), .ZN(n4566) );
  NAND4_X1 U5133 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG2_REG_28__SCAN_IN), .A3(
        REG2_REG_13__SCAN_IN), .A4(DATAI_31_), .ZN(n4564) );
  NAND4_X1 U5134 ( .A1(REG2_REG_17__SCAN_IN), .A2(DATAO_REG_9__SCAN_IN), .A3(
        DATAO_REG_4__SCAN_IN), .A4(DATAO_REG_5__SCAN_IN), .ZN(n4563) );
  NAND4_X1 U5135 ( .A1(n4816), .A2(n4823), .A3(n4832), .A4(n4843), .ZN(n4562)
         );
  NAND4_X1 U5136 ( .A1(REG3_REG_28__SCAN_IN), .A2(DATAI_29_), .A3(
        ADDR_REG_4__SCAN_IN), .A4(ADDR_REG_9__SCAN_IN), .ZN(n4561) );
  NOR4_X1 U5137 ( .A1(n4564), .A2(n4563), .A3(n4562), .A4(n4561), .ZN(n4565)
         );
  NAND4_X1 U5138 ( .A1(REG3_REG_16__SCAN_IN), .A2(DATAO_REG_30__SCAN_IN), .A3(
        n4566), .A4(n4565), .ZN(n4601) );
  NOR4_X1 U5139 ( .A1(n4773), .A2(n4721), .A3(n4717), .A4(REG2_REG_7__SCAN_IN), 
        .ZN(n4599) );
  NOR4_X1 U5140 ( .A1(REG3_REG_6__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        DATAI_7_), .A4(DATAI_6_), .ZN(n4598) );
  NAND4_X1 U5141 ( .A1(REG2_REG_10__SCAN_IN), .A2(DATAO_REG_14__SCAN_IN), .A3(
        ADDR_REG_6__SCAN_IN), .A4(ADDR_REG_2__SCAN_IN), .ZN(n4573) );
  NAND4_X1 U5142 ( .A1(REG0_REG_10__SCAN_IN), .A2(REG3_REG_10__SCAN_IN), .A3(
        DATAI_8_), .A4(n3176), .ZN(n4572) );
  OR4_X1 U5143 ( .A1(REG0_REG_2__SCAN_IN), .A2(REG1_REG_1__SCAN_IN), .A3(
        REG2_REG_1__SCAN_IN), .A4(REG0_REG_1__SCAN_IN), .ZN(n4570) );
  INV_X1 U5144 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4718) );
  NOR4_X1 U5145 ( .A1(REG2_REG_4__SCAN_IN), .A2(REG2_REG_6__SCAN_IN), .A3(
        REG0_REG_8__SCAN_IN), .A4(n4718), .ZN(n4568) );
  INV_X1 U5146 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4745) );
  NOR4_X1 U5147 ( .A1(DATAI_1_), .A2(REG3_REG_0__SCAN_IN), .A3(DATAI_0_), .A4(
        n4745), .ZN(n4567) );
  NAND4_X1 U5148 ( .A1(REG3_REG_2__SCAN_IN), .A2(DATAI_5_), .A3(n4568), .A4(
        n4567), .ZN(n4569) );
  OR4_X1 U5149 ( .A1(n4570), .A2(REG0_REG_5__SCAN_IN), .A3(REG2_REG_5__SCAN_IN), .A4(n4569), .ZN(n4571) );
  NOR3_X1 U5150 ( .A1(n4573), .A2(n4572), .A3(n4571), .ZN(n4597) );
  NAND3_X1 U5151 ( .A1(n4574), .A2(n4794), .A3(n4782), .ZN(n4595) );
  NAND4_X1 U5152 ( .A1(IR_REG_19__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(n4650), .ZN(n4575) );
  NOR3_X1 U5153 ( .A1(D_REG_1__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(n4575), 
        .ZN(n4583) );
  NAND4_X1 U5154 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(n4668), .ZN(n4581) );
  NAND3_X1 U5155 ( .A1(n4576), .A2(IR_REG_13__SCAN_IN), .A3(n2195), .ZN(n4580)
         );
  NAND4_X1 U5156 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n4579) );
  NAND4_X1 U5157 ( .A1(n4577), .A2(IR_REG_26__SCAN_IN), .A3(
        REG1_REG_9__SCAN_IN), .A4(IR_REG_14__SCAN_IN), .ZN(n4578) );
  NOR4_X1 U5158 ( .A1(n4581), .A2(n4580), .A3(n4579), .A4(n4578), .ZN(n4582)
         );
  NAND4_X1 U5159 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .A3(n4583), 
        .A4(n4582), .ZN(n4594) );
  NOR4_X1 U5160 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG2_REG_20__SCAN_IN), .A3(
        REG2_REG_16__SCAN_IN), .A4(REG2_REG_15__SCAN_IN), .ZN(n4586) );
  NOR4_X1 U5161 ( .A1(REG1_REG_15__SCAN_IN), .A2(REG0_REG_13__SCAN_IN), .A3(
        REG1_REG_11__SCAN_IN), .A4(REG2_REG_11__SCAN_IN), .ZN(n4585) );
  NOR4_X1 U5162 ( .A1(REG3_REG_24__SCAN_IN), .A2(DATAI_25_), .A3(
        REG1_REG_19__SCAN_IN), .A4(DATAI_24_), .ZN(n4584) );
  NAND4_X1 U5163 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4593)
         );
  NOR4_X1 U5164 ( .A1(REG0_REG_28__SCAN_IN), .A2(DATAO_REG_29__SCAN_IN), .A3(
        DATAO_REG_21__SCAN_IN), .A4(DATAO_REG_17__SCAN_IN), .ZN(n4591) );
  NOR4_X1 U5165 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_12__SCAN_IN), .A3(
        DATAI_15_), .A4(DATAI_18_), .ZN(n4590) );
  NOR4_X1 U5166 ( .A1(REG1_REG_26__SCAN_IN), .A2(REG2_REG_23__SCAN_IN), .A3(
        REG0_REG_19__SCAN_IN), .A4(REG0_REG_11__SCAN_IN), .ZN(n4589) );
  NOR4_X1 U5167 ( .A1(REG1_REG_27__SCAN_IN), .A2(REG2_REG_26__SCAN_IN), .A3(
        DATAO_REG_11__SCAN_IN), .A4(DATAO_REG_3__SCAN_IN), .ZN(n4588) );
  NAND4_X1 U5168 ( .A1(n4591), .A2(n4590), .A3(n4589), .A4(n4588), .ZN(n4592)
         );
  NOR4_X1 U5169 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(n4596)
         );
  NAND4_X1 U5170 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4600)
         );
  NOR4_X1 U5171 ( .A1(n4603), .A2(n4602), .A3(n4601), .A4(n4600), .ZN(n4604)
         );
  XNOR2_X1 U5172 ( .A(n4605), .B(n4604), .ZN(n4862) );
  INV_X1 U5173 ( .A(DATAI_29_), .ZN(n4607) );
  AOI22_X1 U5174 ( .A1(n4608), .A2(keyinput71), .B1(n4607), .B2(keyinput83), 
        .ZN(n4606) );
  OAI221_X1 U5175 ( .B1(n4608), .B2(keyinput71), .C1(n4607), .C2(keyinput83), 
        .A(n4606), .ZN(n4621) );
  INV_X1 U5176 ( .A(DATAI_25_), .ZN(n4611) );
  AOI22_X1 U5177 ( .A1(n4611), .A2(keyinput69), .B1(n4610), .B2(keyinput5), 
        .ZN(n4609) );
  OAI221_X1 U5178 ( .B1(n4611), .B2(keyinput69), .C1(n4610), .C2(keyinput5), 
        .A(n4609), .ZN(n4620) );
  INV_X1 U5179 ( .A(DATAI_24_), .ZN(n4614) );
  AOI22_X1 U5180 ( .A1(n4614), .A2(keyinput48), .B1(n4613), .B2(keyinput90), 
        .ZN(n4612) );
  OAI221_X1 U5181 ( .B1(n4614), .B2(keyinput48), .C1(n4613), .C2(keyinput90), 
        .A(n4612), .ZN(n4619) );
  AOI22_X1 U5182 ( .A1(n4617), .A2(keyinput38), .B1(n4616), .B2(keyinput32), 
        .ZN(n4615) );
  OAI221_X1 U5183 ( .B1(n4617), .B2(keyinput38), .C1(n4616), .C2(keyinput32), 
        .A(n4615), .ZN(n4618) );
  NOR4_X1 U5184 ( .A1(n4621), .A2(n4620), .A3(n4619), .A4(n4618), .ZN(n4665)
         );
  AOI22_X1 U5185 ( .A1(n4623), .A2(keyinput36), .B1(keyinput21), .B2(n2487), 
        .ZN(n4622) );
  OAI221_X1 U5186 ( .B1(n4623), .B2(keyinput36), .C1(n2487), .C2(keyinput21), 
        .A(n4622), .ZN(n4633) );
  INV_X1 U5187 ( .A(DATAI_7_), .ZN(n4626) );
  INV_X1 U5188 ( .A(DATAI_6_), .ZN(n4625) );
  AOI22_X1 U5189 ( .A1(n4626), .A2(keyinput14), .B1(keyinput57), .B2(n4625), 
        .ZN(n4624) );
  OAI221_X1 U5190 ( .B1(n4626), .B2(keyinput14), .C1(n4625), .C2(keyinput57), 
        .A(n4624), .ZN(n4632) );
  XNOR2_X1 U5191 ( .A(DATAI_5_), .B(keyinput88), .ZN(n4630) );
  XNOR2_X1 U5192 ( .A(DATAI_1_), .B(keyinput39), .ZN(n4629) );
  XNOR2_X1 U5193 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput87), .ZN(n4628) );
  XNOR2_X1 U5194 ( .A(DATAI_0_), .B(keyinput117), .ZN(n4627) );
  NAND4_X1 U5195 ( .A1(n4630), .A2(n4629), .A3(n4628), .A4(n4627), .ZN(n4631)
         );
  NOR3_X1 U5196 ( .A1(n4633), .A2(n4632), .A3(n4631), .ZN(n4664) );
  AOI22_X1 U5197 ( .A1(n4636), .A2(keyinput106), .B1(keyinput43), .B2(n4635), 
        .ZN(n4634) );
  OAI221_X1 U5198 ( .B1(n4636), .B2(keyinput106), .C1(n4635), .C2(keyinput43), 
        .A(n4634), .ZN(n4648) );
  AOI22_X1 U5199 ( .A1(n2662), .A2(keyinput113), .B1(keyinput64), .B2(n4638), 
        .ZN(n4637) );
  OAI221_X1 U5200 ( .B1(n2662), .B2(keyinput113), .C1(n4638), .C2(keyinput64), 
        .A(n4637), .ZN(n4647) );
  AOI22_X1 U5201 ( .A1(n4641), .A2(keyinput75), .B1(keyinput119), .B2(n4640), 
        .ZN(n4639) );
  OAI221_X1 U5202 ( .B1(n4641), .B2(keyinput75), .C1(n4640), .C2(keyinput119), 
        .A(n4639), .ZN(n4646) );
  INV_X1 U5203 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4644) );
  AOI22_X1 U5204 ( .A1(n4644), .A2(keyinput94), .B1(keyinput29), .B2(n4643), 
        .ZN(n4642) );
  OAI221_X1 U5205 ( .B1(n4644), .B2(keyinput94), .C1(n4643), .C2(keyinput29), 
        .A(n4642), .ZN(n4645) );
  NOR4_X1 U5206 ( .A1(n4648), .A2(n4647), .A3(n4646), .A4(n4645), .ZN(n4663)
         );
  AOI22_X1 U5207 ( .A1(n4651), .A2(keyinput41), .B1(keyinput46), .B2(n4650), 
        .ZN(n4649) );
  OAI221_X1 U5208 ( .B1(n4651), .B2(keyinput41), .C1(n4650), .C2(keyinput46), 
        .A(n4649), .ZN(n4661) );
  XNOR2_X1 U5209 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput120), .ZN(n4656) );
  XNOR2_X1 U5210 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput111), .ZN(n4655) );
  XNOR2_X1 U5211 ( .A(IR_REG_7__SCAN_IN), .B(keyinput7), .ZN(n4654) );
  XNOR2_X1 U5212 ( .A(n4652), .B(keyinput61), .ZN(n4653) );
  NAND4_X1 U5213 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4660)
         );
  XNOR2_X1 U5214 ( .A(n2518), .B(keyinput2), .ZN(n4659) );
  XNOR2_X1 U5215 ( .A(n4657), .B(keyinput100), .ZN(n4658) );
  NOR4_X1 U5216 ( .A1(n4661), .A2(n4660), .A3(n4659), .A4(n4658), .ZN(n4662)
         );
  NAND4_X1 U5217 ( .A1(n4665), .A2(n4664), .A3(n4663), .A4(n4662), .ZN(n4860)
         );
  AOI22_X1 U5218 ( .A1(n4667), .A2(keyinput95), .B1(n2740), .B2(keyinput101), 
        .ZN(n4666) );
  OAI221_X1 U5219 ( .B1(n4667), .B2(keyinput95), .C1(n2740), .C2(keyinput101), 
        .A(n4666), .ZN(n4677) );
  XNOR2_X1 U5220 ( .A(n4668), .B(keyinput96), .ZN(n4676) );
  XNOR2_X1 U5221 ( .A(n4669), .B(keyinput3), .ZN(n4675) );
  XNOR2_X1 U5222 ( .A(IR_REG_18__SCAN_IN), .B(keyinput33), .ZN(n4673) );
  XNOR2_X1 U5223 ( .A(IR_REG_17__SCAN_IN), .B(keyinput126), .ZN(n4672) );
  XNOR2_X1 U5224 ( .A(IR_REG_21__SCAN_IN), .B(keyinput81), .ZN(n4671) );
  XNOR2_X1 U5225 ( .A(IR_REG_19__SCAN_IN), .B(keyinput63), .ZN(n4670) );
  NAND4_X1 U5226 ( .A1(n4673), .A2(n4672), .A3(n4671), .A4(n4670), .ZN(n4674)
         );
  NOR4_X1 U5227 ( .A1(n4677), .A2(n4676), .A3(n4675), .A4(n4674), .ZN(n4729)
         );
  AOI22_X1 U5228 ( .A1(n4680), .A2(keyinput47), .B1(n4679), .B2(keyinput93), 
        .ZN(n4678) );
  OAI221_X1 U5229 ( .B1(n4680), .B2(keyinput47), .C1(n4679), .C2(keyinput93), 
        .A(n4678), .ZN(n4693) );
  AOI22_X1 U5230 ( .A1(n4683), .A2(keyinput92), .B1(n4682), .B2(keyinput116), 
        .ZN(n4681) );
  OAI221_X1 U5231 ( .B1(n4683), .B2(keyinput92), .C1(n4682), .C2(keyinput116), 
        .A(n4681), .ZN(n4692) );
  AOI22_X1 U5232 ( .A1(n4686), .A2(keyinput8), .B1(keyinput67), .B2(n4685), 
        .ZN(n4684) );
  OAI221_X1 U5233 ( .B1(n4686), .B2(keyinput8), .C1(n4685), .C2(keyinput67), 
        .A(n4684), .ZN(n4691) );
  AOI22_X1 U5234 ( .A1(n4689), .A2(keyinput20), .B1(n4688), .B2(keyinput34), 
        .ZN(n4687) );
  OAI221_X1 U5235 ( .B1(n4689), .B2(keyinput20), .C1(n4688), .C2(keyinput34), 
        .A(n4687), .ZN(n4690) );
  NOR4_X1 U5236 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4728)
         );
  AOI22_X1 U5237 ( .A1(n4696), .A2(keyinput62), .B1(keyinput28), .B2(n4695), 
        .ZN(n4694) );
  OAI221_X1 U5238 ( .B1(n4696), .B2(keyinput62), .C1(n4695), .C2(keyinput28), 
        .A(n4694), .ZN(n4709) );
  AOI22_X1 U5239 ( .A1(n4699), .A2(keyinput15), .B1(keyinput104), .B2(n4698), 
        .ZN(n4697) );
  OAI221_X1 U5240 ( .B1(n4699), .B2(keyinput15), .C1(n4698), .C2(keyinput104), 
        .A(n4697), .ZN(n4708) );
  AOI22_X1 U5241 ( .A1(n4702), .A2(keyinput72), .B1(keyinput23), .B2(n4701), 
        .ZN(n4700) );
  OAI221_X1 U5242 ( .B1(n4702), .B2(keyinput72), .C1(n4701), .C2(keyinput23), 
        .A(n4700), .ZN(n4707) );
  AOI22_X1 U5243 ( .A1(n4705), .A2(keyinput115), .B1(n4704), .B2(keyinput122), 
        .ZN(n4703) );
  OAI221_X1 U5244 ( .B1(n4705), .B2(keyinput115), .C1(n4704), .C2(keyinput122), 
        .A(n4703), .ZN(n4706) );
  NOR4_X1 U5245 ( .A1(n4709), .A2(n4708), .A3(n4707), .A4(n4706), .ZN(n4727)
         );
  AOI22_X1 U5246 ( .A1(n4712), .A2(keyinput123), .B1(n4711), .B2(keyinput0), 
        .ZN(n4710) );
  OAI221_X1 U5247 ( .B1(n4712), .B2(keyinput123), .C1(n4711), .C2(keyinput0), 
        .A(n4710), .ZN(n4725) );
  INV_X1 U5248 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4715) );
  AOI22_X1 U5249 ( .A1(n4715), .A2(keyinput108), .B1(keyinput109), .B2(n4714), 
        .ZN(n4713) );
  OAI221_X1 U5250 ( .B1(n4715), .B2(keyinput108), .C1(n4714), .C2(keyinput109), 
        .A(n4713), .ZN(n4724) );
  AOI22_X1 U5251 ( .A1(n4718), .A2(keyinput30), .B1(n4717), .B2(keyinput53), 
        .ZN(n4716) );
  OAI221_X1 U5252 ( .B1(n4718), .B2(keyinput30), .C1(n4717), .C2(keyinput53), 
        .A(n4716), .ZN(n4723) );
  AOI22_X1 U5253 ( .A1(n4721), .A2(keyinput1), .B1(keyinput89), .B2(n4720), 
        .ZN(n4719) );
  OAI221_X1 U5254 ( .B1(n4721), .B2(keyinput1), .C1(n4720), .C2(keyinput89), 
        .A(n4719), .ZN(n4722) );
  NOR4_X1 U5255 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .ZN(n4726)
         );
  NAND4_X1 U5256 ( .A1(n4729), .A2(n4728), .A3(n4727), .A4(n4726), .ZN(n4859)
         );
  INV_X1 U5257 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5258 ( .A1(n4732), .A2(keyinput73), .B1(keyinput10), .B2(n4731), 
        .ZN(n4730) );
  OAI221_X1 U5259 ( .B1(n4732), .B2(keyinput73), .C1(n4731), .C2(keyinput10), 
        .A(n4730), .ZN(n4742) );
  AOI22_X1 U5260 ( .A1(n3396), .A2(keyinput77), .B1(n4345), .B2(keyinput51), 
        .ZN(n4733) );
  OAI221_X1 U5261 ( .B1(n3396), .B2(keyinput77), .C1(n4345), .C2(keyinput51), 
        .A(n4733), .ZN(n4741) );
  INV_X1 U5262 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5263 ( .A1(n4736), .A2(keyinput42), .B1(n4735), .B2(keyinput97), 
        .ZN(n4734) );
  OAI221_X1 U5264 ( .B1(n4736), .B2(keyinput42), .C1(n4735), .C2(keyinput97), 
        .A(n4734), .ZN(n4740) );
  AOI22_X1 U5265 ( .A1(n4738), .A2(keyinput24), .B1(keyinput84), .B2(n4306), 
        .ZN(n4737) );
  OAI221_X1 U5266 ( .B1(n4738), .B2(keyinput24), .C1(n4306), .C2(keyinput84), 
        .A(n4737), .ZN(n4739) );
  NOR4_X1 U5267 ( .A1(n4742), .A2(n4741), .A3(n4740), .A4(n4739), .ZN(n4791)
         );
  AOI22_X1 U5268 ( .A1(n4745), .A2(keyinput13), .B1(n4744), .B2(keyinput102), 
        .ZN(n4743) );
  OAI221_X1 U5269 ( .B1(n4745), .B2(keyinput13), .C1(n4744), .C2(keyinput102), 
        .A(n4743), .ZN(n4758) );
  AOI22_X1 U5270 ( .A1(n4748), .A2(keyinput76), .B1(keyinput107), .B2(n4747), 
        .ZN(n4746) );
  OAI221_X1 U5271 ( .B1(n4748), .B2(keyinput76), .C1(n4747), .C2(keyinput107), 
        .A(n4746), .ZN(n4757) );
  INV_X1 U5272 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4750) );
  AOI22_X1 U5273 ( .A1(n4751), .A2(keyinput118), .B1(keyinput11), .B2(n4750), 
        .ZN(n4749) );
  OAI221_X1 U5274 ( .B1(n4751), .B2(keyinput118), .C1(n4750), .C2(keyinput11), 
        .A(n4749), .ZN(n4756) );
  INV_X1 U5275 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4754) );
  AOI22_X1 U5276 ( .A1(n4754), .A2(keyinput40), .B1(n4753), .B2(keyinput56), 
        .ZN(n4752) );
  OAI221_X1 U5277 ( .B1(n4754), .B2(keyinput40), .C1(n4753), .C2(keyinput56), 
        .A(n4752), .ZN(n4755) );
  NOR4_X1 U5278 ( .A1(n4758), .A2(n4757), .A3(n4756), .A4(n4755), .ZN(n4790)
         );
  AOI22_X1 U5279 ( .A1(n3176), .A2(keyinput85), .B1(n4760), .B2(keyinput6), 
        .ZN(n4759) );
  OAI221_X1 U5280 ( .B1(n3176), .B2(keyinput85), .C1(n4760), .C2(keyinput6), 
        .A(n4759), .ZN(n4771) );
  INV_X1 U5281 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4763) );
  AOI22_X1 U5282 ( .A1(n4763), .A2(keyinput112), .B1(n4762), .B2(keyinput103), 
        .ZN(n4761) );
  OAI221_X1 U5283 ( .B1(n4763), .B2(keyinput112), .C1(n4762), .C2(keyinput103), 
        .A(n4761), .ZN(n4770) );
  AOI22_X1 U5284 ( .A1(n4252), .A2(keyinput35), .B1(keyinput74), .B2(n4765), 
        .ZN(n4764) );
  OAI221_X1 U5285 ( .B1(n4252), .B2(keyinput35), .C1(n4765), .C2(keyinput74), 
        .A(n4764), .ZN(n4769) );
  XOR2_X1 U5286 ( .A(n2229), .B(keyinput65), .Z(n4767) );
  XNOR2_X1 U5287 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput121), .ZN(n4766) );
  NAND2_X1 U5288 ( .A1(n4767), .A2(n4766), .ZN(n4768) );
  NOR4_X1 U5289 ( .A1(n4771), .A2(n4770), .A3(n4769), .A4(n4768), .ZN(n4789)
         );
  INV_X1 U5290 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4774) );
  AOI22_X1 U5291 ( .A1(n4774), .A2(keyinput66), .B1(keyinput70), .B2(n4773), 
        .ZN(n4772) );
  OAI221_X1 U5292 ( .B1(n4774), .B2(keyinput66), .C1(n4773), .C2(keyinput70), 
        .A(n4772), .ZN(n4787) );
  AOI22_X1 U5293 ( .A1(n4777), .A2(keyinput80), .B1(keyinput55), .B2(n4776), 
        .ZN(n4775) );
  OAI221_X1 U5294 ( .B1(n4777), .B2(keyinput80), .C1(n4776), .C2(keyinput55), 
        .A(n4775), .ZN(n4786) );
  INV_X1 U5295 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4779) );
  AOI22_X1 U5296 ( .A1(n4780), .A2(keyinput19), .B1(keyinput60), .B2(n4779), 
        .ZN(n4778) );
  OAI221_X1 U5297 ( .B1(n4780), .B2(keyinput19), .C1(n4779), .C2(keyinput60), 
        .A(n4778), .ZN(n4785) );
  INV_X1 U5298 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4783) );
  AOI22_X1 U5299 ( .A1(n4783), .A2(keyinput52), .B1(keyinput125), .B2(n4782), 
        .ZN(n4781) );
  OAI221_X1 U5300 ( .B1(n4783), .B2(keyinput52), .C1(n4782), .C2(keyinput125), 
        .A(n4781), .ZN(n4784) );
  NOR4_X1 U5301 ( .A1(n4787), .A2(n4786), .A3(n4785), .A4(n4784), .ZN(n4788)
         );
  NAND4_X1 U5302 ( .A1(n4791), .A2(n4790), .A3(n4789), .A4(n4788), .ZN(n4858)
         );
  INV_X1 U5303 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4793) );
  AOI22_X1 U5304 ( .A1(n4794), .A2(keyinput127), .B1(n4793), .B2(keyinput78), 
        .ZN(n4792) );
  OAI221_X1 U5305 ( .B1(n4794), .B2(keyinput127), .C1(n4793), .C2(keyinput78), 
        .A(n4792), .ZN(n4805) );
  INV_X1 U5306 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4797) );
  INV_X1 U5307 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4796) );
  AOI22_X1 U5308 ( .A1(n4797), .A2(keyinput59), .B1(keyinput114), .B2(n4796), 
        .ZN(n4795) );
  OAI221_X1 U5309 ( .B1(n4797), .B2(keyinput59), .C1(n4796), .C2(keyinput114), 
        .A(n4795), .ZN(n4804) );
  INV_X1 U5310 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4799) );
  AOI22_X1 U5311 ( .A1(n4029), .A2(keyinput4), .B1(keyinput58), .B2(n4799), 
        .ZN(n4798) );
  OAI221_X1 U5312 ( .B1(n4029), .B2(keyinput4), .C1(n4799), .C2(keyinput58), 
        .A(n4798), .ZN(n4803) );
  AOI22_X1 U5313 ( .A1(n4801), .A2(keyinput18), .B1(n2804), .B2(keyinput37), 
        .ZN(n4800) );
  OAI221_X1 U5314 ( .B1(n4801), .B2(keyinput18), .C1(n2804), .C2(keyinput37), 
        .A(n4800), .ZN(n4802) );
  NOR4_X1 U5315 ( .A1(n4805), .A2(n4804), .A3(n4803), .A4(n4802), .ZN(n4856)
         );
  INV_X1 U5316 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4808) );
  INV_X1 U5317 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4807) );
  AOI22_X1 U5318 ( .A1(n4808), .A2(keyinput45), .B1(n4807), .B2(keyinput99), 
        .ZN(n4806) );
  OAI221_X1 U5319 ( .B1(n4808), .B2(keyinput45), .C1(n4807), .C2(keyinput99), 
        .A(n4806), .ZN(n4821) );
  AOI22_X1 U5320 ( .A1(n4811), .A2(keyinput22), .B1(n4810), .B2(keyinput44), 
        .ZN(n4809) );
  OAI221_X1 U5321 ( .B1(n4811), .B2(keyinput22), .C1(n4810), .C2(keyinput44), 
        .A(n4809), .ZN(n4820) );
  AOI22_X1 U5322 ( .A1(n4814), .A2(keyinput105), .B1(keyinput86), .B2(n4813), 
        .ZN(n4812) );
  OAI221_X1 U5323 ( .B1(n4814), .B2(keyinput105), .C1(n4813), .C2(keyinput86), 
        .A(n4812), .ZN(n4819) );
  AOI22_X1 U5324 ( .A1(n4817), .A2(keyinput31), .B1(keyinput82), .B2(n4816), 
        .ZN(n4815) );
  OAI221_X1 U5325 ( .B1(n4817), .B2(keyinput31), .C1(n4816), .C2(keyinput82), 
        .A(n4815), .ZN(n4818) );
  NOR4_X1 U5326 ( .A1(n4821), .A2(n4820), .A3(n4819), .A4(n4818), .ZN(n4855)
         );
  AOI22_X1 U5327 ( .A1(n4824), .A2(keyinput26), .B1(n4823), .B2(keyinput54), 
        .ZN(n4822) );
  OAI221_X1 U5328 ( .B1(n4824), .B2(keyinput26), .C1(n4823), .C2(keyinput54), 
        .A(n4822), .ZN(n4837) );
  AOI22_X1 U5329 ( .A1(n4827), .A2(keyinput98), .B1(keyinput16), .B2(n4826), 
        .ZN(n4825) );
  OAI221_X1 U5330 ( .B1(n4827), .B2(keyinput98), .C1(n4826), .C2(keyinput16), 
        .A(n4825), .ZN(n4836) );
  AOI22_X1 U5331 ( .A1(n4830), .A2(keyinput12), .B1(keyinput49), .B2(n4829), 
        .ZN(n4828) );
  OAI221_X1 U5332 ( .B1(n4830), .B2(keyinput12), .C1(n4829), .C2(keyinput49), 
        .A(n4828), .ZN(n4835) );
  AOI22_X1 U5333 ( .A1(n4833), .A2(keyinput17), .B1(n4832), .B2(keyinput91), 
        .ZN(n4831) );
  OAI221_X1 U5334 ( .B1(n4833), .B2(keyinput17), .C1(n4832), .C2(keyinput91), 
        .A(n4831), .ZN(n4834) );
  NOR4_X1 U5335 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4854)
         );
  AOI22_X1 U5336 ( .A1(n4840), .A2(keyinput110), .B1(keyinput79), .B2(n4839), 
        .ZN(n4838) );
  OAI221_X1 U5337 ( .B1(n4840), .B2(keyinput110), .C1(n4839), .C2(keyinput79), 
        .A(n4838), .ZN(n4852) );
  AOI22_X1 U5338 ( .A1(n4843), .A2(keyinput50), .B1(n4842), .B2(keyinput9), 
        .ZN(n4841) );
  OAI221_X1 U5339 ( .B1(n4843), .B2(keyinput50), .C1(n4842), .C2(keyinput9), 
        .A(n4841), .ZN(n4851) );
  XOR2_X1 U5340 ( .A(n4844), .B(keyinput124), .Z(n4849) );
  INV_X1 U5341 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4845) );
  XOR2_X1 U5342 ( .A(n4845), .B(keyinput68), .Z(n4848) );
  XNOR2_X1 U5343 ( .A(REG3_REG_6__SCAN_IN), .B(keyinput27), .ZN(n4847) );
  XNOR2_X1 U5344 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput25), .ZN(n4846) );
  NAND4_X1 U5345 ( .A1(n4849), .A2(n4848), .A3(n4847), .A4(n4846), .ZN(n4850)
         );
  NOR3_X1 U5346 ( .A1(n4852), .A2(n4851), .A3(n4850), .ZN(n4853) );
  NAND4_X1 U5347 ( .A1(n4856), .A2(n4855), .A3(n4854), .A4(n4853), .ZN(n4857)
         );
  NOR4_X1 U5348 ( .A1(n4860), .A2(n4859), .A3(n4858), .A4(n4857), .ZN(n4861)
         );
  XNOR2_X1 U5349 ( .A(n4862), .B(n4861), .ZN(U3527) );
  CLKBUF_X2 U2469 ( .A(n3597), .Z(n2153) );
  CLKBUF_X1 U2397 ( .A(n2416), .Z(n2148) );
  CLKBUF_X1 U2398 ( .A(n2416), .Z(n2147) );
endmodule

