

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540;

  CLKBUF_X1 U2248 ( .A(n4242), .Z(n2006) );
  NAND2_X1 U2249 ( .A1(n3972), .A2(n2470), .ZN(n2472) );
  AND2_X1 U2250 ( .A1(n2279), .A2(n2280), .ZN(n3393) );
  CLKBUF_X2 U2251 ( .A(n2293), .Z(n2010) );
  INV_X1 U2252 ( .A(n3210), .ZN(n3152) );
  INV_X1 U2253 ( .A(n2758), .ZN(n3164) );
  AOI21_X1 U2254 ( .B1(n3673), .B2(n3650), .A(n3667), .ZN(n2535) );
  NAND2_X1 U2255 ( .A1(n3430), .A2(n3432), .ZN(n2569) );
  NAND2_X2 U2256 ( .A1(n2255), .A2(n2090), .ZN(n3397) );
  AOI21_X1 U2257 ( .B1(n3351), .B2(n3348), .A(n3347), .ZN(n3200) );
  OR2_X1 U2258 ( .A1(n3041), .A2(n3831), .ZN(n2268) );
  XNOR2_X1 U2259 ( .A(n2268), .B(IR_REG_30__SCAN_IN), .ZN(n4240) );
  NOR2_X1 U2260 ( .A1(n2564), .A2(n2614), .ZN(n4242) );
  OAI22_X2 U2261 ( .A1(n2472), .A2(n2155), .B1(n2157), .B2(n2154), .ZN(n3913)
         );
  OAI22_X2 U2262 ( .A1(n3686), .A2(n2533), .B1(n3847), .B2(n3255), .ZN(n3667)
         );
  AOI21_X1 U2263 ( .B1(n2053), .B2(n2052), .A(n2051), .ZN(n3208) );
  OAI22_X1 U2264 ( .A1(n3200), .A2(n3201), .B1(n3108), .B2(n3107), .ZN(n3291)
         );
  AND2_X1 U2265 ( .A1(n2058), .A2(n2057), .ZN(n3307) );
  NAND2_X1 U2266 ( .A1(n2873), .A2(n2872), .ZN(n2916) );
  NAND2_X1 U2267 ( .A1(n3434), .A2(n3433), .ZN(n3520) );
  CLKBUF_X1 U2268 ( .A(n2726), .Z(n4440) );
  NAND4_X1 U2269 ( .A1(n2307), .A2(n2306), .A3(n2305), .A4(n2304), .ZN(n3557)
         );
  INV_X4 U2270 ( .A(n3209), .ZN(n2110) );
  AND4_X1 U2271 ( .A1(n2276), .A2(n2275), .A3(n2274), .A4(n2273), .ZN(n2726)
         );
  INV_X4 U2272 ( .A(n2729), .ZN(n3154) );
  BUF_X1 U2273 ( .A(n2302), .Z(n2008) );
  BUF_X2 U2274 ( .A(n2293), .Z(n2009) );
  BUF_X1 U2275 ( .A(n2302), .Z(n2007) );
  NAND2_X1 U2276 ( .A1(n4240), .A2(n2020), .ZN(n2302) );
  NAND2_X1 U2277 ( .A1(n4240), .A2(n2280), .ZN(n2293) );
  MUX2_X1 U2278 ( .A(REG1_REG_28__SCAN_IN), .B(n2647), .S(n4540), .Z(n2640) );
  MUX2_X1 U2279 ( .A(REG0_REG_28__SCAN_IN), .B(n2647), .S(n4525), .Z(n2648) );
  AND2_X1 U2280 ( .A1(n2053), .A2(n2033), .ZN(n3359) );
  OR2_X1 U2281 ( .A1(n3648), .A2(n3647), .ZN(n3654) );
  NAND2_X1 U2282 ( .A1(n3143), .A2(n3279), .ZN(n3253) );
  AND2_X1 U2283 ( .A1(n2136), .A2(n2013), .ZN(n3648) );
  AND2_X1 U2284 ( .A1(n2136), .A2(n2034), .ZN(n3646) );
  AND2_X1 U2285 ( .A1(n3841), .A2(n3483), .ZN(n3690) );
  NAND2_X1 U2286 ( .A1(n2591), .A2(n3479), .ZN(n3900) );
  NAND2_X1 U2287 ( .A1(n3291), .A2(n3292), .ZN(n3290) );
  NAND2_X1 U2288 ( .A1(n3089), .A2(n3088), .ZN(n3369) );
  AOI21_X2 U2289 ( .B1(n3307), .B2(n3078), .A(n2021), .ZN(n3172) );
  OAI21_X1 U2290 ( .B1(n2976), .B2(n3460), .A(n3452), .ZN(n3003) );
  NAND2_X1 U2291 ( .A1(n2579), .A2(n3448), .ZN(n2976) );
  AND2_X1 U2292 ( .A1(n2992), .A2(n2066), .ZN(n2993) );
  NAND2_X1 U2293 ( .A1(n2064), .A2(n2108), .ZN(n2991) );
  NOR2_X1 U2294 ( .A1(n2334), .A2(n2172), .ZN(n2171) );
  OR2_X1 U2295 ( .A1(n2772), .A2(n2771), .ZN(n2774) );
  AND4_X1 U2296 ( .A1(n2319), .A2(n2318), .A3(n2317), .A4(n2316), .ZN(n2824)
         );
  NAND2_X2 U2297 ( .A1(n4519), .A2(n2110), .ZN(n2758) );
  NAND4_X1 U2298 ( .A1(n2287), .A2(n2286), .A3(n2285), .A4(n2284), .ZN(n2570)
         );
  AND4_X1 U2299 ( .A1(n2298), .A2(n2297), .A3(n2296), .A4(n2295), .ZN(n2821)
         );
  AND4_X1 U2300 ( .A1(n2347), .A2(n2346), .A3(n2345), .A4(n2344), .ZN(n2970)
         );
  NAND2_X2 U2301 ( .A1(n2781), .A2(n2834), .ZN(n3209) );
  OR2_X1 U2302 ( .A1(n2293), .A2(n2668), .ZN(n2274) );
  INV_X1 U2303 ( .A(n2302), .ZN(n2272) );
  NAND2_X1 U2304 ( .A1(n2267), .A2(n2280), .ZN(n2547) );
  XNOR2_X1 U2305 ( .A(n3573), .B(n2145), .ZN(n4271) );
  NAND2_X2 U2306 ( .A1(n2727), .A2(n2834), .ZN(n3210) );
  NAND2_X1 U2307 ( .A1(n2618), .A2(IR_REG_31__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U2308 ( .A1(n2644), .A2(n4245), .ZN(n2834) );
  AND2_X1 U2309 ( .A1(n2555), .A2(n2561), .ZN(n4245) );
  AND2_X1 U2310 ( .A1(n2236), .A2(n2250), .ZN(n2141) );
  AND2_X1 U2311 ( .A1(n2197), .A2(n2249), .ZN(n2196) );
  NAND4_X1 U2312 ( .A1(n2299), .A2(n2070), .A3(n3776), .A4(n2244), .ZN(n2331)
         );
  NOR2_X1 U2313 ( .A1(IR_REG_22__SCAN_IN), .A2(n2200), .ZN(n2199) );
  AND2_X1 U2314 ( .A1(n2308), .A2(n2067), .ZN(n2070) );
  AND2_X1 U2315 ( .A1(n2069), .A2(n2068), .ZN(n2299) );
  NOR3_X1 U2316 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .A3(
        IR_REG_15__SCAN_IN), .ZN(n2249) );
  INV_X1 U2317 ( .A(IR_REG_3__SCAN_IN), .ZN(n3776) );
  NOR2_X1 U2318 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2375)
         );
  NOR2_X1 U2319 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2100)
         );
  NOR2_X1 U2320 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2245)
         );
  NOR2_X1 U2321 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2246)
         );
  NOR2_X1 U2322 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2247)
         );
  INV_X1 U2323 ( .A(IR_REG_5__SCAN_IN), .ZN(n2244) );
  OR2_X1 U2324 ( .A1(n2009), .A2(n2283), .ZN(n2284) );
  INV_X1 U2325 ( .A(n2020), .ZN(n2280) );
  NOR2_X1 U2326 ( .A1(n2655), .A2(n2633), .ZN(n2708) );
  AND2_X1 U2327 ( .A1(n2252), .A2(n2240), .ZN(n2239) );
  NAND2_X1 U2328 ( .A1(n2103), .A2(n2102), .ZN(n2238) );
  INV_X1 U2329 ( .A(IR_REG_17__SCAN_IN), .ZN(n2103) );
  INV_X1 U2330 ( .A(IR_REG_18__SCAN_IN), .ZN(n2102) );
  XNOR2_X1 U2331 ( .A(n2728), .B(n3210), .ZN(n2763) );
  OAI22_X1 U2332 ( .A1(n4426), .A2(n3209), .B1(n4440), .B2(n2729), .ZN(n2728)
         );
  AOI211_X1 U2333 ( .C1(n3154), .C2(n2570), .A(n2707), .B(n2731), .ZN(n2733)
         );
  AND2_X1 U2334 ( .A1(n3369), .A2(n3263), .ZN(n2227) );
  NAND2_X1 U2335 ( .A1(n3253), .A2(n3251), .ZN(n2053) );
  INV_X1 U2336 ( .A(n2834), .ZN(n2071) );
  OR2_X1 U2337 ( .A1(n2008), .A2(n2292), .ZN(n2298) );
  INV_X2 U2338 ( .A(n2282), .ZN(n3392) );
  OAI21_X1 U2339 ( .B1(n2204), .B2(REG1_REG_1__SCAN_IN), .A(n2143), .ZN(n3564)
         );
  NAND2_X1 U2340 ( .A1(n2204), .A2(REG1_REG_1__SCAN_IN), .ZN(n2143) );
  NAND2_X1 U2341 ( .A1(n2078), .A2(REG1_REG_6__SCAN_IN), .ZN(n2081) );
  INV_X1 U2342 ( .A(n4266), .ZN(n2078) );
  INV_X1 U2343 ( .A(n2207), .ZN(n3593) );
  NOR2_X1 U2344 ( .A1(n3674), .A2(n3696), .ZN(n2533) );
  INV_X1 U2345 ( .A(n2237), .ZN(n2236) );
  AND2_X1 U2346 ( .A1(n3191), .A2(n3192), .ZN(n2107) );
  NAND2_X1 U2347 ( .A1(n2746), .A2(n2211), .ZN(n2210) );
  NAND2_X1 U2348 ( .A1(n4251), .A2(REG1_REG_2__SCAN_IN), .ZN(n2211) );
  NAND2_X1 U2349 ( .A1(n4297), .A2(n3599), .ZN(n3600) );
  INV_X1 U2350 ( .A(n4349), .ZN(n2074) );
  AND2_X1 U2351 ( .A1(n2042), .A2(n3483), .ZN(n2134) );
  NAND2_X1 U2352 ( .A1(n3958), .A2(n3942), .ZN(n2162) );
  NOR2_X1 U2353 ( .A1(n3406), .A2(n2139), .ZN(n2138) );
  INV_X1 U2354 ( .A(n2131), .ZN(n2130) );
  AOI21_X1 U2355 ( .B1(n2131), .B2(n2129), .A(n2128), .ZN(n2127) );
  NOR2_X1 U2356 ( .A1(n3508), .A2(n2132), .ZN(n2131) );
  NAND2_X1 U2357 ( .A1(n3016), .A2(n3458), .ZN(n2133) );
  AND2_X1 U2358 ( .A1(n2366), .A2(n2026), .ZN(n2195) );
  NOR2_X1 U2359 ( .A1(n2169), .A2(n2018), .ZN(n2166) );
  NOR2_X1 U2360 ( .A1(n2171), .A2(n2018), .ZN(n2164) );
  AND2_X1 U2361 ( .A1(n2032), .A2(n3031), .ZN(n2096) );
  INV_X1 U2362 ( .A(n4244), .ZN(n2601) );
  NAND2_X1 U2363 ( .A1(n2014), .A2(n2049), .ZN(n2216) );
  NAND2_X1 U2364 ( .A1(n2049), .A2(n2915), .ZN(n2214) );
  INV_X1 U2365 ( .A(n2109), .ZN(n2108) );
  OAI21_X1 U2366 ( .B1(n2216), .B2(n2215), .A(n2221), .ZN(n2109) );
  NAND2_X1 U2367 ( .A1(n2966), .A2(n2965), .ZN(n2221) );
  NOR2_X1 U2368 ( .A1(n2214), .A2(n2215), .ZN(n2213) );
  INV_X1 U2369 ( .A(n2105), .ZN(n2056) );
  OAI21_X1 U2370 ( .B1(n2107), .B2(n2056), .A(n3326), .ZN(n2055) );
  AND3_X1 U2371 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2336) );
  NAND2_X1 U2372 ( .A1(n2116), .A2(n2124), .ZN(n2115) );
  INV_X1 U2373 ( .A(n2118), .ZN(n2116) );
  OAI21_X1 U2374 ( .B1(n3236), .B2(n2039), .A(n2228), .ZN(n3142) );
  AOI21_X1 U2375 ( .B1(n3131), .B2(n2232), .A(n2229), .ZN(n2228) );
  NAND2_X1 U2376 ( .A1(n2810), .A2(n2807), .ZN(n2873) );
  NOR2_X1 U2377 ( .A1(n2706), .A2(n2111), .ZN(n2732) );
  NOR2_X1 U2378 ( .A1(n2758), .A2(n4417), .ZN(n2111) );
  NAND2_X1 U2379 ( .A1(n2705), .A2(n2704), .ZN(n2706) );
  NAND2_X1 U2380 ( .A1(n3055), .A2(n2106), .ZN(n2105) );
  INV_X1 U2381 ( .A(n3061), .ZN(n2106) );
  AOI21_X1 U2382 ( .B1(n2766), .B2(n2765), .A(n2764), .ZN(n3339) );
  AND2_X1 U2383 ( .A1(n2763), .A2(n2762), .ZN(n2764) );
  NOR2_X1 U2384 ( .A1(n3092), .A2(n3093), .ZN(n2225) );
  AND2_X1 U2385 ( .A1(n2019), .A2(n3098), .ZN(n2059) );
  NAND2_X1 U2386 ( .A1(n2120), .A2(n2121), .ZN(n3089) );
  AND4_X1 U2387 ( .A1(n2486), .A2(n2485), .A3(n2484), .A4(n2483), .ZN(n3521)
         );
  OR2_X1 U2388 ( .A1(n2009), .A2(n2683), .ZN(n2305) );
  NAND2_X1 U2389 ( .A1(n2282), .A2(REG1_REG_1__SCAN_IN), .ZN(n2275) );
  NOR2_X1 U2390 ( .A1(n2620), .A2(n2634), .ZN(n2615) );
  OAI21_X1 U2391 ( .B1(n4251), .B2(n4530), .A(n2083), .ZN(n2748) );
  NAND2_X1 U2392 ( .A1(n4251), .A2(n4530), .ZN(n2083) );
  XNOR2_X1 U2393 ( .A(n2210), .B(n4250), .ZN(n2672) );
  OR2_X1 U2394 ( .A1(n2796), .A2(n2077), .ZN(n2076) );
  AND2_X1 U2395 ( .A1(n2694), .A2(n4249), .ZN(n2077) );
  NAND2_X1 U2396 ( .A1(n2076), .A2(n2075), .ZN(n2209) );
  INV_X1 U2397 ( .A(n2696), .ZN(n2075) );
  AND2_X1 U2398 ( .A1(n2080), .A2(n4275), .ZN(n3597) );
  INV_X1 U2399 ( .A(n4274), .ZN(n2082) );
  NAND2_X1 U2400 ( .A1(n4298), .A2(n4299), .ZN(n4297) );
  XNOR2_X1 U2401 ( .A(n3600), .B(n2142), .ZN(n4311) );
  NAND2_X1 U2402 ( .A1(n4319), .A2(n2043), .ZN(n3603) );
  NAND2_X1 U2403 ( .A1(n4331), .A2(n3582), .ZN(n4343) );
  NAND2_X1 U2404 ( .A1(n4373), .A2(n3587), .ZN(n4381) );
  NAND2_X1 U2405 ( .A1(n4382), .A2(n2152), .ZN(n2151) );
  NAND2_X1 U2406 ( .A1(n4390), .A2(n3985), .ZN(n2152) );
  NAND2_X1 U2407 ( .A1(n3640), .A2(n3639), .ZN(n4092) );
  AND2_X1 U2408 ( .A1(n2552), .A2(n2551), .ZN(n3652) );
  NAND2_X1 U2409 ( .A1(n2174), .A2(n2175), .ZN(n3686) );
  AOI21_X1 U2410 ( .B1(n2177), .B2(n2176), .A(n2037), .ZN(n2175) );
  INV_X1 U2411 ( .A(n3697), .ZN(n3868) );
  AND2_X1 U2412 ( .A1(n3861), .A2(n2592), .ZN(n3883) );
  OR2_X1 U2413 ( .A1(n3993), .A2(n3975), .ZN(n2470) );
  AOI21_X1 U2414 ( .B1(n2011), .B2(n2187), .A(n2036), .ZN(n2183) );
  OR2_X1 U2415 ( .A1(n2428), .A2(n2427), .ZN(n2438) );
  AND2_X1 U2416 ( .A1(n2413), .A2(n2028), .ZN(n2189) );
  AOI21_X1 U2417 ( .B1(n2414), .B2(n2189), .A(n2190), .ZN(n2188) );
  NOR2_X1 U2418 ( .A1(n3550), .A2(n4052), .ZN(n2190) );
  INV_X1 U2419 ( .A(n3553), .ZN(n2978) );
  INV_X1 U2420 ( .A(n2171), .ZN(n2170) );
  OR2_X1 U2421 ( .A1(n2861), .A2(n2856), .ZN(n2893) );
  NAND2_X1 U2422 ( .A1(n2842), .A2(n2301), .ZN(n2817) );
  INV_X1 U2423 ( .A(n4412), .ZN(n4426) );
  NAND2_X1 U2424 ( .A1(n2739), .A2(n2712), .ZN(n4439) );
  NAND2_X1 U2425 ( .A1(n2597), .A2(n3423), .ZN(n4436) );
  AND2_X1 U2426 ( .A1(n2601), .A2(n3496), .ZN(n4432) );
  NOR3_X1 U2427 ( .A1(n3869), .A2(n2095), .A3(n3673), .ZN(n3680) );
  NOR2_X1 U2428 ( .A1(n3869), .A2(n2095), .ZN(n3688) );
  OR2_X1 U2429 ( .A1(n4121), .A2(n3865), .ZN(n3869) );
  NAND2_X1 U2430 ( .A1(n4420), .A2(n4486), .ZN(n4522) );
  NAND2_X1 U2431 ( .A1(n4435), .A2(n2601), .ZN(n4486) );
  NAND2_X1 U2432 ( .A1(n2622), .A2(n2006), .ZN(n2655) );
  NOR2_X1 U2433 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2256)
         );
  NOR2_X1 U2434 ( .A1(n3831), .A2(n2240), .ZN(n2126) );
  NAND2_X1 U2435 ( .A1(n2608), .A2(n2252), .ZN(n2607) );
  XNOR2_X1 U2436 ( .A(n2560), .B(n2559), .ZN(n2644) );
  INV_X1 U2437 ( .A(IR_REG_20__SCAN_IN), .ZN(n2559) );
  OR2_X1 U2438 ( .A1(n2424), .A2(IR_REG_10__SCAN_IN), .ZN(n2398) );
  NAND2_X1 U2439 ( .A1(n2308), .A2(n2299), .ZN(n2309) );
  INV_X1 U2440 ( .A(IR_REG_0__SCAN_IN), .ZN(n2068) );
  INV_X1 U2441 ( .A(n2040), .ZN(n2051) );
  AND2_X1 U2442 ( .A1(n3357), .A2(n2033), .ZN(n2052) );
  INV_X1 U2443 ( .A(n3674), .ZN(n3847) );
  NAND2_X1 U2444 ( .A1(n2734), .A2(n4241), .ZN(n3361) );
  OAI211_X1 U2445 ( .C1(n2010), .C2(n3749), .A(n2270), .B(n2269), .ZN(n3650)
         );
  INV_X1 U2446 ( .A(n2824), .ZN(n3556) );
  NAND2_X1 U2447 ( .A1(n3560), .A2(n3561), .ZN(n3559) );
  AND2_X1 U2448 ( .A1(n2790), .A2(REG1_REG_4__SCAN_IN), .ZN(n2796) );
  INV_X1 U2449 ( .A(n2081), .ZN(n4265) );
  NAND2_X1 U2450 ( .A1(n4336), .A2(n3604), .ZN(n4348) );
  OR2_X1 U2451 ( .A1(n4377), .A2(REG1_REG_16__SCAN_IN), .ZN(n2089) );
  XNOR2_X1 U2452 ( .A(n3608), .B(n3609), .ZN(n4377) );
  OR2_X1 U2453 ( .A1(n4377), .A2(n2087), .ZN(n2086) );
  OR2_X1 U2454 ( .A1(n4386), .A2(REG1_REG_16__SCAN_IN), .ZN(n2087) );
  NAND2_X1 U2455 ( .A1(n3610), .A2(n2085), .ZN(n2084) );
  INV_X1 U2456 ( .A(n4386), .ZN(n2085) );
  NAND2_X1 U2457 ( .A1(n2150), .A2(n4341), .ZN(n2149) );
  NAND2_X1 U2458 ( .A1(n2151), .A2(n4393), .ZN(n2150) );
  AOI21_X1 U2459 ( .B1(n4395), .B2(ADDR_REG_18__SCAN_IN), .A(n4394), .ZN(n2148) );
  NOR2_X1 U2460 ( .A1(n2151), .A2(n4393), .ZN(n4392) );
  OR2_X1 U2461 ( .A1(n4262), .A2(n4241), .ZN(n4401) );
  NAND2_X1 U2462 ( .A1(n4092), .A2(n2099), .ZN(n4098) );
  OR2_X1 U2463 ( .A1(n3640), .A2(n3639), .ZN(n2099) );
  NAND2_X1 U2464 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2277)
         );
  NAND2_X1 U2465 ( .A1(n3170), .A2(n2123), .ZN(n2122) );
  INV_X1 U2466 ( .A(n3169), .ZN(n2123) );
  INV_X1 U2467 ( .A(n3466), .ZN(n2128) );
  INV_X1 U2468 ( .A(n3458), .ZN(n2129) );
  NAND2_X1 U2469 ( .A1(n2202), .A2(n2201), .ZN(n2200) );
  AND2_X1 U2470 ( .A1(n2122), .A2(n2124), .ZN(n2117) );
  INV_X1 U2471 ( .A(n3139), .ZN(n2229) );
  INV_X1 U2472 ( .A(n3131), .ZN(n2230) );
  NAND2_X1 U2473 ( .A1(n2723), .A2(n3154), .ZN(n2705) );
  NAND2_X1 U2474 ( .A1(n3085), .A2(n3169), .ZN(n2121) );
  NOR2_X1 U2475 ( .A1(n3088), .A2(n2119), .ZN(n2118) );
  INV_X1 U2476 ( .A(n2121), .ZN(n2119) );
  INV_X1 U2477 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2402) );
  INV_X1 U2478 ( .A(n2210), .ZN(n2693) );
  NAND2_X1 U2479 ( .A1(n4322), .A2(n2044), .ZN(n3581) );
  NOR2_X1 U2480 ( .A1(n4362), .A2(n2153), .ZN(n3586) );
  AND2_X1 U2481 ( .A1(n3591), .A2(REG2_REG_15__SCAN_IN), .ZN(n2153) );
  NAND2_X1 U2482 ( .A1(n3690), .A2(n3484), .ZN(n2136) );
  INV_X1 U2483 ( .A(n2181), .ZN(n2176) );
  AND2_X1 U2484 ( .A1(n2437), .A2(n2263), .ZN(n2461) );
  NAND2_X1 U2485 ( .A1(n2188), .A2(n2186), .ZN(n2185) );
  INV_X1 U2486 ( .A(n2189), .ZN(n2186) );
  INV_X1 U2487 ( .A(n2188), .ZN(n2187) );
  NOR2_X1 U2488 ( .A1(n2403), .A2(n2402), .ZN(n2401) );
  NAND2_X1 U2489 ( .A1(n3285), .A2(n3255), .ZN(n2095) );
  NAND2_X1 U2490 ( .A1(n4033), .A2(n2045), .ZN(n2098) );
  AND2_X1 U2491 ( .A1(n4015), .A2(n3998), .ZN(n2097) );
  NOR2_X1 U2492 ( .A1(n4076), .A2(n4052), .ZN(n4034) );
  INV_X1 U2493 ( .A(n2990), .ZN(n2065) );
  INV_X1 U2494 ( .A(n2213), .ZN(n2062) );
  NAND2_X1 U2495 ( .A1(n2235), .A2(n2231), .ZN(n3179) );
  NAND2_X1 U2496 ( .A1(n3234), .A2(n3233), .ZN(n2234) );
  NAND2_X1 U2497 ( .A1(n3290), .A2(n2112), .ZN(n2235) );
  NOR2_X1 U2498 ( .A1(n3123), .A2(n2113), .ZN(n2112) );
  INV_X1 U2499 ( .A(n3294), .ZN(n2113) );
  INV_X1 U2500 ( .A(n3884), .ZN(n3893) );
  NAND2_X1 U2501 ( .A1(n3060), .A2(n2107), .ZN(n3190) );
  AND2_X1 U2502 ( .A1(n3105), .A2(n3104), .ZN(n3347) );
  INV_X1 U2503 ( .A(n2091), .ZN(n2090) );
  AND4_X1 U2504 ( .A1(n2516), .A2(n2515), .A3(n2514), .A4(n2513), .ZN(n3239)
         );
  NAND2_X1 U2505 ( .A1(n2747), .A2(n2748), .ZN(n2746) );
  NAND2_X1 U2506 ( .A1(n2751), .A2(n2750), .ZN(n2749) );
  NAND2_X1 U2507 ( .A1(n2209), .A2(n2208), .ZN(n2207) );
  NAND2_X1 U2508 ( .A1(n4248), .A2(REG1_REG_5__SCAN_IN), .ZN(n2208) );
  OR2_X1 U2509 ( .A1(n3570), .A2(n2146), .ZN(n3573) );
  NOR2_X1 U2510 ( .A1(n3571), .A2(n3572), .ZN(n2146) );
  NAND2_X1 U2511 ( .A1(n4292), .A2(n3598), .ZN(n4298) );
  NAND2_X1 U2512 ( .A1(n4300), .A2(n3578), .ZN(n3579) );
  NAND2_X1 U2513 ( .A1(n4310), .A2(n3601), .ZN(n4320) );
  NAND2_X1 U2514 ( .A1(n4320), .A2(n4321), .ZN(n4319) );
  XNOR2_X1 U2515 ( .A(n3581), .B(n2144), .ZN(n4332) );
  NAND2_X1 U2516 ( .A1(n4332), .A2(REG2_REG_12__SCAN_IN), .ZN(n4331) );
  OAI21_X1 U2517 ( .B1(n4336), .B2(n2074), .A(n2072), .ZN(n3605) );
  INV_X1 U2518 ( .A(n2073), .ZN(n2072) );
  OAI21_X1 U2519 ( .B1(n3604), .B2(n2074), .A(n2046), .ZN(n2073) );
  XNOR2_X1 U2520 ( .A(n3586), .B(n3609), .ZN(n4374) );
  NAND2_X1 U2521 ( .A1(n4374), .A2(n2451), .ZN(n4373) );
  NAND2_X1 U2522 ( .A1(n4367), .A2(n2203), .ZN(n3608) );
  NAND2_X1 U2523 ( .A1(n3591), .A2(REG1_REG_15__SCAN_IN), .ZN(n2203) );
  OAI21_X1 U2524 ( .B1(n2467), .B2(n2238), .A(IR_REG_31__SCAN_IN), .ZN(n2557)
         );
  INV_X1 U2525 ( .A(IR_REG_19__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U2526 ( .A1(n2135), .A2(n2024), .ZN(n2596) );
  NAND2_X1 U2527 ( .A1(n3390), .A2(n3629), .ZN(n3621) );
  NOR2_X1 U2528 ( .A1(n2535), .A2(n2534), .ZN(n3656) );
  AND2_X1 U2529 ( .A1(n3700), .A2(n3678), .ZN(n2534) );
  NAND2_X1 U2530 ( .A1(n2494), .A2(REG3_REG_22__SCAN_IN), .ZN(n2512) );
  AND2_X1 U2531 ( .A1(n3397), .A2(DATAI_23_), .ZN(n3865) );
  NAND2_X1 U2532 ( .A1(n2140), .A2(n2016), .ZN(n2591) );
  INV_X1 U2533 ( .A(n2162), .ZN(n2154) );
  NAND2_X1 U2534 ( .A1(n2158), .A2(n2162), .ZN(n2155) );
  AOI21_X1 U2535 ( .B1(n2158), .B2(n2161), .A(n2017), .ZN(n2157) );
  NAND2_X1 U2536 ( .A1(n2140), .A2(n2138), .ZN(n3916) );
  OR2_X1 U2537 ( .A1(n2481), .A2(n3202), .ZN(n2488) );
  NAND2_X1 U2538 ( .A1(n2461), .A2(REG3_REG_18__SCAN_IN), .ZN(n2481) );
  AND4_X1 U2539 ( .A1(n2479), .A2(n2478), .A3(n2477), .A4(n2476), .ZN(n3976)
         );
  NAND2_X1 U2540 ( .A1(n2140), .A2(n3405), .ZN(n3973) );
  NOR2_X1 U2541 ( .A1(n4029), .A2(n3374), .ZN(n2450) );
  INV_X1 U2542 ( .A(n2584), .ZN(n3991) );
  AND4_X1 U2543 ( .A1(n2455), .A2(n2454), .A3(n2453), .A4(n2452), .ZN(n4008)
         );
  INV_X1 U2544 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2427) );
  AND4_X1 U2545 ( .A1(n2433), .A2(n2432), .A3(n2431), .A4(n2430), .ZN(n4042)
         );
  NAND2_X1 U2546 ( .A1(n2133), .A2(n2131), .ZN(n4044) );
  NAND2_X1 U2547 ( .A1(n2133), .A2(n3465), .ZN(n4062) );
  INV_X1 U2548 ( .A(n3331), .ZN(n3064) );
  INV_X1 U2549 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U2550 ( .A1(n3003), .A2(n3457), .ZN(n2580) );
  INV_X1 U2551 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2382) );
  AND4_X1 U2552 ( .A1(n2397), .A2(n2396), .A3(n2395), .A4(n2394), .ZN(n3246)
         );
  AOI21_X1 U2553 ( .B1(n2195), .B2(n2027), .A(n2194), .ZN(n2193) );
  NOR2_X1 U2554 ( .A1(n3032), .A2(n2987), .ZN(n2194) );
  AND2_X1 U2555 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .ZN(
        n2260) );
  NAND2_X1 U2556 ( .A1(n2901), .A2(n3442), .ZN(n2575) );
  NAND2_X1 U2557 ( .A1(n2022), .A2(n2164), .ZN(n2163) );
  OAI21_X1 U2558 ( .B1(n2887), .B2(n2886), .A(n3426), .ZN(n2901) );
  NAND2_X1 U2559 ( .A1(n2781), .A2(n2619), .ZN(n2721) );
  INV_X1 U2560 ( .A(n4455), .ZN(n2619) );
  NAND2_X1 U2561 ( .A1(n4491), .A2(n2836), .ZN(n2861) );
  INV_X1 U2562 ( .A(n3520), .ZN(n2571) );
  AND2_X1 U2563 ( .A1(n4418), .A2(n2291), .ZN(n2843) );
  NAND2_X1 U2564 ( .A1(n2843), .A2(n3520), .ZN(n2842) );
  NAND2_X1 U2565 ( .A1(n4241), .A2(n2712), .ZN(n4416) );
  NAND2_X1 U2566 ( .A1(n4434), .A2(n4426), .ZN(n4425) );
  INV_X1 U2567 ( .A(n2723), .ZN(n4434) );
  NOR2_X1 U2568 ( .A1(n4092), .A2(n4095), .ZN(n4091) );
  AND2_X1 U2569 ( .A1(n4432), .A2(n4246), .ZN(n4413) );
  NOR2_X1 U2570 ( .A1(n3869), .A2(n2092), .ZN(n3657) );
  NAND2_X1 U2571 ( .A1(n2094), .A2(n2093), .ZN(n2092) );
  NOR2_X1 U2572 ( .A1(n3673), .A2(n3649), .ZN(n2094) );
  INV_X1 U2573 ( .A(n2095), .ZN(n2093) );
  INV_X1 U2574 ( .A(n3623), .ZN(n3212) );
  AND2_X1 U2575 ( .A1(n3657), .A2(n3212), .ZN(n3640) );
  NOR2_X1 U2576 ( .A1(n3923), .A2(n3905), .ZN(n3906) );
  OR2_X1 U2577 ( .A1(n3946), .A2(n3112), .ZN(n3923) );
  NOR2_X1 U2578 ( .A1(n2098), .A2(n3957), .ZN(n3963) );
  NAND2_X1 U2579 ( .A1(n3963), .A2(n3947), .ZN(n3946) );
  NAND2_X1 U2580 ( .A1(n4033), .A2(n2097), .ZN(n3997) );
  AND2_X1 U2581 ( .A1(n4034), .A2(n3173), .ZN(n4033) );
  NAND2_X1 U2582 ( .A1(n4033), .A2(n4015), .ZN(n4017) );
  OR2_X1 U2583 ( .A1(n4074), .A2(n4073), .ZN(n4076) );
  NAND2_X1 U2584 ( .A1(n2906), .A2(n2035), .ZN(n3009) );
  NOR2_X1 U2585 ( .A1(n3009), .A2(n3193), .ZN(n3022) );
  NAND2_X1 U2586 ( .A1(n2906), .A2(n2096), .ZN(n3028) );
  AND2_X1 U2587 ( .A1(n2906), .A2(n2902), .ZN(n2955) );
  NOR2_X1 U2588 ( .A1(n2893), .A2(n2892), .ZN(n2906) );
  NOR2_X1 U2589 ( .A1(n4425), .A2(n3343), .ZN(n4491) );
  AND2_X1 U2590 ( .A1(n2832), .A2(n2635), .ZN(n2646) );
  XNOR2_X1 U2591 ( .A(n2568), .B(n2567), .ZN(n2739) );
  NAND2_X1 U2592 ( .A1(n2616), .A2(n2201), .ZN(n2618) );
  NAND2_X1 U2593 ( .A1(n2101), .A2(n2100), .ZN(n2237) );
  INV_X1 U2594 ( .A(n2238), .ZN(n2101) );
  INV_X1 U2595 ( .A(IR_REG_9__SCAN_IN), .ZN(n2379) );
  INV_X1 U2596 ( .A(IR_REG_4__SCAN_IN), .ZN(n2067) );
  CLKBUF_X1 U2597 ( .A(n2331), .Z(n2332) );
  NAND2_X1 U2598 ( .A1(n2217), .A2(n2216), .ZN(n2943) );
  INV_X1 U2599 ( .A(n2214), .ZN(n2212) );
  NAND2_X1 U2600 ( .A1(n2943), .A2(n2942), .ZN(n2967) );
  NAND2_X1 U2601 ( .A1(n3179), .A2(n3131), .ZN(n3182) );
  INV_X1 U2602 ( .A(n3552), .ZN(n3032) );
  NAND2_X1 U2603 ( .A1(n2916), .A2(n2213), .ZN(n2064) );
  OAI21_X1 U2604 ( .B1(n3397), .B2(n2204), .A(n2278), .ZN(n4412) );
  NAND2_X1 U2605 ( .A1(n3397), .A2(DATAI_1_), .ZN(n2278) );
  INV_X1 U2606 ( .A(n2762), .ZN(n2730) );
  NAND2_X1 U2607 ( .A1(n3290), .A2(n3294), .ZN(n3236) );
  AND2_X1 U2608 ( .A1(n3397), .A2(DATAI_21_), .ZN(n3905) );
  INV_X1 U2609 ( .A(n3328), .ZN(n2057) );
  OAI21_X1 U2610 ( .B1(n3060), .B2(n2056), .A(n2054), .ZN(n2058) );
  INV_X1 U2611 ( .A(n2055), .ZN(n2054) );
  NAND2_X1 U2612 ( .A1(n2226), .A2(n2224), .ZN(n3274) );
  INV_X1 U2613 ( .A(n2225), .ZN(n2224) );
  NAND2_X1 U2614 ( .A1(n2019), .A2(n2227), .ZN(n2226) );
  OAI21_X1 U2615 ( .B1(n3397), .B2(n2289), .A(n2288), .ZN(n2723) );
  NAND2_X1 U2616 ( .A1(n3397), .A2(DATAI_0_), .ZN(n2288) );
  INV_X1 U2617 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3297) );
  NAND2_X1 U2618 ( .A1(n2734), .A2(n2739), .ZN(n3363) );
  NAND2_X1 U2619 ( .A1(n2235), .A2(n2234), .ZN(n3318) );
  NAND2_X1 U2620 ( .A1(n3190), .A2(n2105), .ZN(n3330) );
  INV_X1 U2621 ( .A(n3381), .ZN(n3340) );
  NAND2_X1 U2622 ( .A1(n2104), .A2(n2223), .ZN(n3351) );
  NAND2_X1 U2623 ( .A1(n2038), .A2(n3098), .ZN(n2223) );
  NAND2_X1 U2624 ( .A1(n2227), .A2(n2059), .ZN(n2104) );
  AND2_X1 U2625 ( .A1(n2219), .A2(n2222), .ZN(n2938) );
  NAND2_X1 U2626 ( .A1(n2916), .A2(n2915), .ZN(n2219) );
  AND2_X1 U2627 ( .A1(n3091), .A2(n3090), .ZN(n3370) );
  INV_X1 U2628 ( .A(n3362), .ZN(n3375) );
  INV_X1 U2629 ( .A(n3361), .ZN(n3373) );
  INV_X1 U2630 ( .A(n3363), .ZN(n3378) );
  NAND2_X1 U2631 ( .A1(n2540), .A2(n2539), .ZN(n3548) );
  OAI211_X1 U2632 ( .C1(n2009), .C2(n2532), .A(n2531), .B(n2530), .ZN(n3674)
         );
  AND2_X1 U2633 ( .A1(n2522), .A2(n2521), .ZN(n2525) );
  AND4_X1 U2634 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n3919)
         );
  NAND4_X1 U2635 ( .A1(n2493), .A2(n2492), .A3(n2491), .A4(n2490), .ZN(n3943)
         );
  INV_X1 U2636 ( .A(n3521), .ZN(n3958) );
  INV_X1 U2637 ( .A(n3246), .ZN(n4066) );
  INV_X1 U2638 ( .A(n2970), .ZN(n3554) );
  OR2_X1 U2639 ( .A1(n2007), .A2(REG3_REG_3__SCAN_IN), .ZN(n2306) );
  OR2_X1 U2640 ( .A1(n2007), .A2(n2281), .ZN(n2286) );
  NOR2_X1 U2641 ( .A1(n2688), .A2(n2687), .ZN(n3570) );
  INV_X1 U2642 ( .A(n2076), .ZN(n2697) );
  INV_X1 U2643 ( .A(n2209), .ZN(n3592) );
  XNOR2_X1 U2644 ( .A(n2207), .B(n3594), .ZN(n4266) );
  NOR2_X1 U2645 ( .A1(n4265), .A2(n3595), .ZN(n4278) );
  XNOR2_X1 U2646 ( .A(n3597), .B(n4296), .ZN(n4293) );
  NAND2_X1 U2647 ( .A1(n4287), .A2(n3577), .ZN(n4301) );
  NAND2_X1 U2648 ( .A1(n4301), .A2(n4302), .ZN(n4300) );
  XNOR2_X1 U2649 ( .A(n3579), .B(n2142), .ZN(n4313) );
  INV_X1 U2650 ( .A(n4470), .ZN(n4327) );
  XNOR2_X1 U2651 ( .A(n3603), .B(n2144), .ZN(n4337) );
  XNOR2_X1 U2652 ( .A(n2557), .B(n2556), .ZN(n3616) );
  AND2_X1 U2653 ( .A1(n2178), .A2(n2180), .ZN(n3839) );
  NAND2_X1 U2654 ( .A1(n2179), .A2(n2181), .ZN(n2178) );
  NAND2_X1 U2655 ( .A1(n2156), .A2(n2158), .ZN(n3931) );
  NAND2_X1 U2656 ( .A1(n2472), .A2(n2160), .ZN(n2156) );
  NAND2_X1 U2657 ( .A1(n2472), .A2(n2471), .ZN(n3954) );
  NAND2_X1 U2658 ( .A1(n2184), .A2(n2188), .ZN(n4025) );
  NAND2_X1 U2659 ( .A1(n4072), .A2(n2189), .ZN(n2184) );
  NAND2_X1 U2660 ( .A1(n2192), .A2(n2366), .ZN(n2981) );
  OR2_X1 U2661 ( .A1(n3029), .A2(n2027), .ZN(n2192) );
  INV_X1 U2662 ( .A(n4004), .ZN(n4081) );
  NAND2_X1 U2663 ( .A1(n2167), .A2(n2168), .ZN(n2900) );
  OR2_X1 U2664 ( .A1(n2854), .A2(n2170), .ZN(n2167) );
  NAND2_X1 U2665 ( .A1(n2854), .A2(n3526), .ZN(n2173) );
  OR2_X1 U2666 ( .A1(n3965), .A2(n4519), .ZN(n4079) );
  INV_X1 U2667 ( .A(n4055), .ZN(n4442) );
  AND2_X2 U2668 ( .A1(n2646), .A2(n2709), .ZN(n4540) );
  XOR2_X1 U2669 ( .A(n4088), .B(n4091), .Z(n4253) );
  OAI21_X1 U2670 ( .B1(n4098), .B2(n4519), .A(n2023), .ZN(n4184) );
  OR2_X1 U2671 ( .A1(n3680), .A2(n3679), .ZN(n4189) );
  AND2_X2 U2672 ( .A1(n2646), .A2(n2831), .ZN(n4525) );
  INV_X1 U2673 ( .A(IR_REG_29__SCAN_IN), .ZN(n2258) );
  INV_X1 U2674 ( .A(n2739), .ZN(n4241) );
  NAND2_X1 U2675 ( .A1(n2613), .A2(n2612), .ZN(n2614) );
  NAND2_X1 U2676 ( .A1(n3831), .A2(n2240), .ZN(n2612) );
  NAND2_X1 U2677 ( .A1(n2607), .A2(n2126), .ZN(n2613) );
  NAND2_X1 U2678 ( .A1(n2777), .A2(STATE_REG_SCAN_IN), .ZN(n4455) );
  XNOR2_X1 U2679 ( .A(n2562), .B(IR_REG_22__SCAN_IN), .ZN(n4244) );
  INV_X1 U2680 ( .A(n3616), .ZN(n4247) );
  AND2_X1 U2681 ( .A1(n2320), .A2(n2311), .ZN(n4250) );
  OR2_X1 U2682 ( .A1(n2299), .A2(n3831), .ZN(n2300) );
  XNOR2_X1 U2683 ( .A(n3208), .B(n3207), .ZN(n3168) );
  NAND2_X1 U2684 ( .A1(n3565), .A2(n2206), .ZN(n3566) );
  NAND2_X1 U2685 ( .A1(n4348), .A2(n4349), .ZN(n4347) );
  NAND2_X1 U2686 ( .A1(n2084), .A2(n2086), .ZN(n4387) );
  INV_X1 U2687 ( .A(n2147), .ZN(n4400) );
  OAI21_X1 U2688 ( .B1(n4392), .B2(n2149), .A(n2148), .ZN(n2147) );
  NAND2_X1 U2689 ( .A1(U3149), .A2(DATAI_1_), .ZN(n2205) );
  AND2_X1 U2690 ( .A1(n2185), .A2(n4024), .ZN(n2011) );
  AND3_X1 U2691 ( .A1(n2086), .A2(n2084), .A3(n2050), .ZN(n2012) );
  AND2_X1 U2692 ( .A1(n2034), .A2(n3655), .ZN(n2013) );
  OR2_X1 U2693 ( .A1(n2218), .A2(n2220), .ZN(n2014) );
  NOR2_X1 U2694 ( .A1(n2518), .A2(n2031), .ZN(n2177) );
  NAND2_X1 U2695 ( .A1(n3976), .A2(n3962), .ZN(n2015) );
  AND2_X1 U2696 ( .A1(n2138), .A2(n2137), .ZN(n2016) );
  AND2_X1 U2697 ( .A1(n3521), .A2(n3947), .ZN(n2017) );
  NAND2_X1 U2698 ( .A1(n2159), .A2(n2015), .ZN(n2158) );
  INV_X1 U2699 ( .A(n2641), .ZN(n3031) );
  INV_X1 U2700 ( .A(n4424), .ZN(n4058) );
  INV_X1 U2701 ( .A(n3673), .ZN(n3678) );
  AND2_X1 U2702 ( .A1(n3397), .A2(DATAI_26_), .ZN(n3673) );
  AND2_X1 U2703 ( .A1(n3397), .A2(DATAI_25_), .ZN(n3696) );
  AND2_X1 U2704 ( .A1(n2456), .A2(n2448), .ZN(n3591) );
  NOR2_X1 U2705 ( .A1(n2923), .A2(n2892), .ZN(n2018) );
  AND2_X1 U2706 ( .A1(n2114), .A2(n2115), .ZN(n2019) );
  AND3_X1 U2707 ( .A1(n2141), .A2(n2196), .A3(n2198), .ZN(n2554) );
  XOR2_X1 U2708 ( .A(n2259), .B(n2258), .Z(n2020) );
  OR2_X1 U2709 ( .A1(n3083), .A2(n3308), .ZN(n2021) );
  INV_X1 U2710 ( .A(n4519), .ZN(n4512) );
  NAND2_X1 U2711 ( .A1(n4432), .A2(n2644), .ZN(n4519) );
  OR2_X1 U2712 ( .A1(n3555), .A2(n2924), .ZN(n2022) );
  NAND2_X1 U2713 ( .A1(n2554), .A2(n2251), .ZN(n2605) );
  AND2_X1 U2714 ( .A1(n4099), .A2(n4100), .ZN(n2023) );
  OR2_X1 U2715 ( .A1(n2013), .A2(n2595), .ZN(n2024) );
  INV_X1 U2716 ( .A(IR_REG_22__SCAN_IN), .ZN(n2251) );
  OR2_X1 U2717 ( .A1(n2467), .A2(n2237), .ZN(n2025) );
  AND2_X1 U2718 ( .A1(n2554), .A2(n2199), .ZN(n2608) );
  OR2_X1 U2719 ( .A1(n3552), .A2(n2995), .ZN(n2026) );
  AND2_X1 U2720 ( .A1(n3553), .A2(n2641), .ZN(n2027) );
  INV_X1 U2721 ( .A(IR_REG_1__SCAN_IN), .ZN(n2069) );
  NAND2_X1 U2722 ( .A1(n3550), .A2(n4052), .ZN(n2028) );
  AND2_X1 U2723 ( .A1(n2199), .A2(n2239), .ZN(n2029) );
  AND2_X1 U2724 ( .A1(n2089), .A2(n2088), .ZN(n2030) );
  INV_X1 U2725 ( .A(IR_REG_31__SCAN_IN), .ZN(n3831) );
  INV_X1 U2726 ( .A(n3594), .ZN(n2145) );
  INV_X1 U2727 ( .A(n4024), .ZN(n2436) );
  INV_X1 U2728 ( .A(IR_REG_26__SCAN_IN), .ZN(n2240) );
  INV_X1 U2729 ( .A(IR_REG_21__SCAN_IN), .ZN(n2250) );
  AND2_X1 U2730 ( .A1(n3697), .A2(n3848), .ZN(n2031) );
  AOI21_X1 U2731 ( .B1(n3913), .B2(n3498), .A(n3500), .ZN(n3898) );
  AND2_X1 U2732 ( .A1(n2902), .A2(n2951), .ZN(n2032) );
  OAI21_X1 U2733 ( .B1(n4072), .B2(n2414), .A(n2413), .ZN(n4050) );
  OR2_X1 U2734 ( .A1(n3149), .A2(n3148), .ZN(n2033) );
  AOI21_X1 U2735 ( .B1(n3898), .B2(n2503), .A(n2502), .ZN(n3878) );
  INV_X1 U2736 ( .A(n3878), .ZN(n2179) );
  INV_X1 U2737 ( .A(IR_REG_23__SCAN_IN), .ZN(n2201) );
  INV_X1 U2738 ( .A(IR_REG_24__SCAN_IN), .ZN(n2202) );
  AND2_X1 U2739 ( .A1(n3943), .A2(n3924), .ZN(n3409) );
  INV_X1 U2740 ( .A(n3409), .ZN(n2137) );
  INV_X1 U2741 ( .A(n2161), .ZN(n2160) );
  NAND2_X1 U2742 ( .A1(n2471), .A2(n2015), .ZN(n2161) );
  INV_X1 U2743 ( .A(n2232), .ZN(n2231) );
  NAND2_X1 U2744 ( .A1(n2233), .A2(n2234), .ZN(n2232) );
  AND2_X1 U2745 ( .A1(n2594), .A2(n3515), .ZN(n2034) );
  NAND2_X1 U2746 ( .A1(n2120), .A2(n2118), .ZN(n2125) );
  INV_X1 U2747 ( .A(n3993), .ZN(n3352) );
  AND4_X1 U2748 ( .A1(n2466), .A2(n2465), .A3(n2464), .A4(n2463), .ZN(n3993)
         );
  OR2_X1 U2749 ( .A1(n3548), .A2(n3659), .ZN(n3389) );
  AND2_X1 U2750 ( .A1(n2096), .A2(n2987), .ZN(n2035) );
  AND2_X1 U2751 ( .A1(n4042), .A2(n3173), .ZN(n2036) );
  AND2_X1 U2752 ( .A1(n3868), .A2(n3285), .ZN(n2037) );
  OR2_X1 U2753 ( .A1(n3097), .A2(n2225), .ZN(n2038) );
  OR2_X1 U2754 ( .A1(n2230), .A2(n3123), .ZN(n2039) );
  NAND2_X1 U2755 ( .A1(n3159), .A2(n3158), .ZN(n2040) );
  OR2_X1 U2756 ( .A1(n3869), .A2(n3848), .ZN(n2041) );
  AND2_X1 U2757 ( .A1(n3484), .A2(n3389), .ZN(n2042) );
  INV_X1 U2758 ( .A(n2518), .ZN(n2180) );
  INV_X1 U2759 ( .A(IR_REG_27__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U2760 ( .A1(n2833), .A2(n4055), .ZN(n4445) );
  INV_X1 U2761 ( .A(n3602), .ZN(n2144) );
  NAND2_X1 U2762 ( .A1(n2993), .A2(n2994), .ZN(n3060) );
  AOI21_X1 U2763 ( .B1(n2169), .B2(n2171), .A(n2018), .ZN(n2168) );
  INV_X1 U2764 ( .A(n3957), .ZN(n3962) );
  XNOR2_X1 U2765 ( .A(n2606), .B(n2202), .ZN(n2620) );
  NAND2_X1 U2766 ( .A1(n2173), .A2(n2322), .ZN(n2885) );
  INV_X1 U2767 ( .A(n3405), .ZN(n2139) );
  INV_X1 U2768 ( .A(n3465), .ZN(n2132) );
  INV_X1 U2769 ( .A(n3956), .ZN(n2159) );
  NAND2_X1 U2770 ( .A1(n2196), .A2(n2198), .ZN(n2467) );
  OR2_X1 U2771 ( .A1(n4327), .A2(n3808), .ZN(n2043) );
  INV_X1 U2772 ( .A(n2642), .ZN(n3998) );
  OR2_X1 U2773 ( .A1(n4327), .A2(n3024), .ZN(n2044) );
  AND2_X1 U2774 ( .A1(n2097), .A2(n3975), .ZN(n2045) );
  OR2_X1 U2775 ( .A1(n4352), .A2(n3706), .ZN(n2046) );
  OR2_X1 U2776 ( .A1(n2467), .A2(IR_REG_17__SCAN_IN), .ZN(n2047) );
  AND2_X1 U2777 ( .A1(n2906), .A2(n2032), .ZN(n2048) );
  INV_X1 U2778 ( .A(n3649), .ZN(n3659) );
  AND2_X1 U2779 ( .A1(n3397), .A2(DATAI_27_), .ZN(n3649) );
  OR2_X1 U2780 ( .A1(n4262), .A2(n2743), .ZN(n4391) );
  NAND2_X1 U2781 ( .A1(n2921), .A2(n2920), .ZN(n2049) );
  AND2_X1 U2782 ( .A1(n3397), .A2(DATAI_24_), .ZN(n3848) );
  INV_X1 U2783 ( .A(n2222), .ZN(n2220) );
  INV_X1 U2784 ( .A(n4309), .ZN(n2142) );
  NOR2_X1 U2785 ( .A1(n2257), .A2(IR_REG_29__SCAN_IN), .ZN(n3041) );
  OR2_X1 U2786 ( .A1(n4459), .A2(REG1_REG_17__SCAN_IN), .ZN(n2050) );
  INV_X1 U2787 ( .A(n3366), .ZN(n3376) );
  AOI21_X2 U2788 ( .B1(n2783), .B2(n2782), .A(U3149), .ZN(n3366) );
  NAND2_X1 U2789 ( .A1(n2108), .A2(n2065), .ZN(n2063) );
  INV_X1 U2790 ( .A(n2063), .ZN(n2060) );
  NAND2_X1 U2791 ( .A1(n2062), .A2(n2060), .ZN(n2061) );
  OAI211_X1 U2792 ( .C1(n2916), .C2(n2063), .A(n2061), .B(n2989), .ZN(n2066)
         );
  NAND3_X1 U2793 ( .A1(n2299), .A2(n2070), .A3(n3776), .ZN(n2329) );
  NAND2_X2 U2794 ( .A1(n2071), .A2(n2781), .ZN(n2729) );
  XNOR2_X1 U2795 ( .A(n3605), .B(n4466), .ZN(n4359) );
  NAND2_X1 U2796 ( .A1(n2079), .A2(n2081), .ZN(n2080) );
  NOR2_X1 U2797 ( .A1(n3595), .A2(n2082), .ZN(n2079) );
  INV_X1 U2798 ( .A(n2089), .ZN(n4378) );
  INV_X1 U2799 ( .A(n3610), .ZN(n2088) );
  OAI21_X1 U2800 ( .B1(n2652), .B2(IR_REG_28__SCAN_IN), .A(n2254), .ZN(n2091)
         );
  NAND2_X1 U2801 ( .A1(n2253), .A2(IR_REG_31__SCAN_IN), .ZN(n2652) );
  INV_X1 U2802 ( .A(n2098), .ZN(n3982) );
  NAND2_X1 U2803 ( .A1(n3172), .A2(n2117), .ZN(n2114) );
  NAND2_X1 U2804 ( .A1(n3172), .A2(n2122), .ZN(n2120) );
  INV_X1 U2805 ( .A(n2125), .ZN(n3262) );
  INV_X1 U2806 ( .A(n3370), .ZN(n2124) );
  OAI21_X1 U2807 ( .B1(n3016), .B2(n2130), .A(n2127), .ZN(n2581) );
  OAI21_X2 U2808 ( .B1(n2855), .B2(n2574), .A(n3444), .ZN(n2887) );
  NAND2_X1 U2809 ( .A1(n3841), .A2(n2134), .ZN(n2135) );
  NAND2_X1 U2810 ( .A1(n3992), .A2(n3991), .ZN(n2140) );
  INV_X1 U2811 ( .A(n2253), .ZN(n2564) );
  NAND4_X1 U2812 ( .A1(n2141), .A2(n2198), .A3(n2029), .A4(n2196), .ZN(n2253)
         );
  XNOR2_X2 U2813 ( .A(n2277), .B(n2069), .ZN(n2204) );
  XNOR2_X1 U2814 ( .A(n2685), .B(n2799), .ZN(n2791) );
  OAI21_X1 U2815 ( .B1(n2684), .B2(n2683), .A(n2682), .ZN(n2685) );
  NOR2_X1 U2816 ( .A1(n4364), .A2(n4363), .ZN(n4362) );
  NOR2_X1 U2817 ( .A1(n3584), .A2(n4354), .ZN(n4364) );
  NAND3_X1 U2818 ( .A1(n2166), .A2(n2022), .A3(n2854), .ZN(n2165) );
  NAND3_X1 U2819 ( .A1(n2165), .A2(n2163), .A3(n2342), .ZN(n2961) );
  INV_X1 U2820 ( .A(n3526), .ZN(n2169) );
  INV_X1 U2821 ( .A(n2322), .ZN(n2172) );
  NAND2_X1 U2822 ( .A1(n3878), .A2(n2177), .ZN(n2174) );
  NOR2_X1 U2823 ( .A1(n2517), .A2(n3883), .ZN(n2181) );
  NAND2_X1 U2824 ( .A1(n4072), .A2(n2011), .ZN(n2182) );
  NAND2_X1 U2825 ( .A1(n2182), .A2(n2183), .ZN(n4012) );
  NAND2_X1 U2826 ( .A1(n3029), .A2(n2195), .ZN(n2191) );
  NAND2_X1 U2827 ( .A1(n2191), .A2(n2193), .ZN(n3008) );
  NOR2_X1 U2828 ( .A1(n2331), .A2(n2248), .ZN(n2434) );
  INV_X1 U2829 ( .A(n2248), .ZN(n2197) );
  INV_X1 U2830 ( .A(n2331), .ZN(n2198) );
  OR2_X1 U2831 ( .A1(n2204), .A2(n4528), .ZN(n2671) );
  OR2_X1 U2832 ( .A1(n2204), .A2(n2668), .ZN(n2669) );
  OAI21_X1 U2833 ( .B1(n2204), .B2(U3149), .A(n2205), .ZN(U3351) );
  MUX2_X1 U2834 ( .A(n2668), .B(REG2_REG_1__SCAN_IN), .S(n2204), .Z(n3560) );
  INV_X1 U2835 ( .A(n2204), .ZN(n2206) );
  INV_X1 U2836 ( .A(n2942), .ZN(n2215) );
  NAND2_X1 U2837 ( .A1(n2916), .A2(n2212), .ZN(n2217) );
  INV_X1 U2838 ( .A(n2937), .ZN(n2218) );
  NAND2_X1 U2839 ( .A1(n2913), .A2(n2914), .ZN(n2222) );
  INV_X1 U2840 ( .A(n3319), .ZN(n2233) );
  NAND2_X1 U2841 ( .A1(n3906), .A2(n3893), .ZN(n4121) );
  XNOR2_X2 U2842 ( .A(n2300), .B(IR_REG_2__SCAN_IN), .ZN(n4251) );
  OR2_X1 U2843 ( .A1(n2547), .A2(n2271), .ZN(n2276) );
  INV_X1 U2844 ( .A(n2547), .ZN(n3383) );
  NAND2_X1 U2845 ( .A1(n2726), .A2(n4412), .ZN(n3432) );
  AOI22_X2 U2846 ( .A1(n3990), .A2(n2584), .B1(n2642), .B2(n3978), .ZN(n3972)
         );
  NAND2_X1 U2847 ( .A1(n2257), .A2(IR_REG_31__SCAN_IN), .ZN(n2259) );
  OR2_X1 U2848 ( .A1(n3047), .A2(n4238), .ZN(n2241) );
  OR2_X1 U2849 ( .A1(n3047), .A2(n4176), .ZN(n2242) );
  OR2_X1 U2850 ( .A1(n3677), .A2(n3659), .ZN(n2243) );
  INV_X1 U2851 ( .A(IR_REG_30__SCAN_IN), .ZN(n3042) );
  XNOR2_X1 U2852 ( .A(n2268), .B(n3042), .ZN(n2279) );
  NAND2_X1 U2853 ( .A1(n3182), .A2(n3137), .ZN(n3280) );
  INV_X1 U2854 ( .A(IR_REG_0__SCAN_IN), .ZN(n2289) );
  AND2_X1 U2855 ( .A1(n3861), .A2(n3859), .ZN(n3480) );
  AND2_X1 U2856 ( .A1(n3505), .A2(n3840), .ZN(n3483) );
  INV_X1 U2857 ( .A(IR_REG_25__SCAN_IN), .ZN(n2252) );
  AND2_X1 U2858 ( .A1(n3139), .A2(n3140), .ZN(n3137) );
  AND2_X1 U2859 ( .A1(n2487), .A2(REG3_REG_21__SCAN_IN), .ZN(n2494) );
  NOR2_X1 U2860 ( .A1(n2488), .A2(n3297), .ZN(n2487) );
  NOR2_X1 U2861 ( .A1(n2438), .A2(n3824), .ZN(n2437) );
  NAND2_X1 U2862 ( .A1(n3624), .A2(n3623), .ZN(n3625) );
  NAND2_X1 U2863 ( .A1(n2272), .A2(REG3_REG_1__SCAN_IN), .ZN(n2273) );
  AND2_X1 U2864 ( .A1(n3397), .A2(DATAI_22_), .ZN(n3884) );
  NAND2_X1 U2865 ( .A1(n2772), .A2(n2771), .ZN(n2773) );
  AND2_X1 U2866 ( .A1(n2716), .A2(n3542), .ZN(n2734) );
  AND2_X1 U2867 ( .A1(n2546), .A2(n3638), .ZN(n3223) );
  OR2_X1 U2868 ( .A1(n2512), .A2(n3184), .ZN(n2519) );
  OR2_X1 U2869 ( .A1(n3266), .A2(n4015), .ZN(n2449) );
  OR2_X1 U2870 ( .A1(n2392), .A2(n3747), .ZN(n2403) );
  OR2_X1 U2871 ( .A1(n2383), .A2(n2382), .ZN(n2392) );
  INV_X1 U2872 ( .A(n4439), .ZN(n4414) );
  INV_X1 U2873 ( .A(n3631), .ZN(n3627) );
  NAND2_X1 U2874 ( .A1(n2652), .A2(IR_REG_27__SCAN_IN), .ZN(n2255) );
  INV_X1 U2875 ( .A(n2957), .ZN(n2951) );
  INV_X1 U2876 ( .A(n4035), .ZN(n3173) );
  INV_X1 U2877 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3202) );
  INV_X1 U2878 ( .A(n4029), .ZN(n3266) );
  INV_X1 U2879 ( .A(n3848), .ZN(n3285) );
  AND2_X1 U2880 ( .A1(n2809), .A2(n2808), .ZN(n2807) );
  AND2_X1 U2881 ( .A1(n3079), .A2(n3080), .ZN(n3309) );
  AND2_X1 U2882 ( .A1(n2774), .A2(n2773), .ZN(n3338) );
  XNOR2_X1 U2883 ( .A(n2877), .B(n3210), .ZN(n2913) );
  AND2_X1 U2884 ( .A1(n4244), .A2(n4245), .ZN(n2712) );
  OR2_X1 U2885 ( .A1(n2519), .A2(n3284), .ZN(n2527) );
  INV_X1 U2886 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3824) );
  OR2_X1 U2887 ( .A1(n4262), .A2(n4259), .ZN(n4264) );
  AND2_X1 U2888 ( .A1(n3389), .A2(n3488), .ZN(n3655) );
  INV_X1 U2889 ( .A(n3686), .ZN(n3687) );
  NAND2_X1 U2890 ( .A1(n3993), .A2(n3975), .ZN(n2471) );
  INV_X1 U2891 ( .A(n4012), .ZN(n4013) );
  OR2_X1 U2892 ( .A1(n4486), .A2(n4245), .ZN(n2720) );
  INV_X1 U2893 ( .A(n4413), .ZN(n4087) );
  AND2_X1 U2894 ( .A1(n3397), .A2(DATAI_20_), .ZN(n3112) );
  INV_X1 U2895 ( .A(n3374), .ZN(n4015) );
  INV_X1 U2896 ( .A(n4436), .ZN(n4069) );
  NOR2_X1 U2897 ( .A1(n2718), .A2(n2708), .ZN(n2832) );
  INV_X1 U2898 ( .A(n3975), .ZN(n3981) );
  MUX2_X1 U2899 ( .A(n4251), .B(DATAI_2_), .S(n3397), .Z(n3343) );
  NAND2_X1 U2900 ( .A1(n2618), .A2(n2617), .ZN(n2777) );
  INV_X1 U2901 ( .A(n3239), .ZN(n3901) );
  INV_X1 U2902 ( .A(n4391), .ZN(n4341) );
  INV_X1 U2903 ( .A(n4264), .ZN(n4397) );
  INV_X1 U2904 ( .A(n4416), .ZN(n4067) );
  INV_X1 U2905 ( .A(n4420), .ZN(n4437) );
  INV_X1 U2906 ( .A(n4079), .ZN(n4428) );
  OR2_X1 U2907 ( .A1(n2721), .A2(n2720), .ZN(n4055) );
  AND2_X1 U2908 ( .A1(n2639), .A2(n2638), .ZN(n2709) );
  INV_X1 U2909 ( .A(n2709), .ZN(n2831) );
  AND2_X1 U2910 ( .A1(n2381), .A2(n2424), .ZN(n4472) );
  AND2_X1 U2911 ( .A1(n2364), .A2(n2350), .ZN(n3596) );
  AND2_X1 U2912 ( .A1(n2667), .A2(n2662), .ZN(n4395) );
  NAND2_X1 U2913 ( .A1(n2722), .A2(n2714), .ZN(n3381) );
  INV_X1 U2914 ( .A(n3652), .ZN(n3624) );
  OAI211_X1 U2915 ( .C1(n2007), .C2(n3283), .A(n2525), .B(n2524), .ZN(n3697)
         );
  INV_X1 U2916 ( .A(n4008), .ZN(n3978) );
  OR2_X1 U2917 ( .A1(n2781), .A2(n4455), .ZN(n3558) );
  INV_X1 U2918 ( .A(n4459), .ZN(n4390) );
  AND2_X1 U2919 ( .A1(n2884), .A2(n2883), .ZN(n4004) );
  NAND2_X1 U2920 ( .A1(n4540), .A2(n4512), .ZN(n4176) );
  INV_X1 U2921 ( .A(n4540), .ZN(n4538) );
  NAND2_X1 U2922 ( .A1(n4525), .A2(n4512), .ZN(n4238) );
  AND2_X1 U2923 ( .A1(n4500), .A2(n4499), .ZN(n4533) );
  INV_X1 U2924 ( .A(n4452), .ZN(n4454) );
  NAND2_X1 U2925 ( .A1(n2711), .A2(n2655), .ZN(n4452) );
  INV_X1 U2926 ( .A(n3596), .ZN(n4477) );
  INV_X2 U2927 ( .A(n3558), .ZN(U4043) );
  NAND4_X1 U2928 ( .A1(n2375), .A2(n2247), .A3(n2246), .A4(n2245), .ZN(n2248)
         );
  NAND2_X1 U2929 ( .A1(n2565), .A2(IR_REG_28__SCAN_IN), .ZN(n2254) );
  NAND2_X1 U2930 ( .A1(n2564), .A2(n2256), .ZN(n2257) );
  NAND2_X1 U2931 ( .A1(n2336), .A2(REG3_REG_6__SCAN_IN), .ZN(n2356) );
  INV_X1 U2932 ( .A(n2356), .ZN(n2261) );
  NAND2_X1 U2933 ( .A1(n2261), .A2(n2260), .ZN(n2368) );
  INV_X1 U2934 ( .A(n2368), .ZN(n2262) );
  NAND2_X1 U2935 ( .A1(n2262), .A2(REG3_REG_9__SCAN_IN), .ZN(n2383) );
  NAND2_X1 U2936 ( .A1(n2401), .A2(REG3_REG_13__SCAN_IN), .ZN(n2428) );
  AND2_X1 U2937 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2263) );
  INV_X1 U2938 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3184) );
  INV_X1 U2939 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3284) );
  INV_X1 U2940 ( .A(n2527), .ZN(n2264) );
  NAND2_X1 U2941 ( .A1(n2264), .A2(REG3_REG_25__SCAN_IN), .ZN(n2529) );
  INV_X1 U2942 ( .A(n2529), .ZN(n2265) );
  NAND2_X1 U2943 ( .A1(n2265), .A2(REG3_REG_26__SCAN_IN), .ZN(n2545) );
  INV_X1 U2944 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U2945 ( .A1(n2529), .A2(n3744), .ZN(n2266) );
  NAND2_X1 U2946 ( .A1(n2545), .A2(n2266), .ZN(n3360) );
  OR2_X1 U2947 ( .A1(n3360), .A2(n2008), .ZN(n2270) );
  INV_X1 U2948 ( .A(n4240), .ZN(n2267) );
  AND2_X2 U2949 ( .A1(n2279), .A2(n2020), .ZN(n2282) );
  AOI22_X1 U2950 ( .A1(n3383), .A2(REG0_REG_26__SCAN_IN), .B1(n2282), .B2(
        REG1_REG_26__SCAN_IN), .ZN(n2269) );
  INV_X1 U2951 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2271) );
  INV_X1 U2952 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2668) );
  INV_X1 U2953 ( .A(n2726), .ZN(n2290) );
  NAND2_X1 U2954 ( .A1(n2290), .A2(n4426), .ZN(n3430) );
  NAND2_X1 U2955 ( .A1(n3393), .A2(REG0_REG_0__SCAN_IN), .ZN(n2287) );
  INV_X1 U2956 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2281) );
  INV_X1 U2957 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4526) );
  OR2_X1 U2958 ( .A1(n3392), .A2(n4526), .ZN(n2285) );
  INV_X1 U2959 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2283) );
  AND2_X1 U2960 ( .A1(n2570), .A2(n2723), .ZN(n4419) );
  NAND2_X1 U2961 ( .A1(n2569), .A2(n4419), .ZN(n4418) );
  NAND2_X1 U2962 ( .A1(n2290), .A2(n4412), .ZN(n2291) );
  INV_X1 U2963 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2292) );
  NAND2_X1 U2964 ( .A1(n2282), .A2(REG1_REG_2__SCAN_IN), .ZN(n2297) );
  INV_X1 U2965 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2849) );
  OR2_X1 U2966 ( .A1(n2010), .A2(n2849), .ZN(n2296) );
  INV_X1 U2967 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2294) );
  OR2_X1 U2968 ( .A1(n2547), .A2(n2294), .ZN(n2295) );
  INV_X1 U2969 ( .A(n2821), .ZN(n2735) );
  INV_X1 U2970 ( .A(n3343), .ZN(n2767) );
  NAND2_X1 U2971 ( .A1(n2735), .A2(n2767), .ZN(n3434) );
  NAND2_X1 U2972 ( .A1(n2821), .A2(n3343), .ZN(n3433) );
  NAND2_X1 U2973 ( .A1(n2821), .A2(n2767), .ZN(n2301) );
  NAND2_X1 U2974 ( .A1(n2282), .A2(REG1_REG_3__SCAN_IN), .ZN(n2307) );
  INV_X1 U2975 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2683) );
  INV_X1 U2976 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2303) );
  OR2_X1 U2977 ( .A1(n2547), .A2(n2303), .ZN(n2304) );
  INV_X1 U2978 ( .A(IR_REG_2__SCAN_IN), .ZN(n2308) );
  NAND2_X1 U2979 ( .A1(n2309), .A2(IR_REG_31__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U2980 ( .A1(n2310), .A2(n3776), .ZN(n2320) );
  OR2_X1 U2981 ( .A1(n2310), .A2(n3776), .ZN(n2311) );
  MUX2_X1 U2982 ( .A(n4250), .B(DATAI_3_), .S(n3397), .Z(n3437) );
  NOR2_X1 U2983 ( .A1(n3557), .A2(n3437), .ZN(n2313) );
  NAND2_X1 U2984 ( .A1(n3557), .A2(n3437), .ZN(n2312) );
  OAI21_X2 U2985 ( .B1(n2817), .B2(n2313), .A(n2312), .ZN(n2854) );
  NAND2_X1 U2986 ( .A1(n3383), .A2(REG0_REG_4__SCAN_IN), .ZN(n2319) );
  INV_X1 U2987 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2314) );
  OR2_X1 U2988 ( .A1(n3392), .A2(n2314), .ZN(n2318) );
  XNOR2_X1 U2989 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n2864) );
  OR2_X1 U2990 ( .A1(n2007), .A2(n2864), .ZN(n2317) );
  INV_X1 U2991 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2315) );
  OR2_X1 U2992 ( .A1(n2009), .A2(n2315), .ZN(n2316) );
  NAND2_X1 U2993 ( .A1(n2320), .A2(IR_REG_31__SCAN_IN), .ZN(n2321) );
  XNOR2_X1 U2994 ( .A(n2321), .B(IR_REG_4__SCAN_IN), .ZN(n4249) );
  MUX2_X1 U2995 ( .A(n4249), .B(DATAI_4_), .S(n3397), .Z(n2856) );
  NAND2_X1 U2996 ( .A1(n2824), .A2(n2856), .ZN(n3440) );
  INV_X1 U2997 ( .A(n2856), .ZN(n2862) );
  NAND2_X1 U2998 ( .A1(n3556), .A2(n2862), .ZN(n3444) );
  NAND2_X1 U2999 ( .A1(n3440), .A2(n3444), .ZN(n3526) );
  NAND2_X1 U3000 ( .A1(n3556), .A2(n2856), .ZN(n2322) );
  AOI21_X1 U3001 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2323) );
  NOR2_X1 U3002 ( .A1(n2323), .A2(n2336), .ZN(n2895) );
  NAND2_X1 U3003 ( .A1(n2272), .A2(n2895), .ZN(n2328) );
  INV_X1 U3004 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2324) );
  OR2_X1 U3005 ( .A1(n2547), .A2(n2324), .ZN(n2327) );
  INV_X1 U3006 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2695) );
  OR2_X1 U3007 ( .A1(n3392), .A2(n2695), .ZN(n2326) );
  OR2_X1 U3008 ( .A1(n2010), .A2(n3572), .ZN(n2325) );
  NAND4_X1 U3009 ( .A1(n2328), .A2(n2327), .A3(n2326), .A4(n2325), .ZN(n2923)
         );
  NAND2_X1 U3010 ( .A1(n2329), .A2(IR_REG_31__SCAN_IN), .ZN(n2330) );
  MUX2_X1 U3011 ( .A(IR_REG_31__SCAN_IN), .B(n2330), .S(IR_REG_5__SCAN_IN), 
        .Z(n2333) );
  AND2_X1 U3012 ( .A1(n2333), .A2(n2332), .ZN(n4248) );
  MUX2_X1 U3013 ( .A(n4248), .B(DATAI_5_), .S(n3397), .Z(n2892) );
  AND2_X1 U3014 ( .A1(n2923), .A2(n2892), .ZN(n2334) );
  NAND2_X1 U3015 ( .A1(n2282), .A2(REG1_REG_6__SCAN_IN), .ZN(n2340) );
  INV_X1 U3016 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2335) );
  OR2_X1 U3017 ( .A1(n2547), .A2(n2335), .ZN(n2339) );
  OAI21_X1 U3018 ( .B1(n2336), .B2(REG3_REG_6__SCAN_IN), .A(n2356), .ZN(n2926)
         );
  OR2_X1 U3019 ( .A1(n2007), .A2(n2926), .ZN(n2338) );
  INV_X1 U3020 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2908) );
  OR2_X1 U3021 ( .A1(n2009), .A2(n2908), .ZN(n2337) );
  NAND4_X1 U3022 ( .A1(n2340), .A2(n2339), .A3(n2338), .A4(n2337), .ZN(n3555)
         );
  NAND2_X1 U3023 ( .A1(n2332), .A2(IR_REG_31__SCAN_IN), .ZN(n2341) );
  XNOR2_X1 U3024 ( .A(n2341), .B(IR_REG_6__SCAN_IN), .ZN(n3594) );
  MUX2_X1 U3025 ( .A(n3594), .B(DATAI_6_), .S(n3397), .Z(n2924) );
  NAND2_X1 U3026 ( .A1(n3555), .A2(n2924), .ZN(n2342) );
  NAND2_X1 U3027 ( .A1(n3393), .A2(REG0_REG_7__SCAN_IN), .ZN(n2347) );
  OR2_X1 U3028 ( .A1(n3392), .A2(n4536), .ZN(n2346) );
  INV_X1 U3029 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2355) );
  XNOR2_X1 U3030 ( .A(n2356), .B(n2355), .ZN(n2958) );
  OR2_X1 U3031 ( .A1(n2007), .A2(n2958), .ZN(n2345) );
  INV_X1 U3032 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2343) );
  OR2_X1 U3033 ( .A1(n2010), .A2(n2343), .ZN(n2344) );
  OAI21_X1 U3034 ( .B1(n2332), .B2(IR_REG_6__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2349) );
  INV_X1 U3035 ( .A(IR_REG_7__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3036 ( .A1(n2349), .A2(n2348), .ZN(n2364) );
  OR2_X1 U3037 ( .A1(n2349), .A2(n2348), .ZN(n2350) );
  MUX2_X1 U3038 ( .A(n3596), .B(DATAI_7_), .S(n3397), .Z(n2957) );
  NAND2_X1 U3039 ( .A1(n2970), .A2(n2957), .ZN(n2576) );
  NAND2_X1 U3040 ( .A1(n3554), .A2(n2951), .ZN(n3449) );
  NAND2_X1 U3041 ( .A1(n2576), .A2(n3449), .ZN(n3527) );
  NAND2_X1 U3042 ( .A1(n2961), .A2(n3527), .ZN(n2352) );
  NAND2_X1 U3043 ( .A1(n3554), .A2(n2957), .ZN(n2351) );
  NAND2_X1 U3044 ( .A1(n2352), .A2(n2351), .ZN(n3029) );
  NAND2_X1 U3045 ( .A1(n3393), .A2(REG0_REG_8__SCAN_IN), .ZN(n2363) );
  INV_X1 U3046 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2353) );
  OR2_X1 U3047 ( .A1(n3392), .A2(n2353), .ZN(n2362) );
  INV_X1 U3048 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2354) );
  OAI21_X1 U3049 ( .B1(n2356), .B2(n2355), .A(n2354), .ZN(n2357) );
  AND2_X1 U3050 ( .A1(n2368), .A2(n2357), .ZN(n4402) );
  INV_X1 U3051 ( .A(n4402), .ZN(n2358) );
  OR2_X1 U3052 ( .A1(n2008), .A2(n2358), .ZN(n2361) );
  INV_X1 U3053 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2359) );
  OR2_X1 U3054 ( .A1(n2010), .A2(n2359), .ZN(n2360) );
  NAND4_X1 U3055 ( .A1(n2363), .A2(n2362), .A3(n2361), .A4(n2360), .ZN(n3553)
         );
  NAND2_X1 U3056 ( .A1(n2364), .A2(IR_REG_31__SCAN_IN), .ZN(n2365) );
  XNOR2_X1 U3057 ( .A(n2365), .B(IR_REG_8__SCAN_IN), .ZN(n4474) );
  MUX2_X1 U3058 ( .A(n4474), .B(DATAI_8_), .S(n3397), .Z(n2641) );
  NAND2_X1 U3059 ( .A1(n2978), .A2(n3031), .ZN(n2366) );
  NAND2_X1 U3060 ( .A1(n3383), .A2(REG0_REG_9__SCAN_IN), .ZN(n2373) );
  INV_X1 U3061 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2367) );
  OR2_X1 U3062 ( .A1(n3392), .A2(n2367), .ZN(n2372) );
  INV_X1 U3063 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2996) );
  NAND2_X1 U3064 ( .A1(n2368), .A2(n2996), .ZN(n2369) );
  NAND2_X1 U3065 ( .A1(n2383), .A2(n2369), .ZN(n2999) );
  OR2_X1 U3066 ( .A1(n2008), .A2(n2999), .ZN(n2371) );
  INV_X1 U3067 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2983) );
  OR2_X1 U3068 ( .A1(n2009), .A2(n2983), .ZN(n2370) );
  NAND4_X1 U3069 ( .A1(n2373), .A2(n2372), .A3(n2371), .A4(n2370), .ZN(n3552)
         );
  INV_X1 U3070 ( .A(IR_REG_8__SCAN_IN), .ZN(n2374) );
  NAND2_X1 U3071 ( .A1(n2375), .A2(n2374), .ZN(n2376) );
  NOR2_X1 U3072 ( .A1(n2332), .A2(n2376), .ZN(n2380) );
  NOR2_X1 U3073 ( .A1(n2380), .A2(n3831), .ZN(n2377) );
  MUX2_X1 U3074 ( .A(n3831), .B(n2377), .S(IR_REG_9__SCAN_IN), .Z(n2378) );
  INV_X1 U3075 ( .A(n2378), .ZN(n2381) );
  NAND2_X1 U3076 ( .A1(n2380), .A2(n2379), .ZN(n2424) );
  MUX2_X1 U3077 ( .A(n4472), .B(DATAI_9_), .S(n3397), .Z(n2995) );
  INV_X1 U3078 ( .A(n2995), .ZN(n2987) );
  NAND2_X1 U3079 ( .A1(n3383), .A2(REG0_REG_10__SCAN_IN), .ZN(n2388) );
  INV_X1 U3080 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4174) );
  OR2_X1 U3081 ( .A1(n3392), .A2(n4174), .ZN(n2387) );
  NAND2_X1 U3082 ( .A1(n2383), .A2(n2382), .ZN(n2384) );
  NAND2_X1 U3083 ( .A1(n2392), .A2(n2384), .ZN(n3194) );
  OR2_X1 U3084 ( .A1(n2008), .A2(n3194), .ZN(n2386) );
  INV_X1 U3085 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3011) );
  OR2_X1 U3086 ( .A1(n2009), .A2(n3011), .ZN(n2385) );
  NAND4_X1 U3087 ( .A1(n2388), .A2(n2387), .A3(n2386), .A4(n2385), .ZN(n3551)
         );
  NAND2_X1 U3088 ( .A1(n2424), .A2(IR_REG_31__SCAN_IN), .ZN(n2389) );
  XNOR2_X1 U3089 ( .A(n2389), .B(IR_REG_10__SCAN_IN), .ZN(n4309) );
  MUX2_X1 U3090 ( .A(n4309), .B(DATAI_10_), .S(n3397), .Z(n3193) );
  AND2_X1 U3091 ( .A1(n3551), .A2(n3193), .ZN(n2391) );
  INV_X1 U3092 ( .A(n3551), .ZN(n3018) );
  INV_X1 U3093 ( .A(n3193), .ZN(n3004) );
  NAND2_X1 U3094 ( .A1(n3018), .A2(n3004), .ZN(n2390) );
  OAI21_X1 U3095 ( .B1(n3008), .B2(n2391), .A(n2390), .ZN(n3021) );
  INV_X1 U3096 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3796) );
  OR2_X1 U3097 ( .A1(n2547), .A2(n3796), .ZN(n2397) );
  INV_X1 U3098 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3808) );
  OR2_X1 U3099 ( .A1(n3392), .A2(n3808), .ZN(n2396) );
  NAND2_X1 U3100 ( .A1(n2392), .A2(n3747), .ZN(n2393) );
  NAND2_X1 U3101 ( .A1(n2403), .A2(n2393), .ZN(n3332) );
  OR2_X1 U3102 ( .A1(n2007), .A2(n3332), .ZN(n2395) );
  INV_X1 U3103 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3024) );
  OR2_X1 U3104 ( .A1(n2010), .A2(n3024), .ZN(n2394) );
  NAND2_X1 U3105 ( .A1(n2398), .A2(IR_REG_31__SCAN_IN), .ZN(n2410) );
  XNOR2_X1 U3106 ( .A(n2410), .B(IR_REG_11__SCAN_IN), .ZN(n4470) );
  MUX2_X1 U3107 ( .A(n4470), .B(DATAI_11_), .S(n3397), .Z(n3331) );
  NAND2_X1 U3108 ( .A1(n3246), .A2(n3331), .ZN(n3465) );
  NAND2_X1 U3109 ( .A1(n4066), .A2(n3064), .ZN(n3458) );
  NAND2_X1 U3110 ( .A1(n3465), .A2(n3458), .ZN(n3528) );
  NAND2_X1 U3111 ( .A1(n3021), .A2(n3528), .ZN(n2400) );
  NAND2_X1 U3112 ( .A1(n3246), .A2(n3064), .ZN(n2399) );
  NAND2_X1 U3113 ( .A1(n2400), .A2(n2399), .ZN(n4072) );
  NAND2_X1 U3114 ( .A1(n3393), .A2(REG0_REG_12__SCAN_IN), .ZN(n2409) );
  INV_X1 U3115 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4166) );
  OR2_X1 U3116 ( .A1(n3392), .A2(n4166), .ZN(n2408) );
  INV_X1 U3117 ( .A(n2401), .ZN(n2415) );
  NAND2_X1 U3118 ( .A1(n2403), .A2(n2402), .ZN(n2404) );
  NAND2_X1 U3119 ( .A1(n2415), .A2(n2404), .ZN(n3245) );
  OR2_X1 U3120 ( .A1(n2008), .A2(n3245), .ZN(n2407) );
  INV_X1 U3121 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2405) );
  OR2_X1 U3122 ( .A1(n2010), .A2(n2405), .ZN(n2406) );
  NAND4_X1 U3123 ( .A1(n2409), .A2(n2408), .A3(n2407), .A4(n2406), .ZN(n4049)
         );
  INV_X1 U3124 ( .A(IR_REG_11__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3125 ( .A1(n2410), .A2(n2422), .ZN(n2411) );
  NAND2_X1 U3126 ( .A1(n2411), .A2(IR_REG_31__SCAN_IN), .ZN(n2412) );
  XNOR2_X1 U3127 ( .A(n2412), .B(IR_REG_12__SCAN_IN), .ZN(n3602) );
  MUX2_X1 U3128 ( .A(n3602), .B(DATAI_12_), .S(n3397), .Z(n4073) );
  NOR2_X1 U3129 ( .A1(n4049), .A2(n4073), .ZN(n2414) );
  NAND2_X1 U3130 ( .A1(n4049), .A2(n4073), .ZN(n2413) );
  NAND2_X1 U3131 ( .A1(n3393), .A2(REG0_REG_13__SCAN_IN), .ZN(n2420) );
  INV_X1 U3132 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3706) );
  OR2_X1 U3133 ( .A1(n3392), .A2(n3706), .ZN(n2419) );
  INV_X1 U3134 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U3135 ( .A1(n2415), .A2(n3312), .ZN(n2416) );
  NAND2_X1 U3136 ( .A1(n2428), .A2(n2416), .ZN(n4056) );
  OR2_X1 U3137 ( .A1(n2008), .A2(n4056), .ZN(n2418) );
  INV_X1 U3138 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4057) );
  OR2_X1 U3139 ( .A1(n2010), .A2(n4057), .ZN(n2417) );
  NAND4_X1 U3140 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(n3550)
         );
  INV_X1 U3141 ( .A(IR_REG_10__SCAN_IN), .ZN(n3828) );
  INV_X1 U3142 ( .A(IR_REG_12__SCAN_IN), .ZN(n2421) );
  NAND3_X1 U3143 ( .A1(n2422), .A2(n3828), .A3(n2421), .ZN(n2423) );
  OAI21_X1 U3144 ( .B1(n2424), .B2(n2423), .A(IR_REG_31__SCAN_IN), .ZN(n2425)
         );
  XNOR2_X1 U3145 ( .A(n2425), .B(IR_REG_13__SCAN_IN), .ZN(n4467) );
  MUX2_X1 U3146 ( .A(n4467), .B(DATAI_13_), .S(n3397), .Z(n4052) );
  NAND2_X1 U3147 ( .A1(n3393), .A2(REG0_REG_14__SCAN_IN), .ZN(n2433) );
  INV_X1 U31480 ( .A(REG1_REG_14__SCAN_IN), .ZN(n2426) );
  OR2_X1 U31490 ( .A1(n3392), .A2(n2426), .ZN(n2432) );
  NAND2_X1 U3150 ( .A1(n2428), .A2(n2427), .ZN(n2429) );
  NAND2_X1 U3151 ( .A1(n2438), .A2(n2429), .ZN(n4036) );
  OR2_X1 U3152 ( .A1(n2007), .A2(n4036), .ZN(n2431) );
  INV_X1 U3153 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4037) );
  OR2_X1 U3154 ( .A1(n2009), .A2(n4037), .ZN(n2430) );
  OR2_X1 U3155 ( .A1(n2434), .A2(n3831), .ZN(n2435) );
  XNOR2_X1 U3156 ( .A(n2435), .B(IR_REG_14__SCAN_IN), .ZN(n3606) );
  MUX2_X1 U3157 ( .A(n3606), .B(DATAI_14_), .S(n3397), .Z(n4035) );
  NAND2_X1 U3158 ( .A1(n4042), .A2(n4035), .ZN(n4006) );
  INV_X1 U3159 ( .A(n4042), .ZN(n3372) );
  NAND2_X1 U3160 ( .A1(n3372), .A2(n3173), .ZN(n3401) );
  NAND2_X1 U3161 ( .A1(n4006), .A2(n3401), .ZN(n4024) );
  NAND2_X1 U3162 ( .A1(n3383), .A2(REG0_REG_15__SCAN_IN), .ZN(n2443) );
  INV_X1 U3163 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4152) );
  OR2_X1 U3164 ( .A1(n3392), .A2(n4152), .ZN(n2442) );
  INV_X1 U3165 ( .A(n2437), .ZN(n2460) );
  NAND2_X1 U3166 ( .A1(n2438), .A2(n3824), .ZN(n2439) );
  NAND2_X1 U3167 ( .A1(n2460), .A2(n2439), .ZN(n4018) );
  OR2_X1 U3168 ( .A1(n2008), .A2(n4018), .ZN(n2441) );
  INV_X1 U3169 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4019) );
  OR2_X1 U3170 ( .A1(n2009), .A2(n4019), .ZN(n2440) );
  NAND4_X1 U3171 ( .A1(n2443), .A2(n2442), .A3(n2441), .A4(n2440), .ZN(n4029)
         );
  INV_X1 U3172 ( .A(IR_REG_14__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3173 ( .A1(n2434), .A2(n2444), .ZN(n2445) );
  NAND2_X1 U3174 ( .A1(n2445), .A2(IR_REG_31__SCAN_IN), .ZN(n2447) );
  INV_X1 U3175 ( .A(IR_REG_15__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3176 ( .A1(n2447), .A2(n2446), .ZN(n2456) );
  OR2_X1 U3177 ( .A1(n2447), .A2(n2446), .ZN(n2448) );
  MUX2_X1 U3178 ( .A(n3591), .B(DATAI_15_), .S(n3397), .Z(n3374) );
  OAI21_X1 U3179 ( .B1(n4012), .B2(n2450), .A(n2449), .ZN(n3990) );
  NAND2_X1 U3180 ( .A1(n3393), .A2(REG0_REG_16__SCAN_IN), .ZN(n2455) );
  INV_X1 U3181 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4147) );
  OR2_X1 U3182 ( .A1(n3392), .A2(n4147), .ZN(n2454) );
  INV_X1 U3183 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2459) );
  XNOR2_X1 U3184 ( .A(n2460), .B(n2459), .ZN(n3265) );
  OR2_X1 U3185 ( .A1(n2008), .A2(n3265), .ZN(n2453) );
  INV_X1 U3186 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2451) );
  OR2_X1 U3187 ( .A1(n2009), .A2(n2451), .ZN(n2452) );
  NAND2_X1 U3188 ( .A1(n2456), .A2(IR_REG_31__SCAN_IN), .ZN(n2457) );
  XNOR2_X1 U3189 ( .A(n2457), .B(IR_REG_16__SCAN_IN), .ZN(n3609) );
  MUX2_X1 U3190 ( .A(n3609), .B(DATAI_16_), .S(n3397), .Z(n2642) );
  NAND2_X1 U3191 ( .A1(n4008), .A2(n2642), .ZN(n3472) );
  NAND2_X1 U3192 ( .A1(n3978), .A2(n3998), .ZN(n3405) );
  NAND2_X1 U3193 ( .A1(n3472), .A2(n3405), .ZN(n2584) );
  NAND2_X1 U3194 ( .A1(n3393), .A2(REG0_REG_17__SCAN_IN), .ZN(n2466) );
  INV_X1 U3195 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4143) );
  OR2_X1 U3196 ( .A1(n3392), .A2(n4143), .ZN(n2465) );
  INV_X1 U3197 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2458) );
  OAI21_X1 U3198 ( .B1(n2460), .B2(n2459), .A(n2458), .ZN(n2462) );
  INV_X1 U3199 ( .A(n2461), .ZN(n2474) );
  NAND2_X1 U3200 ( .A1(n2462), .A2(n2474), .ZN(n3984) );
  OR2_X1 U3201 ( .A1(n2007), .A2(n3984), .ZN(n2464) );
  INV_X1 U3202 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3985) );
  OR2_X1 U3203 ( .A1(n2010), .A2(n3985), .ZN(n2463) );
  NAND2_X1 U3204 ( .A1(n2467), .A2(IR_REG_31__SCAN_IN), .ZN(n2468) );
  XNOR2_X1 U3205 ( .A(n2468), .B(IR_REG_17__SCAN_IN), .ZN(n4459) );
  INV_X1 U3206 ( .A(DATAI_17_), .ZN(n2469) );
  MUX2_X1 U3207 ( .A(n4390), .B(n2469), .S(n3397), .Z(n3975) );
  NAND2_X1 U3208 ( .A1(n3393), .A2(REG0_REG_18__SCAN_IN), .ZN(n2479) );
  INV_X1 U3209 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3611) );
  OR2_X1 U32100 ( .A1(n3392), .A2(n3611), .ZN(n2478) );
  INV_X1 U32110 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U32120 ( .A1(n2474), .A2(n2473), .ZN(n2475) );
  NAND2_X1 U32130 ( .A1(n2481), .A2(n2475), .ZN(n3966) );
  OR2_X1 U32140 ( .A1(n2007), .A2(n3966), .ZN(n2477) );
  INV_X1 U32150 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3967) );
  OR2_X1 U32160 ( .A1(n2010), .A2(n3967), .ZN(n2476) );
  NAND2_X1 U32170 ( .A1(n2047), .A2(IR_REG_31__SCAN_IN), .ZN(n2480) );
  XNOR2_X1 U32180 ( .A(n2480), .B(IR_REG_18__SCAN_IN), .ZN(n3590) );
  MUX2_X1 U32190 ( .A(n3590), .B(DATAI_18_), .S(n3397), .Z(n3957) );
  NAND2_X1 U32200 ( .A1(n3976), .A2(n3957), .ZN(n3935) );
  INV_X1 U32210 ( .A(n3976), .ZN(n3549) );
  NAND2_X1 U32220 ( .A1(n3549), .A2(n3962), .ZN(n3936) );
  NAND2_X1 U32230 ( .A1(n3935), .A2(n3936), .ZN(n3956) );
  NAND2_X1 U32240 ( .A1(n3393), .A2(REG0_REG_19__SCAN_IN), .ZN(n2486) );
  INV_X1 U32250 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4136) );
  OR2_X1 U32260 ( .A1(n3392), .A2(n4136), .ZN(n2485) );
  NAND2_X1 U32270 ( .A1(n2481), .A2(n3202), .ZN(n2482) );
  NAND2_X1 U32280 ( .A1(n2488), .A2(n2482), .ZN(n3948) );
  OR2_X1 U32290 ( .A1(n2008), .A2(n3948), .ZN(n2484) );
  INV_X1 U32300 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3949) );
  OR2_X1 U32310 ( .A1(n2009), .A2(n3949), .ZN(n2483) );
  INV_X1 U32320 ( .A(DATAI_19_), .ZN(n3771) );
  MUX2_X1 U32330 ( .A(n3616), .B(n3771), .S(n3397), .Z(n3947) );
  INV_X1 U32340 ( .A(n3947), .ZN(n3942) );
  NAND2_X1 U32350 ( .A1(n3393), .A2(REG0_REG_20__SCAN_IN), .ZN(n2493) );
  INV_X1 U32360 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4132) );
  OR2_X1 U32370 ( .A1(n3392), .A2(n4132), .ZN(n2492) );
  INV_X1 U32380 ( .A(n2487), .ZN(n2495) );
  NAND2_X1 U32390 ( .A1(n2488), .A2(n3297), .ZN(n2489) );
  NAND2_X1 U32400 ( .A1(n2495), .A2(n2489), .ZN(n3296) );
  OR2_X1 U32410 ( .A1(n2008), .A2(n3296), .ZN(n2491) );
  INV_X1 U32420 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3825) );
  OR2_X1 U32430 ( .A1(n2009), .A2(n3825), .ZN(n2490) );
  NAND2_X1 U32440 ( .A1(n3943), .A2(n3112), .ZN(n3498) );
  NOR2_X1 U32450 ( .A1(n3943), .A2(n3112), .ZN(n3500) );
  NAND2_X1 U32460 ( .A1(n2282), .A2(REG1_REG_21__SCAN_IN), .ZN(n2501) );
  INV_X1 U32470 ( .A(n2494), .ZN(n2510) );
  INV_X1 U32480 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U32490 ( .A1(n2495), .A2(n3238), .ZN(n2496) );
  NAND2_X1 U32500 ( .A1(n2510), .A2(n2496), .ZN(n3237) );
  OR2_X1 U32510 ( .A1(n2008), .A2(n3237), .ZN(n2500) );
  INV_X1 U32520 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2497) );
  OR2_X1 U32530 ( .A1(n2009), .A2(n2497), .ZN(n2499) );
  INV_X1 U32540 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4204) );
  OR2_X1 U32550 ( .A1(n2547), .A2(n4204), .ZN(n2498) );
  INV_X1 U32560 ( .A(n3905), .ZN(n3119) );
  NAND2_X1 U32570 ( .A1(n3919), .A2(n3119), .ZN(n2503) );
  NOR2_X1 U32580 ( .A1(n3919), .A2(n3119), .ZN(n2502) );
  NAND2_X1 U32590 ( .A1(n2512), .A2(n3184), .ZN(n2504) );
  NAND2_X1 U32600 ( .A1(n2519), .A2(n2504), .ZN(n3872) );
  OR2_X1 U32610 ( .A1(n2007), .A2(n3872), .ZN(n2508) );
  NAND2_X1 U32620 ( .A1(n3393), .A2(REG0_REG_23__SCAN_IN), .ZN(n2507) );
  INV_X1 U32630 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4119) );
  OR2_X1 U32640 ( .A1(n3392), .A2(n4119), .ZN(n2506) );
  INV_X1 U32650 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3873) );
  OR2_X1 U32660 ( .A1(n2010), .A2(n3873), .ZN(n2505) );
  NAND4_X1 U32670 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n3885)
         );
  NOR2_X1 U32680 ( .A1(n3885), .A2(n3865), .ZN(n2517) );
  NAND2_X1 U32690 ( .A1(n3393), .A2(REG0_REG_22__SCAN_IN), .ZN(n2516) );
  INV_X1 U32700 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2509) );
  OR2_X1 U32710 ( .A1(n3392), .A2(n2509), .ZN(n2515) );
  INV_X1 U32720 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U32730 ( .A1(n2510), .A2(n3746), .ZN(n2511) );
  NAND2_X1 U32740 ( .A1(n2512), .A2(n2511), .ZN(n3890) );
  OR2_X1 U32750 ( .A1(n2007), .A2(n3890), .ZN(n2514) );
  INV_X1 U32760 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3891) );
  OR2_X1 U32770 ( .A1(n2010), .A2(n3891), .ZN(n2513) );
  NAND2_X1 U32780 ( .A1(n3239), .A2(n3884), .ZN(n3861) );
  NAND2_X1 U32790 ( .A1(n3901), .A2(n3893), .ZN(n2592) );
  NAND2_X1 U32800 ( .A1(n3901), .A2(n3884), .ZN(n3855) );
  INV_X1 U32810 ( .A(n3885), .ZN(n3320) );
  INV_X1 U32820 ( .A(n3865), .ZN(n3870) );
  OAI22_X1 U32830 ( .A1(n2517), .A2(n3855), .B1(n3320), .B2(n3870), .ZN(n2518)
         );
  NAND2_X1 U32840 ( .A1(n2519), .A2(n3284), .ZN(n2520) );
  NAND2_X1 U32850 ( .A1(n2527), .A2(n2520), .ZN(n3283) );
  NAND2_X1 U32860 ( .A1(n3393), .A2(REG0_REG_24__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32870 ( .A1(n2282), .A2(REG1_REG_24__SCAN_IN), .ZN(n2521) );
  INV_X1 U32880 ( .A(n2010), .ZN(n2523) );
  NAND2_X1 U32890 ( .A1(n2523), .A2(REG2_REG_24__SCAN_IN), .ZN(n2524) );
  INV_X1 U32900 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2532) );
  INV_X1 U32910 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U32920 ( .A1(n2527), .A2(n2526), .ZN(n2528) );
  NAND2_X1 U32930 ( .A1(n2529), .A2(n2528), .ZN(n3257) );
  OR2_X1 U32940 ( .A1(n3257), .A2(n2008), .ZN(n2531) );
  AOI22_X1 U32950 ( .A1(n3393), .A2(REG0_REG_25__SCAN_IN), .B1(n2282), .B2(
        REG1_REG_25__SCAN_IN), .ZN(n2530) );
  INV_X1 U32960 ( .A(n3696), .ZN(n3255) );
  INV_X1 U32970 ( .A(n3650), .ZN(n3700) );
  XNOR2_X1 U32980 ( .A(n2545), .B(REG3_REG_27__SCAN_IN), .ZN(n3660) );
  NAND2_X1 U32990 ( .A1(n3660), .A2(n2272), .ZN(n2540) );
  INV_X1 U33000 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U33010 ( .A1(n3383), .A2(REG0_REG_27__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U33020 ( .A1(n2282), .A2(REG1_REG_27__SCAN_IN), .ZN(n2536) );
  OAI211_X1 U33030 ( .C1(n3661), .C2(n2009), .A(n2537), .B(n2536), .ZN(n2538)
         );
  INV_X1 U33040 ( .A(n2538), .ZN(n2539) );
  OR2_X1 U33050 ( .A1(n3548), .A2(n3649), .ZN(n2541) );
  NAND2_X1 U33060 ( .A1(n3656), .A2(n2541), .ZN(n2542) );
  INV_X1 U33070 ( .A(n3548), .ZN(n3677) );
  NAND2_X1 U33080 ( .A1(n2542), .A2(n2243), .ZN(n3622) );
  INV_X1 U33090 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3750) );
  INV_X1 U33100 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2543) );
  OAI21_X1 U33110 ( .B1(n2545), .B2(n3750), .A(n2543), .ZN(n2546) );
  NAND2_X1 U33120 ( .A1(REG3_REG_28__SCAN_IN), .A2(REG3_REG_27__SCAN_IN), .ZN(
        n2544) );
  OR2_X1 U33130 ( .A1(n2545), .A2(n2544), .ZN(n3638) );
  NAND2_X1 U33140 ( .A1(n3223), .A2(n2272), .ZN(n2552) );
  INV_X1 U33150 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3830) );
  INV_X1 U33160 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3783) );
  OR2_X1 U33170 ( .A1(n2547), .A2(n3783), .ZN(n2549) );
  INV_X1 U33180 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3709) );
  OR2_X1 U33190 ( .A1(n3392), .A2(n3709), .ZN(n2548) );
  OAI211_X1 U33200 ( .C1(n2009), .C2(n3830), .A(n2549), .B(n2548), .ZN(n2550)
         );
  INV_X1 U33210 ( .A(n2550), .ZN(n2551) );
  AND2_X1 U33220 ( .A1(n3397), .A2(DATAI_28_), .ZN(n3623) );
  NAND2_X1 U33230 ( .A1(n3652), .A2(n3623), .ZN(n3390) );
  NAND2_X1 U33240 ( .A1(n3624), .A2(n3212), .ZN(n3629) );
  XNOR2_X1 U33250 ( .A(n3622), .B(n3621), .ZN(n3051) );
  NAND2_X1 U33260 ( .A1(n2025), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  MUX2_X1 U33270 ( .A(n2553), .B(IR_REG_31__SCAN_IN), .S(n2250), .Z(n2555) );
  INV_X1 U33280 ( .A(n2554), .ZN(n2561) );
  NAND2_X1 U33290 ( .A1(n2557), .A2(n2556), .ZN(n2558) );
  NAND2_X1 U33300 ( .A1(n2558), .A2(IR_REG_31__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U33310 ( .A1(n2561), .A2(IR_REG_31__SCAN_IN), .ZN(n2562) );
  XNOR2_X1 U33320 ( .A(n2834), .B(n4244), .ZN(n2563) );
  NAND2_X1 U33330 ( .A1(n2563), .A2(n3616), .ZN(n4420) );
  AND2_X1 U33340 ( .A1(n2644), .A2(n4247), .ZN(n4435) );
  INV_X1 U33350 ( .A(n4522), .ZN(n4507) );
  NAND2_X1 U33360 ( .A1(n2564), .A2(n2565), .ZN(n2566) );
  NAND2_X1 U33370 ( .A1(n2566), .A2(IR_REG_31__SCAN_IN), .ZN(n2568) );
  INV_X1 U33380 ( .A(IR_REG_28__SCAN_IN), .ZN(n2567) );
  INV_X1 U33390 ( .A(n2570), .ZN(n4417) );
  NAND2_X1 U33400 ( .A1(n4417), .A2(n2723), .ZN(n3519) );
  OR2_X1 U33410 ( .A1(n2569), .A2(n3519), .ZN(n4409) );
  NAND2_X1 U33420 ( .A1(n4409), .A2(n3432), .ZN(n2572) );
  NAND2_X1 U33430 ( .A1(n2572), .A2(n2571), .ZN(n2846) );
  NAND2_X1 U33440 ( .A1(n2846), .A2(n3433), .ZN(n2573) );
  XNOR2_X1 U33450 ( .A(n3557), .B(n3437), .ZN(n3522) );
  NAND2_X1 U33460 ( .A1(n2573), .A2(n3522), .ZN(n2820) );
  INV_X1 U33470 ( .A(n3557), .ZN(n3436) );
  NAND2_X1 U33480 ( .A1(n3436), .A2(n3437), .ZN(n3439) );
  NAND2_X1 U33490 ( .A1(n2820), .A2(n3439), .ZN(n2855) );
  INV_X1 U33500 ( .A(n3440), .ZN(n2574) );
  INV_X1 U33510 ( .A(n2892), .ZN(n2888) );
  AND2_X1 U33520 ( .A1(n2923), .A2(n2888), .ZN(n2886) );
  INV_X1 U3353 ( .A(n2923), .ZN(n2874) );
  NAND2_X1 U33540 ( .A1(n2874), .A2(n2892), .ZN(n3426) );
  INV_X1 U3355 ( .A(n2924), .ZN(n2902) );
  NAND2_X1 U3356 ( .A1(n3555), .A2(n2902), .ZN(n3442) );
  INV_X1 U3357 ( .A(n3555), .ZN(n2944) );
  NAND2_X1 U3358 ( .A1(n2944), .A2(n2924), .ZN(n3428) );
  NAND2_X1 U3359 ( .A1(n2575), .A2(n3428), .ZN(n2950) );
  INV_X1 U3360 ( .A(n2576), .ZN(n2577) );
  OR2_X1 U3361 ( .A1(n2950), .A2(n2577), .ZN(n2578) );
  NAND2_X1 U3362 ( .A1(n2578), .A2(n3449), .ZN(n3030) );
  NAND2_X1 U3363 ( .A1(n2978), .A2(n2641), .ZN(n3453) );
  NAND2_X1 U3364 ( .A1(n3030), .A2(n3453), .ZN(n2579) );
  NAND2_X1 U3365 ( .A1(n3553), .A2(n3031), .ZN(n3448) );
  AND2_X1 U3366 ( .A1(n3552), .A2(n2987), .ZN(n3460) );
  NAND2_X1 U3367 ( .A1(n3032), .A2(n2995), .ZN(n3452) );
  NAND2_X1 U3368 ( .A1(n3551), .A2(n3004), .ZN(n3457) );
  NAND2_X1 U3369 ( .A1(n3018), .A2(n3193), .ZN(n3463) );
  NAND2_X1 U3370 ( .A1(n2580), .A2(n3463), .ZN(n3016) );
  INV_X1 U3371 ( .A(n4073), .ZN(n4063) );
  NOR2_X1 U3372 ( .A1(n4049), .A2(n4063), .ZN(n3508) );
  NAND2_X1 U3373 ( .A1(n4049), .A2(n4063), .ZN(n4043) );
  INV_X1 U3374 ( .A(n4052), .ZN(n4041) );
  NAND2_X1 U3375 ( .A1(n3550), .A2(n4041), .ZN(n3506) );
  AND2_X1 U3376 ( .A1(n4043), .A2(n3506), .ZN(n3466) );
  INV_X1 U3377 ( .A(n3550), .ZN(n4064) );
  NAND2_X1 U3378 ( .A1(n4064), .A2(n4052), .ZN(n3507) );
  NAND2_X1 U3379 ( .A1(n2581), .A2(n3507), .ZN(n4027) );
  NAND2_X1 U3380 ( .A1(n4027), .A2(n2436), .ZN(n4026) );
  NAND2_X1 U3381 ( .A1(n3266), .A2(n3374), .ZN(n3468) );
  NAND2_X1 U3382 ( .A1(n4029), .A2(n4015), .ZN(n3402) );
  NAND2_X1 U3383 ( .A1(n3468), .A2(n3402), .ZN(n4014) );
  INV_X1 U3384 ( .A(n4006), .ZN(n3400) );
  NOR2_X1 U3385 ( .A1(n4014), .A2(n3400), .ZN(n2582) );
  NAND2_X1 U3386 ( .A1(n4026), .A2(n2582), .ZN(n2583) );
  NAND2_X1 U3387 ( .A1(n2583), .A2(n3402), .ZN(n3992) );
  NAND2_X1 U3388 ( .A1(n3958), .A2(n3947), .ZN(n2585) );
  AND2_X1 U3389 ( .A1(n3936), .A2(n2585), .ZN(n2586) );
  NAND2_X1 U3390 ( .A1(n3352), .A2(n3975), .ZN(n3932) );
  NAND2_X1 U3391 ( .A1(n2586), .A2(n3932), .ZN(n3406) );
  INV_X1 U3392 ( .A(n3112), .ZN(n3924) );
  NAND2_X1 U3393 ( .A1(n3993), .A2(n3981), .ZN(n3933) );
  NAND2_X1 U3394 ( .A1(n3935), .A2(n3933), .ZN(n2587) );
  NAND2_X1 U3395 ( .A1(n2587), .A2(n2586), .ZN(n2589) );
  NAND2_X1 U3396 ( .A1(n3521), .A2(n3942), .ZN(n2588) );
  NAND2_X1 U3397 ( .A1(n2589), .A2(n2588), .ZN(n3914) );
  NOR2_X1 U3398 ( .A1(n3943), .A2(n3924), .ZN(n2590) );
  OR2_X1 U3399 ( .A1(n3914), .A2(n2590), .ZN(n3407) );
  NAND2_X1 U3400 ( .A1(n3407), .A2(n2137), .ZN(n3479) );
  NAND2_X1 U3401 ( .A1(n3919), .A2(n3905), .ZN(n3859) );
  INV_X1 U3402 ( .A(n3480), .ZN(n2593) );
  NOR2_X1 U3403 ( .A1(n3919), .A2(n3905), .ZN(n3857) );
  NAND2_X1 U3404 ( .A1(n3885), .A2(n3870), .ZN(n3504) );
  NAND2_X1 U3405 ( .A1(n3504), .A2(n2592), .ZN(n3486) );
  AOI21_X1 U3406 ( .B1(n3857), .B2(n3861), .A(n3486), .ZN(n3411) );
  OAI21_X1 U3407 ( .B1(n3900), .B2(n2593), .A(n3411), .ZN(n3841) );
  OR2_X1 U3408 ( .A1(n3697), .A2(n3285), .ZN(n3505) );
  NAND2_X1 U3409 ( .A1(n3320), .A2(n3865), .ZN(n3840) );
  NAND2_X1 U3410 ( .A1(n3700), .A2(n3673), .ZN(n3516) );
  NAND2_X1 U3411 ( .A1(n3847), .A2(n3696), .ZN(n3668) );
  NAND2_X1 U3412 ( .A1(n3516), .A2(n3668), .ZN(n3416) );
  INV_X1 U3413 ( .A(n3416), .ZN(n3484) );
  NAND2_X1 U3414 ( .A1(n3674), .A2(n3255), .ZN(n3503) );
  NAND2_X1 U3415 ( .A1(n3697), .A2(n3285), .ZN(n3691) );
  AND2_X1 U3416 ( .A1(n3503), .A2(n3691), .ZN(n3413) );
  OR2_X1 U3417 ( .A1(n3413), .A2(n3416), .ZN(n2594) );
  NAND2_X1 U3418 ( .A1(n3650), .A2(n3678), .ZN(n3515) );
  NAND2_X1 U3419 ( .A1(n3548), .A2(n3659), .ZN(n3488) );
  INV_X1 U3420 ( .A(n3389), .ZN(n2595) );
  XNOR2_X1 U3421 ( .A(n2596), .B(n3621), .ZN(n2598) );
  NAND2_X1 U3422 ( .A1(n4244), .A2(n4247), .ZN(n2597) );
  INV_X1 U3423 ( .A(n2644), .ZN(n4246) );
  NAND2_X1 U3424 ( .A1(n4245), .A2(n4246), .ZN(n3423) );
  NAND2_X1 U3425 ( .A1(n2598), .A2(n4436), .ZN(n2603) );
  AOI22_X1 U3426 ( .A1(n3393), .A2(REG0_REG_29__SCAN_IN), .B1(n2282), .B2(
        REG1_REG_29__SCAN_IN), .ZN(n2600) );
  INV_X1 U3427 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3641) );
  OR2_X1 U3428 ( .A1(n2009), .A2(n3641), .ZN(n2599) );
  OAI211_X1 U3429 ( .C1(n3638), .C2(n2007), .A(n2600), .B(n2599), .ZN(n3547)
         );
  INV_X1 U3430 ( .A(n4245), .ZN(n3496) );
  AOI22_X1 U3431 ( .A1(n3547), .A2(n4414), .B1(n4413), .B2(n3623), .ZN(n2602)
         );
  OAI211_X1 U3432 ( .C1(n3677), .C2(n4416), .A(n2603), .B(n2602), .ZN(n3049)
         );
  INV_X1 U3433 ( .A(n3049), .ZN(n2604) );
  OAI21_X1 U3434 ( .B1(n3051), .B2(n4507), .A(n2604), .ZN(n2647) );
  NAND2_X1 U3435 ( .A1(n2605), .A2(IR_REG_31__SCAN_IN), .ZN(n2616) );
  INV_X1 U3436 ( .A(n2608), .ZN(n2609) );
  NAND2_X1 U3437 ( .A1(n2609), .A2(IR_REG_31__SCAN_IN), .ZN(n2610) );
  MUX2_X1 U3438 ( .A(IR_REG_31__SCAN_IN), .B(n2610), .S(IR_REG_25__SCAN_IN), 
        .Z(n2611) );
  NAND2_X1 U3439 ( .A1(n2607), .A2(n2611), .ZN(n2634) );
  NAND2_X2 U3440 ( .A1(n2615), .A2(n4242), .ZN(n2781) );
  OR2_X1 U3441 ( .A1(n2616), .A2(n2201), .ZN(n2617) );
  NAND2_X1 U3442 ( .A1(n2644), .A2(n3616), .ZN(n2713) );
  AND2_X1 U3443 ( .A1(n2712), .A2(n2713), .ZN(n2779) );
  OR2_X1 U3444 ( .A1(n2721), .A2(n2779), .ZN(n2718) );
  NAND2_X1 U3445 ( .A1(n2620), .A2(n2634), .ZN(n2621) );
  MUX2_X1 U3446 ( .A(n2620), .B(n2621), .S(B_REG_SCAN_IN), .Z(n2622) );
  INV_X1 U3447 ( .A(D_REG_2__SCAN_IN), .ZN(n4453) );
  INV_X1 U3448 ( .A(D_REG_11__SCAN_IN), .ZN(n4449) );
  INV_X1 U3449 ( .A(D_REG_28__SCAN_IN), .ZN(n4447) );
  NAND3_X1 U3450 ( .A1(n4453), .A2(n4449), .A3(n4447), .ZN(n3807) );
  INV_X1 U3451 ( .A(n3807), .ZN(n2626) );
  NOR3_X1 U3452 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .ZN(n2625) );
  NOR4_X1 U3453 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2624) );
  NOR4_X1 U3454 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2623) );
  AND4_X1 U3455 ( .A1(n2626), .A2(n2625), .A3(n2624), .A4(n2623), .ZN(n2632)
         );
  NOR4_X1 U3456 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2630) );
  NOR4_X1 U3457 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2629) );
  NOR4_X1 U34580 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2628) );
  NOR4_X1 U34590 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2627) );
  AND4_X1 U3460 ( .A1(n2630), .A2(n2629), .A3(n2628), .A4(n2627), .ZN(n2631)
         );
  AND2_X1 U3461 ( .A1(n2632), .A2(n2631), .ZN(n2633) );
  INV_X1 U3462 ( .A(n2634), .ZN(n4243) );
  OAI22_X1 U3463 ( .A1(n2655), .A2(D_REG_1__SCAN_IN), .B1(n2006), .B2(n4243), 
        .ZN(n2829) );
  AND2_X1 U3464 ( .A1(n2829), .A2(n2720), .ZN(n2635) );
  INV_X1 U3465 ( .A(n2655), .ZN(n2636) );
  INV_X1 U3466 ( .A(D_REG_0__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U34670 ( .A1(n2636), .A2(n2658), .ZN(n2639) );
  INV_X1 U3468 ( .A(n2006), .ZN(n2637) );
  NAND2_X1 U34690 ( .A1(n2637), .A2(n2620), .ZN(n2638) );
  INV_X1 U3470 ( .A(n2640), .ZN(n2645) );
  INV_X1 U34710 ( .A(n3437), .ZN(n2836) );
  NAND2_X1 U3472 ( .A1(n3022), .A2(n3064), .ZN(n4074) );
  INV_X1 U34730 ( .A(n3640), .ZN(n2643) );
  OAI21_X1 U3474 ( .B1(n3657), .B2(n3212), .A(n2643), .ZN(n3047) );
  NAND2_X1 U34750 ( .A1(n2645), .A2(n2242), .ZN(U3546) );
  INV_X1 U3476 ( .A(n2648), .ZN(n2649) );
  NAND2_X1 U34770 ( .A1(n2649), .A2(n2241), .ZN(U3514) );
  INV_X2 U3478 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U34790 ( .A(DATAI_24_), .ZN(n2650) );
  MUX2_X1 U3480 ( .A(n2650), .B(n2620), .S(STATE_REG_SCAN_IN), .Z(n2651) );
  INV_X1 U34810 ( .A(n2651), .ZN(U3328) );
  INV_X1 U3482 ( .A(DATAI_27_), .ZN(n2654) );
  XNOR2_X1 U34830 ( .A(n2652), .B(IR_REG_27__SCAN_IN), .ZN(n4259) );
  NAND2_X1 U3484 ( .A1(n4259), .A2(STATE_REG_SCAN_IN), .ZN(n2653) );
  OAI21_X1 U34850 ( .B1(STATE_REG_SCAN_IN), .B2(n2654), .A(n2653), .ZN(U3325)
         );
  INV_X1 U3486 ( .A(n2721), .ZN(n2711) );
  INV_X1 U34870 ( .A(n2620), .ZN(n2656) );
  NOR3_X1 U3488 ( .A1(n2006), .A2(n2656), .A3(n4455), .ZN(n2657) );
  AOI21_X1 U34890 ( .B1(n4452), .B2(n2658), .A(n2657), .ZN(U3458) );
  INV_X1 U3490 ( .A(D_REG_1__SCAN_IN), .ZN(n2660) );
  NOR3_X1 U34910 ( .A1(n2006), .A2(n4243), .A3(n4455), .ZN(n2659) );
  AOI21_X1 U3492 ( .B1(n4452), .B2(n2660), .A(n2659), .ZN(U3459) );
  OR2_X1 U34930 ( .A1(n2777), .A2(U3149), .ZN(n3545) );
  NAND2_X1 U3494 ( .A1(n2721), .A2(n3545), .ZN(n2667) );
  NAND2_X1 U34950 ( .A1(n2777), .A2(n2712), .ZN(n2661) );
  AND2_X1 U3496 ( .A1(n3397), .A2(n2661), .ZN(n2666) );
  INV_X1 U34970 ( .A(n2666), .ZN(n2662) );
  NOR2_X1 U3498 ( .A1(n4395), .A2(U4043), .ZN(U3148) );
  INV_X1 U34990 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n3729) );
  NAND2_X1 U3500 ( .A1(n2290), .A2(U4043), .ZN(n2663) );
  OAI21_X1 U35010 ( .B1(U4043), .B2(n3729), .A(n2663), .ZN(U3551) );
  INV_X1 U3502 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U35030 ( .A1(n4029), .A2(U4043), .ZN(n2664) );
  OAI21_X1 U3504 ( .B1(U4043), .B2(n3732), .A(n2664), .ZN(U3565) );
  INV_X1 U35050 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n3730) );
  NAND2_X1 U35060 ( .A1(n2923), .A2(U4043), .ZN(n2665) );
  OAI21_X1 U35070 ( .B1(U4043), .B2(n3730), .A(n2665), .ZN(U3555) );
  INV_X1 U35080 ( .A(n4250), .ZN(n2692) );
  NAND2_X1 U35090 ( .A1(n2667), .A2(n2666), .ZN(n4262) );
  INV_X1 U35100 ( .A(n4259), .ZN(n2741) );
  OR2_X1 U35110 ( .A1(n2739), .A2(n2741), .ZN(n2743) );
  MUX2_X1 U35120 ( .A(REG2_REG_2__SCAN_IN), .B(n2849), .S(n4251), .Z(n2751) );
  NOR2_X1 U35130 ( .A1(n2289), .A2(n2283), .ZN(n3561) );
  NAND2_X1 U35140 ( .A1(n3559), .A2(n2669), .ZN(n2750) );
  NAND2_X1 U35150 ( .A1(n4251), .A2(REG2_REG_2__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U35160 ( .A1(n2749), .A2(n2670), .ZN(n2681) );
  XNOR2_X1 U35170 ( .A(n2681), .B(n4250), .ZN(n2684) );
  XNOR2_X1 U35180 ( .A(n2684), .B(REG2_REG_3__SCAN_IN), .ZN(n2674) );
  INV_X1 U35190 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4532) );
  INV_X1 U35200 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4530) );
  INV_X1 U35210 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4528) );
  AND2_X1 U35220 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n3563) );
  NAND2_X1 U35230 ( .A1(n3564), .A2(n3563), .ZN(n3562) );
  NAND2_X1 U35240 ( .A1(n3562), .A2(n2671), .ZN(n2747) );
  NOR2_X1 U35250 ( .A1(n2672), .A2(n4532), .ZN(n2690) );
  AOI211_X1 U35260 ( .C1(n4532), .C2(n2672), .A(n2690), .B(n4264), .ZN(n2673)
         );
  AOI21_X1 U35270 ( .B1(n4341), .B2(n2674), .A(n2673), .ZN(n2676) );
  INV_X1 U35280 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2838) );
  NOR2_X1 U35290 ( .A1(STATE_REG_SCAN_IN), .A2(n2838), .ZN(n2784) );
  AOI21_X1 U35300 ( .B1(n4395), .B2(ADDR_REG_3__SCAN_IN), .A(n2784), .ZN(n2675) );
  OAI211_X1 U35310 ( .C1(n2692), .C2(n4401), .A(n2676), .B(n2675), .ZN(U3243)
         );
  INV_X1 U35320 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n3742) );
  INV_X1 U35330 ( .A(n3919), .ZN(n2677) );
  NAND2_X1 U35340 ( .A1(n2677), .A2(U4043), .ZN(n2678) );
  OAI21_X1 U35350 ( .B1(U4043), .B2(n3742), .A(n2678), .ZN(U3571) );
  INV_X1 U35360 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n3805) );
  NAND2_X1 U35370 ( .A1(n3352), .A2(U4043), .ZN(n2679) );
  OAI21_X1 U35380 ( .B1(U4043), .B2(n3805), .A(n2679), .ZN(U3567) );
  INV_X1 U35390 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U35400 ( .A1(n3901), .A2(U4043), .ZN(n2680) );
  OAI21_X1 U35410 ( .B1(U4043), .B2(n3741), .A(n2680), .ZN(U3572) );
  INV_X1 U35420 ( .A(n4248), .ZN(n3571) );
  NAND2_X1 U35430 ( .A1(n2681), .A2(n4250), .ZN(n2682) );
  INV_X1 U35440 ( .A(n4249), .ZN(n2799) );
  AND2_X1 U35450 ( .A1(n2685), .A2(n4249), .ZN(n2686) );
  AOI21_X1 U35460 ( .B1(n2791), .B2(REG2_REG_4__SCAN_IN), .A(n2686), .ZN(n2688) );
  INV_X1 U35470 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3572) );
  MUX2_X1 U35480 ( .A(n3572), .B(REG2_REG_5__SCAN_IN), .S(n4248), .Z(n2687) );
  AOI211_X1 U35490 ( .C1(n2688), .C2(n2687), .A(n3570), .B(n4391), .ZN(n2689)
         );
  INV_X1 U35500 ( .A(n2689), .ZN(n2700) );
  AND2_X1 U35510 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2879) );
  INV_X1 U35520 ( .A(n2690), .ZN(n2691) );
  OAI21_X1 U35530 ( .B1(n2693), .B2(n2692), .A(n2691), .ZN(n2694) );
  XNOR2_X1 U35540 ( .A(n2694), .B(n2799), .ZN(n2790) );
  MUX2_X1 U35550 ( .A(n2695), .B(REG1_REG_5__SCAN_IN), .S(n4248), .Z(n2696) );
  AOI211_X1 U35560 ( .C1(n2697), .C2(n2696), .A(n3592), .B(n4264), .ZN(n2698)
         );
  AOI211_X1 U35570 ( .C1(n4395), .C2(ADDR_REG_5__SCAN_IN), .A(n2879), .B(n2698), .ZN(n2699) );
  OAI211_X1 U35580 ( .C1(n4401), .C2(n3571), .A(n2700), .B(n2699), .ZN(U3245)
         );
  INV_X1 U35590 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n3733) );
  NAND2_X1 U35600 ( .A1(n3372), .A2(U4043), .ZN(n2701) );
  OAI21_X1 U35610 ( .B1(U4043), .B2(n3733), .A(n2701), .ZN(U3564) );
  INV_X1 U35620 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n3735) );
  NAND2_X1 U35630 ( .A1(n3958), .A2(U4043), .ZN(n2702) );
  OAI21_X1 U35640 ( .B1(U4043), .B2(n3735), .A(n2702), .ZN(U3569) );
  INV_X1 U35650 ( .A(n2781), .ZN(n2703) );
  NAND2_X1 U35660 ( .A1(n2703), .A2(IR_REG_0__SCAN_IN), .ZN(n2704) );
  NOR2_X1 U35670 ( .A1(n2781), .A2(n4526), .ZN(n2707) );
  NOR2_X1 U35680 ( .A1(n4434), .A2(n3209), .ZN(n2731) );
  XNOR2_X1 U35690 ( .A(n2732), .B(n2733), .ZN(n2742) );
  NOR2_X1 U35700 ( .A1(n2829), .A2(n2708), .ZN(n2710) );
  NAND2_X1 U35710 ( .A1(n2710), .A2(n2709), .ZN(n2717) );
  INV_X1 U35720 ( .A(n2717), .ZN(n2716) );
  AND2_X1 U35730 ( .A1(n2716), .A2(n2711), .ZN(n2722) );
  AOI21_X1 U35740 ( .B1(n4432), .B2(n2713), .A(n2712), .ZN(n2714) );
  NAND2_X1 U35750 ( .A1(n4244), .A2(n3616), .ZN(n2727) );
  OR2_X1 U35760 ( .A1(n4455), .A2(n2727), .ZN(n2715) );
  NOR2_X1 U35770 ( .A1(n2729), .A2(n2715), .ZN(n3542) );
  NAND2_X1 U35780 ( .A1(n2717), .A2(n2720), .ZN(n2783) );
  INV_X1 U35790 ( .A(n2718), .ZN(n2719) );
  NAND2_X1 U35800 ( .A1(n2783), .A2(n2719), .ZN(n3342) );
  AOI22_X1 U35810 ( .A1(n3378), .A2(n2290), .B1(REG3_REG_0__SCAN_IN), .B2(
        n3342), .ZN(n2725) );
  AOI21_X2 U3582 ( .B1(n2722), .B2(n4413), .A(n4442), .ZN(n3362) );
  NAND2_X1 U3583 ( .A1(n3375), .A2(n2723), .ZN(n2724) );
  OAI211_X1 U3584 ( .C1(n2742), .C2(n3381), .A(n2725), .B(n2724), .ZN(U3229)
         );
  OAI22_X1 U3585 ( .A1(n4440), .A2(n2758), .B1(n2729), .B2(n4426), .ZN(n2762)
         );
  XNOR2_X1 U3586 ( .A(n2763), .B(n2730), .ZN(n2766) );
  OAI22_X1 U3587 ( .A1(n2733), .A2(n2732), .B1(n2731), .B2(n3210), .ZN(n2765)
         );
  XNOR2_X1 U3588 ( .A(n2766), .B(n2765), .ZN(n2738) );
  AOI22_X1 U3589 ( .A1(n3373), .A2(n2570), .B1(REG3_REG_1__SCAN_IN), .B2(n3342), .ZN(n2737) );
  AOI22_X1 U3590 ( .A1(n3375), .A2(n4412), .B1(n3378), .B2(n2735), .ZN(n2736)
         );
  OAI211_X1 U3591 ( .C1(n2738), .C2(n3381), .A(n2737), .B(n2736), .ZN(U3219)
         );
  AND2_X1 U3592 ( .A1(n4259), .A2(n2283), .ZN(n2740) );
  NOR2_X1 U3593 ( .A1(n2740), .A2(n2739), .ZN(n4258) );
  NAND3_X1 U3594 ( .A1(n2742), .A2(n4241), .A3(n2741), .ZN(n2745) );
  INV_X1 U3595 ( .A(n2743), .ZN(n3541) );
  AOI21_X1 U3596 ( .B1(n3541), .B2(n3561), .A(n3558), .ZN(n2744) );
  OAI211_X1 U3597 ( .C1(IR_REG_0__SCAN_IN), .C2(n4258), .A(n2745), .B(n2744), 
        .ZN(n2793) );
  INV_X1 U3598 ( .A(n2793), .ZN(n2757) );
  OAI211_X1 U3599 ( .C1(n2748), .C2(n2747), .A(n4397), .B(n2746), .ZN(n2755)
         );
  OAI211_X1 U3600 ( .C1(n2751), .C2(n2750), .A(n4341), .B(n2749), .ZN(n2754)
         );
  AOI22_X1 U3601 ( .A1(n4395), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2753) );
  INV_X1 U3602 ( .A(n4401), .ZN(n3565) );
  NAND2_X1 U3603 ( .A1(n3565), .A2(n4251), .ZN(n2752) );
  NAND4_X1 U3604 ( .A1(n2755), .A2(n2754), .A3(n2753), .A4(n2752), .ZN(n2756)
         );
  OR2_X1 U3605 ( .A1(n2757), .A2(n2756), .ZN(U3242) );
  OAI22_X1 U3606 ( .A1(n3436), .A2(n2758), .B1(n2729), .B2(n2836), .ZN(n2801)
         );
  NAND2_X1 U3607 ( .A1(n3557), .A2(n3154), .ZN(n2760) );
  NAND2_X1 U3608 ( .A1(n3437), .A2(n2110), .ZN(n2759) );
  NAND2_X1 U3609 ( .A1(n2760), .A2(n2759), .ZN(n2761) );
  XNOR2_X1 U3610 ( .A(n2761), .B(n3210), .ZN(n2800) );
  XOR2_X1 U3611 ( .A(n2801), .B(n2800), .Z(n2776) );
  OAI22_X1 U3612 ( .A1(n2821), .A2(n2729), .B1(n3209), .B2(n2767), .ZN(n2768)
         );
  XNOR2_X1 U3613 ( .A(n2768), .B(n3210), .ZN(n2772) );
  OR2_X1 U3614 ( .A1(n2821), .A2(n2758), .ZN(n2770) );
  NAND2_X1 U3615 ( .A1(n3343), .A2(n3154), .ZN(n2769) );
  NAND2_X1 U3616 ( .A1(n2770), .A2(n2769), .ZN(n2771) );
  NAND2_X1 U3617 ( .A1(n3339), .A2(n3338), .ZN(n3337) );
  NAND2_X1 U3618 ( .A1(n3337), .A2(n2774), .ZN(n2775) );
  NAND2_X1 U3619 ( .A1(n2775), .A2(n2776), .ZN(n2810) );
  OAI21_X1 U3620 ( .B1(n2776), .B2(n2775), .A(n2810), .ZN(n2788) );
  INV_X1 U3621 ( .A(n2777), .ZN(n2778) );
  NOR2_X1 U3622 ( .A1(n2779), .A2(n2778), .ZN(n2780) );
  AND2_X1 U3623 ( .A1(n2781), .A2(n2780), .ZN(n2782) );
  AOI22_X1 U3624 ( .A1(n3375), .A2(n3437), .B1(n3373), .B2(n2735), .ZN(n2786)
         );
  AOI21_X1 U3625 ( .B1(n3378), .B2(n3556), .A(n2784), .ZN(n2785) );
  OAI211_X1 U3626 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3376), .A(n2786), .B(n2785), 
        .ZN(n2787) );
  AOI21_X1 U3627 ( .B1(n2788), .B2(n3340), .A(n2787), .ZN(n2789) );
  INV_X1 U3628 ( .A(n2789), .ZN(U3215) );
  AND2_X1 U3629 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n2812) );
  OAI21_X1 U3630 ( .B1(REG1_REG_4__SCAN_IN), .B2(n2790), .A(n4397), .ZN(n2795)
         );
  XOR2_X1 U3631 ( .A(REG2_REG_4__SCAN_IN), .B(n2791), .Z(n2792) );
  NAND2_X1 U3632 ( .A1(n4341), .A2(n2792), .ZN(n2794) );
  OAI211_X1 U3633 ( .C1(n2796), .C2(n2795), .A(n2794), .B(n2793), .ZN(n2797)
         );
  AOI211_X1 U3634 ( .C1(n4395), .C2(ADDR_REG_4__SCAN_IN), .A(n2812), .B(n2797), 
        .ZN(n2798) );
  OAI21_X1 U3635 ( .B1(n2799), .B2(n4401), .A(n2798), .ZN(U3244) );
  INV_X1 U3636 ( .A(n2800), .ZN(n2803) );
  INV_X1 U3637 ( .A(n2801), .ZN(n2802) );
  NAND2_X1 U3638 ( .A1(n2803), .A2(n2802), .ZN(n2809) );
  OAI22_X1 U3639 ( .A1(n2824), .A2(n2729), .B1(n3209), .B2(n2862), .ZN(n2804)
         );
  XNOR2_X1 U3640 ( .A(n2804), .B(n3152), .ZN(n2869) );
  OR2_X1 U3641 ( .A1(n2824), .A2(n2758), .ZN(n2806) );
  NAND2_X1 U3642 ( .A1(n2856), .A2(n3154), .ZN(n2805) );
  NAND2_X1 U3643 ( .A1(n2806), .A2(n2805), .ZN(n2870) );
  XNOR2_X1 U3644 ( .A(n2869), .B(n2870), .ZN(n2808) );
  NAND2_X1 U3645 ( .A1(n2873), .A2(n3340), .ZN(n2816) );
  AOI21_X1 U3646 ( .B1(n2810), .B2(n2809), .A(n2808), .ZN(n2815) );
  AOI22_X1 U3647 ( .A1(n3375), .A2(n2856), .B1(n3373), .B2(n3557), .ZN(n2814)
         );
  NOR2_X1 U3648 ( .A1(n3376), .A2(n2864), .ZN(n2811) );
  AOI211_X1 U3649 ( .C1(n3378), .C2(n2923), .A(n2812), .B(n2811), .ZN(n2813)
         );
  OAI211_X1 U3650 ( .C1(n2816), .C2(n2815), .A(n2814), .B(n2813), .ZN(U3227)
         );
  INV_X1 U3651 ( .A(n3522), .ZN(n2818) );
  XNOR2_X1 U3652 ( .A(n2817), .B(n2818), .ZN(n4498) );
  NAND2_X1 U3653 ( .A1(n4498), .A2(n4437), .ZN(n2828) );
  NAND3_X1 U3654 ( .A1(n2846), .A2(n3433), .A3(n2818), .ZN(n2819) );
  NAND2_X1 U3655 ( .A1(n2820), .A2(n2819), .ZN(n2826) );
  OR2_X1 U3656 ( .A1(n2821), .A2(n4416), .ZN(n2823) );
  NAND2_X1 U3657 ( .A1(n3437), .A2(n4413), .ZN(n2822) );
  OAI211_X1 U3658 ( .C1(n2824), .C2(n4439), .A(n2823), .B(n2822), .ZN(n2825)
         );
  AOI21_X1 U3659 ( .B1(n2826), .B2(n4436), .A(n2825), .ZN(n2827) );
  AND2_X1 U3660 ( .A1(n2828), .A2(n2827), .ZN(n4500) );
  INV_X1 U3661 ( .A(n2829), .ZN(n2830) );
  NAND3_X1 U3662 ( .A1(n2832), .A2(n2831), .A3(n2830), .ZN(n2833) );
  NOR2_X1 U3663 ( .A1(n2834), .A2(n3616), .ZN(n2835) );
  NAND2_X1 U3664 ( .A1(n4445), .A2(n2835), .ZN(n2884) );
  INV_X1 U3665 ( .A(n2884), .ZN(n4443) );
  INV_X2 U3666 ( .A(n4445), .ZN(n4424) );
  NAND2_X1 U3667 ( .A1(n4058), .A2(n3616), .ZN(n3965) );
  OR2_X1 U3668 ( .A1(n4491), .A2(n2836), .ZN(n2837) );
  NAND2_X1 U3669 ( .A1(n2861), .A2(n2837), .ZN(n4496) );
  AOI22_X1 U3670 ( .A1(n4424), .A2(REG2_REG_3__SCAN_IN), .B1(n4442), .B2(n2838), .ZN(n2839) );
  OAI21_X1 U3671 ( .B1(n4079), .B2(n4496), .A(n2839), .ZN(n2840) );
  AOI21_X1 U3672 ( .B1(n4498), .B2(n4443), .A(n2840), .ZN(n2841) );
  OAI21_X1 U3673 ( .B1(n4500), .B2(n4424), .A(n2841), .ZN(U3287) );
  OAI21_X1 U3674 ( .B1(n2843), .B2(n3520), .A(n2842), .ZN(n4495) );
  INV_X1 U3675 ( .A(n4495), .ZN(n2853) );
  AOI22_X1 U3676 ( .A1(n3557), .A2(n4414), .B1(n3343), .B2(n4413), .ZN(n2844)
         );
  OAI21_X1 U3677 ( .B1(n4440), .B2(n4416), .A(n2844), .ZN(n2848) );
  NAND3_X1 U3678 ( .A1(n3520), .A2(n3432), .A3(n4409), .ZN(n2845) );
  AOI21_X1 U3679 ( .B1(n2846), .B2(n2845), .A(n4069), .ZN(n2847) );
  AOI211_X1 U3680 ( .C1(n4437), .C2(n4495), .A(n2848), .B(n2847), .ZN(n4492)
         );
  MUX2_X1 U3681 ( .A(n2849), .B(n4492), .S(n4445), .Z(n2852) );
  AND2_X1 U3682 ( .A1(n4425), .A2(n3343), .ZN(n4490) );
  NOR3_X1 U3683 ( .A1(n4079), .A2(n4491), .A3(n4490), .ZN(n2850) );
  AOI21_X1 U3684 ( .B1(n4442), .B2(REG3_REG_2__SCAN_IN), .A(n2850), .ZN(n2851)
         );
  OAI211_X1 U3685 ( .C1(n2853), .C2(n2884), .A(n2852), .B(n2851), .ZN(U3288)
         );
  XNOR2_X1 U3686 ( .A(n2854), .B(n3526), .ZN(n2866) );
  XOR2_X1 U3687 ( .A(n3526), .B(n2855), .Z(n2859) );
  AOI22_X1 U3688 ( .A1(n2923), .A2(n4414), .B1(n2856), .B2(n4413), .ZN(n2857)
         );
  OAI21_X1 U3689 ( .B1(n3436), .B2(n4416), .A(n2857), .ZN(n2858) );
  AOI21_X1 U3690 ( .B1(n2859), .B2(n4436), .A(n2858), .ZN(n2860) );
  OAI21_X1 U3691 ( .B1(n4420), .B2(n2866), .A(n2860), .ZN(n4502) );
  INV_X1 U3692 ( .A(n2861), .ZN(n2863) );
  OAI211_X1 U3693 ( .C1(n2863), .C2(n2862), .A(n4512), .B(n2893), .ZN(n4501)
         );
  OAI22_X1 U3694 ( .A1(n4501), .A2(n4247), .B1(n4055), .B2(n2864), .ZN(n2865)
         );
  OAI21_X1 U3695 ( .B1(n4502), .B2(n2865), .A(n4058), .ZN(n2868) );
  INV_X1 U3696 ( .A(n2866), .ZN(n4505) );
  AOI22_X1 U3697 ( .A1(n4505), .A2(n4443), .B1(REG2_REG_4__SCAN_IN), .B2(n4424), .ZN(n2867) );
  NAND2_X1 U3698 ( .A1(n2868), .A2(n2867), .ZN(U3286) );
  INV_X1 U3699 ( .A(n2869), .ZN(n2871) );
  NAND2_X1 U3700 ( .A1(n2871), .A2(n2870), .ZN(n2872) );
  OAI22_X1 U3701 ( .A1(n2874), .A2(n2758), .B1(n2729), .B2(n2888), .ZN(n2914)
         );
  NAND2_X1 U3702 ( .A1(n2923), .A2(n3154), .ZN(n2876) );
  NAND2_X1 U3703 ( .A1(n2892), .A2(n2110), .ZN(n2875) );
  NAND2_X1 U3704 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  XOR2_X1 U3705 ( .A(n2914), .B(n2913), .Z(n2915) );
  XNOR2_X1 U3706 ( .A(n2916), .B(n2915), .ZN(n2882) );
  AOI22_X1 U3707 ( .A1(n3375), .A2(n2892), .B1(n3373), .B2(n3556), .ZN(n2881)
         );
  NOR2_X1 U3708 ( .A1(n3363), .A2(n2944), .ZN(n2878) );
  AOI211_X1 U3709 ( .C1(n2895), .C2(n3366), .A(n2879), .B(n2878), .ZN(n2880)
         );
  OAI211_X1 U3710 ( .C1(n2882), .C2(n3381), .A(n2881), .B(n2880), .ZN(U3224)
         );
  NAND2_X1 U3711 ( .A1(n4058), .A2(n4437), .ZN(n2883) );
  INV_X1 U3712 ( .A(n2886), .ZN(n3443) );
  NAND2_X1 U3713 ( .A1(n3443), .A2(n3426), .ZN(n3529) );
  XNOR2_X1 U3714 ( .A(n2885), .B(n3529), .ZN(n4508) );
  XOR2_X1 U3715 ( .A(n3529), .B(n2887), .Z(n2891) );
  OAI22_X1 U3716 ( .A1(n2944), .A2(n4439), .B1(n4087), .B2(n2888), .ZN(n2889)
         );
  AOI21_X1 U3717 ( .B1(n4067), .B2(n3556), .A(n2889), .ZN(n2890) );
  OAI21_X1 U3718 ( .B1(n2891), .B2(n4069), .A(n2890), .ZN(n4509) );
  NAND2_X1 U3719 ( .A1(n4509), .A2(n4058), .ZN(n2899) );
  AND2_X1 U3720 ( .A1(n2893), .A2(n2892), .ZN(n2894) );
  NOR2_X1 U3721 ( .A1(n2906), .A2(n2894), .ZN(n4511) );
  INV_X1 U3722 ( .A(n2895), .ZN(n2896) );
  OAI22_X1 U3723 ( .A1(n4445), .A2(n3572), .B1(n2896), .B2(n4055), .ZN(n2897)
         );
  AOI21_X1 U3724 ( .B1(n4511), .B2(n4428), .A(n2897), .ZN(n2898) );
  OAI211_X1 U3725 ( .C1(n4004), .C2(n4508), .A(n2899), .B(n2898), .ZN(U3285)
         );
  NAND2_X1 U3726 ( .A1(n3428), .A2(n3442), .ZN(n3525) );
  XNOR2_X1 U3727 ( .A(n2900), .B(n3525), .ZN(n2932) );
  INV_X1 U3728 ( .A(n2932), .ZN(n2912) );
  XNOR2_X1 U3729 ( .A(n2901), .B(n3525), .ZN(n2905) );
  OAI22_X1 U3730 ( .A1(n2970), .A2(n4439), .B1(n4087), .B2(n2902), .ZN(n2903)
         );
  AOI21_X1 U3731 ( .B1(n4067), .B2(n2923), .A(n2903), .ZN(n2904) );
  OAI21_X1 U3732 ( .B1(n2905), .B2(n4069), .A(n2904), .ZN(n2931) );
  NAND2_X1 U3733 ( .A1(n2931), .A2(n4058), .ZN(n2911) );
  INV_X1 U3734 ( .A(n2906), .ZN(n2907) );
  AOI21_X1 U3735 ( .B1(n2924), .B2(n2907), .A(n2955), .ZN(n2934) );
  OAI22_X1 U3736 ( .A1(n4445), .A2(n2908), .B1(n2926), .B2(n4055), .ZN(n2909)
         );
  AOI21_X1 U3737 ( .B1(n2934), .B2(n4428), .A(n2909), .ZN(n2910) );
  OAI211_X1 U3738 ( .C1(n4004), .C2(n2912), .A(n2911), .B(n2910), .ZN(U3284)
         );
  NAND2_X1 U3739 ( .A1(n3555), .A2(n3154), .ZN(n2918) );
  NAND2_X1 U3740 ( .A1(n2924), .A2(n2110), .ZN(n2917) );
  NAND2_X1 U3741 ( .A1(n2918), .A2(n2917), .ZN(n2919) );
  XNOR2_X1 U3742 ( .A(n2919), .B(n3152), .ZN(n2921) );
  AOI22_X1 U3743 ( .A1(n3555), .A2(n3164), .B1(n3154), .B2(n2924), .ZN(n2920)
         );
  OR2_X1 U3744 ( .A1(n2921), .A2(n2920), .ZN(n2937) );
  NAND2_X1 U3745 ( .A1(n2049), .A2(n2937), .ZN(n2922) );
  XNOR2_X1 U3746 ( .A(n2938), .B(n2922), .ZN(n2930) );
  AOI22_X1 U3747 ( .A1(n3375), .A2(n2924), .B1(n3373), .B2(n2923), .ZN(n2929)
         );
  INV_X1 U3748 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2925) );
  NOR2_X1 U3749 ( .A1(STATE_REG_SCAN_IN), .A2(n2925), .ZN(n4268) );
  NOR2_X1 U3750 ( .A1(n3376), .A2(n2926), .ZN(n2927) );
  AOI211_X1 U3751 ( .C1(n3378), .C2(n3554), .A(n4268), .B(n2927), .ZN(n2928)
         );
  OAI211_X1 U3752 ( .C1(n2930), .C2(n3381), .A(n2929), .B(n2928), .ZN(U3236)
         );
  AOI21_X1 U3753 ( .B1(n4522), .B2(n2932), .A(n2931), .ZN(n2936) );
  INV_X1 U3754 ( .A(n4525), .ZN(n4523) );
  INV_X1 U3755 ( .A(n4238), .ZN(n4177) );
  AOI22_X1 U3756 ( .A1(n2934), .A2(n4177), .B1(n4523), .B2(REG0_REG_6__SCAN_IN), .ZN(n2933) );
  OAI21_X1 U3757 ( .B1(n2936), .B2(n4523), .A(n2933), .ZN(U3479) );
  INV_X1 U3758 ( .A(n4176), .ZN(n4084) );
  AOI22_X1 U3759 ( .A1(n2934), .A2(n4084), .B1(n4538), .B2(REG1_REG_6__SCAN_IN), .ZN(n2935) );
  OAI21_X1 U3760 ( .B1(n2936), .B2(n4538), .A(n2935), .ZN(U3524) );
  OR2_X1 U3761 ( .A1(n2970), .A2(n2758), .ZN(n2940) );
  NAND2_X1 U3762 ( .A1(n2957), .A2(n3154), .ZN(n2939) );
  NAND2_X1 U3763 ( .A1(n2940), .A2(n2939), .ZN(n2965) );
  OAI22_X1 U3764 ( .A1(n2970), .A2(n2729), .B1(n3209), .B2(n2951), .ZN(n2941)
         );
  XNOR2_X1 U3765 ( .A(n2941), .B(n3210), .ZN(n2966) );
  XOR2_X1 U3766 ( .A(n2965), .B(n2966), .Z(n2942) );
  OAI211_X1 U3767 ( .C1(n2943), .C2(n2942), .A(n2967), .B(n3340), .ZN(n2949)
         );
  INV_X1 U3768 ( .A(n2958), .ZN(n2947) );
  NAND2_X1 U3769 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n4279) );
  OAI21_X1 U3770 ( .B1(n3363), .B2(n2978), .A(n4279), .ZN(n2946) );
  OAI22_X1 U3771 ( .A1(n3362), .A2(n2951), .B1(n2944), .B2(n3361), .ZN(n2945)
         );
  AOI211_X1 U3772 ( .C1(n2947), .C2(n3366), .A(n2946), .B(n2945), .ZN(n2948)
         );
  NAND2_X1 U3773 ( .A1(n2949), .A2(n2948), .ZN(U3210) );
  XNOR2_X1 U3774 ( .A(n2950), .B(n3527), .ZN(n2954) );
  OAI22_X1 U3775 ( .A1(n2978), .A2(n4439), .B1(n4087), .B2(n2951), .ZN(n2952)
         );
  AOI21_X1 U3776 ( .B1(n4067), .B2(n3555), .A(n2952), .ZN(n2953) );
  OAI21_X1 U3777 ( .B1(n2954), .B2(n4069), .A(n2953), .ZN(n4513) );
  INV_X1 U3778 ( .A(n4513), .ZN(n2964) );
  INV_X1 U3779 ( .A(n2955), .ZN(n2956) );
  AOI211_X1 U3780 ( .C1(n2957), .C2(n2956), .A(n4519), .B(n2048), .ZN(n4514)
         );
  INV_X1 U3781 ( .A(n3965), .ZN(n2960) );
  OAI22_X1 U3782 ( .A1(n4445), .A2(n2343), .B1(n2958), .B2(n4055), .ZN(n2959)
         );
  AOI21_X1 U3783 ( .B1(n4514), .B2(n2960), .A(n2959), .ZN(n2963) );
  XOR2_X1 U3784 ( .A(n2961), .B(n3527), .Z(n4515) );
  NAND2_X1 U3785 ( .A1(n4515), .A2(n4081), .ZN(n2962) );
  OAI211_X1 U3786 ( .C1(n2964), .C2(n4424), .A(n2963), .B(n2962), .ZN(U3283)
         );
  OAI22_X1 U3787 ( .A1(n2978), .A2(n2758), .B1(n2729), .B2(n3031), .ZN(n2990)
         );
  OAI22_X1 U3788 ( .A1(n2978), .A2(n2729), .B1(n3209), .B2(n3031), .ZN(n2968)
         );
  XNOR2_X1 U3789 ( .A(n2968), .B(n3210), .ZN(n2989) );
  XOR2_X1 U3790 ( .A(n2990), .B(n2989), .Z(n2969) );
  XNOR2_X1 U3791 ( .A(n2991), .B(n2969), .ZN(n2974) );
  NAND2_X1 U3792 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4289) );
  OAI21_X1 U3793 ( .B1(n3363), .B2(n3032), .A(n4289), .ZN(n2972) );
  OAI22_X1 U3794 ( .A1(n3362), .A2(n3031), .B1(n2970), .B2(n3361), .ZN(n2971)
         );
  AOI211_X1 U3795 ( .C1(n4402), .C2(n3366), .A(n2972), .B(n2971), .ZN(n2973)
         );
  OAI21_X1 U3796 ( .B1(n2974), .B2(n3381), .A(n2973), .ZN(U3218) );
  INV_X1 U3797 ( .A(n3460), .ZN(n2975) );
  NAND2_X1 U3798 ( .A1(n2975), .A2(n3452), .ZN(n3530) );
  XNOR2_X1 U3799 ( .A(n2976), .B(n3530), .ZN(n2980) );
  AOI22_X1 U3800 ( .A1(n3551), .A2(n4414), .B1(n4413), .B2(n2995), .ZN(n2977)
         );
  OAI21_X1 U3801 ( .B1(n2978), .B2(n4416), .A(n2977), .ZN(n2979) );
  AOI21_X1 U3802 ( .B1(n2980), .B2(n4436), .A(n2979), .ZN(n4517) );
  XNOR2_X1 U3803 ( .A(n2981), .B(n3530), .ZN(n4521) );
  INV_X1 U3804 ( .A(n3028), .ZN(n2982) );
  OAI21_X1 U3805 ( .B1(n2982), .B2(n2987), .A(n3009), .ZN(n4518) );
  NOR2_X1 U3806 ( .A1(n4518), .A2(n4079), .ZN(n2985) );
  OAI22_X1 U3807 ( .A1(n4058), .A2(n2983), .B1(n2999), .B2(n4055), .ZN(n2984)
         );
  AOI211_X1 U3808 ( .C1(n4521), .C2(n4081), .A(n2985), .B(n2984), .ZN(n2986)
         );
  OAI21_X1 U3809 ( .B1(n4424), .B2(n4517), .A(n2986), .ZN(U3281) );
  OAI22_X1 U3810 ( .A1(n3032), .A2(n2758), .B1(n2729), .B2(n2987), .ZN(n3057)
         );
  OAI22_X1 U3811 ( .A1(n3032), .A2(n2729), .B1(n3209), .B2(n2987), .ZN(n2988)
         );
  XNOR2_X1 U3812 ( .A(n2988), .B(n3210), .ZN(n3056) );
  XOR2_X1 U3813 ( .A(n3057), .B(n3056), .Z(n2994) );
  NAND2_X1 U3814 ( .A1(n2991), .A2(n2990), .ZN(n2992) );
  OAI21_X1 U3815 ( .B1(n2994), .B2(n2993), .A(n3060), .ZN(n3001) );
  AOI22_X1 U3816 ( .A1(n3375), .A2(n2995), .B1(n3373), .B2(n3553), .ZN(n2998)
         );
  NOR2_X1 U3817 ( .A1(STATE_REG_SCAN_IN), .A2(n2996), .ZN(n4307) );
  AOI21_X1 U3818 ( .B1(n3378), .B2(n3551), .A(n4307), .ZN(n2997) );
  OAI211_X1 U3819 ( .C1(n3376), .C2(n2999), .A(n2998), .B(n2997), .ZN(n3000)
         );
  AOI21_X1 U3820 ( .B1(n3001), .B2(n3340), .A(n3000), .ZN(n3002) );
  INV_X1 U3821 ( .A(n3002), .ZN(U3228) );
  NAND2_X1 U3822 ( .A1(n3463), .A2(n3457), .ZN(n3511) );
  XNOR2_X1 U3823 ( .A(n3003), .B(n3511), .ZN(n3007) );
  OAI22_X1 U3824 ( .A1(n3246), .A2(n4439), .B1(n4087), .B2(n3004), .ZN(n3005)
         );
  AOI21_X1 U3825 ( .B1(n4067), .B2(n3552), .A(n3005), .ZN(n3006) );
  OAI21_X1 U3826 ( .B1(n3007), .B2(n4069), .A(n3006), .ZN(n4172) );
  INV_X1 U3827 ( .A(n4172), .ZN(n3015) );
  XOR2_X1 U3828 ( .A(n3511), .B(n3008), .Z(n4173) );
  AND2_X1 U3829 ( .A1(n3009), .A2(n3193), .ZN(n3010) );
  OR2_X1 U3830 ( .A1(n3010), .A2(n3022), .ZN(n4239) );
  NOR2_X1 U3831 ( .A1(n4239), .A2(n4079), .ZN(n3013) );
  OAI22_X1 U3832 ( .A1(n4445), .A2(n3011), .B1(n3194), .B2(n4055), .ZN(n3012)
         );
  AOI211_X1 U3833 ( .C1(n4173), .C2(n4081), .A(n3013), .B(n3012), .ZN(n3014)
         );
  OAI21_X1 U3834 ( .B1(n4424), .B2(n3015), .A(n3014), .ZN(U3280) );
  XOR2_X1 U3835 ( .A(n3528), .B(n3016), .Z(n3020) );
  AOI22_X1 U3836 ( .A1(n4049), .A2(n4414), .B1(n3331), .B2(n4413), .ZN(n3017)
         );
  OAI21_X1 U3837 ( .B1(n3018), .B2(n4416), .A(n3017), .ZN(n3019) );
  AOI21_X1 U3838 ( .B1(n3020), .B2(n4436), .A(n3019), .ZN(n4170) );
  XNOR2_X1 U3839 ( .A(n3021), .B(n3528), .ZN(n4168) );
  OR2_X1 U3840 ( .A1(n3022), .A2(n3064), .ZN(n3023) );
  NAND2_X1 U3841 ( .A1(n4074), .A2(n3023), .ZN(n4171) );
  NOR2_X1 U3842 ( .A1(n4171), .A2(n4079), .ZN(n3026) );
  OAI22_X1 U3843 ( .A1(n4445), .A2(n3024), .B1(n3332), .B2(n4055), .ZN(n3025)
         );
  AOI211_X1 U3844 ( .C1(n4168), .C2(n4081), .A(n3026), .B(n3025), .ZN(n3027)
         );
  OAI21_X1 U3845 ( .B1(n4170), .B2(n4424), .A(n3027), .ZN(U3279) );
  OAI21_X1 U3846 ( .B1(n2048), .B2(n3031), .A(n3028), .ZN(n4403) );
  INV_X1 U3847 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3794) );
  INV_X1 U3848 ( .A(n4486), .ZN(n4504) );
  NAND2_X1 U3849 ( .A1(n3453), .A2(n3448), .ZN(n3510) );
  XOR2_X1 U3850 ( .A(n3510), .B(n3029), .Z(n4405) );
  XOR2_X1 U3851 ( .A(n3510), .B(n3030), .Z(n3035) );
  OAI22_X1 U3852 ( .A1(n3032), .A2(n4439), .B1(n4087), .B2(n3031), .ZN(n3033)
         );
  AOI21_X1 U3853 ( .B1(n4067), .B2(n3554), .A(n3033), .ZN(n3034) );
  OAI21_X1 U3854 ( .B1(n3035), .B2(n4069), .A(n3034), .ZN(n3036) );
  AOI21_X1 U3855 ( .B1(n4437), .B2(n4405), .A(n3036), .ZN(n4408) );
  INV_X1 U3856 ( .A(n4408), .ZN(n3037) );
  AOI21_X1 U3857 ( .B1(n4504), .B2(n4405), .A(n3037), .ZN(n3039) );
  MUX2_X1 U3858 ( .A(n3794), .B(n3039), .S(n4525), .Z(n3038) );
  OAI21_X1 U3859 ( .B1(n4403), .B2(n4238), .A(n3038), .ZN(U3483) );
  MUX2_X1 U3860 ( .A(n2353), .B(n3039), .S(n4540), .Z(n3040) );
  OAI21_X1 U3861 ( .B1(n4403), .B2(n4176), .A(n3040), .ZN(U3526) );
  INV_X1 U3862 ( .A(n3041), .ZN(n3045) );
  NAND3_X1 U3863 ( .A1(n3042), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3044) );
  INV_X1 U3864 ( .A(DATAI_31_), .ZN(n3043) );
  OAI22_X1 U3865 ( .A1(n3045), .A2(n3044), .B1(STATE_REG_SCAN_IN), .B2(n3043), 
        .ZN(U3321) );
  AOI22_X1 U3866 ( .A1(n3223), .A2(n4442), .B1(n4424), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n3046) );
  OAI21_X1 U3867 ( .B1(n3047), .B2(n4079), .A(n3046), .ZN(n3048) );
  AOI21_X1 U3868 ( .B1(n3049), .B2(n4058), .A(n3048), .ZN(n3050) );
  OAI21_X1 U3869 ( .B1(n3051), .B2(n4004), .A(n3050), .ZN(U3262) );
  AOI22_X1 U3870 ( .A1(n3551), .A2(n3164), .B1(n3154), .B2(n3193), .ZN(n3061)
         );
  NAND2_X1 U3871 ( .A1(n3551), .A2(n3154), .ZN(n3053) );
  NAND2_X1 U3872 ( .A1(n3193), .A2(n2110), .ZN(n3052) );
  NAND2_X1 U3873 ( .A1(n3053), .A2(n3052), .ZN(n3054) );
  XNOR2_X1 U3874 ( .A(n3054), .B(n3210), .ZN(n3055) );
  XNOR2_X1 U3875 ( .A(n3055), .B(n3061), .ZN(n3191) );
  INV_X1 U3876 ( .A(n3056), .ZN(n3059) );
  INV_X1 U3877 ( .A(n3057), .ZN(n3058) );
  NAND2_X1 U3878 ( .A1(n3059), .A2(n3058), .ZN(n3192) );
  OR2_X1 U3879 ( .A1(n3246), .A2(n2758), .ZN(n3063) );
  NAND2_X1 U3880 ( .A1(n3331), .A2(n3154), .ZN(n3062) );
  AND2_X1 U3881 ( .A1(n3063), .A2(n3062), .ZN(n3066) );
  OAI22_X1 U3882 ( .A1(n3246), .A2(n2729), .B1(n3209), .B2(n3064), .ZN(n3065)
         );
  XNOR2_X1 U3883 ( .A(n3065), .B(n3152), .ZN(n3067) );
  NAND2_X1 U3884 ( .A1(n3066), .A2(n3067), .ZN(n3326) );
  NOR2_X1 U3885 ( .A1(n3067), .A2(n3066), .ZN(n3328) );
  NAND2_X1 U3886 ( .A1(n4049), .A2(n3164), .ZN(n3069) );
  NAND2_X1 U3887 ( .A1(n4073), .A2(n3154), .ZN(n3068) );
  NAND2_X1 U3888 ( .A1(n3069), .A2(n3068), .ZN(n3302) );
  NAND2_X1 U3889 ( .A1(n4049), .A2(n3154), .ZN(n3071) );
  NAND2_X1 U3890 ( .A1(n4073), .A2(n2110), .ZN(n3070) );
  NAND2_X1 U3891 ( .A1(n3071), .A2(n3070), .ZN(n3072) );
  XNOR2_X1 U3892 ( .A(n3072), .B(n3210), .ZN(n3303) );
  NAND2_X1 U3893 ( .A1(n3550), .A2(n3154), .ZN(n3074) );
  NAND2_X1 U3894 ( .A1(n4052), .A2(n2110), .ZN(n3073) );
  NAND2_X1 U3895 ( .A1(n3074), .A2(n3073), .ZN(n3075) );
  XNOR2_X1 U3896 ( .A(n3075), .B(n3210), .ZN(n3079) );
  NAND2_X1 U3897 ( .A1(n3550), .A2(n3164), .ZN(n3077) );
  NAND2_X1 U3898 ( .A1(n4052), .A2(n3154), .ZN(n3076) );
  NAND2_X1 U3899 ( .A1(n3077), .A2(n3076), .ZN(n3080) );
  AOI21_X1 U3900 ( .B1(n3302), .B2(n3303), .A(n3309), .ZN(n3078) );
  NOR3_X1 U3901 ( .A1(n3309), .A2(n3302), .A3(n3303), .ZN(n3083) );
  INV_X1 U3902 ( .A(n3079), .ZN(n3082) );
  INV_X1 U3903 ( .A(n3080), .ZN(n3081) );
  AND2_X1 U3904 ( .A1(n3082), .A2(n3081), .ZN(n3308) );
  OAI22_X1 U3905 ( .A1(n4042), .A2(n2729), .B1(n3209), .B2(n3173), .ZN(n3084)
         );
  XNOR2_X1 U3906 ( .A(n3084), .B(n3210), .ZN(n3085) );
  OAI22_X1 U3907 ( .A1(n4042), .A2(n2758), .B1(n2729), .B2(n3173), .ZN(n3169)
         );
  INV_X1 U3908 ( .A(n3085), .ZN(n3170) );
  OAI22_X1 U3909 ( .A1(n3266), .A2(n2729), .B1(n3209), .B2(n4015), .ZN(n3086)
         );
  XNOR2_X1 U3910 ( .A(n3086), .B(n3210), .ZN(n3088) );
  OAI22_X1 U3911 ( .A1(n4008), .A2(n2758), .B1(n2729), .B2(n3998), .ZN(n3093)
         );
  OAI22_X1 U3912 ( .A1(n4008), .A2(n2729), .B1(n3209), .B2(n3998), .ZN(n3087)
         );
  XNOR2_X1 U3913 ( .A(n3087), .B(n3210), .ZN(n3092) );
  XOR2_X1 U3914 ( .A(n3093), .B(n3092), .Z(n3263) );
  NAND2_X1 U3915 ( .A1(n4029), .A2(n3164), .ZN(n3091) );
  NAND2_X1 U3916 ( .A1(n3374), .A2(n3154), .ZN(n3090) );
  OAI22_X1 U3917 ( .A1(n3993), .A2(n2729), .B1(n3209), .B2(n3975), .ZN(n3094)
         );
  XNOR2_X1 U3918 ( .A(n3094), .B(n3210), .ZN(n3272) );
  OR2_X1 U3919 ( .A1(n3993), .A2(n2758), .ZN(n3096) );
  NAND2_X1 U3920 ( .A1(n3981), .A2(n3154), .ZN(n3095) );
  NAND2_X1 U3921 ( .A1(n3096), .A2(n3095), .ZN(n3271) );
  NOR2_X1 U3922 ( .A1(n3272), .A2(n3271), .ZN(n3097) );
  NAND2_X1 U3923 ( .A1(n3272), .A2(n3271), .ZN(n3098) );
  OAI22_X1 U3924 ( .A1(n3976), .A2(n2729), .B1(n3209), .B2(n3962), .ZN(n3099)
         );
  XNOR2_X1 U3925 ( .A(n3099), .B(n3152), .ZN(n3105) );
  INV_X1 U3926 ( .A(n3105), .ZN(n3103) );
  OR2_X1 U3927 ( .A1(n3976), .A2(n2758), .ZN(n3101) );
  NAND2_X1 U3928 ( .A1(n3957), .A2(n3154), .ZN(n3100) );
  AND2_X1 U3929 ( .A1(n3101), .A2(n3100), .ZN(n3104) );
  INV_X1 U3930 ( .A(n3104), .ZN(n3102) );
  NAND2_X1 U3931 ( .A1(n3103), .A2(n3102), .ZN(n3348) );
  OAI22_X1 U3932 ( .A1(n3521), .A2(n2729), .B1(n3209), .B2(n3947), .ZN(n3106)
         );
  XNOR2_X1 U3933 ( .A(n3106), .B(n3210), .ZN(n3108) );
  OAI22_X1 U3934 ( .A1(n3521), .A2(n2758), .B1(n2729), .B2(n3947), .ZN(n3107)
         );
  XNOR2_X1 U3935 ( .A(n3108), .B(n3107), .ZN(n3201) );
  NAND2_X1 U3936 ( .A1(n3943), .A2(n3154), .ZN(n3110) );
  NAND2_X1 U3937 ( .A1(n2110), .A2(n3112), .ZN(n3109) );
  NAND2_X1 U3938 ( .A1(n3110), .A2(n3109), .ZN(n3111) );
  XNOR2_X1 U3939 ( .A(n3111), .B(n3210), .ZN(n3115) );
  NAND2_X1 U3940 ( .A1(n3943), .A2(n3164), .ZN(n3114) );
  NAND2_X1 U3941 ( .A1(n3154), .A2(n3112), .ZN(n3113) );
  NAND2_X1 U3942 ( .A1(n3114), .A2(n3113), .ZN(n3116) );
  NAND2_X1 U3943 ( .A1(n3115), .A2(n3116), .ZN(n3292) );
  INV_X1 U3944 ( .A(n3115), .ZN(n3118) );
  INV_X1 U3945 ( .A(n3116), .ZN(n3117) );
  NAND2_X1 U3946 ( .A1(n3118), .A2(n3117), .ZN(n3294) );
  OAI22_X1 U3947 ( .A1(n3919), .A2(n2729), .B1(n3209), .B2(n3119), .ZN(n3120)
         );
  XNOR2_X1 U3948 ( .A(n3120), .B(n3210), .ZN(n3234) );
  OR2_X1 U3949 ( .A1(n3919), .A2(n2758), .ZN(n3122) );
  NAND2_X1 U3950 ( .A1(n3154), .A2(n3905), .ZN(n3121) );
  NAND2_X1 U3951 ( .A1(n3122), .A2(n3121), .ZN(n3233) );
  NOR2_X1 U3952 ( .A1(n3234), .A2(n3233), .ZN(n3123) );
  OAI22_X1 U3953 ( .A1(n3239), .A2(n2729), .B1(n3209), .B2(n3893), .ZN(n3124)
         );
  XNOR2_X1 U3954 ( .A(n3124), .B(n3210), .ZN(n3126) );
  OAI22_X1 U3955 ( .A1(n3239), .A2(n2758), .B1(n2729), .B2(n3893), .ZN(n3125)
         );
  XNOR2_X1 U3956 ( .A(n3126), .B(n3125), .ZN(n3319) );
  NOR2_X1 U3957 ( .A1(n3126), .A2(n3125), .ZN(n3181) );
  NAND2_X1 U3958 ( .A1(n3885), .A2(n3154), .ZN(n3128) );
  NAND2_X1 U3959 ( .A1(n2110), .A2(n3865), .ZN(n3127) );
  NAND2_X1 U3960 ( .A1(n3128), .A2(n3127), .ZN(n3129) );
  XNOR2_X1 U3961 ( .A(n3129), .B(n3152), .ZN(n3132) );
  AND2_X1 U3962 ( .A1(n3154), .A2(n3865), .ZN(n3130) );
  AOI21_X1 U3963 ( .B1(n3885), .B2(n3164), .A(n3130), .ZN(n3133) );
  XNOR2_X1 U3964 ( .A(n3132), .B(n3133), .ZN(n3180) );
  NOR2_X1 U3965 ( .A1(n3181), .A2(n3180), .ZN(n3131) );
  INV_X1 U3966 ( .A(n3132), .ZN(n3135) );
  INV_X1 U3967 ( .A(n3133), .ZN(n3134) );
  NAND2_X1 U3968 ( .A1(n3135), .A2(n3134), .ZN(n3139) );
  AND2_X1 U3969 ( .A1(n3154), .A2(n3848), .ZN(n3136) );
  AOI21_X1 U3970 ( .B1(n3697), .B2(n3164), .A(n3136), .ZN(n3140) );
  OAI22_X1 U3971 ( .A1(n3868), .A2(n2729), .B1(n3209), .B2(n3285), .ZN(n3138)
         );
  XNOR2_X1 U3972 ( .A(n3138), .B(n3210), .ZN(n3282) );
  NAND2_X1 U3973 ( .A1(n3280), .A2(n3282), .ZN(n3143) );
  INV_X1 U3974 ( .A(n3140), .ZN(n3141) );
  NAND2_X1 U3975 ( .A1(n3142), .A2(n3141), .ZN(n3279) );
  NAND2_X1 U3976 ( .A1(n3674), .A2(n3154), .ZN(n3145) );
  NAND2_X1 U3977 ( .A1(n2110), .A2(n3696), .ZN(n3144) );
  NAND2_X1 U3978 ( .A1(n3145), .A2(n3144), .ZN(n3146) );
  XNOR2_X1 U3979 ( .A(n3146), .B(n3152), .ZN(n3149) );
  AND2_X1 U3980 ( .A1(n3154), .A2(n3696), .ZN(n3147) );
  AOI21_X1 U3981 ( .B1(n3674), .B2(n3164), .A(n3147), .ZN(n3148) );
  NAND2_X1 U3982 ( .A1(n3149), .A2(n3148), .ZN(n3251) );
  NAND2_X1 U3983 ( .A1(n3650), .A2(n3154), .ZN(n3151) );
  NAND2_X1 U3984 ( .A1(n2110), .A2(n3673), .ZN(n3150) );
  NAND2_X1 U3985 ( .A1(n3151), .A2(n3150), .ZN(n3153) );
  XNOR2_X1 U3986 ( .A(n3153), .B(n3152), .ZN(n3159) );
  INV_X1 U3987 ( .A(n3159), .ZN(n3157) );
  AND2_X1 U3988 ( .A1(n3154), .A2(n3673), .ZN(n3155) );
  AOI21_X1 U3989 ( .B1(n3650), .B2(n3164), .A(n3155), .ZN(n3158) );
  INV_X1 U3990 ( .A(n3158), .ZN(n3156) );
  NAND2_X1 U3991 ( .A1(n3157), .A2(n3156), .ZN(n3357) );
  NAND2_X1 U3992 ( .A1(n3548), .A2(n3154), .ZN(n3161) );
  NAND2_X1 U3993 ( .A1(n2110), .A2(n3649), .ZN(n3160) );
  NAND2_X1 U3994 ( .A1(n3161), .A2(n3160), .ZN(n3162) );
  XNOR2_X1 U3995 ( .A(n3162), .B(n3210), .ZN(n3215) );
  AND2_X1 U3996 ( .A1(n3154), .A2(n3649), .ZN(n3163) );
  AOI21_X1 U3997 ( .B1(n3548), .B2(n3164), .A(n3163), .ZN(n3216) );
  XNOR2_X1 U3998 ( .A(n3215), .B(n3216), .ZN(n3207) );
  OAI22_X1 U3999 ( .A1(n3700), .A2(n3361), .B1(STATE_REG_SCAN_IN), .B2(n3750), 
        .ZN(n3166) );
  OAI22_X1 U4000 ( .A1(n3652), .A2(n3363), .B1(n3362), .B2(n3659), .ZN(n3165)
         );
  AOI211_X1 U4001 ( .C1(n3660), .C2(n3366), .A(n3166), .B(n3165), .ZN(n3167)
         );
  OAI21_X1 U4002 ( .B1(n3168), .B2(n3381), .A(n3167), .ZN(U3211) );
  XNOR2_X1 U4003 ( .A(n3170), .B(n3169), .ZN(n3171) );
  XNOR2_X1 U4004 ( .A(n3172), .B(n3171), .ZN(n3178) );
  INV_X1 U4005 ( .A(n4036), .ZN(n3176) );
  NAND2_X1 U4006 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4353) );
  OAI21_X1 U4007 ( .B1(n3363), .B2(n3266), .A(n4353), .ZN(n3175) );
  OAI22_X1 U4008 ( .A1(n3362), .A2(n3173), .B1(n4064), .B2(n3361), .ZN(n3174)
         );
  AOI211_X1 U4009 ( .C1(n3176), .C2(n3366), .A(n3175), .B(n3174), .ZN(n3177)
         );
  OAI21_X1 U4010 ( .B1(n3178), .B2(n3381), .A(n3177), .ZN(U3212) );
  INV_X1 U4011 ( .A(n3179), .ZN(n3317) );
  OAI21_X1 U4012 ( .B1(n3317), .B2(n3181), .A(n3180), .ZN(n3183) );
  NAND3_X1 U4013 ( .A1(n3183), .A2(n3340), .A3(n3182), .ZN(n3189) );
  INV_X1 U4014 ( .A(n3872), .ZN(n3187) );
  OAI22_X1 U4015 ( .A1(n3361), .A2(n3239), .B1(STATE_REG_SCAN_IN), .B2(n3184), 
        .ZN(n3186) );
  OAI22_X1 U4016 ( .A1(n3362), .A2(n3870), .B1(n3868), .B2(n3363), .ZN(n3185)
         );
  AOI211_X1 U4017 ( .C1(n3187), .C2(n3366), .A(n3186), .B(n3185), .ZN(n3188)
         );
  NAND2_X1 U4018 ( .A1(n3189), .A2(n3188), .ZN(U3213) );
  NAND2_X1 U4019 ( .A1(n3190), .A2(n3340), .ZN(n3199) );
  AOI21_X1 U4020 ( .B1(n3060), .B2(n3192), .A(n3191), .ZN(n3198) );
  AOI22_X1 U4021 ( .A1(n3375), .A2(n3193), .B1(n3373), .B2(n3552), .ZN(n3197)
         );
  AND2_X1 U4022 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n4317) );
  NOR2_X1 U4023 ( .A1(n3376), .A2(n3194), .ZN(n3195) );
  AOI211_X1 U4024 ( .C1(n3378), .C2(n4066), .A(n4317), .B(n3195), .ZN(n3196)
         );
  OAI211_X1 U4025 ( .C1(n3199), .C2(n3198), .A(n3197), .B(n3196), .ZN(U3214)
         );
  XOR2_X1 U4026 ( .A(n3201), .B(n3200), .Z(n3206) );
  AOI22_X1 U4027 ( .A1(n3375), .A2(n3942), .B1(n3373), .B2(n3549), .ZN(n3205)
         );
  NOR2_X1 U4028 ( .A1(n3202), .A2(STATE_REG_SCAN_IN), .ZN(n3614) );
  NOR2_X1 U4029 ( .A1(n3376), .A2(n3948), .ZN(n3203) );
  AOI211_X1 U4030 ( .C1(n3378), .C2(n3943), .A(n3614), .B(n3203), .ZN(n3204)
         );
  OAI211_X1 U4031 ( .C1(n3206), .C2(n3381), .A(n3205), .B(n3204), .ZN(U3216)
         );
  NAND2_X1 U4032 ( .A1(n3208), .A2(n3207), .ZN(n3232) );
  OAI22_X1 U4033 ( .A1(n3652), .A2(n2729), .B1(n3209), .B2(n3212), .ZN(n3211)
         );
  XNOR2_X1 U4034 ( .A(n3211), .B(n3210), .ZN(n3214) );
  OAI22_X1 U4035 ( .A1(n3652), .A2(n2758), .B1(n2729), .B2(n3212), .ZN(n3213)
         );
  XNOR2_X1 U4036 ( .A(n3214), .B(n3213), .ZN(n3219) );
  NAND2_X1 U4037 ( .A1(n3219), .A2(n3340), .ZN(n3231) );
  INV_X1 U4038 ( .A(n3215), .ZN(n3217) );
  NOR2_X1 U4039 ( .A1(n3217), .A2(n3216), .ZN(n3220) );
  NOR3_X1 U4040 ( .A1(n3219), .A2(n3220), .A3(n3381), .ZN(n3218) );
  NAND2_X1 U4041 ( .A1(n3232), .A2(n3218), .ZN(n3230) );
  INV_X1 U4042 ( .A(n3219), .ZN(n3222) );
  INV_X1 U40430 ( .A(n3220), .ZN(n3221) );
  NOR3_X1 U4044 ( .A1(n3222), .A2(n3381), .A3(n3221), .ZN(n3228) );
  INV_X1 U4045 ( .A(n3223), .ZN(n3226) );
  AOI22_X1 U4046 ( .A1(n3375), .A2(n3623), .B1(n3378), .B2(n3547), .ZN(n3225)
         );
  AOI22_X1 U4047 ( .A1(n3548), .A2(n3373), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3224) );
  OAI211_X1 U4048 ( .C1(n3376), .C2(n3226), .A(n3225), .B(n3224), .ZN(n3227)
         );
  NOR2_X1 U4049 ( .A1(n3228), .A2(n3227), .ZN(n3229) );
  OAI211_X1 U4050 ( .C1(n3232), .C2(n3231), .A(n3230), .B(n3229), .ZN(U3217)
         );
  XNOR2_X1 U4051 ( .A(n3234), .B(n3233), .ZN(n3235) );
  XNOR2_X1 U4052 ( .A(n3236), .B(n3235), .ZN(n3243) );
  AOI22_X1 U4053 ( .A1(n3375), .A2(n3905), .B1(n3373), .B2(n3943), .ZN(n3242)
         );
  INV_X1 U4054 ( .A(n3237), .ZN(n3908) );
  OAI22_X1 U4055 ( .A1(n3363), .A2(n3239), .B1(STATE_REG_SCAN_IN), .B2(n3238), 
        .ZN(n3240) );
  AOI21_X1 U4056 ( .B1(n3908), .B2(n3366), .A(n3240), .ZN(n3241) );
  OAI211_X1 U4057 ( .C1(n3243), .C2(n3381), .A(n3242), .B(n3241), .ZN(U3220)
         );
  XNOR2_X1 U4058 ( .A(n3303), .B(n3302), .ZN(n3244) );
  XNOR2_X1 U4059 ( .A(n3307), .B(n3244), .ZN(n3250) );
  INV_X1 U4060 ( .A(n3245), .ZN(n4077) );
  NAND2_X1 U4061 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4333) );
  OAI21_X1 U4062 ( .B1(n3363), .B2(n4064), .A(n4333), .ZN(n3248) );
  OAI22_X1 U4063 ( .A1(n3362), .A2(n4063), .B1(n3246), .B2(n3361), .ZN(n3247)
         );
  AOI211_X1 U4064 ( .C1(n4077), .C2(n3366), .A(n3248), .B(n3247), .ZN(n3249)
         );
  OAI21_X1 U4065 ( .B1(n3250), .B2(n3381), .A(n3249), .ZN(U3221) );
  NAND2_X1 U4066 ( .A1(n2033), .A2(n3251), .ZN(n3252) );
  XNOR2_X1 U4067 ( .A(n3253), .B(n3252), .ZN(n3254) );
  NAND2_X1 U4068 ( .A1(n3254), .A2(n3340), .ZN(n3261) );
  OAI22_X1 U4069 ( .A1(n3362), .A2(n3255), .B1(n3868), .B2(n3361), .ZN(n3256)
         );
  INV_X1 U4070 ( .A(n3256), .ZN(n3260) );
  AOI22_X1 U4071 ( .A1(n3378), .A2(n3650), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3259) );
  INV_X1 U4072 ( .A(n3257), .ZN(n3701) );
  NAND2_X1 U4073 ( .A1(n3366), .A2(n3701), .ZN(n3258) );
  NAND4_X1 U4074 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(U3222)
         );
  AOI21_X1 U4075 ( .B1(n3370), .B2(n3369), .A(n3262), .ZN(n3264) );
  XNOR2_X1 U4076 ( .A(n3264), .B(n3263), .ZN(n3270) );
  INV_X1 U4077 ( .A(n3265), .ZN(n4000) );
  NAND2_X1 U4078 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4372) );
  OAI21_X1 U4079 ( .B1(n3363), .B2(n3993), .A(n4372), .ZN(n3268) );
  OAI22_X1 U4080 ( .A1(n3362), .A2(n3998), .B1(n3266), .B2(n3361), .ZN(n3267)
         );
  AOI211_X1 U4081 ( .C1(n4000), .C2(n3366), .A(n3268), .B(n3267), .ZN(n3269)
         );
  OAI21_X1 U4082 ( .B1(n3270), .B2(n3381), .A(n3269), .ZN(U3223) );
  XNOR2_X1 U4083 ( .A(n3272), .B(n3271), .ZN(n3273) );
  XNOR2_X1 U4084 ( .A(n3274), .B(n3273), .ZN(n3278) );
  AOI22_X1 U4085 ( .A1(n3375), .A2(n3981), .B1(n3373), .B2(n3978), .ZN(n3277)
         );
  AND2_X1 U4086 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4385) );
  NOR2_X1 U4087 ( .A1(n3376), .A2(n3984), .ZN(n3275) );
  AOI211_X1 U4088 ( .C1(n3378), .C2(n3549), .A(n4385), .B(n3275), .ZN(n3276)
         );
  OAI211_X1 U4089 ( .C1(n3278), .C2(n3381), .A(n3277), .B(n3276), .ZN(U3225)
         );
  NAND2_X1 U4090 ( .A1(n3279), .A2(n3280), .ZN(n3281) );
  XOR2_X1 U4091 ( .A(n3282), .B(n3281), .Z(n3289) );
  INV_X1 U4092 ( .A(n3283), .ZN(n3850) );
  OAI22_X1 U4093 ( .A1(n3361), .A2(n3320), .B1(STATE_REG_SCAN_IN), .B2(n3284), 
        .ZN(n3287) );
  OAI22_X1 U4094 ( .A1(n3362), .A2(n3285), .B1(n3847), .B2(n3363), .ZN(n3286)
         );
  AOI211_X1 U4095 ( .C1(n3850), .C2(n3366), .A(n3287), .B(n3286), .ZN(n3288)
         );
  OAI21_X1 U4096 ( .B1(n3289), .B2(n3381), .A(n3288), .ZN(U3226) );
  INV_X1 U4097 ( .A(n3290), .ZN(n3295) );
  AOI21_X1 U4098 ( .B1(n3294), .B2(n3292), .A(n3291), .ZN(n3293) );
  AOI21_X1 U4099 ( .B1(n3295), .B2(n3294), .A(n3293), .ZN(n3301) );
  INV_X1 U4100 ( .A(n3296), .ZN(n3926) );
  OAI22_X1 U4101 ( .A1(n3363), .A2(n3919), .B1(STATE_REG_SCAN_IN), .B2(n3297), 
        .ZN(n3299) );
  OAI22_X1 U4102 ( .A1(n3362), .A2(n3924), .B1(n3521), .B2(n3361), .ZN(n3298)
         );
  AOI211_X1 U4103 ( .C1(n3926), .C2(n3366), .A(n3299), .B(n3298), .ZN(n3300)
         );
  OAI21_X1 U4104 ( .B1(n3301), .B2(n3381), .A(n3300), .ZN(U3230) );
  INV_X1 U4105 ( .A(n3303), .ZN(n3306) );
  INV_X1 U4106 ( .A(n3307), .ZN(n3304) );
  OAI21_X1 U4107 ( .B1(n3304), .B2(n3303), .A(n3302), .ZN(n3305) );
  OAI21_X1 U4108 ( .B1(n3307), .B2(n3306), .A(n3305), .ZN(n3311) );
  NOR2_X1 U4109 ( .A1(n3309), .A2(n3308), .ZN(n3310) );
  XNOR2_X1 U4110 ( .A(n3311), .B(n3310), .ZN(n3316) );
  AOI22_X1 U4111 ( .A1(n3375), .A2(n4052), .B1(n3373), .B2(n4049), .ZN(n3315)
         );
  NOR2_X1 U4112 ( .A1(STATE_REG_SCAN_IN), .A2(n3312), .ZN(n4346) );
  NOR2_X1 U4113 ( .A1(n3376), .A2(n4056), .ZN(n3313) );
  AOI211_X1 U4114 ( .C1(n3378), .C2(n3372), .A(n4346), .B(n3313), .ZN(n3314)
         );
  OAI211_X1 U4115 ( .C1(n3316), .C2(n3381), .A(n3315), .B(n3314), .ZN(U3231)
         );
  AOI21_X1 U4116 ( .B1(n3319), .B2(n3318), .A(n3317), .ZN(n3325) );
  INV_X1 U4117 ( .A(n3890), .ZN(n3323) );
  OAI22_X1 U4118 ( .A1(n3361), .A2(n3919), .B1(STATE_REG_SCAN_IN), .B2(n3746), 
        .ZN(n3322) );
  OAI22_X1 U4119 ( .A1(n3362), .A2(n3893), .B1(n3320), .B2(n3363), .ZN(n3321)
         );
  AOI211_X1 U4120 ( .C1(n3323), .C2(n3366), .A(n3322), .B(n3321), .ZN(n3324)
         );
  OAI21_X1 U4121 ( .B1(n3325), .B2(n3381), .A(n3324), .ZN(U3232) );
  INV_X1 U4122 ( .A(n3326), .ZN(n3327) );
  NOR2_X1 U4123 ( .A1(n3328), .A2(n3327), .ZN(n3329) );
  XNOR2_X1 U4124 ( .A(n3330), .B(n3329), .ZN(n3336) );
  AOI22_X1 U4125 ( .A1(n3375), .A2(n3331), .B1(n3373), .B2(n3551), .ZN(n3335)
         );
  NOR2_X1 U4126 ( .A1(STATE_REG_SCAN_IN), .A2(n3747), .ZN(n4329) );
  NOR2_X1 U4127 ( .A1(n3376), .A2(n3332), .ZN(n3333) );
  AOI211_X1 U4128 ( .C1(n3378), .C2(n4049), .A(n4329), .B(n3333), .ZN(n3334)
         );
  OAI211_X1 U4129 ( .C1(n3336), .C2(n3381), .A(n3335), .B(n3334), .ZN(U3233)
         );
  OAI21_X1 U4130 ( .B1(n3339), .B2(n3338), .A(n3337), .ZN(n3341) );
  NAND2_X1 U4131 ( .A1(n3341), .A2(n3340), .ZN(n3346) );
  AOI22_X1 U4132 ( .A1(n3373), .A2(n2290), .B1(REG3_REG_2__SCAN_IN), .B2(n3342), .ZN(n3345) );
  AOI22_X1 U4133 ( .A1(n3375), .A2(n3343), .B1(n3378), .B2(n3557), .ZN(n3344)
         );
  NAND3_X1 U4134 ( .A1(n3346), .A2(n3345), .A3(n3344), .ZN(U3234) );
  INV_X1 U4135 ( .A(n3347), .ZN(n3349) );
  NAND2_X1 U4136 ( .A1(n3349), .A2(n3348), .ZN(n3350) );
  XNOR2_X1 U4137 ( .A(n3351), .B(n3350), .ZN(n3356) );
  AOI22_X1 U4138 ( .A1(n3375), .A2(n3957), .B1(n3373), .B2(n3352), .ZN(n3355)
         );
  AND2_X1 U4139 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4394) );
  NOR2_X1 U4140 ( .A1(n3376), .A2(n3966), .ZN(n3353) );
  AOI211_X1 U4141 ( .C1(n3378), .C2(n3958), .A(n4394), .B(n3353), .ZN(n3354)
         );
  OAI211_X1 U4142 ( .C1(n3356), .C2(n3381), .A(n3355), .B(n3354), .ZN(U3235)
         );
  NAND2_X1 U4143 ( .A1(n2040), .A2(n3357), .ZN(n3358) );
  XNOR2_X1 U4144 ( .A(n3359), .B(n3358), .ZN(n3368) );
  INV_X1 U4145 ( .A(n3360), .ZN(n3681) );
  OAI22_X1 U4146 ( .A1(n3361), .A2(n3847), .B1(STATE_REG_SCAN_IN), .B2(n3744), 
        .ZN(n3365) );
  OAI22_X1 U4147 ( .A1(n3677), .A2(n3363), .B1(n3362), .B2(n3678), .ZN(n3364)
         );
  AOI211_X1 U4148 ( .C1(n3681), .C2(n3366), .A(n3365), .B(n3364), .ZN(n3367)
         );
  OAI21_X1 U4149 ( .B1(n3368), .B2(n3381), .A(n3367), .ZN(U3237) );
  NAND2_X1 U4150 ( .A1(n2125), .A2(n3369), .ZN(n3371) );
  XNOR2_X1 U4151 ( .A(n3371), .B(n3370), .ZN(n3382) );
  AOI22_X1 U4152 ( .A1(n3375), .A2(n3374), .B1(n3373), .B2(n3372), .ZN(n3380)
         );
  NOR2_X1 U4153 ( .A1(STATE_REG_SCAN_IN), .A2(n3824), .ZN(n4366) );
  NOR2_X1 U4154 ( .A1(n3376), .A2(n4018), .ZN(n3377) );
  AOI211_X1 U4155 ( .C1(n3378), .C2(n3978), .A(n4366), .B(n3377), .ZN(n3379)
         );
  OAI211_X1 U4156 ( .C1(n3382), .C2(n3381), .A(n3380), .B(n3379), .ZN(U3238)
         );
  AND2_X1 U4157 ( .A1(n3397), .A2(DATAI_30_), .ZN(n4095) );
  INV_X1 U4158 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4159 ( .A1(n3383), .A2(REG0_REG_31__SCAN_IN), .ZN(n3386) );
  INV_X1 U4160 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3384) );
  OR2_X1 U4161 ( .A1(n3392), .A2(n3384), .ZN(n3385) );
  OAI211_X1 U4162 ( .C1(n2010), .C2(n3387), .A(n3386), .B(n3385), .ZN(n4086)
         );
  INV_X1 U4163 ( .A(n4086), .ZN(n3421) );
  NAND2_X1 U4164 ( .A1(n3397), .A2(DATAI_29_), .ZN(n3639) );
  INV_X1 U4165 ( .A(n3629), .ZN(n3388) );
  AOI21_X1 U4166 ( .B1(n3547), .B2(n3639), .A(n3388), .ZN(n3489) );
  NAND2_X1 U4167 ( .A1(n3390), .A2(n3389), .ZN(n3630) );
  INV_X1 U4168 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3396) );
  INV_X1 U4169 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3391) );
  OR2_X1 U4170 ( .A1(n3392), .A2(n3391), .ZN(n3395) );
  NAND2_X1 U4171 ( .A1(n3393), .A2(REG0_REG_30__SCAN_IN), .ZN(n3394) );
  OAI211_X1 U4172 ( .C1(n2010), .C2(n3396), .A(n3395), .B(n3394), .ZN(n3634)
         );
  INV_X1 U4173 ( .A(n3634), .ZN(n3399) );
  NAND2_X1 U4174 ( .A1(n3397), .A2(DATAI_31_), .ZN(n4088) );
  INV_X1 U4175 ( .A(n4088), .ZN(n3398) );
  NOR2_X1 U4176 ( .A1(n3421), .A2(n3398), .ZN(n3490) );
  AOI21_X1 U4177 ( .B1(n4095), .B2(n3399), .A(n3490), .ZN(n3497) );
  OAI21_X1 U4178 ( .B1(n3547), .B2(n3639), .A(n3497), .ZN(n3415) );
  AOI21_X1 U4179 ( .B1(n3489), .B2(n3630), .A(n3415), .ZN(n3495) );
  NAND3_X1 U4180 ( .A1(n3489), .A2(n3655), .A3(n3515), .ZN(n3419) );
  INV_X1 U4181 ( .A(n3468), .ZN(n3403) );
  NOR3_X1 U4182 ( .A1(n4027), .A2(n3400), .A3(n3403), .ZN(n3404) );
  AND2_X1 U4183 ( .A1(n3402), .A2(n3401), .ZN(n3454) );
  NOR2_X1 U4184 ( .A1(n3403), .A2(n3454), .ZN(n3474) );
  OAI21_X1 U4185 ( .B1(n3404), .B2(n3474), .A(n3472), .ZN(n3408) );
  NOR2_X1 U4186 ( .A1(n3406), .A2(n2139), .ZN(n3475) );
  AOI21_X1 U4187 ( .B1(n3408), .B2(n3475), .A(n3407), .ZN(n3410) );
  OAI21_X1 U4188 ( .B1(n3410), .B2(n3409), .A(n3480), .ZN(n3412) );
  NAND2_X1 U4189 ( .A1(n3412), .A2(n3411), .ZN(n3414) );
  INV_X1 U4190 ( .A(n3413), .ZN(n3669) );
  AOI21_X1 U4191 ( .B1(n3414), .B2(n3483), .A(n3669), .ZN(n3417) );
  NOR4_X1 U4192 ( .A1(n3417), .A2(n3630), .A3(n3416), .A4(n3415), .ZN(n3418)
         );
  AOI21_X1 U4193 ( .B1(n3495), .B2(n3419), .A(n3418), .ZN(n3420) );
  AOI21_X1 U4194 ( .B1(n4095), .B2(n3421), .A(n3420), .ZN(n3425) );
  INV_X1 U4195 ( .A(n4095), .ZN(n3422) );
  NAND2_X1 U4196 ( .A1(n3634), .A2(n3422), .ZN(n3492) );
  AOI21_X1 U4197 ( .B1(n3492), .B2(n4086), .A(n4088), .ZN(n3424) );
  NOR3_X1 U4198 ( .A1(n3425), .A2(n3424), .A3(n3423), .ZN(n3539) );
  INV_X1 U4199 ( .A(n3442), .ZN(n3427) );
  NOR3_X1 U4200 ( .A1(n3427), .A2(n3474), .A3(n3426), .ZN(n3451) );
  INV_X1 U4201 ( .A(n3428), .ZN(n3429) );
  NOR2_X1 U4202 ( .A1(n3429), .A2(n3527), .ZN(n3447) );
  INV_X1 U4203 ( .A(n3519), .ZN(n4410) );
  NAND2_X1 U4204 ( .A1(n2570), .A2(n4434), .ZN(n3518) );
  OAI211_X1 U4205 ( .C1(n4245), .C2(n4410), .A(n3518), .B(n3430), .ZN(n3431)
         );
  NAND3_X1 U4206 ( .A1(n3433), .A2(n3432), .A3(n3431), .ZN(n3435) );
  OAI211_X1 U4207 ( .C1(n3437), .C2(n3436), .A(n3435), .B(n3434), .ZN(n3438)
         );
  NAND3_X1 U4208 ( .A1(n3440), .A2(n3439), .A3(n3438), .ZN(n3441) );
  NAND4_X1 U4209 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3446)
         );
  INV_X1 U4210 ( .A(n3454), .ZN(n3445) );
  AOI21_X1 U4211 ( .B1(n3447), .B2(n3446), .A(n3445), .ZN(n3450) );
  OAI211_X1 U4212 ( .C1(n3451), .C2(n3450), .A(n3449), .B(n3448), .ZN(n3462)
         );
  INV_X1 U4213 ( .A(n3452), .ZN(n3456) );
  INV_X1 U4214 ( .A(n3453), .ZN(n3455) );
  OAI21_X1 U4215 ( .B1(n3456), .B2(n3455), .A(n3454), .ZN(n3461) );
  AND2_X1 U4216 ( .A1(n3458), .A2(n3457), .ZN(n3459) );
  NAND2_X1 U4217 ( .A1(n3466), .A2(n3459), .ZN(n3464) );
  AOI211_X1 U4218 ( .C1(n3462), .C2(n3461), .A(n3460), .B(n3464), .ZN(n3477)
         );
  INV_X1 U4219 ( .A(n3463), .ZN(n3471) );
  INV_X1 U4220 ( .A(n3464), .ZN(n3470) );
  OAI21_X1 U4221 ( .B1(n2132), .B2(n3508), .A(n3466), .ZN(n3467) );
  NAND4_X1 U4222 ( .A1(n4006), .A2(n3507), .A3(n3468), .A4(n3467), .ZN(n3469)
         );
  AOI21_X1 U4223 ( .B1(n3471), .B2(n3470), .A(n3469), .ZN(n3473) );
  OAI21_X1 U4224 ( .B1(n3474), .B2(n3473), .A(n3472), .ZN(n3476) );
  OAI211_X1 U4225 ( .C1(n3477), .C2(n3476), .A(n3475), .B(n2137), .ZN(n3478)
         );
  AND2_X1 U4226 ( .A1(n3479), .A2(n3478), .ZN(n3481) );
  OAI21_X1 U4227 ( .B1(n3857), .B2(n3481), .A(n3480), .ZN(n3482) );
  INV_X1 U4228 ( .A(n3482), .ZN(n3485) );
  OAI211_X1 U4229 ( .C1(n3486), .C2(n3485), .A(n3484), .B(n3483), .ZN(n3487)
         );
  NAND4_X1 U4230 ( .A1(n3489), .A2(n2034), .A3(n3488), .A4(n3487), .ZN(n3494)
         );
  INV_X1 U4231 ( .A(n3490), .ZN(n3493) );
  OR2_X1 U4232 ( .A1(n4086), .A2(n4088), .ZN(n3491) );
  NAND2_X1 U4233 ( .A1(n3492), .A2(n3491), .ZN(n3501) );
  AOI22_X1 U4234 ( .A1(n3495), .A2(n3494), .B1(n3493), .B2(n3501), .ZN(n3537)
         );
  NAND2_X1 U4235 ( .A1(n3497), .A2(n3496), .ZN(n3502) );
  INV_X1 U4236 ( .A(n3498), .ZN(n3499) );
  NOR2_X1 U4237 ( .A1(n3500), .A2(n3499), .ZN(n3917) );
  NOR4_X1 U4238 ( .A1(n3621), .A2(n3502), .A3(n3917), .A4(n3501), .ZN(n3514)
         );
  NAND2_X1 U4239 ( .A1(n3668), .A2(n3503), .ZN(n3693) );
  NAND2_X1 U4240 ( .A1(n3840), .A2(n3504), .ZN(n3863) );
  NAND2_X1 U4241 ( .A1(n3505), .A2(n3691), .ZN(n3843) );
  NAND2_X1 U4242 ( .A1(n3933), .A2(n3932), .ZN(n3974) );
  NOR4_X1 U4243 ( .A1(n3693), .A2(n3863), .A3(n3843), .A4(n3974), .ZN(n3513)
         );
  NAND2_X1 U4244 ( .A1(n3507), .A2(n3506), .ZN(n4051) );
  INV_X1 U4245 ( .A(n4043), .ZN(n3509) );
  OR2_X1 U4246 ( .A1(n3509), .A2(n3508), .ZN(n4071) );
  NOR4_X1 U4247 ( .A1(n4051), .A2(n4071), .A3(n3511), .A4(n3510), .ZN(n3512)
         );
  NAND4_X1 U4248 ( .A1(n3514), .A2(n3655), .A3(n3513), .A4(n3512), .ZN(n3535)
         );
  NAND2_X1 U4249 ( .A1(n3516), .A2(n3515), .ZN(n3671) );
  INV_X1 U4250 ( .A(n3859), .ZN(n3517) );
  OR2_X1 U4251 ( .A1(n3857), .A2(n3517), .ZN(n3899) );
  NAND2_X1 U4252 ( .A1(n3519), .A2(n3518), .ZN(n4482) );
  NOR4_X1 U4253 ( .A1(n3671), .A2(n3899), .A3(n4014), .A4(n4482), .ZN(n3524)
         );
  INV_X1 U4254 ( .A(n3883), .ZN(n3880) );
  NOR4_X1 U4255 ( .A1(n3520), .A2(n3880), .A3(n4024), .A4(n2569), .ZN(n3523)
         );
  XNOR2_X1 U4256 ( .A(n3521), .B(n3947), .ZN(n3938) );
  NAND4_X1 U4257 ( .A1(n3524), .A2(n3523), .A3(n3522), .A4(n3938), .ZN(n3534)
         );
  XNOR2_X1 U4258 ( .A(n3547), .B(n3639), .ZN(n3631) );
  NOR4_X1 U4259 ( .A1(n3528), .A2(n3527), .A3(n3526), .A4(n3525), .ZN(n3532)
         );
  NOR2_X1 U4260 ( .A1(n3530), .A2(n3529), .ZN(n3531) );
  NAND4_X1 U4261 ( .A1(n3532), .A2(n2159), .A3(n3991), .A4(n3531), .ZN(n3533)
         );
  NOR4_X1 U4262 ( .A1(n3535), .A2(n3534), .A3(n3631), .A4(n3533), .ZN(n3536)
         );
  MUX2_X1 U4263 ( .A(n3537), .B(n3536), .S(n4246), .Z(n3538) );
  NOR2_X1 U4264 ( .A1(n3539), .A2(n3538), .ZN(n3540) );
  XNOR2_X1 U4265 ( .A(n3540), .B(n3616), .ZN(n3546) );
  NAND2_X1 U4266 ( .A1(n3542), .A2(n3541), .ZN(n3543) );
  OAI211_X1 U4267 ( .C1(n4244), .C2(n3545), .A(n3543), .B(B_REG_SCAN_IN), .ZN(
        n3544) );
  OAI21_X1 U4268 ( .B1(n3546), .B2(n3545), .A(n3544), .ZN(U3239) );
  MUX2_X1 U4269 ( .A(DATAO_REG_31__SCAN_IN), .B(n4086), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4270 ( .A(DATAO_REG_30__SCAN_IN), .B(n3634), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4271 ( .A(n3547), .B(DATAO_REG_29__SCAN_IN), .S(n3558), .Z(U3579)
         );
  MUX2_X1 U4272 ( .A(DATAO_REG_28__SCAN_IN), .B(n3624), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4273 ( .A(n3548), .B(DATAO_REG_27__SCAN_IN), .S(n3558), .Z(U3577)
         );
  MUX2_X1 U4274 ( .A(n3650), .B(DATAO_REG_26__SCAN_IN), .S(n3558), .Z(U3576)
         );
  MUX2_X1 U4275 ( .A(n3674), .B(DATAO_REG_25__SCAN_IN), .S(n3558), .Z(U3575)
         );
  MUX2_X1 U4276 ( .A(n3697), .B(DATAO_REG_24__SCAN_IN), .S(n3558), .Z(U3574)
         );
  MUX2_X1 U4277 ( .A(n3885), .B(DATAO_REG_23__SCAN_IN), .S(n3558), .Z(U3573)
         );
  MUX2_X1 U4278 ( .A(n3943), .B(DATAO_REG_20__SCAN_IN), .S(n3558), .Z(U3570)
         );
  MUX2_X1 U4279 ( .A(DATAO_REG_18__SCAN_IN), .B(n3549), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4280 ( .A(DATAO_REG_16__SCAN_IN), .B(n3978), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4281 ( .A(n3550), .B(DATAO_REG_13__SCAN_IN), .S(n3558), .Z(U3563)
         );
  MUX2_X1 U4282 ( .A(n4049), .B(DATAO_REG_12__SCAN_IN), .S(n3558), .Z(U3562)
         );
  MUX2_X1 U4283 ( .A(DATAO_REG_11__SCAN_IN), .B(n4066), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4284 ( .A(n3551), .B(DATAO_REG_10__SCAN_IN), .S(n3558), .Z(U3560)
         );
  MUX2_X1 U4285 ( .A(n3552), .B(DATAO_REG_9__SCAN_IN), .S(n3558), .Z(U3559) );
  MUX2_X1 U4286 ( .A(n3553), .B(DATAO_REG_8__SCAN_IN), .S(n3558), .Z(U3558) );
  MUX2_X1 U4287 ( .A(DATAO_REG_7__SCAN_IN), .B(n3554), .S(U4043), .Z(U3557) );
  MUX2_X1 U4288 ( .A(n3555), .B(DATAO_REG_6__SCAN_IN), .S(n3558), .Z(U3556) );
  MUX2_X1 U4289 ( .A(DATAO_REG_4__SCAN_IN), .B(n3556), .S(U4043), .Z(U3554) );
  MUX2_X1 U4290 ( .A(n3557), .B(DATAO_REG_3__SCAN_IN), .S(n3558), .Z(U3553) );
  MUX2_X1 U4291 ( .A(DATAO_REG_2__SCAN_IN), .B(n2735), .S(U4043), .Z(U3552) );
  MUX2_X1 U4292 ( .A(n2570), .B(DATAO_REG_0__SCAN_IN), .S(n3558), .Z(U3550) );
  OAI211_X1 U4293 ( .C1(n3561), .C2(n3560), .A(n4341), .B(n3559), .ZN(n3569)
         );
  OAI211_X1 U4294 ( .C1(n3564), .C2(n3563), .A(n4397), .B(n3562), .ZN(n3568)
         );
  AOI22_X1 U4295 ( .A1(n4395), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3567) );
  NAND4_X1 U4296 ( .A1(n3569), .A2(n3568), .A3(n3567), .A4(n3566), .ZN(U3241)
         );
  MUX2_X1 U4297 ( .A(n3949), .B(REG2_REG_19__SCAN_IN), .S(n3616), .Z(n3589) );
  INV_X1 U4298 ( .A(n3590), .ZN(n4458) );
  AOI22_X1 U4299 ( .A1(n3590), .A2(n3967), .B1(REG2_REG_18__SCAN_IN), .B2(
        n4458), .ZN(n4393) );
  AOI22_X1 U4300 ( .A1(REG2_REG_17__SCAN_IN), .A2(n4459), .B1(n4390), .B2(
        n3985), .ZN(n4383) );
  INV_X1 U4301 ( .A(n3606), .ZN(n4466) );
  INV_X1 U4302 ( .A(n4467), .ZN(n4352) );
  NOR2_X1 U4303 ( .A1(n4352), .A2(n4057), .ZN(n4340) );
  AOI22_X1 U4304 ( .A1(n4470), .A2(REG2_REG_11__SCAN_IN), .B1(n3024), .B2(
        n4327), .ZN(n4324) );
  NAND2_X1 U4305 ( .A1(n4472), .A2(REG2_REG_9__SCAN_IN), .ZN(n3578) );
  INV_X1 U4306 ( .A(n4472), .ZN(n4305) );
  AOI22_X1 U4307 ( .A1(n4472), .A2(REG2_REG_9__SCAN_IN), .B1(n2983), .B2(n4305), .ZN(n4302) );
  NAND2_X1 U4308 ( .A1(REG2_REG_7__SCAN_IN), .A2(n3596), .ZN(n3575) );
  AOI22_X1 U4309 ( .A1(REG2_REG_7__SCAN_IN), .A2(n3596), .B1(n4477), .B2(n2343), .ZN(n4284) );
  NAND2_X1 U4310 ( .A1(n3594), .A2(n3573), .ZN(n3574) );
  NAND2_X1 U4311 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4271), .ZN(n4270) );
  NAND2_X1 U4312 ( .A1(n3574), .A2(n4270), .ZN(n4283) );
  NAND2_X1 U4313 ( .A1(n4284), .A2(n4283), .ZN(n4282) );
  NAND2_X1 U4314 ( .A1(n3575), .A2(n4282), .ZN(n3576) );
  NAND2_X1 U4315 ( .A1(n4474), .A2(n3576), .ZN(n3577) );
  INV_X1 U4316 ( .A(n4474), .ZN(n4296) );
  XNOR2_X1 U4317 ( .A(n3576), .B(n4296), .ZN(n4288) );
  NAND2_X1 U4318 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4288), .ZN(n4287) );
  NAND2_X1 U4319 ( .A1(n3579), .A2(n4309), .ZN(n3580) );
  NAND2_X1 U4320 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4313), .ZN(n4312) );
  NAND2_X1 U4321 ( .A1(n3580), .A2(n4312), .ZN(n4323) );
  NAND2_X1 U4322 ( .A1(n4324), .A2(n4323), .ZN(n4322) );
  NAND2_X1 U4323 ( .A1(n3602), .A2(n3581), .ZN(n3582) );
  OAI22_X1 U4324 ( .A1(n4340), .A2(n4343), .B1(n4467), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n3583) );
  NOR2_X1 U4325 ( .A1(n4466), .A2(n3583), .ZN(n3584) );
  XOR2_X1 U4326 ( .A(n3606), .B(n3583), .Z(n4355) );
  NOR2_X1 U4327 ( .A1(n4037), .A2(n4355), .ZN(n4354) );
  NAND2_X1 U4328 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3591), .ZN(n3585) );
  OAI21_X1 U4329 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3591), .A(n3585), .ZN(n4363) );
  INV_X1 U4330 ( .A(n3609), .ZN(n4462) );
  NAND2_X1 U4331 ( .A1(n3586), .A2(n4462), .ZN(n3587) );
  NAND2_X1 U4332 ( .A1(n4383), .A2(n4381), .ZN(n4382) );
  AOI21_X1 U4333 ( .B1(n3590), .B2(REG2_REG_18__SCAN_IN), .A(n4392), .ZN(n3588) );
  XOR2_X1 U4334 ( .A(n3589), .B(n3588), .Z(n3620) );
  AOI22_X1 U4335 ( .A1(n3590), .A2(REG1_REG_18__SCAN_IN), .B1(n3611), .B2(
        n4458), .ZN(n4398) );
  INV_X1 U4336 ( .A(n3591), .ZN(n4464) );
  AOI22_X1 U4337 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3591), .B1(n4464), .B2(
        n4152), .ZN(n4369) );
  AOI22_X1 U4338 ( .A1(n4467), .A2(REG1_REG_13__SCAN_IN), .B1(n3706), .B2(
        n4352), .ZN(n4349) );
  AOI22_X1 U4339 ( .A1(n4470), .A2(REG1_REG_11__SCAN_IN), .B1(n3808), .B2(
        n4327), .ZN(n4321) );
  NAND2_X1 U4340 ( .A1(n4472), .A2(REG1_REG_9__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4341 ( .A1(n4472), .A2(REG1_REG_9__SCAN_IN), .B1(n2367), .B2(n4305), .ZN(n4299) );
  NOR2_X1 U4342 ( .A1(n3593), .A2(n2145), .ZN(n3595) );
  INV_X1 U4343 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4267) );
  NAND2_X1 U4344 ( .A1(REG1_REG_7__SCAN_IN), .A2(n3596), .ZN(n4274) );
  INV_X1 U4345 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4536) );
  NAND2_X1 U4346 ( .A1(n4536), .A2(n4477), .ZN(n4275) );
  NAND2_X1 U4347 ( .A1(n4474), .A2(n3597), .ZN(n3598) );
  NAND2_X1 U4348 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4293), .ZN(n4292) );
  NAND2_X1 U4349 ( .A1(n3600), .A2(n4309), .ZN(n3601) );
  NAND2_X1 U4350 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4311), .ZN(n4310) );
  NAND2_X1 U4351 ( .A1(n3602), .A2(n3603), .ZN(n3604) );
  NAND2_X1 U4352 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4337), .ZN(n4336) );
  NAND2_X1 U4353 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  NAND2_X1 U4354 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4359), .ZN(n4358) );
  NAND2_X1 U4355 ( .A1(n3607), .A2(n4358), .ZN(n4368) );
  NAND2_X1 U4356 ( .A1(n4369), .A2(n4368), .ZN(n4367) );
  NOR2_X1 U4357 ( .A1(n3609), .A2(n3608), .ZN(n3610) );
  AOI22_X1 U4358 ( .A1(REG1_REG_17__SCAN_IN), .A2(n4390), .B1(n4459), .B2(
        n4143), .ZN(n4386) );
  NAND2_X1 U4359 ( .A1(n4398), .A2(n2012), .ZN(n4396) );
  OAI21_X1 U4360 ( .B1(n3611), .B2(n4458), .A(n4396), .ZN(n3613) );
  XNOR2_X1 U4361 ( .A(n3616), .B(n4136), .ZN(n3612) );
  XNOR2_X1 U4362 ( .A(n3613), .B(n3612), .ZN(n3618) );
  AOI21_X1 U4363 ( .B1(n4395), .B2(ADDR_REG_19__SCAN_IN), .A(n3614), .ZN(n3615) );
  OAI21_X1 U4364 ( .B1(n4401), .B2(n3616), .A(n3615), .ZN(n3617) );
  AOI21_X1 U4365 ( .B1(n3618), .B2(n4397), .A(n3617), .ZN(n3619) );
  OAI21_X1 U4366 ( .B1(n3620), .B2(n4391), .A(n3619), .ZN(U3259) );
  NAND2_X1 U4367 ( .A1(n3622), .A2(n3621), .ZN(n3626) );
  NAND2_X1 U4368 ( .A1(n3626), .A2(n3625), .ZN(n3628) );
  XNOR2_X1 U4369 ( .A(n3628), .B(n3627), .ZN(n4097) );
  INV_X1 U4370 ( .A(n4097), .ZN(n3645) );
  OAI21_X1 U4371 ( .B1(n3648), .B2(n3630), .A(n3629), .ZN(n3632) );
  XNOR2_X1 U4372 ( .A(n3632), .B(n3631), .ZN(n3637) );
  AOI21_X1 U4373 ( .B1(n4259), .B2(B_REG_SCAN_IN), .A(n4439), .ZN(n4085) );
  INV_X1 U4374 ( .A(n3639), .ZN(n3633) );
  AOI22_X1 U4375 ( .A1(n3634), .A2(n4085), .B1(n4413), .B2(n3633), .ZN(n3635)
         );
  OAI21_X1 U4376 ( .B1(n3652), .B2(n4416), .A(n3635), .ZN(n3636) );
  AOI21_X1 U4377 ( .B1(n3637), .B2(n4436), .A(n3636), .ZN(n4099) );
  OAI21_X1 U4378 ( .B1(n4055), .B2(n3638), .A(n4099), .ZN(n3643) );
  OAI22_X1 U4379 ( .A1(n4098), .A2(n4079), .B1(n3641), .B2(n4445), .ZN(n3642)
         );
  AOI21_X1 U4380 ( .B1(n3643), .B2(n4058), .A(n3642), .ZN(n3644) );
  OAI21_X1 U4381 ( .B1(n3645), .B2(n4004), .A(n3644), .ZN(U3354) );
  NOR2_X1 U4382 ( .A1(n3646), .A2(n3655), .ZN(n3647) );
  AOI22_X1 U4383 ( .A1(n3650), .A2(n4067), .B1(n3649), .B2(n4413), .ZN(n3651)
         );
  OAI21_X1 U4384 ( .B1(n3652), .B2(n4439), .A(n3651), .ZN(n3653) );
  AOI21_X1 U4385 ( .B1(n3654), .B2(n4436), .A(n3653), .ZN(n4102) );
  XNOR2_X1 U4386 ( .A(n3656), .B(n3655), .ZN(n4101) );
  NAND2_X1 U4387 ( .A1(n4101), .A2(n4081), .ZN(n3666) );
  INV_X1 U4388 ( .A(n3657), .ZN(n3658) );
  OAI21_X1 U4389 ( .B1(n3680), .B2(n3659), .A(n3658), .ZN(n4104) );
  INV_X1 U4390 ( .A(n4104), .ZN(n3664) );
  INV_X1 U4391 ( .A(n3660), .ZN(n3662) );
  OAI22_X1 U4392 ( .A1(n3662), .A2(n4055), .B1(n3661), .B2(n4445), .ZN(n3663)
         );
  AOI21_X1 U4393 ( .B1(n3664), .B2(n4428), .A(n3663), .ZN(n3665) );
  OAI211_X1 U4394 ( .C1(n4102), .C2(n4424), .A(n3666), .B(n3665), .ZN(U3263)
         );
  XOR2_X1 U4395 ( .A(n3671), .B(n3667), .Z(n4106) );
  INV_X1 U4396 ( .A(n4106), .ZN(n3685) );
  OAI21_X1 U4397 ( .B1(n3690), .B2(n3669), .A(n3668), .ZN(n3670) );
  XOR2_X1 U4398 ( .A(n3671), .B(n3670), .Z(n3672) );
  NAND2_X1 U4399 ( .A1(n3672), .A2(n4436), .ZN(n3676) );
  AOI22_X1 U4400 ( .A1(n3674), .A2(n4067), .B1(n3673), .B2(n4413), .ZN(n3675)
         );
  OAI211_X1 U4401 ( .C1(n3677), .C2(n4439), .A(n3676), .B(n3675), .ZN(n4105)
         );
  NOR2_X1 U4402 ( .A1(n3688), .A2(n3678), .ZN(n3679) );
  AOI22_X1 U4403 ( .A1(n4424), .A2(REG2_REG_26__SCAN_IN), .B1(n3681), .B2(
        n4442), .ZN(n3682) );
  OAI21_X1 U4404 ( .B1(n4189), .B2(n4079), .A(n3682), .ZN(n3683) );
  AOI21_X1 U4405 ( .B1(n4105), .B2(n4058), .A(n3683), .ZN(n3684) );
  OAI21_X1 U4406 ( .B1(n3685), .B2(n4004), .A(n3684), .ZN(U3264) );
  XOR2_X1 U4407 ( .A(n3693), .B(n3687), .Z(n4110) );
  AND2_X1 U4408 ( .A1(n2041), .A2(n3696), .ZN(n3689) );
  OR2_X1 U4409 ( .A1(n3689), .A2(n3688), .ZN(n4193) );
  INV_X1 U4410 ( .A(n3690), .ZN(n3692) );
  NAND2_X1 U4411 ( .A1(n3692), .A2(n3691), .ZN(n3694) );
  XNOR2_X1 U4412 ( .A(n3694), .B(n3693), .ZN(n3695) );
  NAND2_X1 U4413 ( .A1(n3695), .A2(n4436), .ZN(n3699) );
  AOI22_X1 U4414 ( .A1(n3697), .A2(n4067), .B1(n3696), .B2(n4413), .ZN(n3698)
         );
  OAI211_X1 U4415 ( .C1(n3700), .C2(n4439), .A(n3699), .B(n3698), .ZN(n4109)
         );
  NAND2_X1 U4416 ( .A1(n4109), .A2(n4058), .ZN(n3703) );
  AOI22_X1 U4417 ( .A1(n4424), .A2(REG2_REG_25__SCAN_IN), .B1(n3701), .B2(
        n4442), .ZN(n3702) );
  OAI211_X1 U4418 ( .C1(n4193), .C2(n4079), .A(n3703), .B(n3702), .ZN(n3704)
         );
  AOI21_X1 U4419 ( .B1(n4110), .B2(n4081), .A(n3704), .ZN(n3838) );
  AOI22_X1 U4420 ( .A1(n3706), .A2(keyinput30), .B1(keyinput34), .B2(n4119), 
        .ZN(n3705) );
  OAI221_X1 U4421 ( .B1(n3706), .B2(keyinput30), .C1(n4119), .C2(keyinput34), 
        .A(n3705), .ZN(n3715) );
  INV_X1 U4422 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4423 ( .A1(n3709), .A2(keyinput12), .B1(n3708), .B2(keyinput31), 
        .ZN(n3707) );
  OAI221_X1 U4424 ( .B1(n3709), .B2(keyinput12), .C1(n3708), .C2(keyinput31), 
        .A(n3707), .ZN(n3714) );
  AOI22_X1 U4425 ( .A1(n2668), .A2(keyinput24), .B1(keyinput56), .B2(n2283), 
        .ZN(n3710) );
  OAI221_X1 U4426 ( .B1(n2668), .B2(keyinput24), .C1(n2283), .C2(keyinput56), 
        .A(n3710), .ZN(n3713) );
  AOI22_X1 U4427 ( .A1(n2315), .A2(keyinput62), .B1(n2359), .B2(keyinput17), 
        .ZN(n3711) );
  OAI221_X1 U4428 ( .B1(n2315), .B2(keyinput62), .C1(n2359), .C2(keyinput17), 
        .A(n3711), .ZN(n3712) );
  NOR4_X1 U4429 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3712), .ZN(n3758)
         );
  AOI22_X1 U4430 ( .A1(n3011), .A2(keyinput44), .B1(n4037), .B2(keyinput7), 
        .ZN(n3716) );
  OAI221_X1 U4431 ( .B1(n3011), .B2(keyinput44), .C1(n4037), .C2(keyinput7), 
        .A(n3716), .ZN(n3724) );
  AOI22_X1 U4432 ( .A1(n3825), .A2(keyinput55), .B1(keyinput6), .B2(n2451), 
        .ZN(n3717) );
  OAI221_X1 U4433 ( .B1(n3825), .B2(keyinput55), .C1(n2451), .C2(keyinput6), 
        .A(n3717), .ZN(n3723) );
  AOI22_X1 U4434 ( .A1(n3830), .A2(keyinput3), .B1(n3641), .B2(keyinput28), 
        .ZN(n3718) );
  OAI221_X1 U4435 ( .B1(n3830), .B2(keyinput3), .C1(n3641), .C2(keyinput28), 
        .A(n3718), .ZN(n3722) );
  INV_X1 U4436 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4437 ( .A1(n3387), .A2(keyinput32), .B1(keyinput11), .B2(n3720), 
        .ZN(n3719) );
  OAI221_X1 U4438 ( .B1(n3387), .B2(keyinput32), .C1(n3720), .C2(keyinput11), 
        .A(n3719), .ZN(n3721) );
  NOR4_X1 U4439 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3757)
         );
  INV_X1 U4440 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n3727) );
  INV_X1 U4441 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4442 ( .A1(n3727), .A2(keyinput60), .B1(n3726), .B2(keyinput5), 
        .ZN(n3725) );
  OAI221_X1 U4443 ( .B1(n3727), .B2(keyinput60), .C1(n3726), .C2(keyinput5), 
        .A(n3725), .ZN(n3739) );
  AOI22_X1 U4444 ( .A1(n3730), .A2(keyinput1), .B1(keyinput59), .B2(n3729), 
        .ZN(n3728) );
  OAI221_X1 U4445 ( .B1(n3730), .B2(keyinput1), .C1(n3729), .C2(keyinput59), 
        .A(n3728), .ZN(n3738) );
  AOI22_X1 U4446 ( .A1(n3733), .A2(keyinput36), .B1(keyinput46), .B2(n3732), 
        .ZN(n3731) );
  OAI221_X1 U4447 ( .B1(n3733), .B2(keyinput36), .C1(n3732), .C2(keyinput46), 
        .A(n3731), .ZN(n3737) );
  AOI22_X1 U4448 ( .A1(n3735), .A2(keyinput58), .B1(n3805), .B2(keyinput52), 
        .ZN(n3734) );
  OAI221_X1 U4449 ( .B1(n3735), .B2(keyinput58), .C1(n3805), .C2(keyinput52), 
        .A(n3734), .ZN(n3736) );
  NOR4_X1 U4450 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3756)
         );
  AOI22_X1 U4451 ( .A1(n3742), .A2(keyinput38), .B1(keyinput39), .B2(n3741), 
        .ZN(n3740) );
  OAI221_X1 U4452 ( .B1(n3742), .B2(keyinput38), .C1(n3741), .C2(keyinput39), 
        .A(n3740), .ZN(n3754) );
  AOI22_X1 U4453 ( .A1(n3824), .A2(keyinput19), .B1(keyinput49), .B2(n3744), 
        .ZN(n3743) );
  OAI221_X1 U4454 ( .B1(n3824), .B2(keyinput19), .C1(n3744), .C2(keyinput49), 
        .A(n3743), .ZN(n3753) );
  AOI22_X1 U4455 ( .A1(n3747), .A2(keyinput27), .B1(keyinput43), .B2(n3746), 
        .ZN(n3745) );
  OAI221_X1 U4456 ( .B1(n3747), .B2(keyinput27), .C1(n3746), .C2(keyinput43), 
        .A(n3745), .ZN(n3752) );
  INV_X1 U4457 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4458 ( .A1(n3750), .A2(keyinput54), .B1(keyinput42), .B2(n3749), 
        .ZN(n3748) );
  OAI221_X1 U4459 ( .B1(n3750), .B2(keyinput54), .C1(n3749), .C2(keyinput42), 
        .A(n3748), .ZN(n3751) );
  NOR4_X1 U4460 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(n3755)
         );
  NAND4_X1 U4461 ( .A1(n3758), .A2(n3757), .A3(n3756), .A4(n3755), .ZN(n3769)
         );
  INV_X1 U4462 ( .A(D_REG_7__SCAN_IN), .ZN(n4450) );
  INV_X1 U4463 ( .A(D_REG_5__SCAN_IN), .ZN(n4451) );
  AOI22_X1 U4464 ( .A1(n4450), .A2(keyinput15), .B1(n4451), .B2(keyinput20), 
        .ZN(n3759) );
  OAI221_X1 U4465 ( .B1(n4450), .B2(keyinput15), .C1(n4451), .C2(keyinput20), 
        .A(n3759), .ZN(n3768) );
  XOR2_X1 U4466 ( .A(IR_REG_31__SCAN_IN), .B(keyinput21), .Z(n3762) );
  XOR2_X1 U4467 ( .A(IR_REG_5__SCAN_IN), .B(keyinput8), .Z(n3761) );
  XNOR2_X1 U4468 ( .A(n2250), .B(keyinput35), .ZN(n3760) );
  NOR3_X1 U4469 ( .A1(n3762), .A2(n3761), .A3(n3760), .ZN(n3765) );
  XNOR2_X1 U4470 ( .A(IR_REG_10__SCAN_IN), .B(keyinput26), .ZN(n3764) );
  XNOR2_X1 U4471 ( .A(IR_REG_27__SCAN_IN), .B(keyinput41), .ZN(n3763) );
  NAND3_X1 U4472 ( .A1(n3765), .A2(n3764), .A3(n3763), .ZN(n3767) );
  XNOR2_X1 U4473 ( .A(n4453), .B(keyinput53), .ZN(n3766) );
  NOR4_X1 U4474 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(n3804)
         );
  INV_X1 U4475 ( .A(DATAI_28_), .ZN(n3772) );
  AOI22_X1 U4476 ( .A1(n3772), .A2(keyinput14), .B1(keyinput4), .B2(n3771), 
        .ZN(n3770) );
  OAI221_X1 U4477 ( .B1(n3772), .B2(keyinput14), .C1(n3771), .C2(keyinput4), 
        .A(n3770), .ZN(n3780) );
  INV_X1 U4478 ( .A(DATAI_16_), .ZN(n4461) );
  INV_X1 U4479 ( .A(DATAI_14_), .ZN(n4465) );
  AOI22_X1 U4480 ( .A1(n4461), .A2(keyinput45), .B1(keyinput63), .B2(n4465), 
        .ZN(n3773) );
  OAI221_X1 U4481 ( .B1(n4461), .B2(keyinput45), .C1(n4465), .C2(keyinput63), 
        .A(n3773), .ZN(n3779) );
  INV_X1 U4482 ( .A(DATAI_1_), .ZN(n3809) );
  INV_X1 U4483 ( .A(DATAI_6_), .ZN(n4478) );
  AOI22_X1 U4484 ( .A1(n3809), .A2(keyinput61), .B1(n4478), .B2(keyinput23), 
        .ZN(n3774) );
  OAI221_X1 U4485 ( .B1(n3809), .B2(keyinput61), .C1(n4478), .C2(keyinput23), 
        .A(n3774), .ZN(n3778) );
  AOI22_X1 U4486 ( .A1(n2281), .A2(keyinput29), .B1(n3776), .B2(keyinput33), 
        .ZN(n3775) );
  OAI221_X1 U4487 ( .B1(n2281), .B2(keyinput29), .C1(n3776), .C2(keyinput33), 
        .A(n3775), .ZN(n3777) );
  NOR4_X1 U4488 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3803)
         );
  INV_X1 U4489 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4490 ( .A1(n3783), .A2(keyinput50), .B1(n3782), .B2(keyinput10), 
        .ZN(n3781) );
  OAI221_X1 U4491 ( .B1(n3783), .B2(keyinput50), .C1(n3782), .C2(keyinput10), 
        .A(n3781), .ZN(n3790) );
  INV_X1 U4492 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U4493 ( .A1(n4526), .A2(keyinput16), .B1(keyinput25), .B2(n4180), 
        .ZN(n3784) );
  OAI221_X1 U4494 ( .B1(n4526), .B2(keyinput16), .C1(n4180), .C2(keyinput25), 
        .A(n3784), .ZN(n3789) );
  AOI22_X1 U4495 ( .A1(n4528), .A2(keyinput18), .B1(n4530), .B2(keyinput57), 
        .ZN(n3785) );
  OAI221_X1 U4496 ( .B1(n4528), .B2(keyinput18), .C1(n4530), .C2(keyinput57), 
        .A(n3785), .ZN(n3788) );
  AOI22_X1 U4497 ( .A1(n3808), .A2(keyinput13), .B1(keyinput51), .B2(n2695), 
        .ZN(n3786) );
  OAI221_X1 U4498 ( .B1(n3808), .B2(keyinput13), .C1(n2695), .C2(keyinput51), 
        .A(n3786), .ZN(n3787) );
  NOR4_X1 U4499 ( .A1(n3790), .A2(n3789), .A3(n3788), .A4(n3787), .ZN(n3802)
         );
  INV_X1 U4500 ( .A(D_REG_19__SCAN_IN), .ZN(n4448) );
  AOI22_X1 U4501 ( .A1(n4448), .A2(keyinput0), .B1(keyinput22), .B2(n4449), 
        .ZN(n3791) );
  OAI221_X1 U4502 ( .B1(n4448), .B2(keyinput0), .C1(n4449), .C2(keyinput22), 
        .A(n3791), .ZN(n3800) );
  AOI22_X1 U4503 ( .A1(n2335), .A2(keyinput9), .B1(n4447), .B2(keyinput37), 
        .ZN(n3792) );
  OAI221_X1 U4504 ( .B1(n2335), .B2(keyinput9), .C1(n4447), .C2(keyinput37), 
        .A(n3792), .ZN(n3799) );
  INV_X1 U4505 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4524) );
  AOI22_X1 U4506 ( .A1(n4524), .A2(keyinput2), .B1(keyinput47), .B2(n3794), 
        .ZN(n3793) );
  OAI221_X1 U4507 ( .B1(n4524), .B2(keyinput2), .C1(n3794), .C2(keyinput47), 
        .A(n3793), .ZN(n3798) );
  AOI22_X1 U4508 ( .A1(n3796), .A2(keyinput48), .B1(keyinput40), .B2(n4204), 
        .ZN(n3795) );
  OAI221_X1 U4509 ( .B1(n3796), .B2(keyinput48), .C1(n4204), .C2(keyinput40), 
        .A(n3795), .ZN(n3797) );
  NOR4_X1 U4510 ( .A1(n3800), .A2(n3799), .A3(n3798), .A4(n3797), .ZN(n3801)
         );
  NAND4_X1 U4511 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3836)
         );
  NOR4_X1 U4512 ( .A1(DATAO_REG_1__SCAN_IN), .A2(DATAO_REG_15__SCAN_IN), .A3(
        ADDR_REG_3__SCAN_IN), .A4(n3805), .ZN(n3823) );
  NOR4_X1 U4513 ( .A1(REG0_REG_28__SCAN_IN), .A2(ADDR_REG_15__SCAN_IN), .A3(
        ADDR_REG_0__SCAN_IN), .A4(DATAO_REG_19__SCAN_IN), .ZN(n3822) );
  NAND4_X1 U4514 ( .A1(DATAO_REG_21__SCAN_IN), .A2(DATAO_REG_22__SCAN_IN), 
        .A3(DATAO_REG_14__SCAN_IN), .A4(DATAO_REG_5__SCAN_IN), .ZN(n3806) );
  NOR4_X1 U4515 ( .A1(DATAI_28_), .A2(REG3_REG_27__SCAN_IN), .A3(n3807), .A4(
        n3806), .ZN(n3821) );
  NOR4_X1 U4516 ( .A1(REG2_REG_14__SCAN_IN), .A2(n4461), .A3(n2451), .A4(n4465), .ZN(n3813) );
  NOR4_X1 U4517 ( .A1(REG0_REG_9__SCAN_IN), .A2(REG0_REG_11__SCAN_IN), .A3(
        REG0_REG_8__SCAN_IN), .A4(n3808), .ZN(n3812) );
  NOR4_X1 U4518 ( .A1(REG2_REG_8__SCAN_IN), .A2(REG1_REG_5__SCAN_IN), .A3(
        REG1_REG_2__SCAN_IN), .A4(n2315), .ZN(n3811) );
  NOR4_X1 U4519 ( .A1(REG2_REG_1__SCAN_IN), .A2(REG1_REG_1__SCAN_IN), .A3(
        n3809), .A4(n4526), .ZN(n3810) );
  NAND4_X1 U4520 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3819)
         );
  NAND4_X1 U4521 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        REG0_REG_29__SCAN_IN), .A4(REG0_REG_31__SCAN_IN), .ZN(n3818) );
  NAND4_X1 U4522 ( .A1(REG1_REG_29__SCAN_IN), .A2(REG2_REG_29__SCAN_IN), .A3(
        REG1_REG_28__SCAN_IN), .A4(REG2_REG_31__SCAN_IN), .ZN(n3817) );
  NOR3_X1 U4523 ( .A1(REG0_REG_6__SCAN_IN), .A2(DATAI_6_), .A3(
        REG2_REG_0__SCAN_IN), .ZN(n3815) );
  NOR3_X1 U4524 ( .A1(REG1_REG_13__SCAN_IN), .A2(REG2_REG_10__SCAN_IN), .A3(
        n4119), .ZN(n3814) );
  NAND4_X1 U4525 ( .A1(D_REG_19__SCAN_IN), .A2(REG3_REG_0__SCAN_IN), .A3(n3815), .A4(n3814), .ZN(n3816) );
  NOR4_X1 U4526 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3820)
         );
  NAND4_X1 U4527 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3834)
         );
  NAND4_X1 U4528 ( .A1(REG3_REG_11__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .A3(
        REG3_REG_26__SCAN_IN), .A4(n3824), .ZN(n3827) );
  OR4_X1 U4529 ( .A1(REG2_REG_26__SCAN_IN), .A2(DATAI_19_), .A3(
        REG0_REG_21__SCAN_IN), .A4(n3825), .ZN(n3826) );
  NOR3_X1 U4530 ( .A1(IR_REG_27__SCAN_IN), .A2(n3827), .A3(n3826), .ZN(n3829)
         );
  NAND3_X1 U4531 ( .A1(n3829), .A2(n2250), .A3(n3828), .ZN(n3833) );
  NAND4_X1 U4532 ( .A1(n3831), .A2(n3830), .A3(IR_REG_5__SCAN_IN), .A4(
        IR_REG_3__SCAN_IN), .ZN(n3832) );
  NOR3_X1 U4533 ( .A1(n3834), .A2(n3833), .A3(n3832), .ZN(n3835) );
  XNOR2_X1 U4534 ( .A(n3836), .B(n3835), .ZN(n3837) );
  XNOR2_X1 U4535 ( .A(n3838), .B(n3837), .ZN(U3265) );
  XNOR2_X1 U4536 ( .A(n3839), .B(n3843), .ZN(n4114) );
  INV_X1 U4537 ( .A(n4114), .ZN(n3854) );
  NAND2_X1 U4538 ( .A1(n3841), .A2(n3840), .ZN(n3842) );
  XOR2_X1 U4539 ( .A(n3843), .B(n3842), .Z(n3844) );
  NAND2_X1 U4540 ( .A1(n3844), .A2(n4436), .ZN(n3846) );
  AOI22_X1 U4541 ( .A1(n3885), .A2(n4067), .B1(n4413), .B2(n3848), .ZN(n3845)
         );
  OAI211_X1 U4542 ( .C1(n3847), .C2(n4439), .A(n3846), .B(n3845), .ZN(n4113)
         );
  NAND2_X1 U4543 ( .A1(n3869), .A2(n3848), .ZN(n3849) );
  NAND2_X1 U4544 ( .A1(n2041), .A2(n3849), .ZN(n4197) );
  AOI22_X1 U4545 ( .A1(n4424), .A2(REG2_REG_24__SCAN_IN), .B1(n3850), .B2(
        n4442), .ZN(n3851) );
  OAI21_X1 U4546 ( .B1(n4197), .B2(n4079), .A(n3851), .ZN(n3852) );
  AOI21_X1 U4547 ( .B1(n4113), .B2(n4445), .A(n3852), .ZN(n3853) );
  OAI21_X1 U4548 ( .B1(n3854), .B2(n4004), .A(n3853), .ZN(U3266) );
  OR2_X1 U4549 ( .A1(n3878), .A2(n3883), .ZN(n3879) );
  NAND2_X1 U4550 ( .A1(n3879), .A2(n3855), .ZN(n3856) );
  XOR2_X1 U4551 ( .A(n3863), .B(n3856), .Z(n4118) );
  INV_X1 U4552 ( .A(n4118), .ZN(n3877) );
  INV_X1 U4553 ( .A(n3857), .ZN(n3858) );
  NAND2_X1 U4554 ( .A1(n3900), .A2(n3858), .ZN(n3860) );
  NAND2_X1 U4555 ( .A1(n3860), .A2(n3859), .ZN(n3882) );
  NAND2_X1 U4556 ( .A1(n3882), .A2(n3883), .ZN(n3881) );
  NAND2_X1 U4557 ( .A1(n3881), .A2(n3861), .ZN(n3862) );
  XOR2_X1 U4558 ( .A(n3863), .B(n3862), .Z(n3864) );
  NAND2_X1 U4559 ( .A1(n3864), .A2(n4436), .ZN(n3867) );
  AOI22_X1 U4560 ( .A1(n3901), .A2(n4067), .B1(n4413), .B2(n3865), .ZN(n3866)
         );
  OAI211_X1 U4561 ( .C1(n3868), .C2(n4439), .A(n3867), .B(n3866), .ZN(n4117)
         );
  INV_X1 U4562 ( .A(n4121), .ZN(n3871) );
  OAI21_X1 U4563 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n4201) );
  NOR2_X1 U4564 ( .A1(n4201), .A2(n4079), .ZN(n3875) );
  OAI22_X1 U4565 ( .A1(n4445), .A2(n3873), .B1(n3872), .B2(n4055), .ZN(n3874)
         );
  AOI211_X1 U4566 ( .C1(n4117), .C2(n4058), .A(n3875), .B(n3874), .ZN(n3876)
         );
  OAI21_X1 U4567 ( .B1(n3877), .B2(n4004), .A(n3876), .ZN(U3267) );
  OAI21_X1 U4568 ( .B1(n2179), .B2(n3880), .A(n3879), .ZN(n4125) );
  OAI21_X1 U4569 ( .B1(n3883), .B2(n3882), .A(n3881), .ZN(n3889) );
  NAND2_X1 U4570 ( .A1(n3884), .A2(n4413), .ZN(n3887) );
  NAND2_X1 U4571 ( .A1(n3885), .A2(n4414), .ZN(n3886) );
  OAI211_X1 U4572 ( .C1(n3919), .C2(n4416), .A(n3887), .B(n3886), .ZN(n3888)
         );
  AOI21_X1 U4573 ( .B1(n3889), .B2(n4436), .A(n3888), .ZN(n4124) );
  OAI22_X1 U4574 ( .A1(n4445), .A2(n3891), .B1(n3890), .B2(n4055), .ZN(n3892)
         );
  INV_X1 U4575 ( .A(n3892), .ZN(n3895) );
  OR2_X1 U4576 ( .A1(n3906), .A2(n3893), .ZN(n4122) );
  NAND3_X1 U4577 ( .A1(n4121), .A2(n4122), .A3(n4428), .ZN(n3894) );
  OAI211_X1 U4578 ( .C1(n4124), .C2(n4424), .A(n3895), .B(n3894), .ZN(n3896)
         );
  INV_X1 U4579 ( .A(n3896), .ZN(n3897) );
  OAI21_X1 U4580 ( .B1(n4125), .B2(n4004), .A(n3897), .ZN(U3268) );
  XOR2_X1 U4581 ( .A(n3899), .B(n3898), .Z(n4127) );
  INV_X1 U4582 ( .A(n4127), .ZN(n3912) );
  XNOR2_X1 U4583 ( .A(n3900), .B(n3899), .ZN(n3904) );
  AOI22_X1 U4584 ( .A1(n3901), .A2(n4414), .B1(n4413), .B2(n3905), .ZN(n3903)
         );
  NAND2_X1 U4585 ( .A1(n3943), .A2(n4067), .ZN(n3902) );
  OAI211_X1 U4586 ( .C1(n3904), .C2(n4069), .A(n3903), .B(n3902), .ZN(n4126)
         );
  AND2_X1 U4587 ( .A1(n3923), .A2(n3905), .ZN(n3907) );
  OR2_X1 U4588 ( .A1(n3907), .A2(n3906), .ZN(n4206) );
  AOI22_X1 U4589 ( .A1(n4424), .A2(REG2_REG_21__SCAN_IN), .B1(n3908), .B2(
        n4442), .ZN(n3909) );
  OAI21_X1 U4590 ( .B1(n4206), .B2(n4079), .A(n3909), .ZN(n3910) );
  AOI21_X1 U4591 ( .B1(n4126), .B2(n4445), .A(n3910), .ZN(n3911) );
  OAI21_X1 U4592 ( .B1(n3912), .B2(n4004), .A(n3911), .ZN(U3269) );
  XNOR2_X1 U4593 ( .A(n3913), .B(n3917), .ZN(n4131) );
  INV_X1 U4594 ( .A(n4131), .ZN(n3930) );
  INV_X1 U4595 ( .A(n3914), .ZN(n3915) );
  NAND2_X1 U4596 ( .A1(n3916), .A2(n3915), .ZN(n3918) );
  XNOR2_X1 U4597 ( .A(n3918), .B(n3917), .ZN(n3922) );
  OAI22_X1 U4598 ( .A1(n3919), .A2(n4439), .B1(n4087), .B2(n3924), .ZN(n3920)
         );
  AOI21_X1 U4599 ( .B1(n4067), .B2(n3958), .A(n3920), .ZN(n3921) );
  OAI21_X1 U4600 ( .B1(n3922), .B2(n4069), .A(n3921), .ZN(n4130) );
  INV_X1 U4601 ( .A(n3946), .ZN(n3925) );
  OAI21_X1 U4602 ( .B1(n3925), .B2(n3924), .A(n3923), .ZN(n4210) );
  AOI22_X1 U4603 ( .A1(n4424), .A2(REG2_REG_20__SCAN_IN), .B1(n3926), .B2(
        n4442), .ZN(n3927) );
  OAI21_X1 U4604 ( .B1(n4210), .B2(n4079), .A(n3927), .ZN(n3928) );
  AOI21_X1 U4605 ( .B1(n4130), .B2(n4445), .A(n3928), .ZN(n3929) );
  OAI21_X1 U4606 ( .B1(n3930), .B2(n4004), .A(n3929), .ZN(U3270) );
  XNOR2_X1 U4607 ( .A(n3931), .B(n3938), .ZN(n4135) );
  INV_X1 U4608 ( .A(n4135), .ZN(n3953) );
  INV_X1 U4609 ( .A(n3932), .ZN(n3934) );
  OAI21_X1 U4610 ( .B1(n3973), .B2(n3934), .A(n3933), .ZN(n3955) );
  INV_X1 U4611 ( .A(n3935), .ZN(n3937) );
  OAI21_X1 U4612 ( .B1(n3955), .B2(n3937), .A(n3936), .ZN(n3940) );
  INV_X1 U4613 ( .A(n3938), .ZN(n3939) );
  XNOR2_X1 U4614 ( .A(n3940), .B(n3939), .ZN(n3941) );
  NAND2_X1 U4615 ( .A1(n3941), .A2(n4436), .ZN(n3945) );
  AOI22_X1 U4616 ( .A1(n3943), .A2(n4414), .B1(n4413), .B2(n3942), .ZN(n3944)
         );
  OAI211_X1 U4617 ( .C1(n3976), .C2(n4416), .A(n3945), .B(n3944), .ZN(n4134)
         );
  OAI21_X1 U4618 ( .B1(n3963), .B2(n3947), .A(n3946), .ZN(n4214) );
  NOR2_X1 U4619 ( .A1(n4214), .A2(n4079), .ZN(n3951) );
  OAI22_X1 U4620 ( .A1(n4445), .A2(n3949), .B1(n3948), .B2(n4055), .ZN(n3950)
         );
  AOI211_X1 U4621 ( .C1(n4134), .C2(n4058), .A(n3951), .B(n3950), .ZN(n3952)
         );
  OAI21_X1 U4622 ( .B1(n3953), .B2(n4004), .A(n3952), .ZN(U3271) );
  XOR2_X1 U4623 ( .A(n3956), .B(n3954), .Z(n4140) );
  XOR2_X1 U4624 ( .A(n3956), .B(n3955), .Z(n3961) );
  AOI22_X1 U4625 ( .A1(n3958), .A2(n4414), .B1(n3957), .B2(n4413), .ZN(n3959)
         );
  OAI21_X1 U4626 ( .B1(n3993), .B2(n4416), .A(n3959), .ZN(n3960) );
  AOI21_X1 U4627 ( .B1(n3961), .B2(n4436), .A(n3960), .ZN(n4139) );
  INV_X1 U4628 ( .A(n4139), .ZN(n3970) );
  OAI21_X1 U4629 ( .B1(n3982), .B2(n3962), .A(n4512), .ZN(n3964) );
  OR2_X1 U4630 ( .A1(n3964), .A2(n3963), .ZN(n4138) );
  NOR2_X1 U4631 ( .A1(n4138), .A2(n3965), .ZN(n3969) );
  OAI22_X1 U4632 ( .A1(n4445), .A2(n3967), .B1(n3966), .B2(n4055), .ZN(n3968)
         );
  AOI211_X1 U4633 ( .C1(n3970), .C2(n4058), .A(n3969), .B(n3968), .ZN(n3971)
         );
  OAI21_X1 U4634 ( .B1(n4140), .B2(n4004), .A(n3971), .ZN(U3272) );
  XNOR2_X1 U4635 ( .A(n3972), .B(n3974), .ZN(n4142) );
  INV_X1 U4636 ( .A(n4142), .ZN(n3989) );
  XOR2_X1 U4637 ( .A(n3974), .B(n3973), .Z(n3980) );
  OAI22_X1 U4638 ( .A1(n3976), .A2(n4439), .B1(n4087), .B2(n3975), .ZN(n3977)
         );
  AOI21_X1 U4639 ( .B1(n4067), .B2(n3978), .A(n3977), .ZN(n3979) );
  OAI21_X1 U4640 ( .B1(n3980), .B2(n4069), .A(n3979), .ZN(n4141) );
  AND2_X1 U4641 ( .A1(n3997), .A2(n3981), .ZN(n3983) );
  OR2_X1 U4642 ( .A1(n3983), .A2(n3982), .ZN(n4219) );
  NOR2_X1 U4643 ( .A1(n4219), .A2(n4079), .ZN(n3987) );
  OAI22_X1 U4644 ( .A1(n4445), .A2(n3985), .B1(n3984), .B2(n4055), .ZN(n3986)
         );
  AOI211_X1 U4645 ( .C1(n4141), .C2(n4058), .A(n3987), .B(n3986), .ZN(n3988)
         );
  OAI21_X1 U4646 ( .B1(n3989), .B2(n4004), .A(n3988), .ZN(U3273) );
  XNOR2_X1 U4647 ( .A(n3990), .B(n3991), .ZN(n4146) );
  INV_X1 U4648 ( .A(n4146), .ZN(n4005) );
  XNOR2_X1 U4649 ( .A(n3992), .B(n3991), .ZN(n3996) );
  OAI22_X1 U4650 ( .A1(n3993), .A2(n4439), .B1(n4087), .B2(n3998), .ZN(n3994)
         );
  AOI21_X1 U4651 ( .B1(n4067), .B2(n4029), .A(n3994), .ZN(n3995) );
  OAI21_X1 U4652 ( .B1(n3996), .B2(n4069), .A(n3995), .ZN(n4145) );
  INV_X1 U4653 ( .A(n4017), .ZN(n3999) );
  OAI21_X1 U4654 ( .B1(n3999), .B2(n3998), .A(n3997), .ZN(n4223) );
  AOI22_X1 U4655 ( .A1(n4424), .A2(REG2_REG_16__SCAN_IN), .B1(n4000), .B2(
        n4442), .ZN(n4001) );
  OAI21_X1 U4656 ( .B1(n4223), .B2(n4079), .A(n4001), .ZN(n4002) );
  AOI21_X1 U4657 ( .B1(n4145), .B2(n4058), .A(n4002), .ZN(n4003) );
  OAI21_X1 U4658 ( .B1(n4005), .B2(n4004), .A(n4003), .ZN(U3274) );
  NAND2_X1 U4659 ( .A1(n4026), .A2(n4006), .ZN(n4007) );
  XOR2_X1 U4660 ( .A(n4014), .B(n4007), .Z(n4011) );
  NOR2_X1 U4661 ( .A1(n4042), .A2(n4416), .ZN(n4010) );
  OAI22_X1 U4662 ( .A1(n4008), .A2(n4439), .B1(n4087), .B2(n4015), .ZN(n4009)
         );
  AOI211_X1 U4663 ( .C1(n4011), .C2(n4436), .A(n4010), .B(n4009), .ZN(n4149)
         );
  XOR2_X1 U4664 ( .A(n4014), .B(n4013), .Z(n4151) );
  NAND2_X1 U4665 ( .A1(n4151), .A2(n4081), .ZN(n4023) );
  OR2_X1 U4666 ( .A1(n4033), .A2(n4015), .ZN(n4016) );
  NAND2_X1 U4667 ( .A1(n4017), .A2(n4016), .ZN(n4227) );
  INV_X1 U4668 ( .A(n4227), .ZN(n4021) );
  OAI22_X1 U4669 ( .A1(n4445), .A2(n4019), .B1(n4018), .B2(n4055), .ZN(n4020)
         );
  AOI21_X1 U4670 ( .B1(n4021), .B2(n4428), .A(n4020), .ZN(n4022) );
  OAI211_X1 U4671 ( .C1(n4424), .C2(n4149), .A(n4023), .B(n4022), .ZN(U3275)
         );
  XNOR2_X1 U4672 ( .A(n4025), .B(n4024), .ZN(n4154) );
  OAI21_X1 U4673 ( .B1(n2436), .B2(n4027), .A(n4026), .ZN(n4028) );
  NAND2_X1 U4674 ( .A1(n4028), .A2(n4436), .ZN(n4031) );
  AOI22_X1 U4675 ( .A1(n4029), .A2(n4414), .B1(n4413), .B2(n4035), .ZN(n4030)
         );
  OAI211_X1 U4676 ( .C1(n4064), .C2(n4416), .A(n4031), .B(n4030), .ZN(n4032)
         );
  AOI21_X1 U4677 ( .B1(n4154), .B2(n4437), .A(n4032), .ZN(n4158) );
  INV_X1 U4678 ( .A(n4033), .ZN(n4156) );
  INV_X1 U4679 ( .A(n4034), .ZN(n4054) );
  NAND2_X1 U4680 ( .A1(n4054), .A2(n4035), .ZN(n4155) );
  AND3_X1 U4681 ( .A1(n4156), .A2(n4428), .A3(n4155), .ZN(n4039) );
  OAI22_X1 U4682 ( .A1(n4445), .A2(n4037), .B1(n4036), .B2(n4055), .ZN(n4038)
         );
  AOI211_X1 U4683 ( .C1(n4154), .C2(n4443), .A(n4039), .B(n4038), .ZN(n4040)
         );
  OAI21_X1 U4684 ( .B1(n4158), .B2(n4424), .A(n4040), .ZN(U3276) );
  OAI22_X1 U4685 ( .A1(n4042), .A2(n4439), .B1(n4087), .B2(n4041), .ZN(n4048)
         );
  NAND2_X1 U4686 ( .A1(n4044), .A2(n4043), .ZN(n4045) );
  XOR2_X1 U4687 ( .A(n4051), .B(n4045), .Z(n4046) );
  NOR2_X1 U4688 ( .A1(n4046), .A2(n4069), .ZN(n4047) );
  AOI211_X1 U4689 ( .C1(n4067), .C2(n4049), .A(n4048), .B(n4047), .ZN(n4162)
         );
  XOR2_X1 U4690 ( .A(n4050), .B(n4051), .Z(n4160) );
  NAND2_X1 U4691 ( .A1(n4076), .A2(n4052), .ZN(n4053) );
  NAND2_X1 U4692 ( .A1(n4054), .A2(n4053), .ZN(n4163) );
  NOR2_X1 U4693 ( .A1(n4163), .A2(n4079), .ZN(n4060) );
  OAI22_X1 U4694 ( .A1(n4058), .A2(n4057), .B1(n4056), .B2(n4055), .ZN(n4059)
         );
  AOI211_X1 U4695 ( .C1(n4160), .C2(n4081), .A(n4060), .B(n4059), .ZN(n4061)
         );
  OAI21_X1 U4696 ( .B1(n4162), .B2(n4424), .A(n4061), .ZN(U3277) );
  XNOR2_X1 U4697 ( .A(n4062), .B(n4071), .ZN(n4070) );
  OAI22_X1 U4698 ( .A1(n4064), .A2(n4439), .B1(n4087), .B2(n4063), .ZN(n4065)
         );
  AOI21_X1 U4699 ( .B1(n4067), .B2(n4066), .A(n4065), .ZN(n4068) );
  OAI21_X1 U4700 ( .B1(n4070), .B2(n4069), .A(n4068), .ZN(n4164) );
  INV_X1 U4701 ( .A(n4164), .ZN(n4083) );
  XNOR2_X1 U4702 ( .A(n4072), .B(n4071), .ZN(n4165) );
  NAND2_X1 U4703 ( .A1(n4074), .A2(n4073), .ZN(n4075) );
  NAND2_X1 U4704 ( .A1(n4076), .A2(n4075), .ZN(n4233) );
  AOI22_X1 U4705 ( .A1(n4424), .A2(REG2_REG_12__SCAN_IN), .B1(n4077), .B2(
        n4442), .ZN(n4078) );
  OAI21_X1 U4706 ( .B1(n4233), .B2(n4079), .A(n4078), .ZN(n4080) );
  AOI21_X1 U4707 ( .B1(n4165), .B2(n4081), .A(n4080), .ZN(n4082) );
  OAI21_X1 U4708 ( .B1(n4083), .B2(n4424), .A(n4082), .ZN(U3278) );
  NAND2_X1 U4709 ( .A1(n4253), .A2(n4084), .ZN(n4090) );
  NAND2_X1 U4710 ( .A1(n4086), .A2(n4085), .ZN(n4093) );
  OAI21_X1 U4711 ( .B1(n4088), .B2(n4087), .A(n4093), .ZN(n4252) );
  NAND2_X1 U4712 ( .A1(n4540), .A2(n4252), .ZN(n4089) );
  OAI211_X1 U4713 ( .C1(n4540), .C2(n3384), .A(n4090), .B(n4089), .ZN(U3549)
         );
  AOI21_X1 U4714 ( .B1(n4095), .B2(n4092), .A(n4091), .ZN(n4255) );
  INV_X1 U4715 ( .A(n4255), .ZN(n4183) );
  INV_X1 U4716 ( .A(n4093), .ZN(n4094) );
  AOI21_X1 U4717 ( .B1(n4095), .B2(n4413), .A(n4094), .ZN(n4257) );
  MUX2_X1 U4718 ( .A(n3391), .B(n4257), .S(n4540), .Z(n4096) );
  OAI21_X1 U4719 ( .B1(n4183), .B2(n4176), .A(n4096), .ZN(U3548) );
  NAND2_X1 U4720 ( .A1(n4097), .A2(n4522), .ZN(n4100) );
  MUX2_X1 U4721 ( .A(REG1_REG_29__SCAN_IN), .B(n4184), .S(n4540), .Z(U3547) );
  NAND2_X1 U4722 ( .A1(n4101), .A2(n4522), .ZN(n4103) );
  OAI211_X1 U4723 ( .C1(n4519), .C2(n4104), .A(n4103), .B(n4102), .ZN(n4185)
         );
  MUX2_X1 U4724 ( .A(REG1_REG_27__SCAN_IN), .B(n4185), .S(n4540), .Z(U3545) );
  INV_X1 U4725 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4107) );
  AOI21_X1 U4726 ( .B1(n4106), .B2(n4522), .A(n4105), .ZN(n4186) );
  MUX2_X1 U4727 ( .A(n4107), .B(n4186), .S(n4540), .Z(n4108) );
  OAI21_X1 U4728 ( .B1(n4176), .B2(n4189), .A(n4108), .ZN(U3544) );
  INV_X1 U4729 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4111) );
  AOI21_X1 U4730 ( .B1(n4110), .B2(n4522), .A(n4109), .ZN(n4190) );
  MUX2_X1 U4731 ( .A(n4111), .B(n4190), .S(n4540), .Z(n4112) );
  OAI21_X1 U4732 ( .B1(n4176), .B2(n4193), .A(n4112), .ZN(U3543) );
  INV_X1 U4733 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4115) );
  AOI21_X1 U4734 ( .B1(n4114), .B2(n4522), .A(n4113), .ZN(n4194) );
  MUX2_X1 U4735 ( .A(n4115), .B(n4194), .S(n4540), .Z(n4116) );
  OAI21_X1 U4736 ( .B1(n4176), .B2(n4197), .A(n4116), .ZN(U3542) );
  AOI21_X1 U4737 ( .B1(n4118), .B2(n4522), .A(n4117), .ZN(n4198) );
  MUX2_X1 U4738 ( .A(n4119), .B(n4198), .S(n4540), .Z(n4120) );
  OAI21_X1 U4739 ( .B1(n4176), .B2(n4201), .A(n4120), .ZN(U3541) );
  NAND3_X1 U4740 ( .A1(n4122), .A2(n4512), .A3(n4121), .ZN(n4123) );
  OAI211_X1 U4741 ( .C1(n4125), .C2(n4507), .A(n4124), .B(n4123), .ZN(n4202)
         );
  MUX2_X1 U4742 ( .A(REG1_REG_22__SCAN_IN), .B(n4202), .S(n4540), .Z(U3540) );
  INV_X1 U4743 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4128) );
  AOI21_X1 U4744 ( .B1(n4127), .B2(n4522), .A(n4126), .ZN(n4203) );
  MUX2_X1 U4745 ( .A(n4128), .B(n4203), .S(n4540), .Z(n4129) );
  OAI21_X1 U4746 ( .B1(n4176), .B2(n4206), .A(n4129), .ZN(U3539) );
  AOI21_X1 U4747 ( .B1(n4131), .B2(n4522), .A(n4130), .ZN(n4207) );
  MUX2_X1 U4748 ( .A(n4132), .B(n4207), .S(n4540), .Z(n4133) );
  OAI21_X1 U4749 ( .B1(n4176), .B2(n4210), .A(n4133), .ZN(U3538) );
  AOI21_X1 U4750 ( .B1(n4135), .B2(n4522), .A(n4134), .ZN(n4211) );
  MUX2_X1 U4751 ( .A(n4136), .B(n4211), .S(n4540), .Z(n4137) );
  OAI21_X1 U4752 ( .B1(n4176), .B2(n4214), .A(n4137), .ZN(U3537) );
  OAI211_X1 U4753 ( .C1(n4140), .C2(n4507), .A(n4139), .B(n4138), .ZN(n4215)
         );
  MUX2_X1 U4754 ( .A(REG1_REG_18__SCAN_IN), .B(n4215), .S(n4540), .Z(U3536) );
  AOI21_X1 U4755 ( .B1(n4142), .B2(n4522), .A(n4141), .ZN(n4216) );
  MUX2_X1 U4756 ( .A(n4143), .B(n4216), .S(n4540), .Z(n4144) );
  OAI21_X1 U4757 ( .B1(n4176), .B2(n4219), .A(n4144), .ZN(U3535) );
  AOI21_X1 U4758 ( .B1(n4146), .B2(n4522), .A(n4145), .ZN(n4220) );
  MUX2_X1 U4759 ( .A(n4147), .B(n4220), .S(n4540), .Z(n4148) );
  OAI21_X1 U4760 ( .B1(n4176), .B2(n4223), .A(n4148), .ZN(U3534) );
  INV_X1 U4761 ( .A(n4149), .ZN(n4150) );
  AOI21_X1 U4762 ( .B1(n4522), .B2(n4151), .A(n4150), .ZN(n4224) );
  MUX2_X1 U4763 ( .A(n4152), .B(n4224), .S(n4540), .Z(n4153) );
  OAI21_X1 U4764 ( .B1(n4176), .B2(n4227), .A(n4153), .ZN(U3533) );
  INV_X1 U4765 ( .A(n4154), .ZN(n4159) );
  NAND3_X1 U4766 ( .A1(n4156), .A2(n4512), .A3(n4155), .ZN(n4157) );
  OAI211_X1 U4767 ( .C1(n4159), .C2(n4486), .A(n4158), .B(n4157), .ZN(n4228)
         );
  MUX2_X1 U4768 ( .A(REG1_REG_14__SCAN_IN), .B(n4228), .S(n4540), .Z(U3532) );
  NAND2_X1 U4769 ( .A1(n4160), .A2(n4522), .ZN(n4161) );
  OAI211_X1 U4770 ( .C1(n4519), .C2(n4163), .A(n4162), .B(n4161), .ZN(n4229)
         );
  MUX2_X1 U4771 ( .A(REG1_REG_13__SCAN_IN), .B(n4229), .S(n4540), .Z(U3531) );
  AOI21_X1 U4772 ( .B1(n4522), .B2(n4165), .A(n4164), .ZN(n4230) );
  MUX2_X1 U4773 ( .A(n4166), .B(n4230), .S(n4540), .Z(n4167) );
  OAI21_X1 U4774 ( .B1(n4176), .B2(n4233), .A(n4167), .ZN(U3530) );
  NAND2_X1 U4775 ( .A1(n4168), .A2(n4522), .ZN(n4169) );
  OAI211_X1 U4776 ( .C1(n4519), .C2(n4171), .A(n4170), .B(n4169), .ZN(n4234)
         );
  MUX2_X1 U4777 ( .A(REG1_REG_11__SCAN_IN), .B(n4234), .S(n4540), .Z(U3529) );
  AOI21_X1 U4778 ( .B1(n4173), .B2(n4522), .A(n4172), .ZN(n4235) );
  MUX2_X1 U4779 ( .A(n4174), .B(n4235), .S(n4540), .Z(n4175) );
  OAI21_X1 U4780 ( .B1(n4176), .B2(n4239), .A(n4175), .ZN(U3528) );
  NAND2_X1 U4781 ( .A1(n4253), .A2(n4177), .ZN(n4179) );
  NAND2_X1 U4782 ( .A1(n4525), .A2(n4252), .ZN(n4178) );
  OAI211_X1 U4783 ( .C1(n4525), .C2(n4180), .A(n4179), .B(n4178), .ZN(U3517)
         );
  INV_X1 U4784 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4181) );
  MUX2_X1 U4785 ( .A(n4181), .B(n4257), .S(n4525), .Z(n4182) );
  OAI21_X1 U4786 ( .B1(n4183), .B2(n4238), .A(n4182), .ZN(U3516) );
  MUX2_X1 U4787 ( .A(REG0_REG_29__SCAN_IN), .B(n4184), .S(n4525), .Z(U3515) );
  MUX2_X1 U4788 ( .A(REG0_REG_27__SCAN_IN), .B(n4185), .S(n4525), .Z(U3513) );
  INV_X1 U4789 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4187) );
  MUX2_X1 U4790 ( .A(n4187), .B(n4186), .S(n4525), .Z(n4188) );
  OAI21_X1 U4791 ( .B1(n4189), .B2(n4238), .A(n4188), .ZN(U3512) );
  INV_X1 U4792 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4191) );
  MUX2_X1 U4793 ( .A(n4191), .B(n4190), .S(n4525), .Z(n4192) );
  OAI21_X1 U4794 ( .B1(n4193), .B2(n4238), .A(n4192), .ZN(U3511) );
  INV_X1 U4795 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4195) );
  MUX2_X1 U4796 ( .A(n4195), .B(n4194), .S(n4525), .Z(n4196) );
  OAI21_X1 U4797 ( .B1(n4197), .B2(n4238), .A(n4196), .ZN(U3510) );
  INV_X1 U4798 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4199) );
  MUX2_X1 U4799 ( .A(n4199), .B(n4198), .S(n4525), .Z(n4200) );
  OAI21_X1 U4800 ( .B1(n4201), .B2(n4238), .A(n4200), .ZN(U3509) );
  MUX2_X1 U4801 ( .A(REG0_REG_22__SCAN_IN), .B(n4202), .S(n4525), .Z(U3508) );
  MUX2_X1 U4802 ( .A(n4204), .B(n4203), .S(n4525), .Z(n4205) );
  OAI21_X1 U4803 ( .B1(n4206), .B2(n4238), .A(n4205), .ZN(U3507) );
  INV_X1 U4804 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4208) );
  MUX2_X1 U4805 ( .A(n4208), .B(n4207), .S(n4525), .Z(n4209) );
  OAI21_X1 U4806 ( .B1(n4210), .B2(n4238), .A(n4209), .ZN(U3506) );
  INV_X1 U4807 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4212) );
  MUX2_X1 U4808 ( .A(n4212), .B(n4211), .S(n4525), .Z(n4213) );
  OAI21_X1 U4809 ( .B1(n4214), .B2(n4238), .A(n4213), .ZN(U3505) );
  MUX2_X1 U4810 ( .A(REG0_REG_18__SCAN_IN), .B(n4215), .S(n4525), .Z(U3503) );
  INV_X1 U4811 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4217) );
  MUX2_X1 U4812 ( .A(n4217), .B(n4216), .S(n4525), .Z(n4218) );
  OAI21_X1 U4813 ( .B1(n4219), .B2(n4238), .A(n4218), .ZN(U3501) );
  INV_X1 U4814 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4221) );
  MUX2_X1 U4815 ( .A(n4221), .B(n4220), .S(n4525), .Z(n4222) );
  OAI21_X1 U4816 ( .B1(n4223), .B2(n4238), .A(n4222), .ZN(U3499) );
  INV_X1 U4817 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4225) );
  MUX2_X1 U4818 ( .A(n4225), .B(n4224), .S(n4525), .Z(n4226) );
  OAI21_X1 U4819 ( .B1(n4227), .B2(n4238), .A(n4226), .ZN(U3497) );
  MUX2_X1 U4820 ( .A(REG0_REG_14__SCAN_IN), .B(n4228), .S(n4525), .Z(U3495) );
  MUX2_X1 U4821 ( .A(REG0_REG_13__SCAN_IN), .B(n4229), .S(n4525), .Z(U3493) );
  INV_X1 U4822 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4231) );
  MUX2_X1 U4823 ( .A(n4231), .B(n4230), .S(n4525), .Z(n4232) );
  OAI21_X1 U4824 ( .B1(n4233), .B2(n4238), .A(n4232), .ZN(U3491) );
  MUX2_X1 U4825 ( .A(REG0_REG_11__SCAN_IN), .B(n4234), .S(n4525), .Z(U3489) );
  INV_X1 U4826 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4236) );
  MUX2_X1 U4827 ( .A(n4236), .B(n4235), .S(n4525), .Z(n4237) );
  OAI21_X1 U4828 ( .B1(n4239), .B2(n4238), .A(n4237), .ZN(U3487) );
  MUX2_X1 U4829 ( .A(DATAI_30_), .B(n4240), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4830 ( .A(DATAI_29_), .B(n2020), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4831 ( .A(DATAI_28_), .B(n4241), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4832 ( .A(n2006), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4833 ( .A(n4243), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U4834 ( .A(n4244), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4835 ( .A(n4245), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4836 ( .A(DATAI_20_), .B(n4246), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4837 ( .A(DATAI_19_), .B(n4247), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4838 ( .A(DATAI_10_), .B(n4309), .S(STATE_REG_SCAN_IN), .Z(U3342)
         );
  MUX2_X1 U4839 ( .A(n4248), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4840 ( .A(DATAI_4_), .B(n4249), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4841 ( .A(n4250), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4842 ( .A(n4251), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  AOI22_X1 U4843 ( .A1(n4253), .A2(n4428), .B1(n4445), .B2(n4252), .ZN(n4254)
         );
  OAI21_X1 U4844 ( .B1(n4445), .B2(n3387), .A(n4254), .ZN(U3260) );
  AOI22_X1 U4845 ( .A1(n4255), .A2(n4428), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4424), .ZN(n4256) );
  OAI21_X1 U4846 ( .B1(n4424), .B2(n4257), .A(n4256), .ZN(U3261) );
  OAI21_X1 U4847 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4259), .A(n4258), .ZN(n4260)
         );
  XNOR2_X1 U4848 ( .A(n4260), .B(n2289), .ZN(n4263) );
  AOI22_X1 U4849 ( .A1(n4395), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4261) );
  OAI21_X1 U4850 ( .B1(n4263), .B2(n4262), .A(n4261), .ZN(U3240) );
  AOI211_X1 U4851 ( .C1(n4267), .C2(n4266), .A(n4265), .B(n4264), .ZN(n4269)
         );
  AOI211_X1 U4852 ( .C1(n4395), .C2(ADDR_REG_6__SCAN_IN), .A(n4269), .B(n4268), 
        .ZN(n4273) );
  OAI211_X1 U4853 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4271), .A(n4341), .B(n4270), 
        .ZN(n4272) );
  OAI211_X1 U4854 ( .C1(n4401), .C2(n2145), .A(n4273), .B(n4272), .ZN(U3246)
         );
  NAND2_X1 U4855 ( .A1(n4275), .A2(n4274), .ZN(n4277) );
  OAI21_X1 U4856 ( .B1(n4278), .B2(n4277), .A(n4397), .ZN(n4276) );
  AOI21_X1 U4857 ( .B1(n4278), .B2(n4277), .A(n4276), .ZN(n4281) );
  INV_X1 U4858 ( .A(n4279), .ZN(n4280) );
  AOI211_X1 U4859 ( .C1(n4395), .C2(ADDR_REG_7__SCAN_IN), .A(n4281), .B(n4280), 
        .ZN(n4286) );
  OAI211_X1 U4860 ( .C1(n4284), .C2(n4283), .A(n4341), .B(n4282), .ZN(n4285)
         );
  OAI211_X1 U4861 ( .C1(n4401), .C2(n4477), .A(n4286), .B(n4285), .ZN(U3247)
         );
  OAI211_X1 U4862 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4288), .A(n4341), .B(n4287), 
        .ZN(n4290) );
  NAND2_X1 U4863 ( .A1(n4290), .A2(n4289), .ZN(n4291) );
  AOI21_X1 U4864 ( .B1(n4395), .B2(ADDR_REG_8__SCAN_IN), .A(n4291), .ZN(n4295)
         );
  OAI211_X1 U4865 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4293), .A(n4397), .B(n4292), 
        .ZN(n4294) );
  OAI211_X1 U4866 ( .C1(n4401), .C2(n4296), .A(n4295), .B(n4294), .ZN(U3248)
         );
  OAI211_X1 U4867 ( .C1(n4299), .C2(n4298), .A(n4397), .B(n4297), .ZN(n4304)
         );
  OAI211_X1 U4868 ( .C1(n4302), .C2(n4301), .A(n4341), .B(n4300), .ZN(n4303)
         );
  OAI211_X1 U4869 ( .C1(n4401), .C2(n4305), .A(n4304), .B(n4303), .ZN(n4306)
         );
  AOI211_X1 U4870 ( .C1(n4395), .C2(ADDR_REG_9__SCAN_IN), .A(n4307), .B(n4306), 
        .ZN(n4308) );
  INV_X1 U4871 ( .A(n4308), .ZN(U3249) );
  OAI211_X1 U4872 ( .C1(n4311), .C2(REG1_REG_10__SCAN_IN), .A(n4397), .B(n4310), .ZN(n4315) );
  OAI211_X1 U4873 ( .C1(n4313), .C2(REG2_REG_10__SCAN_IN), .A(n4341), .B(n4312), .ZN(n4314) );
  OAI211_X1 U4874 ( .C1(n4401), .C2(n2142), .A(n4315), .B(n4314), .ZN(n4316)
         );
  AOI211_X1 U4875 ( .C1(n4395), .C2(ADDR_REG_10__SCAN_IN), .A(n4317), .B(n4316), .ZN(n4318) );
  INV_X1 U4876 ( .A(n4318), .ZN(U3250) );
  OAI211_X1 U4877 ( .C1(n4321), .C2(n4320), .A(n4397), .B(n4319), .ZN(n4326)
         );
  OAI211_X1 U4878 ( .C1(n4324), .C2(n4323), .A(n4341), .B(n4322), .ZN(n4325)
         );
  OAI211_X1 U4879 ( .C1(n4401), .C2(n4327), .A(n4326), .B(n4325), .ZN(n4328)
         );
  AOI211_X1 U4880 ( .C1(n4395), .C2(ADDR_REG_11__SCAN_IN), .A(n4329), .B(n4328), .ZN(n4330) );
  INV_X1 U4881 ( .A(n4330), .ZN(U3251) );
  OAI211_X1 U4882 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4332), .A(n4341), .B(n4331), .ZN(n4334) );
  NAND2_X1 U4883 ( .A1(n4334), .A2(n4333), .ZN(n4335) );
  AOI21_X1 U4884 ( .B1(n4395), .B2(ADDR_REG_12__SCAN_IN), .A(n4335), .ZN(n4339) );
  OAI211_X1 U4885 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4337), .A(n4397), .B(n4336), .ZN(n4338) );
  OAI211_X1 U4886 ( .C1(n4401), .C2(n2144), .A(n4339), .B(n4338), .ZN(U3252)
         );
  AOI21_X1 U4887 ( .B1(n4352), .B2(n4057), .A(n4340), .ZN(n4344) );
  OAI21_X1 U4888 ( .B1(n4344), .B2(n4343), .A(n4341), .ZN(n4342) );
  AOI21_X1 U4889 ( .B1(n4344), .B2(n4343), .A(n4342), .ZN(n4345) );
  AOI211_X1 U4890 ( .C1(n4395), .C2(ADDR_REG_13__SCAN_IN), .A(n4346), .B(n4345), .ZN(n4351) );
  OAI211_X1 U4891 ( .C1(n4349), .C2(n4348), .A(n4397), .B(n4347), .ZN(n4350)
         );
  OAI211_X1 U4892 ( .C1(n4401), .C2(n4352), .A(n4351), .B(n4350), .ZN(U3253)
         );
  INV_X1 U4893 ( .A(n4353), .ZN(n4357) );
  AOI211_X1 U4894 ( .C1(n4037), .C2(n4355), .A(n4354), .B(n4391), .ZN(n4356)
         );
  AOI211_X1 U4895 ( .C1(n4395), .C2(ADDR_REG_14__SCAN_IN), .A(n4357), .B(n4356), .ZN(n4361) );
  OAI211_X1 U4896 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4359), .A(n4397), .B(n4358), .ZN(n4360) );
  OAI211_X1 U4897 ( .C1(n4401), .C2(n4466), .A(n4361), .B(n4360), .ZN(U3254)
         );
  AOI211_X1 U4898 ( .C1(n4364), .C2(n4363), .A(n4362), .B(n4391), .ZN(n4365)
         );
  AOI211_X1 U4899 ( .C1(ADDR_REG_15__SCAN_IN), .C2(n4395), .A(n4366), .B(n4365), .ZN(n4371) );
  OAI211_X1 U4900 ( .C1(n4369), .C2(n4368), .A(n4397), .B(n4367), .ZN(n4370)
         );
  OAI211_X1 U4901 ( .C1(n4401), .C2(n4464), .A(n4371), .B(n4370), .ZN(U3255)
         );
  INV_X1 U4902 ( .A(n4372), .ZN(n4376) );
  AOI221_X1 U4903 ( .B1(n4374), .B2(n4373), .C1(n2451), .C2(n4373), .A(n4391), 
        .ZN(n4375) );
  AOI211_X1 U4904 ( .C1(n4395), .C2(ADDR_REG_16__SCAN_IN), .A(n4376), .B(n4375), .ZN(n4380) );
  OAI221_X1 U4905 ( .B1(n4378), .B2(REG1_REG_16__SCAN_IN), .C1(n4378), .C2(
        n4377), .A(n4397), .ZN(n4379) );
  OAI211_X1 U4906 ( .C1(n4401), .C2(n4462), .A(n4380), .B(n4379), .ZN(U3256)
         );
  AOI221_X1 U4907 ( .B1(n4383), .B2(n4382), .C1(n4381), .C2(n4382), .A(n4391), 
        .ZN(n4384) );
  AOI211_X1 U4908 ( .C1(n4395), .C2(ADDR_REG_17__SCAN_IN), .A(n4385), .B(n4384), .ZN(n4389) );
  OAI221_X1 U4909 ( .B1(n4387), .B2(n2030), .C1(n4387), .C2(n4386), .A(n4397), 
        .ZN(n4388) );
  OAI211_X1 U4910 ( .C1(n4401), .C2(n4390), .A(n4389), .B(n4388), .ZN(U3257)
         );
  OAI211_X1 U4911 ( .C1(n4398), .C2(n2012), .A(n4397), .B(n4396), .ZN(n4399)
         );
  OAI211_X1 U4912 ( .C1(n4401), .C2(n4458), .A(n4400), .B(n4399), .ZN(U3258)
         );
  AOI22_X1 U4913 ( .A1(n4402), .A2(n4442), .B1(REG2_REG_8__SCAN_IN), .B2(n4424), .ZN(n4407) );
  INV_X1 U4914 ( .A(n4403), .ZN(n4404) );
  AOI22_X1 U4915 ( .A1(n4405), .A2(n4443), .B1(n4428), .B2(n4404), .ZN(n4406)
         );
  OAI211_X1 U4916 ( .C1(n4424), .C2(n4408), .A(n4407), .B(n4406), .ZN(U3282)
         );
  INV_X1 U4917 ( .A(n2569), .ZN(n4411) );
  OAI21_X1 U4918 ( .B1(n4411), .B2(n4410), .A(n4409), .ZN(n4423) );
  AOI22_X1 U4919 ( .A1(n2735), .A2(n4414), .B1(n4413), .B2(n4412), .ZN(n4415)
         );
  OAI21_X1 U4920 ( .B1(n4417), .B2(n4416), .A(n4415), .ZN(n4422) );
  OAI21_X1 U4921 ( .B1(n2569), .B2(n4419), .A(n4418), .ZN(n4487) );
  NOR2_X1 U4922 ( .A1(n4487), .A2(n4420), .ZN(n4421) );
  AOI211_X1 U4923 ( .C1(n4436), .C2(n4423), .A(n4422), .B(n4421), .ZN(n4484)
         );
  AOI22_X1 U4924 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4442), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4424), .ZN(n4431) );
  INV_X1 U4925 ( .A(n4487), .ZN(n4429) );
  OAI21_X1 U4926 ( .B1(n4426), .B2(n4434), .A(n4425), .ZN(n4485) );
  INV_X1 U4927 ( .A(n4485), .ZN(n4427) );
  AOI22_X1 U4928 ( .A1(n4429), .A2(n4443), .B1(n4428), .B2(n4427), .ZN(n4430)
         );
  OAI211_X1 U4929 ( .C1(n4424), .C2(n4484), .A(n4431), .B(n4430), .ZN(U3289)
         );
  INV_X1 U4930 ( .A(n4432), .ZN(n4433) );
  NOR2_X1 U4931 ( .A1(n4434), .A2(n4433), .ZN(n4481) );
  INV_X1 U4932 ( .A(n4435), .ZN(n4441) );
  OAI21_X1 U4933 ( .B1(n4437), .B2(n4436), .A(n4482), .ZN(n4438) );
  OAI21_X1 U4934 ( .B1(n4440), .B2(n4439), .A(n4438), .ZN(n4480) );
  AOI21_X1 U4935 ( .B1(n4481), .B2(n4441), .A(n4480), .ZN(n4446) );
  AOI22_X1 U4936 ( .A1(n4443), .A2(n4482), .B1(REG3_REG_0__SCAN_IN), .B2(n4442), .ZN(n4444) );
  OAI221_X1 U4937 ( .B1(n4424), .B2(n4446), .C1(n4445), .C2(n2283), .A(n4444), 
        .ZN(U3290) );
  AND2_X1 U4938 ( .A1(D_REG_31__SCAN_IN), .A2(n4452), .ZN(U3291) );
  AND2_X1 U4939 ( .A1(D_REG_30__SCAN_IN), .A2(n4452), .ZN(U3292) );
  AND2_X1 U4940 ( .A1(D_REG_29__SCAN_IN), .A2(n4452), .ZN(U3293) );
  NOR2_X1 U4941 ( .A1(n4454), .A2(n4447), .ZN(U3294) );
  AND2_X1 U4942 ( .A1(D_REG_27__SCAN_IN), .A2(n4452), .ZN(U3295) );
  AND2_X1 U4943 ( .A1(D_REG_26__SCAN_IN), .A2(n4452), .ZN(U3296) );
  AND2_X1 U4944 ( .A1(D_REG_25__SCAN_IN), .A2(n4452), .ZN(U3297) );
  AND2_X1 U4945 ( .A1(D_REG_24__SCAN_IN), .A2(n4452), .ZN(U3298) );
  AND2_X1 U4946 ( .A1(D_REG_23__SCAN_IN), .A2(n4452), .ZN(U3299) );
  AND2_X1 U4947 ( .A1(D_REG_22__SCAN_IN), .A2(n4452), .ZN(U3300) );
  AND2_X1 U4948 ( .A1(D_REG_21__SCAN_IN), .A2(n4452), .ZN(U3301) );
  AND2_X1 U4949 ( .A1(D_REG_20__SCAN_IN), .A2(n4452), .ZN(U3302) );
  NOR2_X1 U4950 ( .A1(n4454), .A2(n4448), .ZN(U3303) );
  AND2_X1 U4951 ( .A1(D_REG_18__SCAN_IN), .A2(n4452), .ZN(U3304) );
  AND2_X1 U4952 ( .A1(D_REG_17__SCAN_IN), .A2(n4452), .ZN(U3305) );
  AND2_X1 U4953 ( .A1(D_REG_16__SCAN_IN), .A2(n4452), .ZN(U3306) );
  AND2_X1 U4954 ( .A1(D_REG_15__SCAN_IN), .A2(n4452), .ZN(U3307) );
  AND2_X1 U4955 ( .A1(D_REG_14__SCAN_IN), .A2(n4452), .ZN(U3308) );
  AND2_X1 U4956 ( .A1(D_REG_13__SCAN_IN), .A2(n4452), .ZN(U3309) );
  AND2_X1 U4957 ( .A1(D_REG_12__SCAN_IN), .A2(n4452), .ZN(U3310) );
  NOR2_X1 U4958 ( .A1(n4454), .A2(n4449), .ZN(U3311) );
  AND2_X1 U4959 ( .A1(D_REG_10__SCAN_IN), .A2(n4452), .ZN(U3312) );
  AND2_X1 U4960 ( .A1(D_REG_9__SCAN_IN), .A2(n4452), .ZN(U3313) );
  AND2_X1 U4961 ( .A1(D_REG_8__SCAN_IN), .A2(n4452), .ZN(U3314) );
  NOR2_X1 U4962 ( .A1(n4454), .A2(n4450), .ZN(U3315) );
  AND2_X1 U4963 ( .A1(D_REG_6__SCAN_IN), .A2(n4452), .ZN(U3316) );
  NOR2_X1 U4964 ( .A1(n4454), .A2(n4451), .ZN(U3317) );
  AND2_X1 U4965 ( .A1(D_REG_4__SCAN_IN), .A2(n4452), .ZN(U3318) );
  AND2_X1 U4966 ( .A1(D_REG_3__SCAN_IN), .A2(n4452), .ZN(U3319) );
  NOR2_X1 U4967 ( .A1(n4454), .A2(n4453), .ZN(U3320) );
  OAI21_X1 U4968 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4455), .ZN(
        n4456) );
  INV_X1 U4969 ( .A(n4456), .ZN(U3329) );
  INV_X1 U4970 ( .A(DATAI_18_), .ZN(n4457) );
  AOI22_X1 U4971 ( .A1(STATE_REG_SCAN_IN), .A2(n4458), .B1(n4457), .B2(U3149), 
        .ZN(U3334) );
  OAI22_X1 U4972 ( .A1(U3149), .A2(n4459), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4460) );
  INV_X1 U4973 ( .A(n4460), .ZN(U3335) );
  AOI22_X1 U4974 ( .A1(STATE_REG_SCAN_IN), .A2(n4462), .B1(n4461), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U4975 ( .A(DATAI_15_), .ZN(n4463) );
  AOI22_X1 U4976 ( .A1(STATE_REG_SCAN_IN), .A2(n4464), .B1(n4463), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U4977 ( .A1(STATE_REG_SCAN_IN), .A2(n4466), .B1(n4465), .B2(U3149), 
        .ZN(U3338) );
  OAI22_X1 U4978 ( .A1(U3149), .A2(n4467), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4468) );
  INV_X1 U4979 ( .A(n4468), .ZN(U3339) );
  INV_X1 U4980 ( .A(DATAI_12_), .ZN(n4469) );
  AOI22_X1 U4981 ( .A1(STATE_REG_SCAN_IN), .A2(n2144), .B1(n4469), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U4982 ( .A1(U3149), .A2(n4470), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4471) );
  INV_X1 U4983 ( .A(n4471), .ZN(U3341) );
  OAI22_X1 U4984 ( .A1(U3149), .A2(n4472), .B1(DATAI_9_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4473) );
  INV_X1 U4985 ( .A(n4473), .ZN(U3343) );
  OAI22_X1 U4986 ( .A1(U3149), .A2(n4474), .B1(DATAI_8_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4475) );
  INV_X1 U4987 ( .A(n4475), .ZN(U3344) );
  INV_X1 U4988 ( .A(DATAI_7_), .ZN(n4476) );
  AOI22_X1 U4989 ( .A1(STATE_REG_SCAN_IN), .A2(n4477), .B1(n4476), .B2(U3149), 
        .ZN(U3345) );
  AOI22_X1 U4990 ( .A1(STATE_REG_SCAN_IN), .A2(n2145), .B1(n4478), .B2(U3149), 
        .ZN(U3346) );
  OAI22_X1 U4991 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4479) );
  INV_X1 U4992 ( .A(n4479), .ZN(U3352) );
  AOI211_X1 U4993 ( .C1(n4504), .C2(n4482), .A(n4481), .B(n4480), .ZN(n4527)
         );
  INV_X1 U4994 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4483) );
  AOI22_X1 U4995 ( .A1(n4525), .A2(n4527), .B1(n4483), .B2(n4523), .ZN(U3467)
         );
  INV_X1 U4996 ( .A(n4484), .ZN(n4489) );
  OAI22_X1 U4997 ( .A1(n4487), .A2(n4486), .B1(n4519), .B2(n4485), .ZN(n4488)
         );
  NOR2_X1 U4998 ( .A1(n4489), .A2(n4488), .ZN(n4529) );
  AOI22_X1 U4999 ( .A1(n4525), .A2(n4529), .B1(n2271), .B2(n4523), .ZN(U3469)
         );
  NOR3_X1 U5000 ( .A1(n4491), .A2(n4490), .A3(n4519), .ZN(n4494) );
  INV_X1 U5001 ( .A(n4492), .ZN(n4493) );
  AOI211_X1 U5002 ( .C1(n4504), .C2(n4495), .A(n4494), .B(n4493), .ZN(n4531)
         );
  AOI22_X1 U5003 ( .A1(n4525), .A2(n4531), .B1(n2294), .B2(n4523), .ZN(U3471)
         );
  NOR2_X1 U5004 ( .A1(n4496), .A2(n4519), .ZN(n4497) );
  AOI21_X1 U5005 ( .B1(n4498), .B2(n4504), .A(n4497), .ZN(n4499) );
  AOI22_X1 U5006 ( .A1(n4525), .A2(n4533), .B1(n2303), .B2(n4523), .ZN(U3473)
         );
  INV_X1 U5007 ( .A(n4501), .ZN(n4503) );
  AOI211_X1 U5008 ( .C1(n4505), .C2(n4504), .A(n4503), .B(n4502), .ZN(n4534)
         );
  INV_X1 U5009 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U5010 ( .A1(n4525), .A2(n4534), .B1(n4506), .B2(n4523), .ZN(U3475)
         );
  NOR2_X1 U5011 ( .A1(n4508), .A2(n4507), .ZN(n4510) );
  AOI211_X1 U5012 ( .C1(n4512), .C2(n4511), .A(n4510), .B(n4509), .ZN(n4535)
         );
  AOI22_X1 U5013 ( .A1(n4525), .A2(n4535), .B1(n2324), .B2(n4523), .ZN(U3477)
         );
  AOI211_X1 U5014 ( .C1(n4515), .C2(n4522), .A(n4514), .B(n4513), .ZN(n4537)
         );
  INV_X1 U5015 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4516) );
  AOI22_X1 U5016 ( .A1(n4525), .A2(n4537), .B1(n4516), .B2(n4523), .ZN(U3481)
         );
  OAI21_X1 U5017 ( .B1(n4519), .B2(n4518), .A(n4517), .ZN(n4520) );
  AOI21_X1 U5018 ( .B1(n4522), .B2(n4521), .A(n4520), .ZN(n4539) );
  AOI22_X1 U5019 ( .A1(n4525), .A2(n4539), .B1(n4524), .B2(n4523), .ZN(U3485)
         );
  AOI22_X1 U5020 ( .A1(n4540), .A2(n4527), .B1(n4526), .B2(n4538), .ZN(U3518)
         );
  AOI22_X1 U5021 ( .A1(n4540), .A2(n4529), .B1(n4528), .B2(n4538), .ZN(U3519)
         );
  AOI22_X1 U5022 ( .A1(n4540), .A2(n4531), .B1(n4530), .B2(n4538), .ZN(U3520)
         );
  AOI22_X1 U5023 ( .A1(n4540), .A2(n4533), .B1(n4532), .B2(n4538), .ZN(U3521)
         );
  AOI22_X1 U5024 ( .A1(n4540), .A2(n4534), .B1(n2314), .B2(n4538), .ZN(U3522)
         );
  AOI22_X1 U5025 ( .A1(n4540), .A2(n4535), .B1(n2695), .B2(n4538), .ZN(U3523)
         );
  AOI22_X1 U5026 ( .A1(n4540), .A2(n4537), .B1(n4536), .B2(n4538), .ZN(U3525)
         );
  AOI22_X1 U5027 ( .A1(n4540), .A2(n4539), .B1(n2367), .B2(n4538), .ZN(U3527)
         );
endmodule

