

module b20_C_AntiSAT_k_128_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4335, n4336, n4337, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259;

  NAND2_X2 U4841 ( .A1(n5131), .A2(n5130), .ZN(n6493) );
  AND2_X2 U4842 ( .A1(n9434), .A2(n5105), .ZN(n5151) );
  BUF_X1 U4843 ( .A(n7800), .Z(n4336) );
  AND2_X1 U4844 ( .A1(n6296), .A2(n8229), .ZN(n8219) );
  NAND2_X1 U4845 ( .A1(n7796), .A2(n4992), .ZN(n5173) );
  INV_X1 U4846 ( .A(n8894), .ZN(n5616) );
  INV_X1 U4847 ( .A(n4342), .ZN(n5500) );
  INV_X1 U4848 ( .A(n8219), .ZN(n8206) );
  INV_X1 U4849 ( .A(n6095), .ZN(n5886) );
  INV_X1 U4850 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4603) );
  INV_X1 U4852 ( .A(n5126), .ZN(n6478) );
  AND2_X1 U4853 ( .A1(n5749), .A2(n7739), .ZN(n5728) );
  INV_X1 U4854 ( .A(n5842), .ZN(n8025) );
  NAND2_X1 U4855 ( .A1(n4706), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U4856 ( .A1(n5711), .A2(n4565), .ZN(n6531) );
  AOI21_X1 U4857 ( .B1(n5468), .B2(n4965), .A(n5467), .ZN(n8952) );
  INV_X1 U4858 ( .A(n8003), .ZN(n9747) );
  XNOR2_X1 U4859 ( .A(n5338), .B(n5337), .ZN(n6577) );
  AND2_X2 U4860 ( .A1(n4743), .A2(n4350), .ZN(n4567) );
  AND4_X2 U4861 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), .ZN(n6303)
         );
  BUF_X4 U4862 ( .A(n5521), .Z(n4335) );
  OAI21_X2 U4863 ( .B1(n5359), .B2(n4878), .A(n4876), .ZN(n5401) );
  NAND2_X2 U4864 ( .A1(n5355), .A2(n5026), .ZN(n5359) );
  XNOR2_X2 U4865 ( .A(n4590), .B(P2_IR_REG_1__SCAN_IN), .ZN(n4592) );
  XNOR2_X2 U4866 ( .A(n4822), .B(n5800), .ZN(n6711) );
  CLKBUF_X1 U4867 ( .A(n7800), .Z(n4337) );
  NAND2_X4 U4868 ( .A1(n4507), .A2(n6299), .ZN(n6412) );
  XNOR2_X2 U4869 ( .A(n5767), .B(n8861), .ZN(n7666) );
  OAI21_X2 U4870 ( .B1(n5424), .B2(n4853), .A(n4851), .ZN(n5514) );
  AOI22_X4 U4871 ( .A1(n9240), .A2(n9242), .B1(n9045), .B2(n9381), .ZN(n9225)
         );
  OAI22_X2 U4872 ( .A1(n6466), .A2(n6465), .B1(n8917), .B2(n9265), .ZN(n9240)
         );
  XNOR2_X2 U4873 ( .A(n5301), .B(n5302), .ZN(n6555) );
  AND2_X4 U4874 ( .A1(n5728), .A2(n6531), .ZN(n5159) );
  XNOR2_X2 U4875 ( .A(n5769), .B(n5768), .ZN(n7654) );
  NAND2_X1 U4876 ( .A1(n7819), .A2(n7815), .ZN(n7954) );
  OR2_X1 U4877 ( .A1(n7303), .A2(n4746), .ZN(n4745) );
  INV_X2 U4879 ( .A(n9752), .ZN(n9754) );
  INV_X1 U4880 ( .A(n9786), .ZN(n7073) );
  INV_X1 U4881 ( .A(n9055), .ZN(n7165) );
  NAND2_X2 U4882 ( .A1(n8894), .A2(n5618), .ZN(n5150) );
  INV_X1 U4883 ( .A(n8357), .ZN(n4615) );
  NAND4_X1 U4884 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(n9932)
         );
  BUF_X2 U4885 ( .A(n5173), .Z(n4342) );
  NAND2_X1 U4886 ( .A1(n5106), .A2(n5109), .ZN(n7800) );
  BUF_X1 U4887 ( .A(n5832), .Z(n4344) );
  BUF_X2 U4888 ( .A(n5828), .Z(n5816) );
  CLKBUF_X2 U4889 ( .A(n6711), .Z(n9912) );
  NAND2_X1 U4890 ( .A1(n4835), .A2(n4833), .ZN(n4997) );
  AND4_X1 U4891 ( .A1(n4566), .A2(n5070), .A3(n5056), .A4(n5074), .ZN(n5057)
         );
  INV_X1 U4892 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5800) );
  NOR2_X1 U4893 ( .A1(n8977), .A2(n4400), .ZN(n8874) );
  AND2_X1 U4894 ( .A1(n6169), .A2(n9928), .ZN(n4639) );
  AND2_X1 U4895 ( .A1(n7802), .A2(n8004), .ZN(n8007) );
  OAI21_X1 U4896 ( .B1(n6255), .B2(n6254), .A(n6253), .ZN(n8026) );
  AND2_X1 U4897 ( .A1(n7979), .A2(n7978), .ZN(n7998) );
  NAND2_X1 U4898 ( .A1(n7931), .A2(n7929), .ZN(n7972) );
  NAND2_X1 U4899 ( .A1(n8969), .A2(n8970), .ZN(n8968) );
  OR2_X1 U4900 ( .A1(n9341), .A2(n6483), .ZN(n7931) );
  NAND2_X1 U4901 ( .A1(n7729), .A2(n7927), .ZN(n9145) );
  NOR2_X1 U4902 ( .A1(n8489), .A2(n8488), .ZN(n8491) );
  XNOR2_X1 U4903 ( .A(n7794), .B(n7793), .ZN(n9426) );
  INV_X1 U4904 ( .A(n7919), .ZN(n7729) );
  NAND2_X1 U4905 ( .A1(n6476), .A2(n6475), .ZN(n9341) );
  AND2_X1 U4906 ( .A1(n9139), .A2(n9038), .ZN(n7919) );
  OAI21_X1 U4907 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n7790) );
  XNOR2_X1 U4908 ( .A(n7659), .B(n7658), .ZN(n7662) );
  INV_X1 U4909 ( .A(n4796), .ZN(n4795) );
  NAND2_X1 U4910 ( .A1(n6116), .A2(n6115), .ZN(n8798) );
  NAND2_X1 U4911 ( .A1(n8330), .A2(n4963), .ZN(n7682) );
  XNOR2_X1 U4912 ( .A(n6257), .B(n6256), .ZN(n8020) );
  NAND2_X1 U4913 ( .A1(n5657), .A2(n5656), .ZN(n9356) );
  NOR2_X1 U4914 ( .A1(n5574), .A2(n4803), .ZN(n4799) );
  XNOR2_X1 U4915 ( .A(n5655), .B(n5654), .ZN(n7614) );
  XNOR2_X1 U4916 ( .A(n6134), .B(n6133), .ZN(n7624) );
  AND2_X1 U4917 ( .A1(n7911), .A2(n7910), .ZN(n9199) );
  NAND2_X1 U4918 ( .A1(n8235), .A2(n8234), .ZN(n8233) );
  AOI21_X1 U4919 ( .B1(n5673), .B2(n5672), .A(n5671), .ZN(n6134) );
  NAND3_X1 U4920 ( .A1(n4777), .A2(n4776), .A3(n4372), .ZN(n7515) );
  NAND2_X1 U4921 ( .A1(n7504), .A2(n4427), .ZN(n7568) );
  NAND2_X1 U4922 ( .A1(n5583), .A2(n5582), .ZN(n9371) );
  OR2_X1 U4923 ( .A1(n8391), .A2(n8392), .ZN(n4720) );
  NAND2_X1 U4924 ( .A1(n7506), .A2(n7505), .ZN(n7504) );
  OAI21_X1 U4925 ( .B1(n7535), .B2(n4692), .A(n4694), .ZN(n6224) );
  AND2_X1 U4926 ( .A1(n7763), .A2(n7761), .ZN(n9299) );
  NAND2_X1 U4927 ( .A1(n4778), .A2(n4781), .ZN(n4776) );
  AND2_X1 U4928 ( .A1(n9697), .A2(n7748), .ZN(n9680) );
  XNOR2_X1 U4929 ( .A(n5599), .B(n5598), .ZN(n6078) );
  NAND2_X1 U4930 ( .A1(n5540), .A2(n5539), .ZN(n9381) );
  OAI21_X1 U4931 ( .B1(n4781), .B2(n4370), .A(n4780), .ZN(n4779) );
  OR2_X1 U4932 ( .A1(n8673), .A2(n8658), .ZN(n8166) );
  OR2_X1 U4933 ( .A1(n8769), .A2(n8636), .ZN(n8168) );
  NAND2_X1 U4934 ( .A1(n6027), .A2(n6026), .ZN(n8673) );
  NAND2_X1 U4935 ( .A1(n6041), .A2(n6040), .ZN(n8769) );
  NAND2_X1 U4936 ( .A1(n5936), .A2(n5935), .ZN(n7538) );
  NAND2_X1 U4937 ( .A1(n5472), .A2(n5471), .ZN(n9323) );
  NAND2_X1 U4938 ( .A1(n5431), .A2(n5430), .ZN(n9512) );
  NAND2_X1 U4939 ( .A1(n5992), .A2(n5991), .ZN(n8848) );
  NAND2_X1 U4940 ( .A1(n4849), .A2(n4847), .ZN(n5535) );
  NAND2_X1 U4941 ( .A1(n5445), .A2(n5444), .ZN(n9402) );
  AND2_X1 U4942 ( .A1(n7861), .A2(n7874), .ZN(n7960) );
  NAND2_X1 U4943 ( .A1(n7521), .A2(n7558), .ZN(n7874) );
  AND2_X1 U4944 ( .A1(n7852), .A2(n7748), .ZN(n9699) );
  NAND2_X1 U4945 ( .A1(n5963), .A2(n5962), .ZN(n8855) );
  NAND2_X1 U4946 ( .A1(n5039), .A2(n5040), .ZN(n5424) );
  AND2_X1 U4947 ( .A1(n5410), .A2(n5409), .ZN(n9839) );
  NAND3_X1 U4948 ( .A1(n4751), .A2(n5210), .A3(n5230), .ZN(n6897) );
  AND2_X1 U4949 ( .A1(n7219), .A2(n7834), .ZN(n7832) );
  NAND2_X1 U4950 ( .A1(n5364), .A2(n5363), .ZN(n9818) );
  NAND2_X1 U4951 ( .A1(n6849), .A2(n6850), .ZN(n4751) );
  AND2_X1 U4952 ( .A1(n5884), .A2(n5883), .ZN(n7244) );
  INV_X1 U4953 ( .A(n6519), .ZN(n9721) );
  NAND2_X1 U4954 ( .A1(n5359), .A2(n5027), .ZN(n5338) );
  NAND2_X1 U4955 ( .A1(n5274), .A2(n4561), .ZN(n6519) );
  INV_X1 U4956 ( .A(n4562), .ZN(n4561) );
  NAND2_X1 U4957 ( .A1(n5272), .A2(n5273), .ZN(n6542) );
  AND2_X1 U4958 ( .A1(n8091), .A2(n8097), .ZN(n8038) );
  NAND2_X1 U4959 ( .A1(n5271), .A2(n5270), .ZN(n5273) );
  AND3_X2 U4960 ( .A1(n6248), .A2(n6835), .A3(n6836), .ZN(n10008) );
  AND3_X2 U4961 ( .A1(n5169), .A2(n4892), .A3(n5170), .ZN(n6851) );
  NAND4_X1 U4962 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n9052)
         );
  INV_X2 U4964 ( .A(n5618), .ZN(n8896) );
  OAI211_X1 U4965 ( .C1(n7796), .C2(n9537), .A(n5143), .B(n5142), .ZN(n6429)
         );
  INV_X2 U4966 ( .A(n6300), .ZN(n4339) );
  OR2_X2 U4967 ( .A1(n6489), .A2(n5097), .ZN(n5618) );
  OR2_X1 U4968 ( .A1(n5404), .A2(n6549), .ZN(n5142) );
  NAND3_X1 U4969 ( .A1(n4367), .A2(n5801), .A3(n4614), .ZN(n9948) );
  NOR2_X1 U4970 ( .A1(n4844), .A2(n4840), .ZN(n4839) );
  AOI21_X1 U4971 ( .B1(n4843), .B2(n4845), .A(n4402), .ZN(n4842) );
  INV_X2 U4972 ( .A(n4337), .ZN(n4345) );
  INV_X2 U4973 ( .A(n4336), .ZN(n4340) );
  NAND2_X1 U4974 ( .A1(n6154), .A2(n6153), .ZN(n7201) );
  OR2_X1 U4975 ( .A1(n5816), .A2(n5793), .ZN(n5796) );
  CLKBUF_X1 U4976 ( .A(n5790), .Z(n6028) );
  AND2_X1 U4977 ( .A1(n5016), .A2(n5015), .ZN(n5286) );
  NAND2_X1 U4978 ( .A1(n5094), .A2(n4563), .ZN(n8003) );
  NOR2_X1 U4979 ( .A1(n5302), .A2(n4846), .ZN(n4845) );
  XNOR2_X1 U4980 ( .A(n6179), .B(n6178), .ZN(n6189) );
  INV_X2 U4981 ( .A(n8530), .ZN(n8503) );
  XNOR2_X1 U4982 ( .A(n6038), .B(n6037), .ZN(n8539) );
  XNOR2_X1 U4983 ( .A(n4707), .B(P1_IR_REG_27__SCAN_IN), .ZN(n7626) );
  INV_X1 U4984 ( .A(n5720), .ZN(n7739) );
  XNOR2_X1 U4985 ( .A(n5777), .B(n4954), .ZN(n6165) );
  NAND2_X1 U4986 ( .A1(n5064), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5083) );
  NAND2_X2 U4987 ( .A1(n7795), .A2(P2_U3151), .ZN(n8019) );
  OR2_X1 U4988 ( .A1(n5766), .A2(n4603), .ZN(n6205) );
  AND2_X1 U4989 ( .A1(n5898), .A2(n4952), .ZN(n5766) );
  INV_X1 U4990 ( .A(n4997), .ZN(n4992) );
  NOR2_X1 U4991 ( .A1(n4742), .A2(n5058), .ZN(n5081) );
  NAND2_X1 U4992 ( .A1(n5823), .A2(n5822), .ZN(n6799) );
  CLKBUF_X3 U4993 ( .A(n4997), .Z(n4346) );
  OR2_X1 U4994 ( .A1(n5764), .A2(n5763), .ZN(n4961) );
  AND2_X1 U4995 ( .A1(n5051), .A2(n4917), .ZN(n4350) );
  AND2_X1 U4996 ( .A1(n4756), .A2(n4754), .ZN(n4740) );
  AND3_X1 U4997 ( .A1(n5132), .A2(n5050), .A3(n5054), .ZN(n4743) );
  INV_X1 U4998 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5713) );
  INV_X1 U4999 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5091) );
  INV_X1 U5000 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5073) );
  INV_X1 U5001 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5070) );
  INV_X4 U5002 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U5003 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4756) );
  NOR2_X1 U5004 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4754) );
  INV_X1 U5005 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4834) );
  NOR2_X1 U5006 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4753) );
  NOR2_X1 U5007 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4755) );
  INV_X4 U5008 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5009 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5799) );
  INV_X1 U5010 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5756) );
  INV_X1 U5011 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5838) );
  NOR2_X1 U5012 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4464) );
  INV_X1 U5013 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6021) );
  NOR2_X1 U5014 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6016) );
  NOR2_X1 U5015 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5760) );
  NOR2_X1 U5016 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5761) );
  OAI21_X1 U5017 ( .B1(n8913), .B2(n4799), .A(n4795), .ZN(n5597) );
  AOI21_X2 U5018 ( .B1(n6518), .B2(n9702), .A(n6517), .ZN(n9343) );
  NOR2_X1 U5019 ( .A1(n9202), .A2(n6510), .ZN(n9191) );
  OAI21_X1 U5020 ( .B1(n9202), .B2(n4712), .A(n4711), .ZN(n9177) );
  AND2_X2 U5021 ( .A1(n9434), .A2(n5109), .ZN(n5521) );
  OAI22_X2 U5022 ( .A1(n9727), .A2(n9726), .B1(n9740), .B2(n6493), .ZN(n6780)
         );
  BUF_X2 U5023 ( .A(n5173), .Z(n4341) );
  NAND2_X2 U5024 ( .A1(n6165), .A2(n6166), .ZN(n5827) );
  OAI21_X2 U5025 ( .B1(n7639), .B2(n6455), .A(n6456), .ZN(n7627) );
  OAI21_X1 U5026 ( .B1(n9429), .B2(n5100), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5101) );
  XNOR2_X2 U5027 ( .A(n6484), .B(n7972), .ZN(n9344) );
  OAI21_X2 U5028 ( .B1(n9139), .B2(n6516), .A(n9137), .ZN(n6484) );
  NAND2_X1 U5029 ( .A1(n5770), .A2(n7666), .ZN(n5832) );
  OAI22_X2 U5030 ( .A1(n7538), .A2(n5948), .B1(n8349), .B2(n7547), .ZN(n7598)
         );
  AOI22_X2 U5031 ( .A1(n9272), .A2(n6464), .B1(n8972), .B2(n9392), .ZN(n9257)
         );
  AOI21_X2 U5032 ( .B1(n9291), .B2(n6463), .A(n6462), .ZN(n9272) );
  NAND2_X2 U5033 ( .A1(n6454), .A2(n6453), .ZN(n7639) );
  AND2_X2 U5034 ( .A1(n5896), .A2(n5757), .ZN(n5898) );
  NOR2_X2 U5035 ( .A1(n4463), .A2(n4460), .ZN(n5896) );
  OAI21_X2 U5036 ( .B1(n7454), .B2(n5923), .A(n5922), .ZN(n7336) );
  OAI22_X2 U5037 ( .A1(n7266), .A2(n5912), .B1(n8352), .B2(n9980), .ZN(n7454)
         );
  INV_X1 U5038 ( .A(n5016), .ZN(n4846) );
  AND2_X1 U5039 ( .A1(n6298), .A2(n6297), .ZN(n6299) );
  NAND2_X1 U5040 ( .A1(n6295), .A2(n6294), .ZN(n4507) );
  NOR2_X1 U5041 ( .A1(n7201), .A2(n6296), .ZN(n6294) );
  NAND2_X1 U5042 ( .A1(n9927), .A2(n5862), .ZN(n4642) );
  NAND2_X1 U5043 ( .A1(n5096), .A2(n8003), .ZN(n5727) );
  INV_X1 U5044 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U5045 ( .A1(n4377), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U5046 ( .A1(n8001), .A2(n5749), .ZN(n4528) );
  INV_X1 U5047 ( .A(n7319), .ZN(n5096) );
  NAND2_X1 U5048 ( .A1(n4458), .A2(n4457), .ZN(n8089) );
  NAND2_X1 U5049 ( .A1(n8127), .A2(n4448), .ZN(n8124) );
  NAND2_X1 U5050 ( .A1(n7875), .A2(n7874), .ZN(n4548) );
  NAND2_X1 U5051 ( .A1(n8192), .A2(n8206), .ZN(n4456) );
  NAND2_X1 U5052 ( .A1(n8191), .A2(n8219), .ZN(n4454) );
  AOI21_X1 U5053 ( .B1(n8209), .B2(n8208), .A(n8207), .ZN(n8214) );
  NOR2_X1 U5054 ( .A1(n4857), .A2(n5494), .ZN(n4855) );
  INV_X1 U5055 ( .A(n5491), .ZN(n5494) );
  NAND2_X1 U5056 ( .A1(n5045), .A2(n5044), .ZN(n5048) );
  NOR2_X1 U5057 ( .A1(n4889), .A2(n4887), .ZN(n4886) );
  NAND2_X1 U5058 ( .A1(n5403), .A2(n4890), .ZN(n4888) );
  AND2_X1 U5059 ( .A1(n5035), .A2(n4891), .ZN(n4890) );
  NAND2_X1 U5060 ( .A1(n5114), .A2(SI_14_), .ZN(n4891) );
  NOR2_X1 U5061 ( .A1(n7042), .A2(n4829), .ZN(n7045) );
  OR2_X1 U5062 ( .A1(n7301), .A2(n7300), .ZN(n7302) );
  INV_X1 U5063 ( .A(n7443), .ZN(n4748) );
  NOR2_X1 U5064 ( .A1(n6081), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4570) );
  INV_X1 U5065 ( .A(n5812), .ZN(n4629) );
  NAND2_X1 U5066 ( .A1(n4628), .A2(n5812), .ZN(n4627) );
  INV_X1 U5067 ( .A(n5803), .ZN(n4628) );
  NAND2_X1 U5068 ( .A1(n6303), .A2(n6300), .ZN(n8081) );
  OR2_X1 U5069 ( .A1(n8803), .A2(n8285), .ZN(n6232) );
  OR2_X1 U5070 ( .A1(n4621), .A2(n4620), .ZN(n4619) );
  OR2_X1 U5071 ( .A1(n8848), .A2(n8334), .ZN(n8153) );
  XNOR2_X1 U5072 ( .A(n5779), .B(n5778), .ZN(n6166) );
  NAND2_X1 U5073 ( .A1(n6183), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5779) );
  NOR2_X1 U5074 ( .A1(n4357), .A2(n7418), .ZN(n4784) );
  OR2_X1 U5075 ( .A1(n5336), .A2(n7418), .ZN(n4785) );
  OR2_X1 U5076 ( .A1(n4964), .A2(n5645), .ZN(n4763) );
  INV_X1 U5077 ( .A(n9171), .ZN(n4896) );
  NAND2_X1 U5078 ( .A1(n9371), .A2(n9043), .ZN(n4929) );
  NAND2_X1 U5079 ( .A1(n4380), .A2(n5057), .ZN(n5058) );
  NAND2_X1 U5080 ( .A1(n5029), .A2(SI_12_), .ZN(n5030) );
  NOR2_X1 U5081 ( .A1(n5337), .A2(n4884), .ZN(n4883) );
  INV_X1 U5082 ( .A(n5027), .ZN(n4884) );
  XNOR2_X1 U5083 ( .A(n5020), .B(SI_9_), .ZN(n5317) );
  INV_X1 U5084 ( .A(n5286), .ZN(n4843) );
  INV_X1 U5085 ( .A(n4845), .ZN(n4844) );
  INV_X1 U5086 ( .A(n5816), .ZN(n6160) );
  NAND2_X1 U5087 ( .A1(n4574), .A2(n4573), .ZN(n5942) );
  INV_X1 U5088 ( .A(n6028), .ZN(n6046) );
  OAI21_X1 U5089 ( .B1(n7302), .B2(n7373), .A(n7358), .ZN(n7303) );
  INV_X1 U5090 ( .A(n8361), .ZN(n4651) );
  NOR2_X1 U5091 ( .A1(n8433), .A2(n8419), .ZN(n8456) );
  OAI21_X1 U5092 ( .B1(n8508), .B2(n8507), .A(n9913), .ZN(n4655) );
  AND2_X1 U5093 ( .A1(n4385), .A2(n6011), .ZN(n4626) );
  OR2_X1 U5094 ( .A1(n6052), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U5095 ( .A1(n5879), .A2(n5878), .ZN(n7239) );
  AND2_X1 U5096 ( .A1(n4389), .A2(n5863), .ZN(n4641) );
  NAND2_X1 U5097 ( .A1(n6218), .A2(n8037), .ZN(n6959) );
  OR2_X1 U5098 ( .A1(n7547), .A2(n7569), .ZN(n8133) );
  INV_X1 U5099 ( .A(n5824), .ZN(n6039) );
  NAND2_X1 U5100 ( .A1(n5776), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5777) );
  AND2_X1 U5101 ( .A1(n5898), .A2(n4348), .ZN(n4643) );
  NAND2_X1 U5102 ( .A1(n4599), .A2(n4598), .ZN(n6152) );
  AOI21_X1 U5103 ( .B1(n4601), .B2(n4603), .A(n4603), .ZN(n4599) );
  NAND2_X1 U5104 ( .A1(n6024), .A2(n4601), .ZN(n4598) );
  NOR2_X1 U5105 ( .A1(n5723), .A2(n5728), .ZN(n5112) );
  INV_X1 U5106 ( .A(n8962), .ZN(n4766) );
  OR2_X1 U5107 ( .A1(n9332), .A2(n9125), .ZN(n8004) );
  NAND2_X1 U5108 ( .A1(n4567), .A2(n5053), .ZN(n5442) );
  AND2_X1 U5109 ( .A1(n5600), .A2(n5581), .ZN(n5598) );
  INV_X1 U5110 ( .A(n5827), .ZN(n6535) );
  INV_X1 U5111 ( .A(n6380), .ZN(n6383) );
  INV_X1 U5112 ( .A(n8222), .ZN(n4872) );
  NAND2_X1 U5113 ( .A1(n4596), .A2(n8221), .ZN(n4595) );
  NOR2_X1 U5114 ( .A1(n8468), .A2(n10071), .ZN(n8488) );
  NAND2_X1 U5115 ( .A1(n4523), .A2(n4526), .ZN(n4522) );
  NOR2_X1 U5116 ( .A1(n8015), .A2(n5749), .ZN(n4526) );
  NAND2_X1 U5117 ( .A1(n4375), .A2(n7998), .ZN(n4523) );
  INV_X1 U5118 ( .A(n4525), .ZN(n4524) );
  OAI21_X1 U5119 ( .B1(n4527), .B2(n8010), .A(n5732), .ZN(n4525) );
  OAI211_X1 U5120 ( .C1(n4447), .C2(n4452), .A(n4451), .B(n4446), .ZN(n8127)
         );
  NAND2_X1 U5121 ( .A1(n8122), .A2(n8206), .ZN(n4446) );
  OAI21_X1 U5122 ( .B1(n4353), .B2(n4399), .A(n8145), .ZN(n4610) );
  NAND2_X1 U5123 ( .A1(n4548), .A2(n4547), .ZN(n4546) );
  INV_X1 U5124 ( .A(n7877), .ZN(n4552) );
  NAND2_X1 U5125 ( .A1(n7878), .A2(n7879), .ZN(n4544) );
  INV_X1 U5126 ( .A(n7901), .ZN(n4560) );
  OAI21_X1 U5127 ( .B1(n7906), .B2(n7905), .A(n4557), .ZN(n4556) );
  AND2_X1 U5128 ( .A1(n9224), .A2(n4361), .ZN(n4557) );
  INV_X1 U5129 ( .A(n5425), .ZN(n5041) );
  NAND2_X1 U5130 ( .A1(n4453), .A2(n4604), .ZN(n8209) );
  AND2_X1 U5131 ( .A1(n4605), .A2(n8205), .ZN(n4604) );
  NAND2_X1 U5132 ( .A1(n4406), .A2(n8210), .ZN(n4582) );
  MUX2_X1 U5133 ( .A(n8212), .B(n8211), .S(n8219), .Z(n8213) );
  AND2_X1 U5134 ( .A1(n8500), .A2(n4644), .ZN(n8505) );
  NAND2_X1 U5135 ( .A1(n8502), .A2(n8501), .ZN(n4644) );
  OAI21_X1 U5136 ( .B1(n6188), .B2(P2_D_REG_0__SCAN_IN), .A(n6583), .ZN(n6293)
         );
  OR2_X1 U5137 ( .A1(n8842), .A2(n8321), .ZN(n8165) );
  INV_X1 U5138 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5054) );
  NOR2_X1 U5139 ( .A1(n5041), .A2(SI_16_), .ZN(n5043) );
  NAND3_X1 U5140 ( .A1(n9122), .A2(n4837), .A3(n4836), .ZN(n4835) );
  INV_X1 U5141 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4836) );
  OR2_X1 U5142 ( .A1(n6363), .A2(n8623), .ZN(n6364) );
  XNOR2_X1 U5143 ( .A(n6412), .B(n6986), .ZN(n6310) );
  AOI21_X1 U5144 ( .B1(n6317), .B2(n6318), .A(n4388), .ZN(n4491) );
  INV_X1 U5145 ( .A(n6874), .ZN(n4723) );
  AND2_X1 U5146 ( .A1(n6870), .A2(n6869), .ZN(n6871) );
  AND2_X1 U5147 ( .A1(n7039), .A2(n7044), .ZN(n7040) );
  AND2_X1 U5148 ( .A1(n5757), .A2(n5758), .ZN(n4613) );
  OAI21_X1 U5149 ( .B1(n4820), .B2(n7376), .A(n4819), .ZN(n7483) );
  NAND2_X1 U5150 ( .A1(n7432), .A2(n4821), .ZN(n4819) );
  OR2_X1 U5151 ( .A1(n7375), .A2(n7379), .ZN(n4820) );
  OR2_X1 U5152 ( .A1(n4649), .A2(n8398), .ZN(n4647) );
  OR2_X1 U5153 ( .A1(n8360), .A2(n4648), .ZN(n4646) );
  NAND2_X1 U5154 ( .A1(n4651), .A2(n8363), .ZN(n4648) );
  NOR2_X1 U5155 ( .A1(n8505), .A2(n8504), .ZN(n8529) );
  AND2_X1 U5156 ( .A1(n5953), .A2(n4577), .ZN(n4576) );
  INV_X1 U5157 ( .A(n5955), .ZN(n5954) );
  NOR2_X1 U5158 ( .A1(n5916), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n4574) );
  INV_X1 U5159 ( .A(n8352), .ZN(n6220) );
  NAND2_X1 U5160 ( .A1(n7201), .A2(n8539), .ZN(n6297) );
  NOR2_X1 U5161 ( .A1(n4679), .A2(n4678), .ZN(n4677) );
  INV_X1 U5162 ( .A(n8195), .ZN(n4678) );
  NOR2_X1 U5163 ( .A1(n4680), .A2(n8196), .ZN(n4679) );
  OR2_X1 U5164 ( .A1(n8738), .A2(n7713), .ZN(n8203) );
  OR2_X1 U5165 ( .A1(n8798), .A2(n8557), .ZN(n8195) );
  OR2_X1 U5166 ( .A1(n8831), .A2(n8659), .ZN(n8169) );
  OR2_X1 U5167 ( .A1(n8825), .A2(n8637), .ZN(n8178) );
  INV_X1 U5168 ( .A(n5983), .ZN(n4620) );
  NAND2_X1 U5169 ( .A1(n4697), .A2(n8138), .ZN(n4695) );
  OR2_X1 U5170 ( .A1(n7606), .A2(n8348), .ZN(n7596) );
  INV_X1 U5171 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5778) );
  NOR3_X1 U5172 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n5765) );
  AND2_X1 U5173 ( .A1(n5157), .A2(n5156), .ZN(n5163) );
  AND2_X1 U5174 ( .A1(n5553), .A2(n4802), .ZN(n4801) );
  INV_X1 U5175 ( .A(n5574), .ZN(n4802) );
  INV_X1 U5176 ( .A(n6531), .ZN(n5723) );
  OR2_X1 U5177 ( .A1(n7924), .A2(n4538), .ZN(n4537) );
  NAND2_X1 U5178 ( .A1(n7780), .A2(n4539), .ZN(n4538) );
  NOR2_X1 U5179 ( .A1(n7972), .A2(n4534), .ZN(n4533) );
  NAND2_X1 U5180 ( .A1(n4536), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U5181 ( .A1(n7919), .A2(n7937), .ZN(n4535) );
  NAND2_X1 U5182 ( .A1(n7918), .A2(n7917), .ZN(n4543) );
  NOR2_X1 U5183 ( .A1(n7919), .A2(n4542), .ZN(n4541) );
  NAND2_X1 U5184 ( .A1(n7930), .A2(n7937), .ZN(n7935) );
  OR2_X1 U5185 ( .A1(n6741), .A2(n4381), .ZN(n4494) );
  INV_X1 U5186 ( .A(n6636), .ZN(n4498) );
  AND2_X1 U5187 ( .A1(n4661), .A2(n4660), .ZN(n9453) );
  NAND2_X1 U5188 ( .A1(n6638), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4660) );
  OR2_X1 U5189 ( .A1(n9341), .A2(n9346), .ZN(n4793) );
  OAI21_X1 U5190 ( .B1(n4711), .B2(n7971), .A(n7769), .ZN(n4710) );
  INV_X1 U5191 ( .A(n4712), .ZN(n4487) );
  AND2_X1 U5192 ( .A1(n4811), .A2(n9207), .ZN(n4810) );
  NOR2_X1 U5193 ( .A1(n9371), .A2(n9376), .ZN(n4811) );
  OR2_X1 U5194 ( .A1(n9371), .A2(n8980), .ZN(n7902) );
  NOR2_X1 U5195 ( .A1(n9267), .A2(n9381), .ZN(n9226) );
  OR2_X1 U5196 ( .A1(n9381), .A2(n8982), .ZN(n7903) );
  OR2_X1 U5197 ( .A1(n9323), .A2(n9512), .ZN(n4816) );
  INV_X1 U5198 ( .A(n7874), .ZN(n4737) );
  INV_X1 U5199 ( .A(n4808), .ZN(n4807) );
  NAND2_X1 U5200 ( .A1(n9780), .A2(n9774), .ZN(n4808) );
  OAI22_X1 U5201 ( .A1(n6542), .A2(n5404), .B1(n7796), .B2(n9565), .ZN(n4562)
         );
  INV_X1 U5202 ( .A(n5670), .ZN(n5671) );
  AND2_X1 U5203 ( .A1(n6135), .A2(n5677), .ZN(n6133) );
  INV_X1 U5204 ( .A(n4861), .ZN(n5624) );
  AOI21_X1 U5205 ( .B1(n5558), .B2(n4865), .A(n4862), .ZN(n4861) );
  NAND2_X1 U5206 ( .A1(n4863), .A2(n5600), .ZN(n4862) );
  NAND2_X1 U5207 ( .A1(n4865), .A2(n4867), .ZN(n4863) );
  AND2_X1 U5208 ( .A1(n5625), .A2(n5604), .ZN(n5623) );
  NAND2_X1 U5209 ( .A1(n4871), .A2(n5556), .ZN(n4870) );
  INV_X1 U5210 ( .A(n5576), .ZN(n4871) );
  AOI21_X1 U5211 ( .B1(n4403), .B2(n4851), .A(n4848), .ZN(n4847) );
  INV_X1 U5212 ( .A(n5512), .ZN(n4848) );
  NOR2_X1 U5213 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5086) );
  NOR2_X1 U5214 ( .A1(n5469), .A2(n4860), .ZN(n4859) );
  OAI21_X1 U5215 ( .B1(n5469), .B2(n4858), .A(n5048), .ZN(n4857) );
  NAND2_X1 U5216 ( .A1(n5043), .A2(n5042), .ZN(n4858) );
  INV_X1 U5217 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U5218 ( .A1(n5031), .A2(SI_13_), .ZN(n5035) );
  INV_X1 U5219 ( .A(n5317), .ZN(n4840) );
  XNOR2_X1 U5220 ( .A(n5017), .B(SI_8_), .ZN(n5302) );
  INV_X1 U5221 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4666) );
  AOI21_X1 U5222 ( .B1(n7708), .B2(n4363), .A(n4937), .ZN(n4936) );
  NOR2_X1 U5223 ( .A1(n7708), .A2(n8557), .ZN(n4938) );
  INV_X1 U5224 ( .A(n4491), .ZN(n4490) );
  OAI211_X1 U5225 ( .C1(n4507), .C2(n6300), .A(n4505), .B(n4503), .ZN(n6301)
         );
  NAND2_X1 U5226 ( .A1(n4339), .A2(n4506), .ZN(n4505) );
  NAND2_X1 U5227 ( .A1(n4507), .A2(n4504), .ZN(n4503) );
  NAND2_X1 U5228 ( .A1(n7682), .A2(n7681), .ZN(n4951) );
  AND2_X1 U5229 ( .A1(n7721), .A2(n6371), .ZN(n8278) );
  NAND2_X1 U5230 ( .A1(n7190), .A2(n6332), .ZN(n6333) );
  INV_X1 U5231 ( .A(n6412), .ZN(n6375) );
  XNOR2_X1 U5232 ( .A(n9948), .B(n6412), .ZN(n6307) );
  NAND2_X1 U5233 ( .A1(n4492), .A2(n4491), .ZN(n6933) );
  OR2_X1 U5234 ( .A1(n4873), .A2(n4467), .ZN(n4466) );
  NAND2_X1 U5235 ( .A1(n8217), .A2(n8219), .ZN(n4467) );
  NAND2_X1 U5236 ( .A1(n8032), .A2(n8215), .ZN(n4701) );
  OAI21_X1 U5237 ( .B1(n8026), .B2(n4703), .A(n4391), .ZN(n4702) );
  INV_X1 U5238 ( .A(n8033), .ZN(n4703) );
  AND4_X1 U5239 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n8238)
         );
  AND4_X1 U5240 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n7510)
         );
  OR2_X1 U5241 ( .A1(n5816), .A2(n5907), .ZN(n5908) );
  NAND2_X1 U5242 ( .A1(n4823), .A2(n4827), .ZN(n4824) );
  INV_X1 U5243 ( .A(n6707), .ZN(n4823) );
  XNOR2_X1 U5244 ( .A(n6870), .B(n6861), .ZN(n6802) );
  OAI21_X1 U5245 ( .B1(n6798), .B2(n4405), .A(n4583), .ZN(n7042) );
  NAND2_X1 U5246 ( .A1(n4969), .A2(n4828), .ZN(n4583) );
  INV_X1 U5247 ( .A(n6868), .ZN(n4828) );
  INV_X1 U5248 ( .A(n4727), .ZN(n4726) );
  INV_X1 U5249 ( .A(n7040), .ZN(n4728) );
  OR2_X1 U5250 ( .A1(n7303), .A2(n5902), .ZN(n4747) );
  NAND2_X1 U5251 ( .A1(n4748), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4746) );
  NAND2_X1 U5252 ( .A1(n7360), .A2(n4748), .ZN(n4744) );
  XNOR2_X1 U5253 ( .A(n7483), .B(n7486), .ZN(n4585) );
  NOR2_X1 U5254 ( .A1(n8358), .A2(n8365), .ZN(n4649) );
  NAND2_X1 U5255 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  INV_X1 U5256 ( .A(n8393), .ZN(n4719) );
  NOR2_X1 U5257 ( .A1(n8456), .A2(n8457), .ZN(n8460) );
  OR2_X1 U5258 ( .A1(n8460), .A2(n8459), .ZN(n4818) );
  NAND2_X1 U5259 ( .A1(n6105), .A2(n6104), .ZN(n6117) );
  INV_X1 U5260 ( .A(n6106), .ZN(n6105) );
  INV_X1 U5261 ( .A(n6062), .ZN(n6061) );
  AOI21_X1 U5262 ( .B1(n4689), .B2(n4368), .A(n4688), .ZN(n4687) );
  INV_X1 U5263 ( .A(n8168), .ZN(n4688) );
  NAND2_X1 U5264 ( .A1(n6004), .A2(n4366), .ZN(n6052) );
  INV_X1 U5265 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4578) );
  OR2_X1 U5266 ( .A1(n5993), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6005) );
  INV_X1 U5267 ( .A(n8349), .ZN(n7569) );
  OR2_X1 U5268 ( .A1(n9980), .A2(n6220), .ZN(n8113) );
  NAND2_X1 U5269 ( .A1(n5904), .A2(n5903), .ZN(n5916) );
  INV_X1 U5270 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5903) );
  INV_X1 U5271 ( .A(n5905), .ZN(n5904) );
  OR2_X1 U5272 ( .A1(n5888), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5905) );
  AND4_X1 U5273 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n9924)
         );
  OR2_X1 U5274 ( .A1(n5790), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U5275 ( .A1(n6263), .A2(n6262), .ZN(n6283) );
  NOR2_X1 U5276 ( .A1(n4638), .A2(n4636), .ZN(n4635) );
  NAND2_X1 U5277 ( .A1(n6170), .A2(n9995), .ZN(n4636) );
  NAND2_X1 U5278 ( .A1(n8578), .A2(n8585), .ZN(n6114) );
  NOR2_X1 U5279 ( .A1(n8198), .A2(n4681), .ZN(n4680) );
  INV_X1 U5280 ( .A(n8189), .ZN(n4681) );
  OR2_X1 U5281 ( .A1(n8809), .A2(n8248), .ZN(n8189) );
  NAND2_X1 U5282 ( .A1(n4624), .A2(n4623), .ZN(n8622) );
  NOR2_X1 U5283 ( .A1(n4625), .A2(n4390), .ZN(n4623) );
  NOR2_X1 U5284 ( .A1(n4690), .A2(n6057), .ZN(n4689) );
  INV_X1 U5285 ( .A(n4379), .ZN(n4690) );
  NOR2_X1 U5286 ( .A1(n5984), .A2(n4622), .ZN(n4621) );
  INV_X1 U5287 ( .A(n5971), .ZN(n4622) );
  AND2_X1 U5288 ( .A1(n8147), .A2(n8694), .ZN(n8146) );
  INV_X1 U5289 ( .A(n8049), .ZN(n8142) );
  NAND2_X1 U5290 ( .A1(n4698), .A2(n8133), .ZN(n4697) );
  INV_X1 U5291 ( .A(n8139), .ZN(n4698) );
  INV_X1 U5292 ( .A(n8720), .ZN(n9933) );
  INV_X1 U5293 ( .A(n8718), .ZN(n9930) );
  NOR2_X1 U5294 ( .A1(n7535), .A2(n8136), .ZN(n4699) );
  NAND2_X1 U5295 ( .A1(n8072), .A2(n7318), .ZN(n9989) );
  NAND2_X1 U5296 ( .A1(n5758), .A2(n4517), .ZN(n4516) );
  INV_X1 U5297 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4517) );
  AND2_X1 U5298 ( .A1(n5765), .A2(n4705), .ZN(n4348) );
  INV_X1 U5299 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4705) );
  INV_X1 U5300 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5768) );
  INV_X1 U5301 ( .A(n6166), .ZN(n8530) );
  NAND2_X1 U5302 ( .A1(n6024), .A2(n4374), .ZN(n4600) );
  INV_X1 U5303 ( .A(n4602), .ZN(n4601) );
  OAI21_X1 U5304 ( .B1(n4374), .B2(n4603), .A(n6151), .ZN(n4602) );
  INV_X1 U5305 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4462) );
  OR2_X1 U5306 ( .A1(n5858), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5880) );
  NOR2_X1 U5307 ( .A1(n5820), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5839) );
  OR2_X1 U5308 ( .A1(n5799), .A2(n4603), .ZN(n4822) );
  AND2_X1 U5309 ( .A1(n8962), .A2(n5596), .ZN(n8870) );
  NOR2_X1 U5310 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  INV_X1 U5311 ( .A(n4779), .ZN(n4778) );
  INV_X1 U5312 ( .A(n7464), .ZN(n4780) );
  NAND2_X1 U5313 ( .A1(n8913), .A2(n4801), .ZN(n4800) );
  NAND2_X1 U5314 ( .A1(n8913), .A2(n5553), .ZN(n4794) );
  NAND2_X1 U5315 ( .A1(n7078), .A2(n7080), .ZN(n4752) );
  NAND2_X1 U5316 ( .A1(n5258), .A2(n5257), .ZN(n7077) );
  AND2_X1 U5317 ( .A1(n5231), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5259) );
  INV_X1 U5318 ( .A(n4763), .ZN(n4762) );
  AOI21_X1 U5319 ( .B1(n4765), .B2(n4763), .A(n4359), .ZN(n4761) );
  AND2_X1 U5320 ( .A1(n5111), .A2(n5110), .ZN(n8886) );
  NOR2_X1 U5321 ( .A1(n9489), .A2(n9490), .ZN(n9491) );
  NAND2_X1 U5322 ( .A1(n4670), .A2(n4669), .ZN(n9089) );
  AOI21_X1 U5323 ( .B1(n4371), .B2(n9634), .A(n9082), .ZN(n4669) );
  OR2_X1 U5324 ( .A1(n9635), .A2(n9634), .ZN(n4671) );
  INV_X1 U5325 ( .A(n4792), .ZN(n4787) );
  NOR2_X1 U5326 ( .A1(n9135), .A2(n4793), .ZN(n4792) );
  NOR2_X1 U5327 ( .A1(n9352), .A2(n4973), .ZN(n9159) );
  NAND2_X1 U5328 ( .A1(n9356), .A2(n9040), .ZN(n4893) );
  NAND2_X1 U5329 ( .A1(n9017), .A2(n7776), .ZN(n4895) );
  OR2_X1 U5330 ( .A1(n9184), .A2(n9356), .ZN(n4973) );
  AOI21_X1 U5331 ( .B1(n4369), .B2(n9234), .A(n4732), .ZN(n4731) );
  INV_X1 U5332 ( .A(n7908), .ZN(n4732) );
  NOR2_X1 U5333 ( .A1(n6468), .A2(n4925), .ZN(n4924) );
  INV_X1 U5334 ( .A(n4929), .ZN(n4925) );
  NAND2_X1 U5335 ( .A1(n4409), .A2(n4929), .ZN(n4923) );
  AND2_X1 U5336 ( .A1(n9215), .A2(n8980), .ZN(n4930) );
  INV_X1 U5337 ( .A(n6467), .ZN(n4926) );
  AND2_X1 U5338 ( .A1(n7902), .A2(n7908), .ZN(n9218) );
  OR2_X1 U5339 ( .A1(n9233), .A2(n9234), .ZN(n4734) );
  NOR2_X1 U5340 ( .A1(n9386), .A2(n9278), .ZN(n6465) );
  NAND2_X1 U5341 ( .A1(n7757), .A2(n4488), .ZN(n4713) );
  OR2_X1 U5342 ( .A1(n9328), .A2(n4716), .ZN(n4488) );
  NAND2_X1 U5343 ( .A1(n7629), .A2(n7630), .ZN(n7628) );
  NAND2_X1 U5344 ( .A1(n7757), .A2(n7760), .ZN(n9328) );
  INV_X1 U5345 ( .A(n7960), .ZN(n7398) );
  AND2_X1 U5346 ( .A1(n5391), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5411) );
  OR3_X1 U5347 ( .A1(n9707), .A2(n9818), .A3(n4343), .ZN(n9708) );
  AOI21_X1 U5348 ( .B1(n7278), .B2(n4901), .A(n4397), .ZN(n4900) );
  INV_X1 U5349 ( .A(n9008), .ZN(n9309) );
  NAND2_X1 U5350 ( .A1(n6512), .A2(n8005), .ZN(n9702) );
  NAND2_X1 U5351 ( .A1(n6778), .A2(n7822), .ZN(n4749) );
  AND2_X1 U5352 ( .A1(n9763), .A2(n5749), .ZN(n9734) );
  INV_X1 U5353 ( .A(n9006), .ZN(n9311) );
  OR2_X1 U5354 ( .A1(n6485), .A2(n9423), .ZN(n9334) );
  INV_X1 U5355 ( .A(n7565), .ZN(n5711) );
  NAND2_X1 U5356 ( .A1(n6569), .A2(n5718), .ZN(n9423) );
  AND2_X1 U5357 ( .A1(n6531), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5718) );
  XNOR2_X1 U5358 ( .A(n5101), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5106) );
  INV_X1 U5359 ( .A(n9429), .ZN(n5098) );
  NAND2_X1 U5360 ( .A1(n5081), .A2(n5060), .ZN(n5064) );
  INV_X1 U5361 ( .A(n4870), .ZN(n4869) );
  OAI21_X1 U5362 ( .B1(n4870), .B2(n4868), .A(n5575), .ZN(n4867) );
  INV_X1 U5363 ( .A(n5557), .ZN(n4868) );
  NAND2_X1 U5364 ( .A1(n4771), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5714) );
  AND2_X1 U5365 ( .A1(n4774), .A2(n5074), .ZN(n4772) );
  NAND2_X1 U5366 ( .A1(n5469), .A2(n4860), .ZN(n4478) );
  OR2_X1 U5367 ( .A1(n5039), .A2(n4481), .ZN(n4477) );
  OR2_X1 U5368 ( .A1(n4384), .A2(n4481), .ZN(n4480) );
  INV_X1 U5369 ( .A(n5038), .ZN(n5441) );
  AND2_X1 U5370 ( .A1(n4753), .A2(n4755), .ZN(n4738) );
  NAND2_X1 U5371 ( .A1(n5052), .A2(n4350), .ZN(n4918) );
  INV_X1 U5372 ( .A(n4877), .ZN(n4876) );
  OAI21_X1 U5373 ( .B1(n4883), .B2(n4878), .A(n5030), .ZN(n4877) );
  INV_X1 U5374 ( .A(n4879), .ZN(n4878) );
  OAI21_X1 U5375 ( .B1(n5029), .B2(SI_12_), .A(n5030), .ZN(n5383) );
  NOR2_X1 U5376 ( .A1(n5383), .A2(n4882), .ZN(n4879) );
  NAND2_X1 U5377 ( .A1(n5359), .A2(n4883), .ZN(n4880) );
  OAI21_X1 U5378 ( .B1(n5287), .B2(n4844), .A(n4842), .ZN(n5316) );
  NAND2_X1 U5379 ( .A1(n5238), .A2(n5006), .ZN(n5271) );
  AND2_X1 U5380 ( .A1(n5132), .A2(n5050), .ZN(n5052) );
  NAND2_X1 U5381 ( .A1(n4995), .A2(n5174), .ZN(n5178) );
  AND2_X1 U5382 ( .A1(n6934), .A2(n6324), .ZN(n7056) );
  NOR2_X1 U5383 ( .A1(n4944), .A2(n4943), .ZN(n4942) );
  OAI21_X1 U5384 ( .B1(n4945), .B2(n4943), .A(n4941), .ZN(n4940) );
  INV_X1 U5385 ( .A(n8254), .ZN(n4943) );
  NAND2_X1 U5386 ( .A1(n6138), .A2(n6137), .ZN(n8547) );
  INV_X1 U5387 ( .A(n8315), .ZN(n8327) );
  NAND2_X1 U5388 ( .A1(n6132), .A2(n6131), .ZN(n8571) );
  OR2_X1 U5389 ( .A1(n5790), .A2(n5791), .ZN(n5798) );
  OR2_X1 U5390 ( .A1(n5886), .A2(n5794), .ZN(n5795) );
  OR2_X1 U5391 ( .A1(n5828), .A2(n6955), .ZN(n5774) );
  NAND2_X1 U5392 ( .A1(n4592), .A2(n4373), .ZN(n4591) );
  NAND2_X1 U5393 ( .A1(n4652), .A2(n4651), .ZN(n4650) );
  INV_X1 U5394 ( .A(n4718), .ZN(n8416) );
  INV_X1 U5395 ( .A(n4708), .ZN(n8487) );
  INV_X1 U5396 ( .A(n8514), .ZN(n4653) );
  NAND2_X1 U5397 ( .A1(n4655), .A2(n8528), .ZN(n4654) );
  NAND2_X1 U5398 ( .A1(n8512), .A2(n8511), .ZN(n4656) );
  OAI21_X1 U5399 ( .B1(n8499), .B2(n8498), .A(n8497), .ZN(n8515) );
  AND2_X1 U5400 ( .A1(n4637), .A2(n4633), .ZN(n6249) );
  NOR2_X1 U5401 ( .A1(n4638), .A2(n4634), .ZN(n4633) );
  INV_X1 U5402 ( .A(n6170), .ZN(n4634) );
  AOI21_X1 U5403 ( .B1(n9426), .B2(n8025), .A(n8024), .ZN(n8786) );
  INV_X1 U5404 ( .A(n6283), .ZN(n7689) );
  INV_X1 U5405 ( .A(n4635), .ZN(n4632) );
  NAND2_X1 U5406 ( .A1(n6080), .A2(n6079), .ZN(n8815) );
  NAND2_X1 U5407 ( .A1(n5940), .A2(n5939), .ZN(n7547) );
  OR2_X1 U5408 ( .A1(n9997), .A2(n9989), .ZN(n8834) );
  AND2_X1 U5409 ( .A1(n5434), .A2(n5433), .ZN(n9026) );
  AOI21_X1 U5410 ( .B1(n4524), .B2(n4527), .A(n4444), .ZN(n4520) );
  OAI211_X1 U5411 ( .C1(n7943), .C2(n7942), .A(n8004), .B(n7941), .ZN(n8002)
         );
  OR2_X1 U5412 ( .A1(n6648), .A2(n8012), .ZN(n9649) );
  NAND2_X1 U5413 ( .A1(n8086), .A2(n4459), .ZN(n4458) );
  AND2_X1 U5414 ( .A1(n8097), .A2(n8206), .ZN(n4459) );
  INV_X1 U5415 ( .A(n7828), .ZN(n4531) );
  NOR2_X1 U5416 ( .A1(n4450), .A2(n4449), .ZN(n4448) );
  INV_X1 U5417 ( .A(n8128), .ZN(n4450) );
  INV_X1 U5418 ( .A(n8123), .ZN(n4449) );
  NAND2_X1 U5419 ( .A1(n4553), .A2(n7843), .ZN(n7851) );
  NAND2_X1 U5420 ( .A1(n4611), .A2(n8146), .ZN(n8156) );
  INV_X1 U5421 ( .A(n4610), .ZN(n4609) );
  INV_X1 U5422 ( .A(n7873), .ZN(n4547) );
  NAND2_X1 U5423 ( .A1(n4550), .A2(n4549), .ZN(n7875) );
  NAND2_X1 U5424 ( .A1(n7860), .A2(n7932), .ZN(n4549) );
  NAND2_X1 U5425 ( .A1(n7859), .A2(n7937), .ZN(n4550) );
  INV_X1 U5426 ( .A(n8181), .ZN(n4608) );
  AND2_X1 U5427 ( .A1(n8613), .A2(n8180), .ZN(n4607) );
  AND2_X1 U5428 ( .A1(n4545), .A2(n4544), .ZN(n7880) );
  NAND2_X1 U5429 ( .A1(n8202), .A2(n8201), .ZN(n4606) );
  INV_X1 U5430 ( .A(n4606), .ZN(n4455) );
  OR2_X1 U5431 ( .A1(n4606), .A2(n8193), .ZN(n4605) );
  OAI211_X1 U5432 ( .C1(n4559), .C2(n4558), .A(n7907), .B(n4556), .ZN(n7909)
         );
  AOI21_X1 U5433 ( .B1(n7906), .B2(n4472), .A(n4560), .ZN(n4559) );
  INV_X1 U5434 ( .A(n5513), .ZN(n4850) );
  NOR2_X1 U5435 ( .A1(n8368), .A2(n4956), .ZN(n4589) );
  AND2_X1 U5436 ( .A1(n6638), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4500) );
  AND2_X1 U5437 ( .A1(n9286), .A2(n8972), .ZN(n7893) );
  INV_X1 U5438 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5056) );
  INV_X1 U5439 ( .A(n4866), .ZN(n4865) );
  OAI21_X1 U5440 ( .B1(n4867), .B2(n4869), .A(n5598), .ZN(n4866) );
  NAND2_X1 U5441 ( .A1(n5497), .A2(n5496), .ZN(n5512) );
  NOR2_X1 U5442 ( .A1(n5114), .A2(SI_14_), .ZN(n4889) );
  NOR2_X1 U5443 ( .A1(n6374), .A2(n8579), .ZN(n4937) );
  INV_X1 U5444 ( .A(n6299), .ZN(n4506) );
  AOI21_X1 U5445 ( .B1(n4950), .B2(n4948), .A(n8313), .ZN(n4947) );
  INV_X1 U5446 ( .A(n7681), .ZN(n4948) );
  INV_X1 U5447 ( .A(n8213), .ZN(n4874) );
  NAND2_X1 U5448 ( .A1(n8214), .A2(n4406), .ZN(n4875) );
  NAND2_X1 U5449 ( .A1(n6706), .A2(n6707), .ZN(n6756) );
  AND2_X1 U5450 ( .A1(n4584), .A2(n6869), .ZN(n4969) );
  NAND2_X1 U5451 ( .A1(n4589), .A2(n8387), .ZN(n8369) );
  OR2_X1 U5452 ( .A1(n8379), .A2(n8378), .ZN(n8381) );
  NAND2_X1 U5453 ( .A1(n8369), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4832) );
  AOI21_X1 U5454 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8431), .A(n8430), .ZN(
        n8454) );
  AND2_X1 U5455 ( .A1(n4818), .A2(n4593), .ZN(n8492) );
  NAND2_X1 U5456 ( .A1(n8471), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4593) );
  OR2_X1 U5457 ( .A1(n6283), .A2(n6264), .ZN(n8033) );
  AND2_X1 U5458 ( .A1(n6003), .A2(n4580), .ZN(n4579) );
  INV_X1 U5459 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4580) );
  INV_X1 U5460 ( .A(n6005), .ZN(n6004) );
  NAND2_X1 U5461 ( .A1(n8356), .A2(n9954), .ZN(n8091) );
  OR2_X1 U5462 ( .A1(n5816), .A2(n6984), .ZN(n5804) );
  AND2_X1 U5463 ( .A1(n6190), .A2(n6580), .ZN(n6244) );
  INV_X1 U5464 ( .A(n8555), .ZN(n6266) );
  OR2_X1 U5465 ( .A1(n8815), .A2(n6368), .ZN(n8183) );
  NAND2_X1 U5466 ( .A1(n4642), .A2(n5863), .ZN(n7209) );
  NAND2_X1 U5467 ( .A1(n6216), .A2(n6215), .ZN(n6944) );
  AND2_X1 U5468 ( .A1(n6022), .A2(n6021), .ZN(n6023) );
  AND2_X1 U5469 ( .A1(n6020), .A2(n6019), .ZN(n6022) );
  INV_X1 U5470 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4461) );
  INV_X1 U5471 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5757) );
  OR2_X1 U5472 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  OAI21_X1 U5473 ( .B1(n4801), .B2(n8979), .A(n4797), .ZN(n4796) );
  NAND2_X1 U5474 ( .A1(n4798), .A2(n5574), .ZN(n4797) );
  INV_X1 U5475 ( .A(n5553), .ZN(n4798) );
  AND2_X1 U5476 ( .A1(n4663), .A2(n4662), .ZN(n9556) );
  NAND2_X1 U5477 ( .A1(n6634), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4662) );
  INV_X1 U5478 ( .A(n9545), .ZN(n4499) );
  INV_X1 U5479 ( .A(n4495), .ZN(n9460) );
  AOI22_X1 U5480 ( .A1(n9545), .A2(n4497), .B1(n9560), .B2(n4496), .ZN(n4495)
         );
  NOR2_X1 U5481 ( .A1(n4500), .A2(n4498), .ZN(n4497) );
  INV_X1 U5482 ( .A(n4500), .ZN(n4496) );
  NOR2_X1 U5483 ( .A1(n9460), .A2(n9459), .ZN(n9461) );
  OR2_X1 U5484 ( .A1(n9571), .A2(n4440), .ZN(n9573) );
  NAND2_X1 U5485 ( .A1(n9076), .A2(n4658), .ZN(n9590) );
  OR2_X1 U5486 ( .A1(n9077), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4658) );
  NOR2_X1 U5487 ( .A1(n9591), .A2(n9590), .ZN(n9592) );
  NAND2_X1 U5488 ( .A1(n9062), .A2(n9063), .ZN(n9596) );
  NOR2_X1 U5489 ( .A1(n9596), .A2(n9597), .ZN(n9598) );
  NOR2_X1 U5490 ( .A1(n9592), .A2(n4657), .ZN(n9610) );
  AND2_X1 U5491 ( .A1(n9589), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4657) );
  NOR2_X1 U5492 ( .A1(n9610), .A2(n9611), .ZN(n9612) );
  NOR2_X1 U5493 ( .A1(n9598), .A2(n4510), .ZN(n9617) );
  AND2_X1 U5494 ( .A1(n9589), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5495 ( .A1(n7925), .A2(n7917), .ZN(n7970) );
  NAND2_X1 U5496 ( .A1(n4923), .A2(n4922), .ZN(n4919) );
  INV_X1 U5497 ( .A(n4924), .ZN(n4922) );
  NAND2_X1 U5498 ( .A1(n9259), .A2(n4472), .ZN(n7983) );
  INV_X1 U5499 ( .A(n7893), .ZN(n7765) );
  INV_X1 U5500 ( .A(n7872), .ZN(n4716) );
  AND2_X1 U5501 ( .A1(n7757), .A2(n7630), .ZN(n4715) );
  NAND2_X1 U5502 ( .A1(n9833), .A2(n4358), .ZN(n4768) );
  NOR2_X1 U5503 ( .A1(n7960), .A2(n4907), .ZN(n4906) );
  INV_X1 U5504 ( .A(n9667), .ZN(n4907) );
  INV_X1 U5505 ( .A(n6451), .ZN(n4908) );
  NOR2_X1 U5506 ( .A1(n4902), .A2(n4899), .ZN(n4898) );
  INV_X1 U5507 ( .A(n7278), .ZN(n4902) );
  INV_X1 U5508 ( .A(n6439), .ZN(n4901) );
  NAND2_X1 U5509 ( .A1(n4750), .A2(n4749), .ZN(n7741) );
  AND2_X1 U5510 ( .A1(n4387), .A2(n7821), .ZN(n4750) );
  INV_X1 U5511 ( .A(n7812), .ZN(n7827) );
  NOR2_X1 U5512 ( .A1(n7737), .A2(n9735), .ZN(n7945) );
  AND2_X1 U5513 ( .A1(n4753), .A2(n5132), .ZN(n4739) );
  AND4_X1 U5514 ( .A1(n4755), .A2(n5050), .A3(n5054), .A4(n5059), .ZN(n4741)
         );
  INV_X1 U5515 ( .A(n4855), .ZN(n4853) );
  AOI21_X1 U5516 ( .B1(n4855), .B2(n4852), .A(n4432), .ZN(n4851) );
  INV_X1 U5517 ( .A(n4859), .ZN(n4852) );
  INV_X1 U5518 ( .A(n5043), .ZN(n4483) );
  NAND2_X1 U5519 ( .A1(n4482), .A2(n5042), .ZN(n4481) );
  INV_X1 U5520 ( .A(n5469), .ZN(n4482) );
  NAND2_X1 U5521 ( .A1(n4888), .A2(n4885), .ZN(n5038) );
  INV_X1 U5522 ( .A(n4889), .ZN(n4885) );
  OR2_X1 U5523 ( .A1(n5303), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5342) );
  OAI21_X1 U5524 ( .B1(n7795), .B2(n4977), .A(n4976), .ZN(n4980) );
  INV_X1 U5525 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U5526 ( .A1(n4998), .A2(SI_3_), .ZN(n5000) );
  OAI211_X1 U5527 ( .C1(n4835), .C2(n4476), .A(n4475), .B(n4474), .ZN(n4985)
         );
  INV_X1 U5528 ( .A(n8253), .ZN(n4941) );
  INV_X1 U5529 ( .A(n4947), .ZN(n4944) );
  AOI21_X1 U5530 ( .B1(n4947), .B2(n4949), .A(n4946), .ZN(n4945) );
  INV_X1 U5531 ( .A(n8312), .ZN(n4946) );
  INV_X1 U5532 ( .A(n4950), .ZN(n4949) );
  AND2_X1 U5533 ( .A1(n8269), .A2(n4383), .ZN(n4950) );
  NAND2_X1 U5534 ( .A1(n8356), .A2(n6311), .ZN(n6881) );
  AND2_X1 U5535 ( .A1(n8261), .A2(n6358), .ZN(n8291) );
  INV_X1 U5536 ( .A(n6301), .ZN(n6302) );
  NAND2_X1 U5537 ( .A1(n4939), .A2(n4945), .ZN(n8311) );
  NAND2_X1 U5538 ( .A1(n7682), .A2(n4947), .ZN(n4939) );
  INV_X1 U5539 ( .A(n6559), .ZN(n6401) );
  OR2_X1 U5540 ( .A1(n5816), .A2(n6794), .ZN(n5836) );
  XNOR2_X1 U5541 ( .A(n6693), .B(n6714), .ZN(n9885) );
  OR2_X1 U5542 ( .A1(n9894), .A2(n6955), .ZN(n9892) );
  OAI21_X1 U5543 ( .B1(n6711), .B2(n5792), .A(n4730), .ZN(n9902) );
  NAND2_X1 U5544 ( .A1(n4826), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6758) );
  INV_X1 U5545 ( .A(n6756), .ZN(n4826) );
  OR2_X1 U5546 ( .A1(n6753), .A2(n10000), .ZN(n6755) );
  AND2_X1 U5547 ( .A1(n6802), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6872) );
  XNOR2_X1 U5548 ( .A(n4584), .B(n6869), .ZN(n6798) );
  OR2_X1 U5549 ( .A1(n6798), .A2(n6794), .ZN(n4831) );
  INV_X1 U5550 ( .A(n4969), .ZN(n4830) );
  NAND2_X1 U5551 ( .A1(n4722), .A2(n4721), .ZN(n7038) );
  NAND2_X1 U5552 ( .A1(n6871), .A2(n4723), .ZN(n4721) );
  NAND2_X1 U5553 ( .A1(n6802), .A2(n4393), .ZN(n4722) );
  NAND2_X1 U5554 ( .A1(n7045), .A2(n7044), .ZN(n7046) );
  OR2_X1 U5555 ( .A1(n7040), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U5556 ( .A1(n4729), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4725) );
  OR2_X1 U5557 ( .A1(n7040), .A2(n5864), .ZN(n4727) );
  NOR2_X1 U5558 ( .A1(n7287), .A2(n7286), .ZN(n7372) );
  AND2_X1 U5559 ( .A1(n7299), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7286) );
  NOR2_X1 U5560 ( .A1(n7372), .A2(n7374), .ZN(n7375) );
  AND2_X1 U5561 ( .A1(n4587), .A2(n4586), .ZN(n7488) );
  NAND2_X1 U5562 ( .A1(n7485), .A2(n7486), .ZN(n4586) );
  NOR2_X1 U5563 ( .A1(n8406), .A2(n4832), .ZN(n8405) );
  NAND2_X1 U5564 ( .A1(n4588), .A2(n8369), .ZN(n8370) );
  AND2_X1 U5565 ( .A1(n4646), .A2(n4435), .ZN(n8422) );
  INV_X1 U5566 ( .A(n8400), .ZN(n4645) );
  NAND2_X1 U5567 ( .A1(n4646), .A2(n4647), .ZN(n8399) );
  AND2_X1 U5568 ( .A1(n4588), .A2(n4832), .ZN(n8409) );
  XNOR2_X1 U5569 ( .A(n8454), .B(n8455), .ZN(n8433) );
  AND2_X1 U5570 ( .A1(n4718), .A2(n4717), .ZN(n8439) );
  NAND2_X1 U5571 ( .A1(n8431), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4717) );
  NOR2_X1 U5572 ( .A1(n8445), .A2(n8444), .ZN(n8478) );
  XNOR2_X1 U5573 ( .A(n8492), .B(n8501), .ZN(n8472) );
  NOR2_X1 U5574 ( .A1(n8472), .A2(n8689), .ZN(n8493) );
  NAND2_X1 U5575 ( .A1(n8482), .A2(n8481), .ZN(n8500) );
  OR2_X1 U5576 ( .A1(n8467), .A2(n4709), .ZN(n4708) );
  AND2_X1 U5577 ( .A1(n8471), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U5578 ( .A1(n8506), .A2(n8527), .ZN(n8508) );
  NAND2_X1 U5579 ( .A1(n4570), .A2(n6092), .ZN(n6106) );
  INV_X1 U5580 ( .A(n4570), .ZN(n6093) );
  OR2_X1 U5581 ( .A1(n6071), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6081) );
  AND2_X1 U5582 ( .A1(n8169), .A2(n8173), .ZN(n8640) );
  AND3_X1 U5583 ( .A1(n6066), .A2(n6065), .A3(n6064), .ZN(n8637) );
  NAND2_X1 U5584 ( .A1(n6004), .A2(n4579), .ZN(n6044) );
  NAND2_X1 U5585 ( .A1(n6012), .A2(n6011), .ZN(n8630) );
  NAND2_X1 U5586 ( .A1(n6004), .A2(n6003), .ZN(n6029) );
  NAND2_X1 U5587 ( .A1(n5954), .A2(n4364), .ZN(n5993) );
  INV_X1 U5588 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U5589 ( .A1(n5954), .A2(n4576), .ZN(n5977) );
  NAND2_X1 U5590 ( .A1(n4572), .A2(n5941), .ZN(n5955) );
  INV_X1 U5591 ( .A(n5942), .ZN(n4572) );
  NAND2_X1 U5592 ( .A1(n5954), .A2(n5953), .ZN(n5964) );
  INV_X1 U5593 ( .A(n8351), .ZN(n7339) );
  INV_X1 U5594 ( .A(n4574), .ZN(n5928) );
  NAND2_X1 U5595 ( .A1(n4684), .A2(n8108), .ZN(n4683) );
  INV_X1 U5596 ( .A(n8114), .ZN(n4684) );
  NAND2_X1 U5597 ( .A1(n5866), .A2(n5865), .ZN(n5888) );
  INV_X1 U5598 ( .A(n5867), .ZN(n5866) );
  AND2_X1 U5599 ( .A1(n4630), .A2(n5847), .ZN(n5848) );
  NAND2_X1 U5600 ( .A1(n6982), .A2(n5812), .ZN(n7092) );
  NAND2_X1 U5601 ( .A1(n5813), .A2(n6985), .ZN(n5830) );
  NAND2_X1 U5602 ( .A1(n8719), .A2(n6986), .ZN(n8097) );
  NAND2_X1 U5603 ( .A1(n8724), .A2(n5803), .ZN(n6982) );
  INV_X1 U5604 ( .A(n8082), .ZN(n8722) );
  OR2_X1 U5605 ( .A1(n6840), .A2(n6236), .ZN(n8717) );
  AOI21_X1 U5606 ( .B1(n4677), .B2(n8196), .A(n4675), .ZN(n4674) );
  INV_X1 U5607 ( .A(n8197), .ZN(n4675) );
  NAND2_X1 U5608 ( .A1(n6124), .A2(n6123), .ZN(n8738) );
  OAI21_X1 U5609 ( .B1(n8604), .B2(n6088), .A(n6089), .ZN(n8589) );
  AND3_X1 U5610 ( .A1(n6056), .A2(n6055), .A3(n6054), .ZN(n8659) );
  OR2_X1 U5611 ( .A1(n8206), .A2(n6390), .ZN(n8720) );
  OR2_X1 U5612 ( .A1(n8206), .A2(n6167), .ZN(n8718) );
  AOI21_X1 U5613 ( .B1(n4352), .B2(n4620), .A(n4392), .ZN(n4617) );
  AND2_X1 U5614 ( .A1(n4695), .A2(n8143), .ZN(n4694) );
  OR2_X1 U5615 ( .A1(n8140), .A2(n8136), .ZN(n4692) );
  AND2_X1 U5616 ( .A1(n6537), .A2(n6584), .ZN(n6559) );
  AND2_X1 U5617 ( .A1(n6184), .A2(n6183), .ZN(n6187) );
  NAND2_X1 U5618 ( .A1(n5766), .A2(n5765), .ZN(n6181) );
  NAND2_X1 U5619 ( .A1(n6024), .A2(n6023), .ZN(n6150) );
  OR2_X1 U5620 ( .A1(n5475), .A2(n5107), .ZN(n5503) );
  NAND2_X1 U5621 ( .A1(n5282), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U5622 ( .A1(n8968), .A2(n5531), .ZN(n8914) );
  AND2_X1 U5623 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5231) );
  AND2_X1 U5624 ( .A1(n8925), .A2(n5622), .ZN(n8960) );
  NAND2_X1 U5625 ( .A1(n5163), .A2(n5158), .ZN(n6657) );
  AND2_X1 U5626 ( .A1(n5518), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5541) );
  NOR2_X1 U5627 ( .A1(n5503), .A2(n8885), .ZN(n5518) );
  OAI21_X1 U5628 ( .B1(n4783), .B2(n4785), .A(n4396), .ZN(n4781) );
  INV_X1 U5629 ( .A(n5382), .ZN(n4783) );
  OR2_X1 U5630 ( .A1(n5565), .A2(n8983), .ZN(n5584) );
  NAND2_X1 U5631 ( .A1(n7323), .A2(n4784), .ZN(n4782) );
  INV_X1 U5632 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7588) );
  XNOR2_X1 U5633 ( .A(n5146), .B(n8894), .ZN(n5165) );
  NAND3_X1 U5634 ( .A1(n4752), .A2(n7077), .A3(n5278), .ZN(n7149) );
  INV_X1 U5635 ( .A(n7152), .ZN(n5278) );
  AND2_X1 U5636 ( .A1(n5259), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5282) );
  INV_X1 U5637 ( .A(n9039), .ZN(n9007) );
  NAND2_X1 U5638 ( .A1(n5411), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5447) );
  AOI21_X1 U5639 ( .B1(n4540), .B2(n4532), .A(n7936), .ZN(n7939) );
  NAND2_X1 U5640 ( .A1(n4543), .A2(n4541), .ZN(n4540) );
  AND2_X1 U5641 ( .A1(n4537), .A2(n4533), .ZN(n4532) );
  AND3_X1 U5642 ( .A1(n5545), .A2(n5544), .A3(n5543), .ZN(n8982) );
  AND2_X1 U5643 ( .A1(n5285), .A2(n5284), .ZN(n7330) );
  NOR2_X1 U5644 ( .A1(n9530), .A2(n4513), .ZN(n9531) );
  NAND2_X1 U5645 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n4513) );
  OR2_X1 U5646 ( .A1(n9473), .A2(n9472), .ZN(n9474) );
  INV_X1 U5647 ( .A(n4494), .ZN(n9478) );
  NAND2_X1 U5648 ( .A1(n4494), .A2(n4493), .ZN(n9479) );
  INV_X1 U5649 ( .A(n9477), .ZN(n4493) );
  AND2_X1 U5650 ( .A1(n9474), .A2(n4659), .ZN(n6670) );
  NAND2_X1 U5651 ( .A1(n6629), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4659) );
  NOR2_X1 U5652 ( .A1(n4499), .A2(n4498), .ZN(n9559) );
  NOR2_X1 U5653 ( .A1(n9455), .A2(n4425), .ZN(n9489) );
  NOR2_X1 U5654 ( .A1(n9495), .A2(n9496), .ZN(n9497) );
  NOR2_X1 U5655 ( .A1(n9491), .A2(n4664), .ZN(n6621) );
  AND2_X1 U5656 ( .A1(n6644), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U5657 ( .A1(n6621), .A2(n6622), .ZN(n6995) );
  NAND2_X1 U5658 ( .A1(n6999), .A2(n4511), .ZN(n9443) );
  OR2_X1 U5659 ( .A1(n7000), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4511) );
  AND2_X1 U5660 ( .A1(n9573), .A2(n4672), .ZN(n6996) );
  NAND2_X1 U5661 ( .A1(n9570), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U5662 ( .A1(n7005), .A2(n7004), .ZN(n9062) );
  NOR2_X1 U5663 ( .A1(n9631), .A2(n9632), .ZN(n9630) );
  AND2_X1 U5664 ( .A1(n9089), .A2(n9088), .ZN(n9091) );
  OR2_X1 U5665 ( .A1(n9645), .A2(n9646), .ZN(n9642) );
  OR2_X1 U5666 ( .A1(n9650), .A2(n9651), .ZN(n9647) );
  XNOR2_X1 U5667 ( .A(n4502), .B(n4501), .ZN(n9114) );
  INV_X1 U5668 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U5669 ( .A1(n9642), .A2(n9111), .ZN(n4502) );
  INV_X1 U5670 ( .A(n4793), .ZN(n4791) );
  AND2_X1 U5671 ( .A1(n6477), .A2(n5741), .ZN(n8902) );
  INV_X1 U5672 ( .A(n4484), .ZN(n9166) );
  NAND2_X1 U5673 ( .A1(n9176), .A2(n4487), .ZN(n4486) );
  INV_X1 U5674 ( .A(n4710), .ZN(n4485) );
  INV_X1 U5675 ( .A(n7970), .ZN(n9165) );
  NAND2_X1 U5676 ( .A1(n9190), .A2(n7734), .ZN(n4711) );
  NAND2_X1 U5677 ( .A1(n7911), .A2(n7734), .ZN(n4712) );
  NOR2_X1 U5678 ( .A1(n9188), .A2(n9009), .ZN(n6471) );
  AND2_X1 U5679 ( .A1(n4810), .A2(n9188), .ZN(n4809) );
  NAND2_X1 U5680 ( .A1(n9226), .A2(n4811), .ZN(n9211) );
  NAND2_X1 U5681 ( .A1(n9226), .A2(n6520), .ZN(n9227) );
  NAND2_X1 U5682 ( .A1(n9274), .A2(n7765), .ZN(n9259) );
  NOR2_X1 U5683 ( .A1(n7640), .A2(n4813), .ZN(n9282) );
  NAND2_X1 U5684 ( .A1(n4815), .A2(n4814), .ZN(n4813) );
  INV_X1 U5685 ( .A(n4816), .ZN(n4815) );
  NOR2_X1 U5686 ( .A1(n9397), .A2(n9286), .ZN(n4814) );
  NAND2_X1 U5687 ( .A1(n9275), .A2(n9276), .ZN(n9274) );
  AND2_X1 U5688 ( .A1(n7764), .A2(n7765), .ZN(n9276) );
  NOR3_X1 U5689 ( .A1(n7640), .A2(n4816), .A3(n9397), .ZN(n9293) );
  NOR2_X1 U5690 ( .A1(n7640), .A2(n4816), .ZN(n9319) );
  NAND2_X1 U5691 ( .A1(n4408), .A2(n7865), .ZN(n4736) );
  OR2_X1 U5692 ( .A1(n4347), .A2(n9402), .ZN(n7640) );
  AND2_X1 U5693 ( .A1(n5728), .A2(n9747), .ZN(n6489) );
  NAND2_X1 U5694 ( .A1(n7392), .A2(n7874), .ZN(n7525) );
  NAND2_X1 U5695 ( .A1(n9660), .A2(n7751), .ZN(n7390) );
  NAND2_X1 U5696 ( .A1(n6507), .A2(n7960), .ZN(n7392) );
  NOR2_X1 U5697 ( .A1(n5367), .A2(n7588), .ZN(n5391) );
  NOR3_X1 U5698 ( .A1(n9708), .A2(n9665), .A3(n9691), .ZN(n9669) );
  NOR2_X1 U5699 ( .A1(n9708), .A2(n9691), .ZN(n9687) );
  NOR2_X1 U5700 ( .A1(n6499), .A2(n6500), .ZN(n6506) );
  INV_X1 U5701 ( .A(n7747), .ZN(n6505) );
  INV_X1 U5702 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7499) );
  AND2_X1 U5703 ( .A1(n5310), .A2(n5309), .ZN(n7426) );
  NAND2_X1 U5704 ( .A1(n7227), .A2(n9809), .ZN(n9707) );
  AND2_X1 U5705 ( .A1(n7253), .A2(n9802), .ZN(n7227) );
  AOI21_X1 U5706 ( .B1(n7954), .B2(n4914), .A(n4398), .ZN(n4913) );
  INV_X1 U5707 ( .A(n6436), .ZN(n4914) );
  NOR2_X1 U5708 ( .A1(n9733), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U5709 ( .A1(n7741), .A2(n7823), .ZN(n7813) );
  NOR2_X1 U5710 ( .A1(n9733), .A2(n9786), .ZN(n4806) );
  OR2_X1 U5711 ( .A1(n9733), .A2(n6784), .ZN(n6923) );
  OR2_X1 U5712 ( .A1(n7980), .A2(n5737), .ZN(n9008) );
  OR2_X1 U5713 ( .A1(n7980), .A2(n6647), .ZN(n9006) );
  INV_X1 U5714 ( .A(n7182), .ZN(n9802) );
  AND2_X1 U5715 ( .A1(n9763), .A2(n8008), .ZN(n9787) );
  INV_X1 U5716 ( .A(n9740), .ZN(n9767) );
  INV_X1 U5717 ( .A(n9787), .ZN(n9846) );
  AND2_X1 U5718 ( .A1(n7319), .A2(n5720), .ZN(n9763) );
  AND2_X1 U5719 ( .A1(n7529), .A2(n9765), .ZN(n9791) );
  XNOR2_X1 U5720 ( .A(n7790), .B(n7789), .ZN(n7783) );
  INV_X1 U5721 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5099) );
  NOR2_X1 U5722 ( .A1(n4775), .A2(n5071), .ZN(n4774) );
  NAND2_X1 U5723 ( .A1(n5073), .A2(n5066), .ZN(n4775) );
  NOR2_X1 U5724 ( .A1(n5088), .A2(n5087), .ZN(n4564) );
  NAND2_X1 U5725 ( .A1(n5470), .A2(n5070), .ZN(n5088) );
  NAND2_X1 U5726 ( .A1(n4856), .A2(n4854), .ZN(n5495) );
  INV_X1 U5727 ( .A(n4857), .ZN(n4854) );
  NAND2_X1 U5728 ( .A1(n5403), .A2(n5035), .ZN(n5113) );
  AND2_X1 U5729 ( .A1(n5035), .A2(n5034), .ZN(n5400) );
  OAI21_X1 U5730 ( .B1(n4842), .B2(n4840), .A(n4404), .ZN(n4838) );
  NAND2_X1 U5731 ( .A1(n5289), .A2(n5016), .ZN(n5301) );
  AND2_X1 U5732 ( .A1(n5011), .A2(n5010), .ZN(n5270) );
  AND2_X1 U5733 ( .A1(n5006), .A2(n5005), .ZN(n5239) );
  NAND2_X1 U5734 ( .A1(n5198), .A2(n5000), .ZN(n5222) );
  AND3_X1 U5735 ( .A1(n4667), .A2(n5133), .A3(n4665), .ZN(n6626) );
  NAND2_X1 U5736 ( .A1(n4407), .A2(P1_IR_REG_1__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U5737 ( .A1(n4666), .A2(n5360), .ZN(n4665) );
  AND4_X1 U5738 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(n8658)
         );
  NAND2_X1 U5739 ( .A1(n4490), .A2(n4935), .ZN(n4489) );
  AOI21_X1 U5740 ( .B1(n6932), .B2(n4935), .A(n4356), .ZN(n4933) );
  NAND2_X1 U5741 ( .A1(n7402), .A2(n6336), .ZN(n7506) );
  NAND2_X1 U5742 ( .A1(n4354), .A2(n4428), .ZN(n4514) );
  NAND2_X1 U5743 ( .A1(n8244), .A2(n4386), .ZN(n4515) );
  AND2_X1 U5744 ( .A1(n4951), .A2(n4950), .ZN(n8314) );
  AND2_X1 U5745 ( .A1(n4951), .A2(n4383), .ZN(n8270) );
  NAND2_X1 U5746 ( .A1(n6329), .A2(n6328), .ZN(n7192) );
  AND3_X1 U5747 ( .A1(n6049), .A2(n6048), .A3(n6047), .ZN(n8636) );
  NAND2_X1 U5748 ( .A1(n6070), .A2(n6069), .ZN(n8756) );
  NAND2_X1 U5749 ( .A1(n7401), .A2(n7403), .ZN(n7402) );
  AND2_X1 U5750 ( .A1(n6389), .A2(n6390), .ZN(n8318) );
  NAND2_X1 U5751 ( .A1(n6379), .A2(n6378), .ZN(n8315) );
  OR2_X1 U5752 ( .A1(n6391), .A2(n6390), .ZN(n8320) );
  NAND2_X1 U5753 ( .A1(n6321), .A2(n6320), .ZN(n6934) );
  INV_X1 U5754 ( .A(n8318), .ZN(n8335) );
  NAND2_X1 U5755 ( .A1(n6387), .A2(n9936), .ZN(n8250) );
  NAND2_X1 U5756 ( .A1(n7719), .A2(n6374), .ZN(n7710) );
  NAND2_X1 U5757 ( .A1(n8233), .A2(n4429), .ZN(n8330) );
  NAND2_X1 U5758 ( .A1(n8233), .A2(n6342), .ZN(n8329) );
  INV_X1 U5759 ( .A(n8320), .ZN(n8338) );
  AOI21_X1 U5760 ( .B1(n4702), .B2(n4700), .A(n4955), .ZN(n8063) );
  AND2_X1 U5761 ( .A1(n8061), .A2(n4701), .ZN(n4700) );
  XNOR2_X1 U5762 ( .A(n6155), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8229) );
  INV_X1 U5763 ( .A(n8248), .ZN(n8605) );
  NAND4_X1 U5764 ( .A1(n5911), .A2(n5910), .A3(n5909), .A4(n5908), .ZN(n8352)
         );
  OR2_X1 U5765 ( .A1(n6537), .A2(n6536), .ZN(n8507) );
  NAND2_X1 U5766 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4590) );
  NAND2_X1 U5767 ( .A1(n6711), .A2(n5793), .ZN(n6702) );
  AOI21_X1 U5768 ( .B1(n6699), .B2(n6698), .A(n6750), .ZN(n6701) );
  NAND2_X1 U5769 ( .A1(n4825), .A2(n4824), .ZN(n6797) );
  AOI21_X1 U5770 ( .B1(n7036), .B2(n7035), .A(n7034), .ZN(n7119) );
  NAND2_X1 U5771 ( .A1(n4349), .A2(n4728), .ZN(n4975) );
  INV_X1 U5772 ( .A(n4747), .ZN(n7359) );
  NAND2_X1 U5773 ( .A1(n4745), .A2(n4744), .ZN(n7442) );
  NOR2_X1 U5774 ( .A1(n7376), .A2(n7375), .ZN(n7433) );
  XNOR2_X1 U5775 ( .A(n8439), .B(n8455), .ZN(n8417) );
  NOR2_X1 U5776 ( .A1(n8443), .A2(n8442), .ZN(n8467) );
  OR2_X1 U5777 ( .A1(P2_U3150), .A2(n6604), .ZN(n9899) );
  INV_X1 U5778 ( .A(n4818), .ZN(n8470) );
  XNOR2_X1 U5779 ( .A(n4708), .B(n8480), .ZN(n8468) );
  NOR2_X1 U5780 ( .A1(n8525), .A2(n8524), .ZN(n8526) );
  NAND2_X1 U5781 ( .A1(n6118), .A2(n6126), .ZN(n8574) );
  OR2_X1 U5782 ( .A1(n9989), .A2(n8222), .ZN(n8709) );
  NAND2_X1 U5783 ( .A1(n5915), .A2(n5914), .ZN(n9986) );
  NAND2_X1 U5784 ( .A1(n5901), .A2(n5900), .ZN(n9980) );
  NAND2_X1 U5785 ( .A1(n6219), .A2(n8071), .ZN(n7207) );
  NAND2_X1 U5786 ( .A1(n6959), .A2(n8092), .ZN(n7089) );
  INV_X1 U5787 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6985) );
  OR2_X1 U5788 ( .A1(n5824), .A2(n4982), .ZN(n4614) );
  NAND2_X1 U5789 ( .A1(n6386), .A2(n6559), .ZN(n9936) );
  INV_X1 U5790 ( .A(n9989), .ZN(n9987) );
  INV_X1 U5791 ( .A(n9936), .ZN(n8729) );
  NAND2_X1 U5792 ( .A1(n4676), .A2(n8194), .ZN(n8568) );
  NAND2_X1 U5793 ( .A1(n6231), .A2(n4680), .ZN(n4676) );
  NAND2_X1 U5794 ( .A1(n6103), .A2(n6102), .ZN(n8803) );
  NAND2_X1 U5795 ( .A1(n6231), .A2(n8189), .ZN(n8584) );
  NAND2_X1 U5796 ( .A1(n6091), .A2(n6090), .ZN(n8809) );
  NAND2_X1 U5797 ( .A1(n6060), .A2(n6059), .ZN(n8825) );
  NAND2_X1 U5798 ( .A1(n6051), .A2(n6050), .ZN(n8831) );
  NAND2_X1 U5799 ( .A1(n4691), .A2(n4689), .ZN(n8648) );
  AND2_X1 U5800 ( .A1(n4691), .A2(n4379), .ZN(n8649) );
  OR2_X1 U5801 ( .A1(n8674), .A2(n4368), .ZN(n4691) );
  NAND2_X1 U5802 ( .A1(n6002), .A2(n6001), .ZN(n8842) );
  NAND2_X1 U5803 ( .A1(n4618), .A2(n5983), .ZN(n8698) );
  NAND2_X1 U5804 ( .A1(n5972), .A2(n4621), .ZN(n4618) );
  NAND2_X1 U5805 ( .A1(n5976), .A2(n5975), .ZN(n8326) );
  NAND2_X1 U5806 ( .A1(n5972), .A2(n5971), .ZN(n7696) );
  NAND2_X1 U5807 ( .A1(n4693), .A2(n8138), .ZN(n7617) );
  OR2_X1 U5808 ( .A1(n4699), .A2(n4697), .ZN(n4693) );
  NAND2_X1 U5809 ( .A1(n5952), .A2(n5951), .ZN(n7606) );
  OR2_X1 U5810 ( .A1(n4699), .A2(n4696), .ZN(n7597) );
  INV_X1 U5811 ( .A(n8133), .ZN(n4696) );
  INV_X1 U5812 ( .A(n4699), .ZN(n7536) );
  AND2_X1 U5813 ( .A1(n6533), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6584) );
  NAND2_X1 U5814 ( .A1(n8860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5767) );
  AND2_X1 U5815 ( .A1(n4348), .A2(n4953), .ZN(n4704) );
  INV_X1 U5816 ( .A(n6187), .ZN(n7622) );
  INV_X1 U5817 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10086) );
  INV_X1 U5818 ( .A(n6296), .ZN(n8072) );
  NAND2_X1 U5819 ( .A1(n4597), .A2(n4601), .ZN(n6154) );
  OR2_X1 U5820 ( .A1(n6024), .A2(n4603), .ZN(n4597) );
  INV_X1 U5821 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6943) );
  INV_X1 U5822 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U5823 ( .A1(n5859), .A2(n5880), .ZN(n7043) );
  INV_X1 U5824 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4977) );
  AND2_X1 U5825 ( .A1(n7615), .A2(n7576), .ZN(n4565) );
  XNOR2_X1 U5826 ( .A(n5717), .B(n5716), .ZN(n6569) );
  NAND2_X1 U5827 ( .A1(n4759), .A2(n5695), .ZN(n4758) );
  NAND2_X1 U5828 ( .A1(n4761), .A2(n4762), .ZN(n4759) );
  AOI21_X1 U5829 ( .B1(n7323), .B2(n4370), .A(n4781), .ZN(n7463) );
  INV_X1 U5830 ( .A(n4760), .ZN(n9002) );
  OR2_X1 U5831 ( .A1(n5466), .A2(n5465), .ZN(n5467) );
  INV_X1 U5832 ( .A(n6895), .ZN(n5230) );
  NAND2_X1 U5833 ( .A1(n4751), .A2(n5210), .ZN(n6896) );
  AOI22_X1 U5834 ( .A1(n5500), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6568), .B2(
        n7000), .ZN(n5321) );
  AND2_X1 U5835 ( .A1(n5517), .A2(n5516), .ZN(n9265) );
  AND2_X1 U5836 ( .A1(n5394), .A2(n5393), .ZN(n7585) );
  AND2_X1 U5837 ( .A1(n8869), .A2(n4416), .ZN(n8977) );
  NAND2_X1 U5838 ( .A1(n4752), .A2(n7077), .ZN(n7151) );
  NAND2_X1 U5839 ( .A1(n5736), .A2(n5735), .ZN(n9030) );
  NAND4_X1 U5840 ( .A1(n5236), .A2(n5235), .A3(n5234), .A4(n5233), .ZN(n9056)
         );
  NAND2_X1 U5841 ( .A1(n9479), .A2(n6631), .ZN(n6674) );
  NAND2_X1 U5842 ( .A1(n6674), .A2(n6675), .ZN(n6673) );
  NOR2_X1 U5843 ( .A1(n9497), .A2(n4512), .ZN(n6645) );
  AND2_X1 U5844 ( .A1(n6644), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5845 ( .A1(n6645), .A2(n6646), .ZN(n6999) );
  OR2_X1 U5846 ( .A1(n9630), .A2(n4508), .ZN(n9094) );
  NAND2_X1 U5847 ( .A1(n4509), .A2(n9070), .ZN(n4508) );
  INV_X1 U5848 ( .A(n9068), .ZN(n4509) );
  AND2_X1 U5849 ( .A1(n4671), .A2(n4371), .ZN(n9083) );
  OAI21_X1 U5850 ( .B1(n9114), .B2(n9644), .A(n9625), .ZN(n9115) );
  NAND2_X1 U5851 ( .A1(n4787), .A2(n9332), .ZN(n4786) );
  NOR2_X1 U5852 ( .A1(n9343), .A2(n9754), .ZN(n6529) );
  NOR2_X1 U5853 ( .A1(n9191), .A2(n9190), .ZN(n9189) );
  NAND2_X1 U5854 ( .A1(n4921), .A2(n4923), .ZN(n9197) );
  NAND2_X1 U5855 ( .A1(n9225), .A2(n4924), .ZN(n4921) );
  NAND2_X1 U5856 ( .A1(n4734), .A2(n4369), .ZN(n9216) );
  AND2_X1 U5857 ( .A1(n4734), .A2(n7730), .ZN(n9217) );
  NAND2_X1 U5858 ( .A1(n4927), .A2(n6467), .ZN(n9210) );
  NAND2_X1 U5859 ( .A1(n9225), .A2(n4928), .ZN(n4927) );
  INV_X1 U5860 ( .A(n9265), .ZN(n9386) );
  NAND2_X1 U5861 ( .A1(n7628), .A2(n7872), .ZN(n9308) );
  NAND2_X1 U5862 ( .A1(n6940), .A2(n7782), .ZN(n5472) );
  NAND2_X1 U5863 ( .A1(n9666), .A2(n9667), .ZN(n4909) );
  NAND2_X1 U5864 ( .A1(n7225), .A2(n7226), .ZN(n4903) );
  NAND2_X1 U5865 ( .A1(n6969), .A2(n6970), .ZN(n4915) );
  OR2_X1 U5866 ( .A1(n7261), .A2(n9423), .ZN(n9315) );
  NAND2_X1 U5867 ( .A1(n4749), .A2(n7821), .ZN(n6917) );
  OR2_X1 U5868 ( .A1(n6521), .A2(n9747), .ZN(n9694) );
  INV_X1 U5869 ( .A(n9694), .ZN(n9738) );
  INV_X1 U5870 ( .A(n9720), .ZN(n9739) );
  INV_X1 U5871 ( .A(n9315), .ZN(n9749) );
  AND2_X2 U5872 ( .A1(n9336), .A2(n9335), .ZN(n10233) );
  AND2_X1 U5873 ( .A1(n4932), .A2(n5059), .ZN(n4931) );
  NOR2_X1 U5874 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(n5063), .ZN(n4932) );
  OAI21_X1 U5875 ( .B1(n7790), .B2(n7789), .A(n7788), .ZN(n7794) );
  NAND2_X1 U5876 ( .A1(n5083), .A2(n5065), .ZN(n4707) );
  XNOR2_X1 U5877 ( .A(n5083), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7615) );
  INV_X1 U5878 ( .A(n4864), .ZN(n5599) );
  XNOR2_X1 U5879 ( .A(n5714), .B(n5713), .ZN(n7319) );
  NOR2_X1 U5880 ( .A1(n5071), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4773) );
  INV_X1 U5881 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6858) );
  NOR2_X1 U5882 ( .A1(n4916), .A2(n4918), .ZN(n5116) );
  INV_X1 U5883 ( .A(n5053), .ZN(n4916) );
  NAND2_X1 U5884 ( .A1(n4880), .A2(n4879), .ZN(n5385) );
  NAND2_X1 U5885 ( .A1(n4880), .A2(n4881), .ZN(n5384) );
  INV_X1 U5886 ( .A(n6626), .ZN(n9537) );
  NAND2_X1 U5887 ( .A1(n4650), .A2(n8359), .ZN(n8366) );
  INV_X1 U5888 ( .A(n4720), .ZN(n8394) );
  AOI21_X1 U5889 ( .B1(n8515), .B2(n9919), .A(n4594), .ZN(n8516) );
  NAND2_X1 U5890 ( .A1(n4656), .A2(n4394), .ZN(n4594) );
  AND2_X1 U5891 ( .A1(n4637), .A2(n6168), .ZN(n8553) );
  INV_X1 U5892 ( .A(n6285), .ZN(n6286) );
  OAI22_X1 U5893 ( .A1(n7689), .A2(n8737), .B1(n10008), .B2(n6284), .ZN(n6285)
         );
  OR2_X1 U5894 ( .A1(n8550), .A2(n8783), .ZN(n6251) );
  INV_X1 U5895 ( .A(n6290), .ZN(n6291) );
  OAI21_X1 U5896 ( .B1(n7689), .B2(n8834), .A(n6289), .ZN(n6290) );
  OR2_X1 U5897 ( .A1(n8550), .A2(n8858), .ZN(n6237) );
  NAND2_X1 U5898 ( .A1(n9997), .A2(n6212), .ZN(n4640) );
  OAI211_X1 U5899 ( .C1(n4522), .C2(n7999), .A(n4521), .B(n4518), .ZN(P1_U3242) );
  NAND2_X1 U5900 ( .A1(n8011), .A2(n4524), .ZN(n4521) );
  INV_X1 U5901 ( .A(n4519), .ZN(n4518) );
  OR3_X1 U5902 ( .A1(n9708), .A2(n4768), .A3(n7560), .ZN(n4347) );
  OR2_X1 U5903 ( .A1(n7039), .A2(n7044), .ZN(n4349) );
  AND2_X1 U5904 ( .A1(n9188), .A2(n9041), .ZN(n7921) );
  AND2_X1 U5905 ( .A1(n5069), .A2(n5068), .ZN(n9297) );
  INV_X1 U5906 ( .A(n9297), .ZN(n9397) );
  INV_X1 U5907 ( .A(n5150), .ZN(n5524) );
  INV_X2 U5908 ( .A(n5524), .ZN(n5244) );
  OR2_X1 U5909 ( .A1(n8640), .A2(n8632), .ZN(n4351) );
  AND2_X1 U5910 ( .A1(n8697), .A2(n4619), .ZN(n4352) );
  OR2_X1 U5911 ( .A1(n8142), .A2(n8141), .ZN(n4353) );
  OR2_X1 U5912 ( .A1(n7722), .A2(n7721), .ZN(n4354) );
  OR2_X1 U5913 ( .A1(n5937), .A2(n4961), .ZN(n4355) );
  AND2_X1 U5914 ( .A1(n6325), .A2(n7141), .ZN(n4356) );
  NOR2_X1 U5915 ( .A1(n7322), .A2(n7327), .ZN(n4357) );
  AND2_X1 U5916 ( .A1(n9839), .A2(n4769), .ZN(n4358) );
  NAND2_X1 U5917 ( .A1(n4794), .A2(n5574), .ZN(n8869) );
  INV_X1 U5918 ( .A(n7948), .ZN(n6970) );
  AND2_X1 U5919 ( .A1(n7816), .A2(n7814), .ZN(n7948) );
  NAND2_X1 U5920 ( .A1(n9001), .A2(n9004), .ZN(n4359) );
  NOR2_X1 U5921 ( .A1(n8040), .A2(n4685), .ZN(n4360) );
  AND2_X1 U5922 ( .A1(n7904), .A2(n7937), .ZN(n4361) );
  AND2_X1 U5923 ( .A1(n5632), .A2(n5631), .ZN(n9188) );
  INV_X1 U5924 ( .A(n9188), .ZN(n9361) );
  AND2_X1 U5925 ( .A1(n4953), .A2(n5768), .ZN(n4362) );
  INV_X1 U5926 ( .A(n8557), .ZN(n8579) );
  NAND2_X1 U5927 ( .A1(n6374), .A2(n8579), .ZN(n4363) );
  AND2_X1 U5928 ( .A1(n4576), .A2(n4575), .ZN(n4364) );
  AND2_X1 U5929 ( .A1(n4806), .A2(n4807), .ZN(n4365) );
  NAND2_X1 U5930 ( .A1(n5390), .A2(n5389), .ZN(n9665) );
  NOR2_X1 U5931 ( .A1(n9708), .A2(n4768), .ZN(n4767) );
  AND2_X1 U5932 ( .A1(n4579), .A2(n4578), .ZN(n4366) );
  XNOR2_X1 U5933 ( .A(n5077), .B(n5073), .ZN(n5749) );
  XNOR2_X1 U5934 ( .A(n6152), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6296) );
  OR2_X1 U5935 ( .A1(n5827), .A2(n9912), .ZN(n4367) );
  OR2_X1 U5936 ( .A1(n8675), .A2(n6227), .ZN(n4368) );
  OR2_X1 U5937 ( .A1(n9376), .A2(n8918), .ZN(n7730) );
  NAND2_X1 U5938 ( .A1(n5827), .A2(n4992), .ZN(n5842) );
  AND4_X1 U5939 ( .A1(n4958), .A2(n5819), .A3(n5818), .A4(n5817), .ZN(n6312)
         );
  INV_X1 U5940 ( .A(n5159), .ZN(n5546) );
  AND2_X1 U5941 ( .A1(n9218), .A2(n7730), .ZN(n4369) );
  NAND2_X1 U5942 ( .A1(n5052), .A2(n5051), .ZN(n5218) );
  AND2_X1 U5943 ( .A1(n5382), .A2(n4784), .ZN(n4370) );
  NAND4_X1 U5944 ( .A1(n5798), .A2(n5797), .A3(n5796), .A4(n5795), .ZN(n8357)
         );
  AOI21_X1 U5945 ( .B1(n8872), .B2(n4761), .A(n4758), .ZN(n4757) );
  OR2_X1 U5946 ( .A1(n9080), .A2(n9079), .ZN(n4371) );
  OR2_X1 U5947 ( .A1(n5399), .A2(n5398), .ZN(n4372) );
  NAND2_X1 U5948 ( .A1(n6712), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4373) );
  AND2_X1 U5949 ( .A1(n6023), .A2(n6037), .ZN(n4374) );
  OR2_X2 U5950 ( .A1(n7997), .A2(n9747), .ZN(n4375) );
  AND4_X1 U5951 ( .A1(n5787), .A2(n5786), .A3(n5785), .A4(n5784), .ZN(n4376)
         );
  OR2_X1 U5952 ( .A1(n8009), .A2(n8008), .ZN(n4377) );
  NAND2_X1 U5953 ( .A1(n5564), .A2(n5563), .ZN(n9376) );
  OR2_X1 U5954 ( .A1(n9207), .A2(n8928), .ZN(n4378) );
  OR2_X1 U5955 ( .A1(n6227), .A2(n8676), .ZN(n4379) );
  NAND2_X1 U5956 ( .A1(n7797), .A2(n7796), .ZN(n9332) );
  INV_X1 U5957 ( .A(n9332), .ZN(n4790) );
  INV_X1 U5958 ( .A(n6499), .ZN(n7744) );
  INV_X1 U5959 ( .A(n6869), .ZN(n6861) );
  OR2_X1 U5960 ( .A1(n5841), .A2(n5840), .ZN(n6869) );
  AOI21_X1 U5961 ( .B1(n7783), .B2(n8025), .A(n7668), .ZN(n8027) );
  INV_X1 U5962 ( .A(n8071), .ZN(n4685) );
  AND4_X1 U5963 ( .A1(n5055), .A2(n5713), .A3(n5073), .A4(n5091), .ZN(n4380)
         );
  AND2_X1 U5964 ( .A1(n6628), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4381) );
  OR3_X1 U5965 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U5966 ( .A1(n6347), .A2(n8686), .ZN(n4383) );
  AND2_X1 U5967 ( .A1(n5040), .A2(n4483), .ZN(n4384) );
  NOR2_X1 U5968 ( .A1(n8631), .A2(n8640), .ZN(n4385) );
  AND2_X1 U5969 ( .A1(n7903), .A2(n9241), .ZN(n4472) );
  AND2_X1 U5970 ( .A1(n8277), .A2(n4354), .ZN(n4386) );
  OR2_X1 U5971 ( .A1(n9058), .A2(n9780), .ZN(n4387) );
  NAND2_X1 U5972 ( .A1(n7785), .A2(n7784), .ZN(n9135) );
  NAND2_X1 U5973 ( .A1(n5799), .A2(n5800), .ZN(n5808) );
  INV_X1 U5974 ( .A(n5052), .ZN(n5216) );
  AND2_X1 U5975 ( .A1(n6319), .A2(n6963), .ZN(n4388) );
  NAND2_X1 U5976 ( .A1(n9931), .A2(n7216), .ZN(n4389) );
  INV_X1 U5977 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5360) );
  NOR2_X1 U5978 ( .A1(n8831), .A2(n8624), .ZN(n4390) );
  AND2_X1 U5979 ( .A1(n5502), .A2(n5501), .ZN(n9392) );
  INV_X1 U5980 ( .A(n9392), .ZN(n9286) );
  NOR2_X1 U5981 ( .A1(n8030), .A2(n8212), .ZN(n4391) );
  AND2_X1 U5982 ( .A1(n8848), .A2(n8686), .ZN(n4392) );
  INV_X1 U5983 ( .A(n6932), .ZN(n6320) );
  AND2_X1 U5984 ( .A1(n4723), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4393) );
  INV_X1 U5985 ( .A(n6468), .ZN(n4928) );
  NOR2_X1 U5986 ( .A1(n6520), .A2(n8918), .ZN(n6468) );
  AND2_X1 U5987 ( .A1(n4654), .A2(n4653), .ZN(n4394) );
  INV_X1 U5988 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6037) );
  AND2_X1 U5989 ( .A1(n9839), .A2(n7558), .ZN(n4395) );
  NOR2_X1 U5990 ( .A1(n5381), .A2(n5380), .ZN(n4396) );
  NOR2_X1 U5991 ( .A1(n4343), .A2(n9052), .ZN(n4397) );
  AND2_X1 U5992 ( .A1(n7165), .A2(n9721), .ZN(n4398) );
  AND2_X1 U5993 ( .A1(n8134), .A2(n8135), .ZN(n4399) );
  INV_X1 U5994 ( .A(n6708), .ZN(n4827) );
  INV_X1 U5995 ( .A(n4882), .ZN(n4881) );
  NOR2_X1 U5996 ( .A1(n5028), .A2(SI_11_), .ZN(n4882) );
  XNOR2_X1 U5997 ( .A(n7662), .B(SI_29_), .ZN(n6474) );
  OR2_X1 U5998 ( .A1(n8871), .A2(n8870), .ZN(n4400) );
  AND2_X1 U5999 ( .A1(n4600), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4401) );
  AND4_X1 U6000 ( .A1(n5807), .A2(n5806), .A3(n5805), .A4(n5804), .ZN(n8719)
         );
  INV_X1 U6001 ( .A(n8719), .ZN(n8356) );
  INV_X1 U6002 ( .A(n9780), .ZN(n6926) );
  AND3_X1 U6003 ( .A1(n5203), .A2(n5202), .A3(n5201), .ZN(n9780) );
  AND2_X1 U6004 ( .A1(n5019), .A2(n5018), .ZN(n4402) );
  AND2_X1 U6005 ( .A1(n4853), .A2(n4850), .ZN(n4403) );
  OR2_X1 U6006 ( .A1(n5021), .A2(SI_9_), .ZN(n4404) );
  OR2_X1 U6007 ( .A1(n6868), .A2(n6794), .ZN(n4405) );
  AND2_X1 U6008 ( .A1(n8033), .A2(n8029), .ZN(n4406) );
  NAND2_X1 U6009 ( .A1(n5783), .A2(n5782), .ZN(n6300) );
  AND2_X1 U6010 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4407) );
  INV_X1 U6011 ( .A(n4765), .ZN(n4764) );
  OR2_X1 U6012 ( .A1(n4964), .A2(n4766), .ZN(n4765) );
  OR2_X1 U6013 ( .A1(n7963), .A2(n4737), .ZN(n4408) );
  OR2_X1 U6014 ( .A1(n4930), .A2(n4926), .ZN(n4409) );
  INV_X1 U6015 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5758) );
  AND2_X1 U6016 ( .A1(n4851), .A2(n4850), .ZN(n4410) );
  AND2_X1 U6017 ( .A1(n8168), .A2(n8170), .ZN(n8654) );
  AND2_X1 U6018 ( .A1(n4792), .A2(n4790), .ZN(n4411) );
  INV_X1 U6019 ( .A(n7127), .ZN(n4729) );
  AND3_X1 U6020 ( .A1(n8167), .A2(n8166), .A3(n8165), .ZN(n4412) );
  INV_X1 U6021 ( .A(n9346), .ZN(n9139) );
  NAND2_X1 U6022 ( .A1(n6428), .A2(n6427), .ZN(n9346) );
  AND2_X1 U6023 ( .A1(n7960), .A2(n7865), .ZN(n4413) );
  OR2_X1 U6024 ( .A1(n4353), .A2(n8136), .ZN(n4414) );
  AND2_X1 U6025 ( .A1(n4959), .A2(n8092), .ZN(n4415) );
  INV_X1 U6026 ( .A(n9224), .ZN(n9234) );
  AND2_X1 U6027 ( .A1(n7730), .A2(n7770), .ZN(n9224) );
  AND2_X1 U6028 ( .A1(n4800), .A2(n4803), .ZN(n4416) );
  AND2_X1 U6029 ( .A1(n6330), .A2(n6328), .ZN(n4417) );
  OR2_X1 U6030 ( .A1(n9352), .A2(n9007), .ZN(n7925) );
  NAND2_X1 U6031 ( .A1(n6799), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4418) );
  INV_X1 U6032 ( .A(n6265), .ZN(n6158) );
  AND2_X1 U6033 ( .A1(n4613), .A2(n4612), .ZN(n4419) );
  AND2_X1 U6034 ( .A1(n4360), .A2(n8108), .ZN(n4420) );
  AND2_X1 U6035 ( .A1(n4919), .A2(n4378), .ZN(n4421) );
  INV_X1 U6036 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5074) );
  AND2_X1 U6037 ( .A1(n5778), .A2(n4954), .ZN(n4953) );
  AND2_X1 U6038 ( .A1(n4827), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4422) );
  OR2_X1 U6039 ( .A1(n8209), .A2(n4582), .ZN(n4423) );
  INV_X1 U6040 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4566) );
  INV_X1 U6041 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U6042 ( .A1(n4782), .A2(n4785), .ZN(n7496) );
  NAND2_X1 U6043 ( .A1(n4897), .A2(n4900), .ZN(n9673) );
  INV_X1 U6044 ( .A(n4592), .ZN(n6714) );
  NOR2_X1 U6045 ( .A1(n9293), .A2(n9292), .ZN(n4424) );
  INV_X1 U6046 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4476) );
  AND2_X1 U6047 ( .A1(n6641), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4425) );
  NOR2_X1 U6048 ( .A1(n4589), .A2(n8387), .ZN(n8406) );
  INV_X1 U6049 ( .A(n8406), .ZN(n4588) );
  INV_X1 U6050 ( .A(n5042), .ZN(n4860) );
  OR2_X1 U6051 ( .A1(n7447), .A2(n7361), .ZN(n4426) );
  INV_X1 U6052 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4954) );
  INV_X1 U6053 ( .A(n8979), .ZN(n4803) );
  NAND2_X1 U6054 ( .A1(n5896), .A2(n4613), .ZN(n5937) );
  NOR2_X1 U6055 ( .A1(n5949), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U6056 ( .A1(n9226), .A2(n4810), .ZN(n4812) );
  INV_X1 U6057 ( .A(n7560), .ZN(n9847) );
  NAND2_X1 U6058 ( .A1(n5119), .A2(n5118), .ZN(n7560) );
  NAND2_X1 U6059 ( .A1(n5679), .A2(n5678), .ZN(n9352) );
  OR2_X1 U6060 ( .A1(n6338), .A2(n7569), .ZN(n4427) );
  NAND2_X1 U6061 ( .A1(n8278), .A2(n6372), .ZN(n4428) );
  AND2_X1 U6062 ( .A1(n6343), .A2(n6342), .ZN(n4429) );
  AND2_X1 U6063 ( .A1(n4650), .A2(n4649), .ZN(n4430) );
  INV_X1 U6064 ( .A(n4351), .ZN(n4625) );
  INV_X1 U6065 ( .A(n4571), .ZN(n6126) );
  NOR2_X1 U6066 ( .A1(n6117), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n4571) );
  NAND2_X1 U6067 ( .A1(n6017), .A2(n6019), .ZN(n4431) );
  AND2_X1 U6068 ( .A1(n5493), .A2(SI_18_), .ZN(n4432) );
  AND2_X1 U6069 ( .A1(n6473), .A2(n9007), .ZN(n4433) );
  NAND2_X1 U6070 ( .A1(n5606), .A2(n5605), .ZN(n9367) );
  INV_X1 U6071 ( .A(n4817), .ZN(n9318) );
  NOR2_X1 U6072 ( .A1(n7640), .A2(n9512), .ZN(n4817) );
  INV_X1 U6073 ( .A(n9665), .ZN(n9833) );
  AND2_X1 U6074 ( .A1(n4624), .A2(n4351), .ZN(n4434) );
  AND2_X1 U6075 ( .A1(n4647), .A2(n4645), .ZN(n4435) );
  INV_X1 U6076 ( .A(n7379), .ZN(n4821) );
  NOR2_X1 U6077 ( .A1(n7447), .A2(n7459), .ZN(n7379) );
  NAND2_X1 U6078 ( .A1(n5322), .A2(n5321), .ZN(n9706) );
  INV_X1 U6079 ( .A(n4343), .ZN(n4569) );
  AOI21_X1 U6080 ( .B1(n8574), .B2(n6046), .A(n6121), .ZN(n8557) );
  INV_X1 U6081 ( .A(n9691), .ZN(n4769) );
  INV_X1 U6082 ( .A(n7226), .ZN(n4899) );
  NAND2_X1 U6083 ( .A1(n6219), .A2(n4360), .ZN(n7206) );
  AND2_X1 U6084 ( .A1(n7055), .A2(n6324), .ZN(n4935) );
  OAI211_X1 U6085 ( .C1(n4492), .C2(n4934), .A(n4933), .B(n4489), .ZN(n7135)
         );
  NAND2_X1 U6086 ( .A1(n4915), .A2(n6436), .ZN(n7248) );
  AND2_X1 U6087 ( .A1(n7149), .A2(n5281), .ZN(n7161) );
  NAND2_X1 U6088 ( .A1(n4903), .A2(n6439), .ZN(n7277) );
  NAND2_X1 U6089 ( .A1(n4909), .A2(n6451), .ZN(n7397) );
  NAND2_X1 U6090 ( .A1(n6934), .A2(n4935), .ZN(n7054) );
  NOR2_X1 U6091 ( .A1(n7433), .A2(n7432), .ZN(n4436) );
  AND2_X1 U6092 ( .A1(n4747), .A2(n7358), .ZN(n4437) );
  INV_X1 U6093 ( .A(n4767), .ZN(n4770) );
  AND2_X1 U6094 ( .A1(n4726), .A2(n4349), .ZN(n4438) );
  INV_X1 U6095 ( .A(n6168), .ZN(n4638) );
  INV_X1 U6096 ( .A(SI_15_), .ZN(n4887) );
  OR2_X1 U6097 ( .A1(n4808), .A2(n9733), .ZN(n4439) );
  XOR2_X1 U6098 ( .A(n9570), .B(n6993), .Z(n4440) );
  NOR2_X1 U6099 ( .A1(n6872), .A2(n6871), .ZN(n4441) );
  OR2_X1 U6100 ( .A1(n9559), .A2(n9560), .ZN(n4442) );
  AND2_X1 U6101 ( .A1(n4727), .A2(n4349), .ZN(n4443) );
  OR2_X1 U6102 ( .A1(n9542), .A2(n9541), .ZN(n4663) );
  NOR2_X1 U6103 ( .A1(n8014), .A2(n8013), .ZN(n4444) );
  OR2_X1 U6104 ( .A1(n9556), .A2(n9555), .ZN(n4661) );
  INV_X1 U6105 ( .A(n9774), .ZN(n6784) );
  AND2_X1 U6106 ( .A1(n4831), .A2(n4830), .ZN(n4445) );
  INV_X1 U6107 ( .A(n5749), .ZN(n8000) );
  INV_X1 U6108 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n4573) );
  INV_X1 U6109 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4581) );
  INV_X1 U6110 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4577) );
  INV_X1 U6111 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4837) );
  NAND2_X1 U6112 ( .A1(n7925), .A2(n7932), .ZN(n4542) );
  NAND2_X1 U6113 ( .A1(n7928), .A2(n7932), .ZN(n4536) );
  AOI21_X1 U6114 ( .B1(n7926), .B2(n7925), .A(n7932), .ZN(n4539) );
  NOR2_X1 U6115 ( .A1(n7876), .A2(n7932), .ZN(n4551) );
  AND2_X1 U6116 ( .A1(n7819), .A2(n7932), .ZN(n4530) );
  NAND2_X1 U6117 ( .A1(n4920), .A2(n4421), .ZN(n6470) );
  INV_X1 U6118 ( .A(n5287), .ZN(n4841) );
  NAND2_X1 U6119 ( .A1(n4896), .A2(n4895), .ZN(n4894) );
  NAND2_X1 U6120 ( .A1(n5195), .A2(n4999), .ZN(n5198) );
  OAI22_X1 U6121 ( .A1(n6472), .A2(n6471), .B1(n9361), .B2(n9041), .ZN(n9171)
         );
  NAND2_X1 U6122 ( .A1(n5401), .A2(n5400), .ZN(n5403) );
  NAND2_X1 U6123 ( .A1(n7627), .A2(n6457), .ZN(n6461) );
  NOR2_X1 U6124 ( .A1(n8105), .A2(n8206), .ZN(n4447) );
  NAND2_X1 U6125 ( .A1(n8121), .A2(n8219), .ZN(n4451) );
  OAI211_X1 U6126 ( .C1(n8106), .C2(n8219), .A(n8111), .B(n8112), .ZN(n4452)
         );
  NAND3_X1 U6127 ( .A1(n5898), .A2(n4952), .A3(n4348), .ZN(n6183) );
  NAND4_X1 U6128 ( .A1(n5898), .A2(n4952), .A3(n4348), .A4(n4362), .ZN(n8860)
         );
  NAND3_X1 U6129 ( .A1(n4456), .A2(n4455), .A3(n4454), .ZN(n4453) );
  NAND3_X1 U6130 ( .A1(n8087), .A2(n8091), .A3(n8219), .ZN(n4457) );
  NAND2_X2 U6131 ( .A1(n4615), .A2(n9948), .ZN(n8086) );
  NAND4_X1 U6132 ( .A1(n5756), .A2(n5800), .A3(n5780), .A4(n6712), .ZN(n5820)
         );
  NAND4_X1 U6133 ( .A1(n5756), .A2(n5838), .A3(n4462), .A4(n4461), .ZN(n4460)
         );
  NAND4_X1 U6134 ( .A1(n4464), .A2(n5800), .A3(n5780), .A4(n6712), .ZN(n4463)
         );
  NAND3_X1 U6135 ( .A1(n4466), .A2(n4465), .A3(n8220), .ZN(n4596) );
  NAND3_X1 U6136 ( .A1(n4873), .A2(n8217), .A3(n8218), .ZN(n4465) );
  NAND2_X1 U6137 ( .A1(n4412), .A2(n8176), .ZN(n4469) );
  NAND2_X1 U6138 ( .A1(n8163), .A2(n8176), .ZN(n4468) );
  NAND3_X1 U6139 ( .A1(n4469), .A2(n4468), .A3(n4608), .ZN(n4471) );
  NAND2_X1 U6140 ( .A1(n4470), .A2(n8182), .ZN(n8188) );
  NAND2_X1 U6141 ( .A1(n4471), .A2(n4607), .ZN(n4470) );
  NAND2_X2 U6142 ( .A1(n5273), .A2(n5011), .ZN(n5287) );
  NAND2_X2 U6143 ( .A1(n7983), .A2(n7904), .ZN(n9233) );
  INV_X1 U6144 ( .A(n4833), .ZN(n4473) );
  NAND2_X1 U6145 ( .A1(n4473), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4474) );
  NAND3_X1 U6146 ( .A1(n4835), .A2(n4833), .A3(P1_DATAO_REG_2__SCAN_IN), .ZN(
        n4475) );
  INV_X1 U6147 ( .A(n4985), .ZN(n4984) );
  NAND2_X1 U6148 ( .A1(n5178), .A2(n4996), .ZN(n5195) );
  NAND4_X1 U6149 ( .A1(n4480), .A2(n4479), .A3(n4478), .A4(n4477), .ZN(n6940)
         );
  NAND3_X1 U6150 ( .A1(n4384), .A2(n5469), .A3(n5039), .ZN(n4479) );
  OAI21_X2 U6151 ( .B1(n9202), .B2(n4486), .A(n4485), .ZN(n4484) );
  NOR2_X2 U6152 ( .A1(n9198), .A2(n7969), .ZN(n9202) );
  NAND2_X2 U6153 ( .A1(n4733), .A2(n4731), .ZN(n9198) );
  NAND2_X1 U6154 ( .A1(n6822), .A2(n6317), .ZN(n4492) );
  OAI21_X1 U6155 ( .B1(n6822), .B2(n6318), .A(n6317), .ZN(n6908) );
  INV_X1 U6156 ( .A(n6933), .ZN(n6321) );
  NOR2_X1 U6157 ( .A1(n4339), .A2(n4506), .ZN(n4504) );
  XNOR2_X1 U6158 ( .A(n9067), .B(n9079), .ZN(n9631) );
  NOR2_X1 U6159 ( .A1(n9630), .A2(n9068), .ZN(n9071) );
  AOI21_X2 U6160 ( .B1(n7682), .B2(n4942), .A(n4940), .ZN(n8293) );
  MUX2_X1 U6161 ( .A(n6624), .B(P1_REG1_REG_1__SCAN_IN), .S(n6626), .Z(n9530)
         );
  NAND2_X1 U6162 ( .A1(n8244), .A2(n8277), .ZN(n7720) );
  NAND2_X2 U6163 ( .A1(n4515), .A2(n4514), .ZN(n7719) );
  NOR2_X2 U6164 ( .A1(n4961), .A2(n4516), .ZN(n4952) );
  OAI21_X2 U6165 ( .B1(n4522), .B2(n4375), .A(n4520), .ZN(n4519) );
  OAI211_X1 U6166 ( .C1(n7932), .C2(n7819), .A(n4529), .B(n7818), .ZN(n7820)
         );
  NAND2_X1 U6167 ( .A1(n4530), .A2(n4531), .ZN(n4529) );
  AND2_X1 U6168 ( .A1(n7815), .A2(n7814), .ZN(n7828) );
  NAND3_X1 U6169 ( .A1(n4552), .A2(n4551), .A3(n4546), .ZN(n4545) );
  AOI21_X1 U6170 ( .B1(n7851), .B2(n7850), .A(n7849), .ZN(n7856) );
  NAND2_X1 U6171 ( .A1(n4555), .A2(n4554), .ZN(n4553) );
  INV_X1 U6172 ( .A(n7838), .ZN(n4554) );
  NAND4_X1 U6173 ( .A1(n7831), .A2(n7833), .A3(n7830), .A4(n7832), .ZN(n4555)
         );
  NAND3_X1 U6174 ( .A1(n9224), .A2(n7932), .A3(n7902), .ZN(n4558) );
  NOR2_X1 U6175 ( .A1(n4564), .A2(n5093), .ZN(n4563) );
  NAND2_X2 U6176 ( .A1(n8914), .A2(n8915), .ZN(n8913) );
  AND3_X2 U6177 ( .A1(n4567), .A2(n5053), .A3(n4566), .ZN(n5427) );
  NAND2_X1 U6178 ( .A1(n5427), .A2(n4773), .ZN(n5076) );
  XNOR2_X1 U6179 ( .A(n4568), .B(n8894), .ZN(n5332) );
  OAI21_X1 U6180 ( .B1(n5524), .B2(n4569), .A(n5329), .ZN(n4568) );
  NAND3_X1 U6181 ( .A1(n5813), .A2(n5829), .A3(n6985), .ZN(n5850) );
  NAND4_X1 U6182 ( .A1(n5813), .A2(n6985), .A3(n5829), .A4(n4581), .ZN(n5867)
         );
  NAND3_X1 U6183 ( .A1(n4824), .A2(n4418), .A3(n4825), .ZN(n4584) );
  NAND3_X1 U6184 ( .A1(n4422), .A2(n6707), .A3(n6706), .ZN(n4825) );
  NAND2_X1 U6185 ( .A1(n4585), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4587) );
  INV_X1 U6186 ( .A(n4585), .ZN(n7380) );
  INV_X1 U6187 ( .A(n4587), .ZN(n7484) );
  NAND2_X1 U6188 ( .A1(n6703), .A2(n4591), .ZN(n9894) );
  OAI21_X1 U6189 ( .B1(n4596), .B2(n4872), .A(n4595), .ZN(n8223) );
  OAI21_X1 U6190 ( .B1(n8137), .B2(n4414), .A(n4609), .ZN(n4611) );
  NAND2_X1 U6191 ( .A1(n5896), .A2(n4419), .ZN(n5949) );
  INV_X1 U6192 ( .A(n9948), .ZN(n6733) );
  NAND2_X1 U6193 ( .A1(n5972), .A2(n4352), .ZN(n4616) );
  NAND2_X1 U6194 ( .A1(n4616), .A2(n4617), .ZN(n8685) );
  NAND2_X1 U6195 ( .A1(n6012), .A2(n4626), .ZN(n4624) );
  OAI211_X1 U6196 ( .C1(n8724), .C2(n4629), .A(n5845), .B(n4627), .ZN(n4630)
         );
  NAND2_X1 U6197 ( .A1(n4639), .A2(n6265), .ZN(n4637) );
  NAND2_X1 U6198 ( .A1(n6158), .A2(n4635), .ZN(n4631) );
  OAI211_X1 U6199 ( .C1(n4639), .C2(n4632), .A(n4631), .B(n4640), .ZN(n6238)
         );
  OAI22_X2 U6200 ( .A1(n8589), .A2(n6101), .B1(n8605), .B2(n8809), .ZN(n8578)
         );
  NAND2_X1 U6201 ( .A1(n4642), .A2(n4641), .ZN(n5879) );
  NAND3_X1 U6202 ( .A1(n4643), .A2(n4952), .A3(n5778), .ZN(n5776) );
  INV_X1 U6203 ( .A(n8360), .ZN(n4652) );
  NAND2_X1 U6204 ( .A1(n9884), .A2(n9885), .ZN(n9883) );
  MUX2_X1 U6205 ( .A(n6692), .B(n6955), .S(n8530), .Z(n6693) );
  MUX2_X1 U6206 ( .A(n4668), .B(P1_REG2_REG_1__SCAN_IN), .S(n6626), .Z(n9524)
         );
  NAND2_X1 U6207 ( .A1(n4371), .A2(n9635), .ZN(n4670) );
  XNOR2_X1 U6208 ( .A(n9080), .B(n9079), .ZN(n9635) );
  INV_X1 U6209 ( .A(n4671), .ZN(n9633) );
  INV_X1 U6210 ( .A(n7654), .ZN(n5770) );
  NAND2_X1 U6211 ( .A1(n5885), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U6212 ( .A1(n6231), .A2(n4677), .ZN(n4673) );
  NAND2_X1 U6213 ( .A1(n4673), .A2(n4674), .ZN(n8561) );
  NAND2_X1 U6214 ( .A1(n6219), .A2(n4420), .ZN(n4682) );
  NAND2_X1 U6215 ( .A1(n4682), .A2(n4683), .ZN(n7265) );
  NAND2_X1 U6216 ( .A1(n8674), .A2(n4689), .ZN(n4686) );
  NAND2_X1 U6217 ( .A1(n4686), .A2(n4687), .ZN(n8642) );
  NAND2_X1 U6218 ( .A1(n6959), .A2(n4415), .ZN(n9923) );
  NAND2_X1 U6219 ( .A1(n5766), .A2(n4704), .ZN(n4706) );
  NAND2_X2 U6220 ( .A1(n7796), .A2(n7795), .ZN(n5404) );
  NAND2_X2 U6221 ( .A1(n7626), .A2(n5737), .ZN(n7796) );
  NAND2_X1 U6222 ( .A1(n7629), .A2(n4715), .ZN(n4714) );
  NAND2_X1 U6223 ( .A1(n4714), .A2(n4713), .ZN(n9300) );
  OAI21_X1 U6224 ( .B1(n4349), .B2(n7127), .A(n4724), .ZN(n7301) );
  NAND2_X1 U6225 ( .A1(n6711), .A2(n5792), .ZN(n4730) );
  NAND2_X1 U6226 ( .A1(n9901), .A2(n9902), .ZN(n9900) );
  NAND2_X1 U6227 ( .A1(n9900), .A2(n6716), .ZN(n6717) );
  NAND2_X1 U6228 ( .A1(n9233), .A2(n4369), .ZN(n4733) );
  INV_X1 U6229 ( .A(n4734), .ZN(n9232) );
  NAND2_X1 U6230 ( .A1(n6507), .A2(n4413), .ZN(n4735) );
  NAND2_X1 U6231 ( .A1(n4735), .A2(n4736), .ZN(n7645) );
  AND2_X1 U6232 ( .A1(n4740), .A2(n4738), .ZN(n5053) );
  NAND4_X1 U6233 ( .A1(n4741), .A2(n4740), .A3(n4739), .A4(n4350), .ZN(n4742)
         );
  NOR2_X2 U6234 ( .A1(n5442), .A2(n5058), .ZN(n5078) );
  NAND3_X1 U6235 ( .A1(n4745), .A2(n4744), .A3(n4426), .ZN(n7362) );
  OAI21_X1 U6236 ( .B1(n8872), .B2(n4762), .A(n4761), .ZN(n9003) );
  INV_X1 U6237 ( .A(n4757), .ZN(n8901) );
  AOI21_X1 U6238 ( .B1(n8872), .B2(n4764), .A(n4762), .ZN(n4760) );
  NAND2_X1 U6239 ( .A1(n8872), .A2(n8962), .ZN(n8924) );
  NAND2_X1 U6240 ( .A1(n5427), .A2(n4774), .ZN(n5095) );
  NAND2_X1 U6241 ( .A1(n5427), .A2(n4772), .ZN(n4771) );
  NAND2_X1 U6242 ( .A1(n5427), .A2(n5066), .ZN(n5072) );
  NAND2_X1 U6243 ( .A1(n4778), .A2(n7323), .ZN(n4777) );
  AND2_X1 U6244 ( .A1(n9159), .A2(n4791), .ZN(n9131) );
  OR2_X1 U6245 ( .A1(n9159), .A2(n4790), .ZN(n4788) );
  NAND2_X1 U6246 ( .A1(n9159), .A2(n9139), .ZN(n9141) );
  NAND2_X1 U6247 ( .A1(n9159), .A2(n4792), .ZN(n9130) );
  NAND3_X1 U6248 ( .A1(n4789), .A2(n4788), .A3(n4786), .ZN(n9123) );
  NAND2_X1 U6249 ( .A1(n9159), .A2(n4411), .ZN(n4789) );
  NAND2_X1 U6250 ( .A1(n8869), .A2(n4800), .ZN(n8978) );
  NAND2_X1 U6251 ( .A1(n4807), .A2(n4804), .ZN(n7252) );
  NAND2_X1 U6252 ( .A1(n9795), .A2(n7073), .ZN(n4805) );
  NAND2_X1 U6253 ( .A1(n9226), .A2(n4809), .ZN(n9184) );
  INV_X1 U6254 ( .A(n4812), .ZN(n9204) );
  INV_X1 U6255 ( .A(n4831), .ZN(n6866) );
  AND2_X1 U6256 ( .A1(n7043), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4829) );
  NAND3_X1 U6257 ( .A1(n4834), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4833) );
  INV_X2 U6258 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9122) );
  NAND2_X1 U6259 ( .A1(n5287), .A2(n5286), .ZN(n5289) );
  AOI21_X2 U6260 ( .B1(n4841), .B2(n4839), .A(n4838), .ZN(n5355) );
  NAND2_X1 U6261 ( .A1(n5424), .A2(n4410), .ZN(n4849) );
  NAND2_X1 U6262 ( .A1(n5424), .A2(n4859), .ZN(n4856) );
  AOI21_X1 U6263 ( .B1(n5558), .B2(n4869), .A(n4867), .ZN(n4864) );
  OAI21_X1 U6264 ( .B1(n5558), .B2(n5557), .A(n5556), .ZN(n5577) );
  NAND3_X1 U6265 ( .A1(n4423), .A2(n4875), .A3(n4874), .ZN(n4873) );
  NAND2_X1 U6266 ( .A1(n4888), .A2(n4886), .ZN(n5037) );
  AND2_X1 U6267 ( .A1(n5171), .A2(n5172), .ZN(n4892) );
  NAND2_X2 U6268 ( .A1(n7822), .A2(n7821), .ZN(n7949) );
  NAND2_X1 U6269 ( .A1(n6851), .A2(n6784), .ZN(n7821) );
  NAND2_X2 U6270 ( .A1(n9059), .A2(n9774), .ZN(n7822) );
  INV_X2 U6271 ( .A(n6851), .ZN(n9059) );
  AOI21_X2 U6272 ( .B1(n9156), .B2(n7970), .A(n4433), .ZN(n9138) );
  AND2_X2 U6273 ( .A1(n4894), .A2(n4893), .ZN(n9156) );
  NAND2_X1 U6274 ( .A1(n7225), .A2(n4898), .ZN(n4897) );
  NAND2_X1 U6275 ( .A1(n4905), .A2(n4904), .ZN(n7524) );
  AOI21_X1 U6276 ( .B1(n7398), .B2(n4908), .A(n4395), .ZN(n4904) );
  NAND2_X1 U6277 ( .A1(n9666), .A2(n4906), .ZN(n4905) );
  NAND2_X1 U6278 ( .A1(n6969), .A2(n4910), .ZN(n4912) );
  NOR2_X1 U6279 ( .A1(n7948), .A2(n4911), .ZN(n4910) );
  INV_X1 U6280 ( .A(n7954), .ZN(n4911) );
  NAND2_X1 U6281 ( .A1(n4912), .A2(n4913), .ZN(n7178) );
  INV_X1 U6282 ( .A(n4918), .ZN(n5265) );
  NAND2_X1 U6283 ( .A1(n6469), .A2(n4923), .ZN(n4920) );
  NAND2_X1 U6284 ( .A1(n5078), .A2(n4931), .ZN(n9429) );
  NAND2_X1 U6285 ( .A1(n6329), .A2(n4417), .ZN(n7190) );
  NAND3_X1 U6286 ( .A1(n6367), .A2(n8277), .A3(n6368), .ZN(n8244) );
  NAND2_X1 U6287 ( .A1(n6367), .A2(n8277), .ZN(n8243) );
  INV_X1 U6288 ( .A(n4935), .ZN(n4934) );
  OAI21_X2 U6289 ( .B1(n7719), .B2(n4938), .A(n4936), .ZN(n6380) );
  NOR2_X1 U6290 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  AOI21_X2 U6291 ( .B1(n6122), .B2(n4972), .A(n4971), .ZN(n8554) );
  NAND2_X1 U6292 ( .A1(n5095), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5075) );
  OR2_X1 U6293 ( .A1(n9376), .A2(n9044), .ZN(n6467) );
  NAND2_X1 U6294 ( .A1(n4335), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6295 ( .A1(n6493), .A2(n5159), .ZN(n5145) );
  NAND2_X1 U6296 ( .A1(n6281), .A2(n6280), .ZN(n7688) );
  INV_X1 U6297 ( .A(n6279), .ZN(n6280) );
  OAI21_X1 U6298 ( .B1(n6711), .B2(n5793), .A(n6702), .ZN(n9917) );
  NAND2_X1 U6299 ( .A1(n5106), .A2(n5105), .ZN(n5126) );
  INV_X1 U6300 ( .A(n9226), .ZN(n9247) );
  INV_X1 U6301 ( .A(n5106), .ZN(n9434) );
  AOI21_X2 U6302 ( .B1(n9949), .B2(n6282), .A(n7688), .ZN(n6292) );
  NAND2_X1 U6303 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  OAI21_X1 U6304 ( .B1(n5535), .B2(n5534), .A(n5533), .ZN(n5537) );
  INV_X1 U6305 ( .A(n4376), .ZN(n6946) );
  OAI21_X1 U6306 ( .B1(n6278), .B2(n8717), .A(n6277), .ZN(n6279) );
  NAND2_X1 U6307 ( .A1(n5771), .A2(n7654), .ZN(n5828) );
  XNOR2_X1 U6308 ( .A(n8026), .B(n4406), .ZN(n6278) );
  AOI22_X2 U6309 ( .A1(n7568), .A2(n6340), .B1(n6339), .B2(n8348), .ZN(n8235)
         );
  OAI222_X1 U6310 ( .A1(P2_U3151), .A2(n7666), .B1(n8017), .B2(n9435), .C1(
        n7667), .C2(n8019), .ZN(P2_U3265) );
  NOR2_X1 U6311 ( .A1(n8060), .A2(n8059), .ZN(n4955) );
  INV_X1 U6312 ( .A(n10008), .ZN(n6287) );
  NOR2_X1 U6313 ( .A1(n8377), .A2(n8367), .ZN(n4956) );
  AND3_X1 U6314 ( .A1(n6422), .A2(n6421), .A3(n8315), .ZN(n4957) );
  INV_X2 U6315 ( .A(n9997), .ZN(n9995) );
  NAND2_X1 U6316 ( .A1(n6095), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n4958) );
  OR2_X1 U6317 ( .A1(n9932), .A2(n9959), .ZN(n4959) );
  OR2_X1 U6318 ( .A1(n9344), .A2(n9307), .ZN(n4960) );
  NAND2_X1 U6319 ( .A1(n6112), .A2(n6111), .ZN(n8590) );
  INV_X1 U6320 ( .A(n8590), .ZN(n8285) );
  NOR2_X1 U6321 ( .A1(n5411), .A2(n5392), .ZN(n4962) );
  INV_X1 U6322 ( .A(n9928), .ZN(n6157) );
  OR2_X1 U6323 ( .A1(n6346), .A2(n6345), .ZN(n4963) );
  NOR2_X1 U6324 ( .A1(n5644), .A2(n8925), .ZN(n4964) );
  AND2_X1 U6325 ( .A1(n4966), .A2(n5460), .ZN(n4965) );
  OR2_X1 U6326 ( .A1(n8940), .A2(n8939), .ZN(n4966) );
  NAND2_X1 U6327 ( .A1(n6312), .A2(n7105), .ZN(n4967) );
  NOR2_X1 U6328 ( .A1(n5609), .A2(n5633), .ZN(n4968) );
  INV_X1 U6329 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4982) );
  OR2_X1 U6330 ( .A1(n7908), .A2(n7932), .ZN(n4970) );
  AND2_X1 U6331 ( .A1(n8798), .A2(n8579), .ZN(n4971) );
  OR2_X1 U6332 ( .A1(n8798), .A2(n8579), .ZN(n4972) );
  OAI21_X1 U6333 ( .B1(n7239), .B2(n5895), .A(n5894), .ZN(n7266) );
  AND2_X1 U6334 ( .A1(n4988), .A2(n4987), .ZN(n4974) );
  AND2_X1 U6335 ( .A1(n9315), .A2(n5751), .ZN(n9034) );
  INV_X1 U6336 ( .A(n9034), .ZN(n5752) );
  AND2_X1 U6337 ( .A1(n7922), .A2(n7734), .ZN(n7916) );
  AOI211_X1 U6338 ( .C1(n7923), .C2(n7922), .A(n7921), .B(n7920), .ZN(n7924)
         );
  INV_X1 U6339 ( .A(n7931), .ZN(n7933) );
  INV_X1 U6340 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U6341 ( .A1(n7933), .A2(n7932), .ZN(n7934) );
  NAND2_X1 U6342 ( .A1(n7935), .A2(n7934), .ZN(n7936) );
  OR2_X1 U6343 ( .A1(n6705), .A2(n6762), .ZN(n6706) );
  INV_X1 U6344 ( .A(n8591), .ZN(n6368) );
  NAND2_X1 U6345 ( .A1(n6213), .A2(n6948), .ZN(n6947) );
  NAND2_X1 U6346 ( .A1(n4346), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4976) );
  OR2_X1 U6347 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  INV_X1 U6348 ( .A(n6848), .ZN(n6214) );
  AND2_X1 U6349 ( .A1(n8101), .A2(n9922), .ZN(n8096) );
  NOR2_X1 U6350 ( .A1(n5608), .A2(n5607), .ZN(n5633) );
  INV_X1 U6351 ( .A(n7819), .ZN(n6500) );
  NOR2_X1 U6352 ( .A1(n7252), .A2(n6519), .ZN(n7253) );
  NAND2_X1 U6353 ( .A1(n7154), .A2(n6971), .ZN(n7816) );
  INV_X1 U6354 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5060) );
  INV_X1 U6355 ( .A(n5554), .ZN(n5555) );
  INV_X1 U6356 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5066) );
  INV_X1 U6357 ( .A(n7403), .ZN(n6335) );
  NAND2_X1 U6358 ( .A1(n6366), .A2(n6365), .ZN(n8277) );
  NAND2_X1 U6359 ( .A1(n6373), .A2(n8285), .ZN(n6374) );
  NAND2_X1 U6360 ( .A1(n7047), .A2(n7046), .ZN(n7048) );
  INV_X1 U6361 ( .A(n7373), .ZN(n7374) );
  INV_X1 U6362 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5306) );
  OAI21_X1 U6363 ( .B1(n8008), .B2(n5096), .A(n6531), .ZN(n5097) );
  OR2_X1 U6364 ( .A1(n5584), .A2(n8875), .ZN(n5608) );
  OR2_X1 U6365 ( .A1(n5126), .A2(n5125), .ZN(n5129) );
  INV_X1 U6366 ( .A(n9376), .ZN(n6520) );
  OR2_X1 U6367 ( .A1(n7659), .A2(n7658), .ZN(n7660) );
  INV_X1 U6368 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5059) );
  INV_X1 U6369 ( .A(n5427), .ZN(n5428) );
  OR2_X1 U6370 ( .A1(n5387), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5388) );
  INV_X1 U6371 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U6372 ( .A1(n6335), .A2(n8350), .ZN(n6336) );
  INV_X1 U6373 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5829) );
  INV_X1 U6374 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5813) );
  AOI22_X1 U6375 ( .A1(n7347), .A2(n7348), .B1(n7339), .B2(n6334), .ZN(n7401)
         );
  INV_X1 U6376 ( .A(n8571), .ZN(n7713) );
  INV_X1 U6377 ( .A(n8539), .ZN(n8062) );
  NAND2_X1 U6378 ( .A1(n9892), .A2(n6703), .ZN(n9916) );
  OR2_X1 U6379 ( .A1(n6139), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7678) );
  NAND2_X1 U6380 ( .A1(n6061), .A2(n10077), .ZN(n6071) );
  AND2_X1 U6381 ( .A1(n7201), .A2(n8062), .ZN(n8222) );
  AND2_X1 U6382 ( .A1(n8219), .A2(n8221), .ZN(n6840) );
  NAND2_X1 U6383 ( .A1(n8222), .A2(n7318), .ZN(n9982) );
  NAND2_X1 U6384 ( .A1(n6177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6179) );
  AND2_X1 U6385 ( .A1(n5696), .A2(n5697), .ZN(n5695) );
  AND2_X1 U6386 ( .A1(n6655), .A2(n5164), .ZN(n6768) );
  NOR2_X1 U6387 ( .A1(n5448), .A2(n10167), .ZN(n5473) );
  OR3_X1 U6388 ( .A1(n5447), .A2(n9023), .A3(n5446), .ZN(n5448) );
  INV_X1 U6389 ( .A(n7796), .ZN(n6568) );
  OR2_X1 U6390 ( .A1(n5365), .A2(n7499), .ZN(n5367) );
  INV_X1 U6391 ( .A(n9324), .ZN(n7630) );
  INV_X1 U6392 ( .A(n9702), .ZN(n9759) );
  AND2_X1 U6393 ( .A1(n5669), .A2(n5630), .ZN(n5649) );
  XNOR2_X1 U6394 ( .A(n5028), .B(SI_11_), .ZN(n5337) );
  AND2_X1 U6395 ( .A1(n4981), .A2(n5001), .ZN(n5221) );
  NAND2_X1 U6396 ( .A1(n6405), .A2(n6404), .ZN(n8323) );
  AND2_X1 U6397 ( .A1(n6100), .A2(n6099), .ZN(n8248) );
  INV_X1 U6398 ( .A(n9899), .ZN(n9905) );
  INV_X1 U6399 ( .A(n8509), .ZN(n9906) );
  INV_X1 U6400 ( .A(n9913), .ZN(n9891) );
  AND2_X1 U6401 ( .A1(n8113), .A2(n8118), .ZN(n8045) );
  INV_X1 U6402 ( .A(n9939), .ZN(n8705) );
  INV_X1 U6403 ( .A(n8737), .ZN(n8780) );
  AND2_X1 U6404 ( .A1(n6395), .A2(n6242), .ZN(n6835) );
  INV_X1 U6405 ( .A(n8177), .ZN(n8613) );
  INV_X1 U6406 ( .A(n8150), .ZN(n8684) );
  INV_X1 U6407 ( .A(n8834), .ZN(n8854) );
  NAND2_X1 U6408 ( .A1(n8717), .A2(n9982), .ZN(n9994) );
  AND2_X1 U6409 ( .A1(n5999), .A2(n5990), .ZN(n8450) );
  INV_X1 U6410 ( .A(n9839), .ZN(n7521) );
  INV_X1 U6411 ( .A(n8959), .ZN(n9014) );
  AND2_X1 U6412 ( .A1(n5746), .A2(n5722), .ZN(n9021) );
  AND2_X1 U6413 ( .A1(n5572), .A2(n5571), .ZN(n8918) );
  OR2_X1 U6414 ( .A1(n6648), .A2(n6663), .ZN(n9644) );
  INV_X1 U6415 ( .A(n9644), .ZN(n9112) );
  INV_X1 U6416 ( .A(n7971), .ZN(n9176) );
  INV_X1 U6417 ( .A(n7962), .ZN(n7644) );
  INV_X1 U6418 ( .A(n9307), .ZN(n9715) );
  INV_X1 U6419 ( .A(n9135), .ZN(n9339) );
  INV_X1 U6420 ( .A(n9791), .ZN(n9842) );
  AND2_X1 U6421 ( .A1(n7261), .A2(n7260), .ZN(n9336) );
  XNOR2_X1 U6422 ( .A(n5075), .B(n5074), .ZN(n5720) );
  INV_X1 U6423 ( .A(n8323), .ZN(n8333) );
  NAND2_X1 U6424 ( .A1(n6145), .A2(n6144), .ZN(n8555) );
  NAND2_X1 U6425 ( .A1(n6087), .A2(n6086), .ZN(n8591) );
  INV_X1 U6426 ( .A(n8238), .ZN(n8348) );
  INV_X1 U6427 ( .A(n9919), .ZN(n9896) );
  INV_X1 U6428 ( .A(n8733), .ZN(n8713) );
  NAND2_X1 U6429 ( .A1(n8733), .A2(n6981), .ZN(n9943) );
  NAND2_X1 U6430 ( .A1(n6839), .A2(n8728), .ZN(n9939) );
  NAND2_X1 U6431 ( .A1(n10008), .A2(n9994), .ZN(n8783) );
  OR2_X1 U6432 ( .A1(n9997), .A2(n9965), .ZN(n8858) );
  AND3_X1 U6433 ( .A1(n9970), .A2(n9969), .A3(n9968), .ZN(n10003) );
  AND2_X1 U6434 ( .A1(n6211), .A2(n6210), .ZN(n9997) );
  AND2_X1 U6435 ( .A1(n6559), .A2(n6188), .ZN(n6579) );
  INV_X1 U6436 ( .A(n8229), .ZN(n7318) );
  INV_X1 U6437 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6856) );
  INV_X1 U6438 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6573) );
  INV_X1 U6439 ( .A(n9030), .ZN(n9012) );
  INV_X1 U6440 ( .A(n9021), .ZN(n8999) );
  OR2_X1 U6441 ( .A1(n6648), .A2(n6647), .ZN(n9625) );
  INV_X1 U6442 ( .A(n9522), .ZN(n9659) );
  AND2_X1 U6443 ( .A1(n9686), .A2(n6492), .ZN(n9307) );
  NAND2_X1 U6444 ( .A1(n6521), .A2(n9315), .ZN(n9752) );
  INV_X1 U6445 ( .A(n10233), .ZN(n9878) );
  INV_X1 U6446 ( .A(n9854), .ZN(n9852) );
  AND2_X2 U6447 ( .A1(n9336), .A2(n7263), .ZN(n9854) );
  OR2_X1 U6448 ( .A1(n9423), .A2(n9422), .ZN(n9756) );
  INV_X1 U6449 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6941) );
  INV_X1 U6450 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6565) );
  OR2_X1 U6451 ( .A1(n5269), .A2(n5268), .ZN(n9565) );
  INV_X1 U6452 ( .A(n8507), .ZN(P2_U3893) );
  AND2_X1 U6453 ( .A1(n6569), .A2(n6532), .ZN(P1_U3973) );
  NAND2_X1 U6454 ( .A1(n4960), .A2(n6530), .ZN(P1_U3356) );
  INV_X4 U6455 ( .A(n4992), .ZN(n7795) );
  INV_X1 U6456 ( .A(n4980), .ZN(n4979) );
  INV_X1 U6457 ( .A(SI_4_), .ZN(n4978) );
  NAND2_X1 U6458 ( .A1(n4979), .A2(n4978), .ZN(n4981) );
  NAND2_X1 U6459 ( .A1(n4980), .A2(SI_4_), .ZN(n5001) );
  INV_X1 U6460 ( .A(SI_2_), .ZN(n4983) );
  NAND2_X1 U6461 ( .A1(n4984), .A2(n4983), .ZN(n4986) );
  NAND2_X1 U6462 ( .A1(n4985), .A2(SI_2_), .ZN(n4996) );
  NAND2_X1 U6463 ( .A1(n4986), .A2(n4996), .ZN(n5176) );
  INV_X1 U6464 ( .A(n5176), .ZN(n4995) );
  OAI211_X1 U6465 ( .C1(SI_1_), .C2(P2_DATAO_REG_1__SCAN_IN), .A(SI_0_), .B(
        P2_DATAO_REG_0__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6466 ( .A1(SI_1_), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4987) );
  OR2_X1 U6467 ( .A1(n4992), .A2(n4974), .ZN(n4994) );
  OAI211_X1 U6468 ( .C1(SI_1_), .C2(P1_DATAO_REG_1__SCAN_IN), .A(SI_0_), .B(
        P1_DATAO_REG_0__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U6469 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U6470 ( .A1(n4990), .A2(n4989), .ZN(n4991) );
  NAND2_X1 U6471 ( .A1(n4992), .A2(n4991), .ZN(n4993) );
  NAND2_X1 U6472 ( .A1(n4994), .A2(n4993), .ZN(n5174) );
  MUX2_X1 U6473 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4346), .Z(n4998) );
  OAI21_X1 U6474 ( .B1(n4998), .B2(SI_3_), .A(n5000), .ZN(n5196) );
  INV_X1 U6475 ( .A(n5196), .ZN(n4999) );
  NAND2_X1 U6476 ( .A1(n5221), .A2(n5222), .ZN(n5220) );
  NAND2_X1 U6477 ( .A1(n5220), .A2(n5001), .ZN(n5240) );
  MUX2_X1 U6478 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7795), .Z(n5002) );
  NAND2_X1 U6479 ( .A1(n5002), .A2(SI_5_), .ZN(n5006) );
  INV_X1 U6480 ( .A(n5002), .ZN(n5004) );
  INV_X1 U6481 ( .A(SI_5_), .ZN(n5003) );
  NAND2_X1 U6482 ( .A1(n5004), .A2(n5003), .ZN(n5005) );
  NAND2_X1 U6483 ( .A1(n5240), .A2(n5239), .ZN(n5238) );
  MUX2_X1 U6484 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7795), .Z(n5007) );
  NAND2_X1 U6485 ( .A1(n5007), .A2(SI_6_), .ZN(n5011) );
  INV_X1 U6486 ( .A(n5007), .ZN(n5009) );
  INV_X1 U6487 ( .A(SI_6_), .ZN(n5008) );
  NAND2_X1 U6488 ( .A1(n5009), .A2(n5008), .ZN(n5010) );
  MUX2_X1 U6489 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7795), .Z(n5012) );
  NAND2_X1 U6490 ( .A1(n5012), .A2(SI_7_), .ZN(n5016) );
  INV_X1 U6491 ( .A(n5012), .ZN(n5014) );
  INV_X1 U6492 ( .A(SI_7_), .ZN(n5013) );
  NAND2_X1 U6493 ( .A1(n5014), .A2(n5013), .ZN(n5015) );
  MUX2_X1 U6494 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n4346), .Z(n5017) );
  INV_X1 U6495 ( .A(n5017), .ZN(n5019) );
  INV_X1 U6496 ( .A(SI_8_), .ZN(n5018) );
  MUX2_X1 U6497 ( .A(n6573), .B(n6565), .S(n4346), .Z(n5020) );
  INV_X1 U6498 ( .A(n5020), .ZN(n5021) );
  MUX2_X1 U6499 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7795), .Z(n5022) );
  NAND2_X1 U6500 ( .A1(n5022), .A2(SI_10_), .ZN(n5027) );
  INV_X1 U6501 ( .A(n5022), .ZN(n5024) );
  INV_X1 U6502 ( .A(SI_10_), .ZN(n5023) );
  NAND2_X1 U6503 ( .A1(n5024), .A2(n5023), .ZN(n5025) );
  NAND2_X1 U6504 ( .A1(n5027), .A2(n5025), .ZN(n5356) );
  INV_X1 U6505 ( .A(n5356), .ZN(n5026) );
  MUX2_X1 U6506 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4346), .Z(n5028) );
  MUX2_X1 U6507 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4346), .Z(n5029) );
  MUX2_X1 U6508 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4346), .Z(n5031) );
  INV_X1 U6509 ( .A(n5031), .ZN(n5033) );
  INV_X1 U6510 ( .A(SI_13_), .ZN(n5032) );
  NAND2_X1 U6511 ( .A1(n5033), .A2(n5032), .ZN(n5034) );
  MUX2_X1 U6512 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4346), .Z(n5114) );
  MUX2_X1 U6513 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7795), .Z(n5439) );
  INV_X1 U6514 ( .A(n5439), .ZN(n5036) );
  NAND2_X1 U6515 ( .A1(n5037), .A2(n5036), .ZN(n5040) );
  NAND2_X1 U6516 ( .A1(n5038), .A2(n4887), .ZN(n5039) );
  MUX2_X1 U6517 ( .A(n6856), .B(n6858), .S(n4346), .Z(n5425) );
  NAND2_X1 U6518 ( .A1(n5041), .A2(SI_16_), .ZN(n5042) );
  MUX2_X1 U6519 ( .A(n6943), .B(n6941), .S(n7795), .Z(n5045) );
  INV_X1 U6520 ( .A(SI_17_), .ZN(n5044) );
  INV_X1 U6521 ( .A(n5045), .ZN(n5046) );
  NAND2_X1 U6522 ( .A1(n5046), .A2(SI_17_), .ZN(n5047) );
  NAND2_X1 U6523 ( .A1(n5048), .A2(n5047), .ZN(n5469) );
  INV_X1 U6524 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7063) );
  INV_X1 U6525 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5049) );
  MUX2_X1 U6526 ( .A(n7063), .B(n5049), .S(n7795), .Z(n5492) );
  XNOR2_X1 U6527 ( .A(n5492), .B(SI_18_), .ZN(n5491) );
  XNOR2_X1 U6528 ( .A(n5495), .B(n5491), .ZN(n7012) );
  NOR2_X4 U6529 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5132) );
  NOR2_X2 U6530 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5050) );
  NOR2_X1 U6531 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5055) );
  INV_X1 U6532 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5062) );
  INV_X1 U6533 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6534 ( .A1(n5062), .A2(n5061), .ZN(n5063) );
  OR2_X2 U6535 ( .A1(n5098), .A2(n5360), .ZN(n5103) );
  XNOR2_X2 U6536 ( .A(n5103), .B(n5099), .ZN(n5737) );
  NAND2_X1 U6537 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n5065) );
  INV_X2 U6538 ( .A(n5404), .ZN(n7782) );
  NAND2_X1 U6539 ( .A1(n7012), .A2(n7782), .ZN(n5069) );
  NAND2_X1 U6540 ( .A1(n5072), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6541 ( .A1(n5088), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5067) );
  XNOR2_X1 U6542 ( .A(n5067), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9654) );
  AOI22_X1 U6543 ( .A1(n5500), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6568), .B2(
        n9654), .ZN(n5068) );
  NAND2_X1 U6544 ( .A1(n5086), .A2(n5070), .ZN(n5071) );
  NAND2_X1 U6545 ( .A1(n5076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5077) );
  INV_X1 U6546 ( .A(n5078), .ZN(n5079) );
  NAND2_X1 U6547 ( .A1(n5079), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5080) );
  MUX2_X1 U6548 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5080), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5082) );
  INV_X1 U6549 ( .A(n5081), .ZN(n5084) );
  NAND2_X1 U6550 ( .A1(n5082), .A2(n5084), .ZN(n7565) );
  NAND2_X1 U6551 ( .A1(n5084), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5085) );
  XNOR2_X1 U6552 ( .A(n5085), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7576) );
  NAND3_X1 U6553 ( .A1(n5088), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n5094) );
  INV_X1 U6554 ( .A(n5086), .ZN(n5087) );
  NAND2_X1 U6555 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n5089) );
  NAND2_X1 U6556 ( .A1(n5089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5090) );
  OAI21_X1 U6557 ( .B1(n5091), .B2(P1_IR_REG_31__SCAN_IN), .A(n5090), .ZN(
        n5092) );
  INV_X1 U6558 ( .A(n5092), .ZN(n5093) );
  NAND2_X1 U6559 ( .A1(n5749), .A2(n8003), .ZN(n8008) );
  INV_X1 U6560 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U6561 ( .A1(n5099), .A2(n9427), .ZN(n5100) );
  NAND2_X1 U6562 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5102) );
  NAND2_X1 U6563 ( .A1(n5103), .A2(n5102), .ZN(n5104) );
  XNOR2_X2 U6564 ( .A(n5104), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5109) );
  INV_X1 U6565 ( .A(n5109), .ZN(n5105) );
  AOI22_X1 U6566 ( .A1(n4340), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n5520), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5111) );
  NOR2_X2 U6567 ( .A1(n5307), .A2(n5306), .ZN(n5323) );
  NAND2_X1 U6568 ( .A1(n5323), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5365) );
  INV_X1 U6569 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9023) );
  INV_X1 U6570 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5446) );
  INV_X1 U6571 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10167) );
  NAND2_X1 U6572 ( .A1(n5473), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5475) );
  INV_X1 U6573 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6574 ( .A1(n5475), .A2(n5107), .ZN(n5108) );
  AND2_X1 U6575 ( .A1(n5503), .A2(n5108), .ZN(n9294) );
  AOI22_X1 U6576 ( .A1(n6478), .A2(n9294), .B1(n5521), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5110) );
  INV_X1 U6577 ( .A(n8886), .ZN(n9312) );
  AOI22_X1 U6578 ( .A1(n9397), .A2(n5159), .B1(n8896), .B2(n9312), .ZN(n8991)
         );
  NAND2_X4 U6579 ( .A1(n5727), .A2(n5112), .ZN(n8894) );
  XNOR2_X1 U6580 ( .A(n5114), .B(SI_14_), .ZN(n5115) );
  XNOR2_X1 U6581 ( .A(n5113), .B(n5115), .ZN(n6680) );
  NAND2_X1 U6582 ( .A1(n6680), .A2(n7782), .ZN(n5119) );
  OR2_X1 U6583 ( .A1(n5116), .A2(n5360), .ZN(n5117) );
  XNOR2_X1 U6584 ( .A(n5117), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9609) );
  AOI22_X1 U6585 ( .A1(n5500), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6568), .B2(
        n9609), .ZN(n5118) );
  INV_X2 U6586 ( .A(n5126), .ZN(n5450) );
  XNOR2_X1 U6587 ( .A(n5447), .B(P1_REG3_REG_14__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U6588 ( .A1(n5450), .A2(n7555), .ZN(n5123) );
  NAND2_X1 U6589 ( .A1(n4340), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6590 ( .A1(n4335), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6591 ( .A1(n5520), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5120) );
  NAND4_X1 U6592 ( .A1(n5123), .A2(n5122), .A3(n5121), .A4(n5120), .ZN(n9047)
         );
  AOI22_X1 U6593 ( .A1(n7560), .A2(n5244), .B1(n5159), .B2(n9047), .ZN(n5124)
         );
  XOR2_X1 U6594 ( .A(n8894), .B(n5124), .Z(n5421) );
  INV_X1 U6595 ( .A(n5421), .ZN(n7552) );
  INV_X1 U6596 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6597 ( .A1(n5521), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6598 ( .A1(n5151), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5127) );
  AND3_X1 U6599 ( .A1(n5129), .A2(n5128), .A3(n5127), .ZN(n5131) );
  NAND2_X1 U6600 ( .A1(n4340), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5130) );
  INV_X1 U6601 ( .A(n5132), .ZN(n5133) );
  INV_X1 U6602 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6587) );
  OR2_X1 U6603 ( .A1(n5173), .A2(n6587), .ZN(n5143) );
  MUX2_X1 U6604 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n7795), .Z(n5134) );
  NAND2_X1 U6605 ( .A1(n5134), .A2(SI_0_), .ZN(n5136) );
  INV_X1 U6606 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6550) );
  MUX2_X1 U6607 ( .A(n6550), .B(n6587), .S(n7795), .Z(n5135) );
  XNOR2_X1 U6608 ( .A(n5136), .B(n5135), .ZN(n5138) );
  INV_X1 U6609 ( .A(SI_1_), .ZN(n5137) );
  NAND2_X1 U6610 ( .A1(n5138), .A2(n5137), .ZN(n5141) );
  INV_X1 U6611 ( .A(n5138), .ZN(n5139) );
  NAND2_X1 U6612 ( .A1(n5139), .A2(SI_1_), .ZN(n5140) );
  NAND2_X1 U6613 ( .A1(n5141), .A2(n5140), .ZN(n6549) );
  NAND2_X1 U6614 ( .A1(n5150), .A2(n6429), .ZN(n5144) );
  NAND2_X1 U6615 ( .A1(n5145), .A2(n5144), .ZN(n5146) );
  AND2_X1 U6616 ( .A1(n6429), .A2(n5159), .ZN(n5147) );
  AOI21_X1 U6617 ( .B1(n6493), .B2(n8896), .A(n5147), .ZN(n5166) );
  XNOR2_X1 U6618 ( .A(n5165), .B(n5166), .ZN(n6769) );
  INV_X1 U6619 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U6620 ( .A1(n7795), .A2(SI_0_), .ZN(n5149) );
  INV_X1 U6621 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5148) );
  XNOR2_X1 U6622 ( .A(n5149), .B(n5148), .ZN(n9439) );
  MUX2_X1 U6623 ( .A(n6625), .B(n9439), .S(n7796), .Z(n9735) );
  INV_X1 U6624 ( .A(n9735), .ZN(n9762) );
  NAND2_X1 U6625 ( .A1(n9762), .A2(n5150), .ZN(n5157) );
  NAND2_X1 U6626 ( .A1(n5450), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6627 ( .A1(n4345), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6628 ( .A1(n5151), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U6629 ( .A1(n5521), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5152) );
  NAND4_X2 U6630 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n7737)
         );
  NAND2_X1 U6631 ( .A1(n7737), .A2(n5159), .ZN(n5156) );
  NAND2_X1 U6632 ( .A1(n5723), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6633 ( .A1(n7737), .A2(n8896), .ZN(n5162) );
  OAI22_X1 U6634 ( .A1(n9735), .A2(n5546), .B1(n6531), .B2(n6625), .ZN(n5160)
         );
  INV_X1 U6635 ( .A(n5160), .ZN(n5161) );
  NAND2_X1 U6636 ( .A1(n5162), .A2(n5161), .ZN(n6656) );
  NAND2_X1 U6637 ( .A1(n6657), .A2(n6656), .ZN(n6655) );
  NAND2_X1 U6638 ( .A1(n5163), .A2(n5616), .ZN(n5164) );
  NAND2_X1 U6639 ( .A1(n6769), .A2(n6768), .ZN(n6767) );
  INV_X1 U6640 ( .A(n5165), .ZN(n5167) );
  NAND2_X1 U6641 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  NAND2_X1 U6642 ( .A1(n6767), .A2(n5168), .ZN(n6813) );
  NAND2_X1 U6643 ( .A1(n4340), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6644 ( .A1(n5450), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6645 ( .A1(n5151), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6646 ( .A1(n4335), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6647 ( .A1(n9059), .A2(n5159), .ZN(n5184) );
  OR2_X1 U6648 ( .A1(n4341), .A2(n4476), .ZN(n5182) );
  INV_X1 U6649 ( .A(n5174), .ZN(n5175) );
  NAND2_X1 U6650 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  NAND2_X1 U6651 ( .A1(n5178), .A2(n5177), .ZN(n6553) );
  OR2_X1 U6652 ( .A1(n5404), .A2(n6553), .ZN(n5181) );
  OR2_X1 U6653 ( .A1(n5132), .A2(n5360), .ZN(n5179) );
  XNOR2_X1 U6654 ( .A(n5179), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6628) );
  INV_X1 U6655 ( .A(n6628), .ZN(n6745) );
  OR2_X1 U6656 ( .A1(n7796), .A2(n6745), .ZN(n5180) );
  AND3_X2 U6657 ( .A1(n5182), .A2(n5181), .A3(n5180), .ZN(n9774) );
  NAND2_X1 U6658 ( .A1(n6784), .A2(n5150), .ZN(n5183) );
  NAND2_X1 U6659 ( .A1(n5184), .A2(n5183), .ZN(n5185) );
  XNOR2_X1 U6660 ( .A(n5185), .B(n8894), .ZN(n5186) );
  AOI22_X1 U6661 ( .A1(n9059), .A2(n8896), .B1(n6784), .B2(n5159), .ZN(n5187)
         );
  XNOR2_X1 U6662 ( .A(n5186), .B(n5187), .ZN(n6814) );
  NAND2_X1 U6663 ( .A1(n6813), .A2(n6814), .ZN(n5190) );
  INV_X1 U6664 ( .A(n5186), .ZN(n5188) );
  NAND2_X1 U6665 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  NAND2_X1 U6666 ( .A1(n5190), .A2(n5189), .ZN(n6849) );
  INV_X1 U6667 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6925) );
  NAND2_X1 U6668 ( .A1(n5450), .A2(n6925), .ZN(n5194) );
  NAND2_X1 U6669 ( .A1(n4345), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6670 ( .A1(n5151), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6671 ( .A1(n4335), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5191) );
  NAND4_X2 U6672 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), .ZN(n9058)
         );
  NAND2_X1 U6673 ( .A1(n9058), .A2(n5159), .ZN(n5205) );
  INV_X1 U6674 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6541) );
  OR2_X1 U6675 ( .A1(n4341), .A2(n6541), .ZN(n5203) );
  INV_X1 U6676 ( .A(n5195), .ZN(n5197) );
  NAND2_X1 U6677 ( .A1(n5197), .A2(n5196), .ZN(n5199) );
  NAND2_X1 U6678 ( .A1(n5199), .A2(n5198), .ZN(n6552) );
  OR2_X1 U6679 ( .A1(n5404), .A2(n6552), .ZN(n5202) );
  NAND2_X1 U6680 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4382), .ZN(n5200) );
  XNOR2_X1 U6681 ( .A(n5200), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6629) );
  INV_X1 U6682 ( .A(n6629), .ZN(n9484) );
  OR2_X1 U6683 ( .A1(n7796), .A2(n9484), .ZN(n5201) );
  NAND2_X1 U6684 ( .A1(n6926), .A2(n5150), .ZN(n5204) );
  NAND2_X1 U6685 ( .A1(n5205), .A2(n5204), .ZN(n5206) );
  XNOR2_X1 U6686 ( .A(n5206), .B(n8894), .ZN(n5207) );
  AOI22_X1 U6687 ( .A1(n9058), .A2(n8896), .B1(n6926), .B2(n5159), .ZN(n5208)
         );
  XNOR2_X1 U6688 ( .A(n5207), .B(n5208), .ZN(n6850) );
  INV_X1 U6689 ( .A(n5207), .ZN(n5209) );
  NAND2_X1 U6690 ( .A1(n5209), .A2(n5208), .ZN(n5210) );
  NOR2_X1 U6691 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5211) );
  NOR2_X1 U6692 ( .A1(n5231), .A2(n5211), .ZN(n6894) );
  NAND2_X1 U6693 ( .A1(n5450), .A2(n6894), .ZN(n5215) );
  NAND2_X1 U6694 ( .A1(n4345), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6695 ( .A1(n4335), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6696 ( .A1(n5151), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5212) );
  NAND4_X1 U6697 ( .A1(n5215), .A2(n5214), .A3(n5213), .A4(n5212), .ZN(n9057)
         );
  NAND2_X1 U6698 ( .A1(n9057), .A2(n5159), .ZN(n5227) );
  NAND2_X1 U6699 ( .A1(n5216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5217) );
  MUX2_X1 U6700 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5217), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5219) );
  NAND2_X1 U6701 ( .A1(n5219), .A2(n5218), .ZN(n6678) );
  INV_X1 U6702 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6538) );
  OR2_X1 U6703 ( .A1(n4342), .A2(n6538), .ZN(n5225) );
  OR2_X1 U6704 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  NAND2_X1 U6705 ( .A1(n5220), .A2(n5223), .ZN(n6554) );
  OR2_X1 U6706 ( .A1(n5404), .A2(n6554), .ZN(n5224) );
  OAI211_X1 U6707 ( .C1(n7796), .C2(n6678), .A(n5225), .B(n5224), .ZN(n9786)
         );
  NAND2_X1 U6708 ( .A1(n5244), .A2(n9786), .ZN(n5226) );
  NAND2_X1 U6709 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  XNOR2_X1 U6710 ( .A(n5228), .B(n5616), .ZN(n5248) );
  AND2_X1 U6711 ( .A1(n9786), .A2(n5159), .ZN(n5229) );
  AOI21_X1 U6712 ( .B1(n9057), .B2(n8896), .A(n5229), .ZN(n5249) );
  XNOR2_X1 U6713 ( .A(n5248), .B(n5249), .ZN(n6895) );
  NOR2_X1 U6714 ( .A1(n5231), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5232) );
  NOR2_X1 U6715 ( .A1(n5259), .A2(n5232), .ZN(n7084) );
  NAND2_X1 U6716 ( .A1(n5450), .A2(n7084), .ZN(n5236) );
  NAND2_X1 U6717 ( .A1(n4345), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6718 ( .A1(n5151), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6719 ( .A1(n4335), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6720 ( .A1(n9056), .A2(n5159), .ZN(n5246) );
  NAND2_X1 U6721 ( .A1(n5218), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5237) );
  XNOR2_X1 U6722 ( .A(n5237), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6634) );
  INV_X1 U6723 ( .A(n6634), .ZN(n9551) );
  OR2_X1 U6724 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NAND2_X1 U6725 ( .A1(n5238), .A2(n5241), .ZN(n6544) );
  OR2_X1 U6726 ( .A1(n5404), .A2(n6544), .ZN(n5243) );
  INV_X1 U6727 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6539) );
  OR2_X1 U6728 ( .A1(n4341), .A2(n6539), .ZN(n5242) );
  OAI211_X1 U6729 ( .C1(n7796), .C2(n9551), .A(n5243), .B(n5242), .ZN(n6971)
         );
  NAND2_X1 U6730 ( .A1(n5244), .A2(n6971), .ZN(n5245) );
  NAND2_X1 U6731 ( .A1(n5246), .A2(n5245), .ZN(n5247) );
  XNOR2_X1 U6732 ( .A(n5247), .B(n8894), .ZN(n5257) );
  INV_X1 U6733 ( .A(n5257), .ZN(n5252) );
  INV_X1 U6734 ( .A(n5248), .ZN(n5251) );
  INV_X1 U6735 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6736 ( .A1(n5251), .A2(n5250), .ZN(n5256) );
  AND2_X1 U6737 ( .A1(n5252), .A2(n5256), .ZN(n5253) );
  NAND2_X1 U6738 ( .A1(n6897), .A2(n5253), .ZN(n7078) );
  NAND2_X1 U6739 ( .A1(n9056), .A2(n8896), .ZN(n5255) );
  NAND2_X1 U6740 ( .A1(n6971), .A2(n5159), .ZN(n5254) );
  NAND2_X1 U6741 ( .A1(n5255), .A2(n5254), .ZN(n7080) );
  NAND2_X1 U6742 ( .A1(n6897), .A2(n5256), .ZN(n5258) );
  NOR2_X1 U6743 ( .A1(n5259), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5260) );
  NOR2_X1 U6744 ( .A1(n5282), .A2(n5260), .ZN(n9718) );
  NAND2_X1 U6745 ( .A1(n6478), .A2(n9718), .ZN(n5264) );
  NAND2_X1 U6746 ( .A1(n4345), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6747 ( .A1(n4335), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6748 ( .A1(n5151), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5261) );
  NAND4_X1 U6749 ( .A1(n5264), .A2(n5263), .A3(n5262), .A4(n5261), .ZN(n9055)
         );
  NAND2_X1 U6750 ( .A1(n9055), .A2(n5159), .ZN(n5276) );
  NOR2_X1 U6751 ( .A1(n5265), .A2(n5360), .ZN(n5266) );
  MUX2_X1 U6752 ( .A(n5360), .B(n5266), .S(P1_IR_REG_6__SCAN_IN), .Z(n5269) );
  INV_X1 U6753 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6754 ( .A1(n5265), .A2(n5267), .ZN(n5303) );
  INV_X1 U6755 ( .A(n5303), .ZN(n5268) );
  OR2_X1 U6756 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  INV_X1 U6757 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6540) );
  OR2_X1 U6758 ( .A1(n4342), .A2(n6540), .ZN(n5274) );
  NAND2_X1 U6759 ( .A1(n5244), .A2(n6519), .ZN(n5275) );
  NAND2_X1 U6760 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  XNOR2_X1 U6761 ( .A(n5277), .B(n5616), .ZN(n5280) );
  AOI22_X1 U6762 ( .A1(n9055), .A2(n8896), .B1(n5159), .B2(n6519), .ZN(n5279)
         );
  XNOR2_X1 U6763 ( .A(n5280), .B(n5279), .ZN(n7152) );
  NAND2_X1 U6764 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  AOI22_X1 U6765 ( .A1(n4345), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n5151), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n5285) );
  OAI21_X1 U6766 ( .B1(n5282), .B2(P1_REG3_REG_7__SCAN_IN), .A(n5307), .ZN(
        n5283) );
  INV_X1 U6767 ( .A(n5283), .ZN(n7181) );
  AOI22_X1 U6768 ( .A1(n6478), .A2(n7181), .B1(n4335), .B2(
        P1_REG0_REG_7__SCAN_IN), .ZN(n5284) );
  OR2_X1 U6769 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  NAND2_X1 U6770 ( .A1(n5289), .A2(n5288), .ZN(n6547) );
  OR2_X1 U6771 ( .A1(n6547), .A2(n5404), .ZN(n5292) );
  NAND2_X1 U6772 ( .A1(n5303), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5290) );
  XNOR2_X1 U6773 ( .A(n5290), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U6774 ( .A1(n5500), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6568), .B2(
        n6641), .ZN(n5291) );
  NAND2_X1 U6775 ( .A1(n5292), .A2(n5291), .ZN(n7182) );
  NAND2_X1 U6776 ( .A1(n7182), .A2(n5244), .ZN(n5293) );
  OAI21_X1 U6777 ( .B1(n7330), .B2(n5546), .A(n5293), .ZN(n5294) );
  XNOR2_X1 U6778 ( .A(n5294), .B(n8894), .ZN(n7163) );
  INV_X1 U6779 ( .A(n7163), .ZN(n5298) );
  OR2_X1 U6780 ( .A1(n7330), .A2(n5618), .ZN(n5296) );
  NAND2_X1 U6781 ( .A1(n7182), .A2(n5159), .ZN(n5295) );
  NAND2_X1 U6782 ( .A1(n5296), .A2(n5295), .ZN(n7162) );
  INV_X1 U6783 ( .A(n7162), .ZN(n5297) );
  NAND2_X1 U6784 ( .A1(n5298), .A2(n5297), .ZN(n5300) );
  AND2_X1 U6785 ( .A1(n7163), .A2(n7162), .ZN(n5299) );
  AOI21_X2 U6786 ( .B1(n7161), .B2(n5300), .A(n5299), .ZN(n7323) );
  NAND2_X1 U6787 ( .A1(n6555), .A2(n7782), .ZN(n5305) );
  NAND2_X1 U6788 ( .A1(n5342), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5318) );
  XNOR2_X1 U6789 ( .A(n5318), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6644) );
  AOI22_X1 U6790 ( .A1(n5500), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6568), .B2(
        n6644), .ZN(n5304) );
  NAND2_X1 U6791 ( .A1(n5305), .A2(n5304), .ZN(n7228) );
  NAND2_X1 U6792 ( .A1(n7228), .A2(n5244), .ZN(n5312) );
  AOI22_X1 U6793 ( .A1(n4345), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n5151), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n5310) );
  AND2_X1 U6794 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  NOR2_X1 U6795 ( .A1(n5323), .A2(n5308), .ZN(n7333) );
  AOI22_X1 U6796 ( .A1(n5450), .A2(n7333), .B1(n5521), .B2(
        P1_REG0_REG_8__SCAN_IN), .ZN(n5309) );
  OR2_X1 U6797 ( .A1(n7426), .A2(n5546), .ZN(n5311) );
  NAND2_X1 U6798 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  XNOR2_X1 U6799 ( .A(n5313), .B(n5616), .ZN(n7322) );
  NAND2_X1 U6800 ( .A1(n7228), .A2(n5159), .ZN(n5315) );
  OR2_X1 U6801 ( .A1(n7426), .A2(n5618), .ZN(n5314) );
  AND2_X1 U6802 ( .A1(n5315), .A2(n5314), .ZN(n7327) );
  XNOR2_X1 U6803 ( .A(n5316), .B(n5317), .ZN(n6564) );
  NAND2_X1 U6804 ( .A1(n6564), .A2(n7782), .ZN(n5322) );
  INV_X1 U6805 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6806 ( .A1(n5318), .A2(n5340), .ZN(n5319) );
  NAND2_X1 U6807 ( .A1(n5319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5320) );
  XNOR2_X1 U6808 ( .A(n5320), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7000) );
  OR2_X1 U6809 ( .A1(n5323), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5324) );
  AND2_X1 U6810 ( .A1(n5365), .A2(n5324), .ZN(n7428) );
  NAND2_X1 U6811 ( .A1(n5450), .A2(n7428), .ZN(n5328) );
  NAND2_X1 U6812 ( .A1(n4345), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6813 ( .A1(n5151), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6814 ( .A1(n9052), .A2(n5159), .ZN(n5329) );
  NAND2_X1 U6815 ( .A1(n4343), .A2(n5159), .ZN(n5331) );
  NAND2_X1 U6816 ( .A1(n9052), .A2(n8896), .ZN(n5330) );
  NAND2_X1 U6817 ( .A1(n5331), .A2(n5330), .ZN(n5333) );
  NOR2_X1 U6818 ( .A1(n5332), .A2(n5333), .ZN(n7417) );
  AOI21_X1 U6819 ( .B1(n7322), .B2(n7327), .A(n7417), .ZN(n5336) );
  INV_X1 U6820 ( .A(n5332), .ZN(n5335) );
  INV_X1 U6821 ( .A(n5333), .ZN(n5334) );
  NOR2_X1 U6822 ( .A1(n5335), .A2(n5334), .ZN(n7418) );
  NAND2_X1 U6823 ( .A1(n6577), .A2(n7782), .ZN(n5346) );
  INV_X1 U6824 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6825 ( .A1(n5340), .A2(n5339), .ZN(n5341) );
  NOR2_X1 U6826 ( .A1(n5342), .A2(n5341), .ZN(n5361) );
  INV_X1 U6827 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6828 ( .A1(n5361), .A2(n5343), .ZN(n5387) );
  NAND2_X1 U6829 ( .A1(n5387), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5344) );
  XNOR2_X1 U6830 ( .A(n5344), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9570) );
  AOI22_X1 U6831 ( .A1(n5500), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6568), .B2(
        n9570), .ZN(n5345) );
  NAND2_X2 U6832 ( .A1(n5346), .A2(n5345), .ZN(n9691) );
  AND2_X1 U6833 ( .A1(n5367), .A2(n7588), .ZN(n5347) );
  NOR2_X1 U6834 ( .A1(n5391), .A2(n5347), .ZN(n9690) );
  NAND2_X1 U6835 ( .A1(n5450), .A2(n9690), .ZN(n5351) );
  NAND2_X1 U6836 ( .A1(n4345), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6837 ( .A1(n5151), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6838 ( .A1(n5521), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5348) );
  NAND4_X1 U6839 ( .A1(n5351), .A2(n5350), .A3(n5349), .A4(n5348), .ZN(n9050)
         );
  AOI22_X1 U6840 ( .A1(n9691), .A2(n5244), .B1(n5159), .B2(n9050), .ZN(n5352)
         );
  XOR2_X1 U6841 ( .A(n8894), .B(n5352), .Z(n7581) );
  NAND2_X1 U6842 ( .A1(n9691), .A2(n5159), .ZN(n5354) );
  NAND2_X1 U6843 ( .A1(n9050), .A2(n8896), .ZN(n5353) );
  NAND2_X1 U6844 ( .A1(n5354), .A2(n5353), .ZN(n7582) );
  INV_X1 U6845 ( .A(n5355), .ZN(n5357) );
  NAND2_X1 U6846 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  NAND2_X1 U6847 ( .A1(n5359), .A2(n5358), .ZN(n6566) );
  OR2_X1 U6848 ( .A1(n6566), .A2(n5404), .ZN(n5364) );
  OR2_X1 U6849 ( .A1(n5361), .A2(n5360), .ZN(n5362) );
  XNOR2_X1 U6850 ( .A(n5362), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9449) );
  AOI22_X1 U6851 ( .A1(n5500), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6568), .B2(
        n9449), .ZN(n5363) );
  NAND2_X1 U6852 ( .A1(n9818), .A2(n5244), .ZN(n5373) );
  NAND2_X1 U6853 ( .A1(n5365), .A2(n7499), .ZN(n5366) );
  AND2_X1 U6854 ( .A1(n5367), .A2(n5366), .ZN(n9704) );
  NAND2_X1 U6855 ( .A1(n5450), .A2(n9704), .ZN(n5371) );
  NAND2_X1 U6856 ( .A1(n4340), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6857 ( .A1(n4335), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6858 ( .A1(n5151), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5368) );
  NAND4_X1 U6859 ( .A1(n5371), .A2(n5370), .A3(n5369), .A4(n5368), .ZN(n9051)
         );
  NAND2_X1 U6860 ( .A1(n9051), .A2(n5159), .ZN(n5372) );
  NAND2_X1 U6861 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  XNOR2_X1 U6862 ( .A(n5374), .B(n5616), .ZN(n7580) );
  INV_X1 U6863 ( .A(n7580), .ZN(n5377) );
  NAND2_X1 U6864 ( .A1(n9818), .A2(n5159), .ZN(n5376) );
  NAND2_X1 U6865 ( .A1(n9051), .A2(n8896), .ZN(n5375) );
  AND2_X1 U6866 ( .A1(n5376), .A2(n5375), .ZN(n5378) );
  INV_X1 U6867 ( .A(n5378), .ZN(n7498) );
  AOI22_X1 U6868 ( .A1(n7581), .A2(n7582), .B1(n5377), .B2(n7498), .ZN(n5382)
         );
  NAND2_X1 U6869 ( .A1(n7580), .A2(n5378), .ZN(n5379) );
  AOI21_X1 U6870 ( .B1(n7582), .B2(n5379), .A(n7581), .ZN(n5381) );
  NOR2_X1 U6871 ( .A1(n5379), .A2(n7582), .ZN(n5380) );
  NAND2_X1 U6872 ( .A1(n5384), .A2(n5383), .ZN(n5386) );
  NAND2_X1 U6873 ( .A1(n5386), .A2(n5385), .ZN(n6592) );
  OR2_X1 U6874 ( .A1(n6592), .A2(n5404), .ZN(n5390) );
  NAND2_X1 U6875 ( .A1(n5388), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5406) );
  XNOR2_X1 U6876 ( .A(n5406), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9077) );
  AOI22_X1 U6877 ( .A1(n5500), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6568), .B2(
        n9077), .ZN(n5389) );
  NAND2_X1 U6878 ( .A1(n9665), .A2(n5244), .ZN(n5396) );
  AOI22_X1 U6879 ( .A1(n4345), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n5151), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n5394) );
  NOR2_X1 U6880 ( .A1(n5391), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5392) );
  AOI22_X1 U6881 ( .A1(n5450), .A2(n4962), .B1(n4335), .B2(
        P1_REG0_REG_12__SCAN_IN), .ZN(n5393) );
  OR2_X1 U6882 ( .A1(n7585), .A2(n5546), .ZN(n5395) );
  NAND2_X1 U6883 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  XNOR2_X1 U6884 ( .A(n5397), .B(n8894), .ZN(n5399) );
  OAI22_X1 U6885 ( .A1(n9833), .A2(n5546), .B1(n7585), .B2(n5618), .ZN(n5398)
         );
  XNOR2_X1 U6886 ( .A(n5399), .B(n5398), .ZN(n7464) );
  OR2_X1 U6887 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  NAND2_X1 U6888 ( .A1(n5403), .A2(n5402), .ZN(n6613) );
  OR2_X1 U6889 ( .A1(n6613), .A2(n5404), .ZN(n5410) );
  INV_X1 U6890 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6891 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  NAND2_X1 U6892 ( .A1(n5407), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5408) );
  XNOR2_X1 U6893 ( .A(n5408), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9589) );
  AOI22_X1 U6894 ( .A1(n5500), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6568), .B2(
        n9589), .ZN(n5409) );
  OR2_X1 U6895 ( .A1(n5411), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5412) );
  AND2_X1 U6896 ( .A1(n5447), .A2(n5412), .ZN(n7517) );
  NAND2_X1 U6897 ( .A1(n6478), .A2(n7517), .ZN(n5416) );
  NAND2_X1 U6898 ( .A1(n4345), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6899 ( .A1(n5521), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6900 ( .A1(n5520), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5413) );
  NAND4_X1 U6901 ( .A1(n5416), .A2(n5415), .A3(n5414), .A4(n5413), .ZN(n9048)
         );
  AOI22_X1 U6902 ( .A1(n7521), .A2(n5244), .B1(n5159), .B2(n9048), .ZN(n5417)
         );
  XNOR2_X1 U6903 ( .A(n5417), .B(n8894), .ZN(n5419) );
  INV_X1 U6904 ( .A(n9048), .ZN(n7558) );
  OAI22_X1 U6905 ( .A1(n9839), .A2(n5546), .B1(n7558), .B2(n5618), .ZN(n5418)
         );
  XNOR2_X1 U6906 ( .A(n5419), .B(n5418), .ZN(n7516) );
  INV_X1 U6907 ( .A(n5418), .ZN(n5420) );
  AOI22_X2 U6908 ( .A1(n7515), .A2(n7516), .B1(n5420), .B2(n5419), .ZN(n7554)
         );
  INV_X1 U6909 ( .A(n7554), .ZN(n5423) );
  INV_X1 U6910 ( .A(n9047), .ZN(n9024) );
  OAI22_X1 U6911 ( .A1(n9847), .A2(n5546), .B1(n9024), .B2(n5618), .ZN(n7551)
         );
  AOI21_X1 U6912 ( .B1(n7554), .B2(n5421), .A(n7551), .ZN(n5422) );
  AOI21_X1 U6913 ( .B1(n7552), .B2(n5423), .A(n5422), .ZN(n8936) );
  INV_X1 U6914 ( .A(n8936), .ZN(n5468) );
  XNOR2_X1 U6915 ( .A(n5425), .B(SI_16_), .ZN(n5426) );
  XNOR2_X1 U6916 ( .A(n5424), .B(n5426), .ZN(n6855) );
  NAND2_X1 U6917 ( .A1(n6855), .A2(n7782), .ZN(n5431) );
  NAND2_X1 U6918 ( .A1(n5428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5429) );
  XNOR2_X1 U6919 ( .A(n5429), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9095) );
  AOI22_X1 U6920 ( .A1(n5500), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6568), .B2(
        n9095), .ZN(n5430) );
  NAND2_X1 U6921 ( .A1(n9512), .A2(n5244), .ZN(n5436) );
  AND2_X1 U6922 ( .A1(n5448), .A2(n10167), .ZN(n5432) );
  NOR2_X1 U6923 ( .A1(n5473), .A2(n5432), .ZN(n8946) );
  AOI22_X1 U6924 ( .A1(n6478), .A2(n8946), .B1(n5520), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n5434) );
  AOI22_X1 U6925 ( .A1(n4340), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n5521), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5433) );
  OR2_X1 U6926 ( .A1(n9026), .A2(n5546), .ZN(n5435) );
  NAND2_X1 U6927 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  XNOR2_X1 U6928 ( .A(n5437), .B(n5616), .ZN(n8940) );
  NOR2_X1 U6929 ( .A1(n9026), .A2(n5618), .ZN(n5438) );
  AOI21_X1 U6930 ( .B1(n9512), .B2(n5159), .A(n5438), .ZN(n8939) );
  XNOR2_X1 U6931 ( .A(n5439), .B(SI_15_), .ZN(n5440) );
  XNOR2_X1 U6932 ( .A(n5441), .B(n5440), .ZN(n6775) );
  NAND2_X1 U6933 ( .A1(n6775), .A2(n7782), .ZN(n5445) );
  NAND2_X1 U6934 ( .A1(n5442), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5443) );
  XNOR2_X1 U6935 ( .A(n5443), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9638) );
  AOI22_X1 U6936 ( .A1(n5500), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6568), .B2(
        n9638), .ZN(n5444) );
  NAND2_X1 U6937 ( .A1(n9402), .A2(n5244), .ZN(n5456) );
  OAI21_X1 U6938 ( .B1(n5447), .B2(n5446), .A(n9023), .ZN(n5449) );
  AND2_X1 U6939 ( .A1(n5449), .A2(n5448), .ZN(n9031) );
  NAND2_X1 U6940 ( .A1(n5450), .A2(n9031), .ZN(n5454) );
  NAND2_X1 U6941 ( .A1(n4345), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6942 ( .A1(n5520), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6943 ( .A1(n4335), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5451) );
  NAND4_X1 U6944 ( .A1(n5454), .A2(n5453), .A3(n5452), .A4(n5451), .ZN(n9046)
         );
  NAND2_X1 U6945 ( .A1(n9046), .A2(n5159), .ZN(n5455) );
  NAND2_X1 U6946 ( .A1(n5456), .A2(n5455), .ZN(n5457) );
  XNOR2_X1 U6947 ( .A(n5457), .B(n8894), .ZN(n8938) );
  NAND2_X1 U6948 ( .A1(n9402), .A2(n5159), .ZN(n5459) );
  NAND2_X1 U6949 ( .A1(n9046), .A2(n8896), .ZN(n5458) );
  NAND2_X1 U6950 ( .A1(n5459), .A2(n5458), .ZN(n5461) );
  NAND2_X1 U6951 ( .A1(n8938), .A2(n5461), .ZN(n5460) );
  INV_X1 U6952 ( .A(n8939), .ZN(n5463) );
  INV_X1 U6953 ( .A(n8938), .ZN(n8937) );
  INV_X1 U6954 ( .A(n5461), .ZN(n9020) );
  NAND2_X1 U6955 ( .A1(n8937), .A2(n9020), .ZN(n5464) );
  INV_X1 U6956 ( .A(n8940), .ZN(n5462) );
  AOI21_X1 U6957 ( .B1(n5463), .B2(n5464), .A(n5462), .ZN(n5466) );
  XNOR2_X1 U6958 ( .A(n5470), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9110) );
  AOI22_X1 U6959 ( .A1(n5500), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6568), .B2(
        n9110), .ZN(n5471) );
  NAND2_X1 U6960 ( .A1(n9323), .A2(n5150), .ZN(n5481) );
  OR2_X1 U6961 ( .A1(n5473), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5474) );
  AND2_X1 U6962 ( .A1(n5475), .A2(n5474), .ZN(n9314) );
  NAND2_X1 U6963 ( .A1(n6478), .A2(n9314), .ZN(n5479) );
  NAND2_X1 U6964 ( .A1(n4340), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U6965 ( .A1(n4335), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6966 ( .A1(n5520), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5476) );
  NAND4_X1 U6967 ( .A1(n5479), .A2(n5478), .A3(n5477), .A4(n5476), .ZN(n9301)
         );
  NAND2_X1 U6968 ( .A1(n9301), .A2(n5159), .ZN(n5480) );
  NAND2_X1 U6969 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  XNOR2_X1 U6970 ( .A(n5482), .B(n5616), .ZN(n5485) );
  AND2_X1 U6971 ( .A1(n9301), .A2(n8896), .ZN(n5483) );
  AOI21_X1 U6972 ( .B1(n9323), .B2(n5159), .A(n5483), .ZN(n5484) );
  NOR2_X1 U6973 ( .A1(n5485), .A2(n5484), .ZN(n5486) );
  AOI21_X1 U6974 ( .B1(n5485), .B2(n5484), .A(n5486), .ZN(n8951) );
  NAND2_X1 U6975 ( .A1(n8952), .A2(n8951), .ZN(n8950) );
  INV_X1 U6976 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U6977 ( .A1(n8950), .A2(n5487), .ZN(n5490) );
  OAI22_X1 U6978 ( .A1(n9297), .A2(n5524), .B1(n8886), .B2(n5546), .ZN(n5488)
         );
  XNOR2_X1 U6979 ( .A(n5488), .B(n8894), .ZN(n5489) );
  NAND2_X1 U6980 ( .A1(n5490), .A2(n5489), .ZN(n8989) );
  NOR2_X1 U6981 ( .A1(n5490), .A2(n5489), .ZN(n8988) );
  AOI21_X2 U6982 ( .B1(n8991), .B2(n8989), .A(n8988), .ZN(n8884) );
  INV_X1 U6983 ( .A(n5492), .ZN(n5493) );
  INV_X1 U6984 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7160) );
  INV_X1 U6985 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7728) );
  MUX2_X1 U6986 ( .A(n7160), .B(n7728), .S(n7795), .Z(n5497) );
  INV_X1 U6987 ( .A(SI_19_), .ZN(n5496) );
  INV_X1 U6988 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U6989 ( .A1(n5498), .A2(SI_19_), .ZN(n5499) );
  NAND2_X1 U6990 ( .A1(n5512), .A2(n5499), .ZN(n5513) );
  XNOR2_X1 U6991 ( .A(n5514), .B(n5513), .ZN(n7159) );
  NAND2_X1 U6992 ( .A1(n7159), .A2(n7782), .ZN(n5502) );
  AOI22_X1 U6993 ( .A1(n5500), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9747), .B2(
        n6568), .ZN(n5501) );
  INV_X1 U6994 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8885) );
  AND2_X1 U6995 ( .A1(n5503), .A2(n8885), .ZN(n5504) );
  OR2_X1 U6996 ( .A1(n5504), .A2(n5518), .ZN(n9283) );
  AOI22_X1 U6997 ( .A1(n4345), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n5520), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U6998 ( .A1(n4335), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5505) );
  OAI211_X1 U6999 ( .C1(n9283), .C2(n5126), .A(n5506), .B(n5505), .ZN(n9302)
         );
  INV_X1 U7000 ( .A(n9302), .ZN(n8972) );
  OAI22_X1 U7001 ( .A1(n9392), .A2(n5524), .B1(n8972), .B2(n5546), .ZN(n5507)
         );
  XNOR2_X1 U7002 ( .A(n5507), .B(n5616), .ZN(n5511) );
  OR2_X1 U7003 ( .A1(n9392), .A2(n5546), .ZN(n5509) );
  NAND2_X1 U7004 ( .A1(n9302), .A2(n8896), .ZN(n5508) );
  AND2_X1 U7005 ( .A1(n5509), .A2(n5508), .ZN(n5510) );
  NOR2_X1 U7006 ( .A1(n5511), .A2(n5510), .ZN(n8882) );
  NAND2_X1 U7007 ( .A1(n5511), .A2(n5510), .ZN(n8880) );
  OAI21_X1 U7008 ( .B1(n8884), .B2(n8882), .A(n8880), .ZN(n8969) );
  MUX2_X1 U7009 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7795), .Z(n5532) );
  INV_X1 U7010 ( .A(SI_20_), .ZN(n5534) );
  XNOR2_X1 U7011 ( .A(n5532), .B(n5534), .ZN(n5515) );
  XNOR2_X1 U7012 ( .A(n5535), .B(n5515), .ZN(n7188) );
  NAND2_X1 U7013 ( .A1(n7188), .A2(n7782), .ZN(n5517) );
  INV_X1 U7014 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7189) );
  OR2_X1 U7015 ( .A1(n4341), .A2(n7189), .ZN(n5516) );
  NOR2_X1 U7016 ( .A1(n5518), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5519) );
  OR2_X1 U7017 ( .A1(n5541), .A2(n5519), .ZN(n9262) );
  AOI22_X1 U7018 ( .A1(n4345), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n5520), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7019 ( .A1(n4335), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5522) );
  OAI211_X1 U7020 ( .C1(n9262), .C2(n5126), .A(n5523), .B(n5522), .ZN(n9278)
         );
  INV_X1 U7021 ( .A(n9278), .ZN(n8917) );
  OAI22_X1 U7022 ( .A1(n9265), .A2(n5524), .B1(n8917), .B2(n5546), .ZN(n5525)
         );
  XNOR2_X1 U7023 ( .A(n5525), .B(n8894), .ZN(n5529) );
  OR2_X1 U7024 ( .A1(n9265), .A2(n5546), .ZN(n5527) );
  NAND2_X1 U7025 ( .A1(n9278), .A2(n8896), .ZN(n5526) );
  NAND2_X1 U7026 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  NOR2_X1 U7027 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  AOI21_X1 U7028 ( .B1(n5529), .B2(n5528), .A(n5530), .ZN(n8970) );
  INV_X1 U7029 ( .A(n5530), .ZN(n5531) );
  INV_X1 U7030 ( .A(n5532), .ZN(n5533) );
  NAND2_X1 U7031 ( .A1(n5537), .A2(n5536), .ZN(n5558) );
  INV_X1 U7032 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7235) );
  INV_X1 U7033 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7205) );
  MUX2_X1 U7034 ( .A(n7235), .B(n7205), .S(n7795), .Z(n5554) );
  XNOR2_X1 U7035 ( .A(n5554), .B(SI_21_), .ZN(n5538) );
  XNOR2_X1 U7036 ( .A(n5558), .B(n5538), .ZN(n7204) );
  NAND2_X1 U7037 ( .A1(n7204), .A2(n7782), .ZN(n5540) );
  OR2_X1 U7038 ( .A1(n4341), .A2(n7205), .ZN(n5539) );
  NAND2_X1 U7039 ( .A1(n9381), .A2(n5150), .ZN(n5548) );
  NAND2_X1 U7040 ( .A1(n5541), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5565) );
  OR2_X1 U7041 ( .A1(n5541), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5542) );
  AND2_X1 U7042 ( .A1(n5565), .A2(n5542), .ZN(n9249) );
  NAND2_X1 U7043 ( .A1(n9249), .A2(n6478), .ZN(n5545) );
  AOI22_X1 U7044 ( .A1(n5520), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5521), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7045 ( .A1(n4340), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5543) );
  OR2_X1 U7046 ( .A1(n8982), .A2(n5546), .ZN(n5547) );
  NAND2_X1 U7047 ( .A1(n5548), .A2(n5547), .ZN(n5549) );
  XNOR2_X1 U7048 ( .A(n5549), .B(n8894), .ZN(n5552) );
  INV_X1 U7049 ( .A(n8982), .ZN(n9045) );
  AOI22_X1 U7050 ( .A1(n9381), .A2(n5159), .B1(n8896), .B2(n9045), .ZN(n5550)
         );
  XNOR2_X1 U7051 ( .A(n5552), .B(n5550), .ZN(n8915) );
  INV_X1 U7052 ( .A(n5550), .ZN(n5551) );
  NOR2_X1 U7053 ( .A1(n5555), .A2(SI_21_), .ZN(n5557) );
  NAND2_X1 U7054 ( .A1(n5555), .A2(SI_21_), .ZN(n5556) );
  INV_X1 U7055 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7321) );
  MUX2_X1 U7056 ( .A(n10086), .B(n7321), .S(n7795), .Z(n5560) );
  INV_X1 U7057 ( .A(SI_22_), .ZN(n5559) );
  NAND2_X1 U7058 ( .A1(n5560), .A2(n5559), .ZN(n5575) );
  INV_X1 U7059 ( .A(n5560), .ZN(n5561) );
  NAND2_X1 U7060 ( .A1(n5561), .A2(SI_22_), .ZN(n5562) );
  NAND2_X1 U7061 ( .A1(n5575), .A2(n5562), .ZN(n5576) );
  XNOR2_X1 U7062 ( .A(n5577), .B(n5576), .ZN(n7317) );
  NAND2_X1 U7063 ( .A1(n7317), .A2(n7782), .ZN(n5564) );
  OR2_X1 U7064 ( .A1(n4342), .A2(n7321), .ZN(n5563) );
  INV_X1 U7065 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U7066 ( .A1(n5565), .A2(n8983), .ZN(n5566) );
  NAND2_X1 U7067 ( .A1(n5584), .A2(n5566), .ZN(n9229) );
  OR2_X1 U7068 ( .A1(n9229), .A2(n5126), .ZN(n5572) );
  INV_X1 U7069 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7070 ( .A1(n4335), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7071 ( .A1(n5520), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5567) );
  OAI211_X1 U7072 ( .C1(n5569), .C2(n4337), .A(n5568), .B(n5567), .ZN(n5570)
         );
  INV_X1 U7073 ( .A(n5570), .ZN(n5571) );
  INV_X1 U7074 ( .A(n8918), .ZN(n9044) );
  AOI22_X1 U7075 ( .A1(n9376), .A2(n5150), .B1(n5159), .B2(n9044), .ZN(n5573)
         );
  XNOR2_X1 U7076 ( .A(n5573), .B(n8894), .ZN(n5574) );
  OAI22_X1 U7077 ( .A1(n6520), .A2(n5546), .B1(n8918), .B2(n5618), .ZN(n8979)
         );
  INV_X1 U7078 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7413) );
  INV_X1 U7079 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7416) );
  MUX2_X1 U7080 ( .A(n7413), .B(n7416), .S(n7795), .Z(n5579) );
  INV_X1 U7081 ( .A(SI_23_), .ZN(n5578) );
  NAND2_X1 U7082 ( .A1(n5579), .A2(n5578), .ZN(n5600) );
  INV_X1 U7083 ( .A(n5579), .ZN(n5580) );
  NAND2_X1 U7084 ( .A1(n5580), .A2(SI_23_), .ZN(n5581) );
  NAND2_X1 U7085 ( .A1(n6078), .A2(n7782), .ZN(n5583) );
  OR2_X1 U7086 ( .A1(n4341), .A2(n7416), .ZN(n5582) );
  NAND2_X1 U7087 ( .A1(n9371), .A2(n5150), .ZN(n5591) );
  INV_X1 U7088 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U7089 ( .A1(n5584), .A2(n8875), .ZN(n5585) );
  AND2_X1 U7090 ( .A1(n5608), .A2(n5585), .ZN(n9213) );
  INV_X1 U7091 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7092 ( .A1(n5520), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7093 ( .A1(n4335), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5586) );
  OAI211_X1 U7094 ( .C1(n4337), .C2(n5588), .A(n5587), .B(n5586), .ZN(n5589)
         );
  AOI21_X1 U7095 ( .B1(n9213), .B2(n6478), .A(n5589), .ZN(n8980) );
  OR2_X1 U7096 ( .A1(n8980), .A2(n5546), .ZN(n5590) );
  NAND2_X1 U7097 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  XNOR2_X1 U7098 ( .A(n5592), .B(n5616), .ZN(n5595) );
  NOR2_X1 U7099 ( .A1(n8980), .A2(n5618), .ZN(n5593) );
  AOI21_X1 U7100 ( .B1(n9371), .B2(n5159), .A(n5593), .ZN(n5594) );
  NAND2_X1 U7101 ( .A1(n5595), .A2(n5594), .ZN(n8962) );
  OR2_X1 U7102 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  NAND2_X2 U7103 ( .A1(n5597), .A2(n8870), .ZN(n8872) );
  INV_X1 U7104 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10055) );
  INV_X1 U7105 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7564) );
  MUX2_X1 U7106 ( .A(n10055), .B(n7564), .S(n7795), .Z(n5602) );
  INV_X1 U7107 ( .A(SI_24_), .ZN(n5601) );
  NAND2_X1 U7108 ( .A1(n5602), .A2(n5601), .ZN(n5625) );
  INV_X1 U7109 ( .A(n5602), .ZN(n5603) );
  NAND2_X1 U7110 ( .A1(n5603), .A2(SI_24_), .ZN(n5604) );
  XNOR2_X1 U7111 ( .A(n5624), .B(n5623), .ZN(n7563) );
  NAND2_X1 U7112 ( .A1(n7563), .A2(n7782), .ZN(n5606) );
  OR2_X1 U7113 ( .A1(n4342), .A2(n7564), .ZN(n5605) );
  NAND2_X1 U7114 ( .A1(n9367), .A2(n5150), .ZN(n5615) );
  INV_X1 U7115 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5607) );
  AND2_X1 U7116 ( .A1(n5608), .A2(n5607), .ZN(n5609) );
  INV_X1 U7117 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7118 ( .A1(n5520), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7119 ( .A1(n4335), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U7120 ( .C1(n4336), .C2(n5612), .A(n5611), .B(n5610), .ZN(n5613)
         );
  AOI21_X1 U7121 ( .B1(n4968), .B2(n6478), .A(n5613), .ZN(n8928) );
  OR2_X1 U7122 ( .A1(n8928), .A2(n5546), .ZN(n5614) );
  NAND2_X1 U7123 ( .A1(n5615), .A2(n5614), .ZN(n5617) );
  XNOR2_X1 U7124 ( .A(n5617), .B(n5616), .ZN(n5621) );
  NOR2_X1 U7125 ( .A1(n8928), .A2(n5618), .ZN(n5619) );
  AOI21_X1 U7126 ( .B1(n9367), .B2(n5159), .A(n5619), .ZN(n5620) );
  NAND2_X1 U7127 ( .A1(n5621), .A2(n5620), .ZN(n8925) );
  OR2_X1 U7128 ( .A1(n5621), .A2(n5620), .ZN(n5622) );
  NAND2_X1 U7129 ( .A1(n5624), .A2(n5623), .ZN(n5626) );
  NAND2_X1 U7130 ( .A1(n5626), .A2(n5625), .ZN(n5650) );
  INV_X1 U7131 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7594) );
  INV_X1 U7132 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7577) );
  MUX2_X1 U7133 ( .A(n7594), .B(n7577), .S(n7795), .Z(n5628) );
  INV_X1 U7134 ( .A(SI_25_), .ZN(n5627) );
  NAND2_X1 U7135 ( .A1(n5628), .A2(n5627), .ZN(n5669) );
  INV_X1 U7136 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U7137 ( .A1(n5629), .A2(SI_25_), .ZN(n5630) );
  XNOR2_X1 U7138 ( .A(n5650), .B(n5649), .ZN(n7575) );
  NAND2_X1 U7139 ( .A1(n7575), .A2(n7782), .ZN(n5632) );
  OR2_X1 U7140 ( .A1(n4342), .A2(n7577), .ZN(n5631) );
  OR2_X1 U7141 ( .A1(n5633), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7142 ( .A1(n5633), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5659) );
  AND2_X1 U7143 ( .A1(n5634), .A2(n5659), .ZN(n9186) );
  NAND2_X1 U7144 ( .A1(n9186), .A2(n6478), .ZN(n5640) );
  INV_X1 U7145 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7146 ( .A1(n5521), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7147 ( .A1(n5520), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5635) );
  OAI211_X1 U7148 ( .C1(n5637), .C2(n4336), .A(n5636), .B(n5635), .ZN(n5638)
         );
  INV_X1 U7149 ( .A(n5638), .ZN(n5639) );
  NAND2_X1 U7150 ( .A1(n5640), .A2(n5639), .ZN(n9041) );
  AOI22_X1 U7151 ( .A1(n9361), .A2(n5150), .B1(n5159), .B2(n9041), .ZN(n5641)
         );
  XNOR2_X1 U7152 ( .A(n5641), .B(n8894), .ZN(n5648) );
  OR2_X1 U7153 ( .A1(n9188), .A2(n5546), .ZN(n5643) );
  NAND2_X1 U7154 ( .A1(n9041), .A2(n8896), .ZN(n5642) );
  NAND2_X1 U7155 ( .A1(n5643), .A2(n5642), .ZN(n5646) );
  XNOR2_X1 U7156 ( .A(n5648), .B(n5646), .ZN(n8927) );
  AND2_X1 U7157 ( .A1(n8960), .A2(n8927), .ZN(n5645) );
  INV_X1 U7158 ( .A(n8927), .ZN(n5644) );
  INV_X1 U7159 ( .A(n5646), .ZN(n5647) );
  NAND2_X1 U7160 ( .A1(n5648), .A2(n5647), .ZN(n9001) );
  NAND2_X1 U7161 ( .A1(n5650), .A2(n5649), .ZN(n5673) );
  NAND2_X1 U7162 ( .A1(n5673), .A2(n5669), .ZN(n5655) );
  INV_X1 U7163 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10218) );
  INV_X1 U7164 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10169) );
  MUX2_X1 U7165 ( .A(n10218), .B(n10169), .S(n7795), .Z(n5652) );
  INV_X1 U7166 ( .A(SI_26_), .ZN(n5651) );
  NAND2_X1 U7167 ( .A1(n5652), .A2(n5651), .ZN(n5668) );
  INV_X1 U7168 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U7169 ( .A1(n5653), .A2(SI_26_), .ZN(n5670) );
  AND2_X1 U7170 ( .A1(n5668), .A2(n5670), .ZN(n5654) );
  NAND2_X1 U7171 ( .A1(n7614), .A2(n7782), .ZN(n5657) );
  OR2_X1 U7172 ( .A1(n4341), .A2(n10169), .ZN(n5656) );
  NAND2_X1 U7173 ( .A1(n9356), .A2(n5150), .ZN(n5665) );
  INV_X1 U7174 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9011) );
  INV_X1 U7175 ( .A(n5659), .ZN(n5658) );
  NAND2_X1 U7176 ( .A1(n5658), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5680) );
  INV_X1 U7177 ( .A(n5680), .ZN(n5738) );
  AOI21_X1 U7178 ( .B1(n9011), .B2(n5659), .A(n5738), .ZN(n9010) );
  NAND2_X1 U7179 ( .A1(n6478), .A2(n9010), .ZN(n5663) );
  NAND2_X1 U7180 ( .A1(n4340), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7181 ( .A1(n4335), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7182 ( .A1(n5520), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5660) );
  NAND4_X1 U7183 ( .A1(n5663), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n9040)
         );
  NAND2_X1 U7184 ( .A1(n9040), .A2(n5159), .ZN(n5664) );
  NAND2_X1 U7185 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  XNOR2_X1 U7186 ( .A(n5666), .B(n8894), .ZN(n5694) );
  AND2_X1 U7187 ( .A1(n9040), .A2(n8896), .ZN(n5667) );
  AOI21_X1 U7188 ( .B1(n9356), .B2(n5159), .A(n5667), .ZN(n5692) );
  XNOR2_X1 U7189 ( .A(n5694), .B(n5692), .ZN(n9004) );
  AND2_X1 U7190 ( .A1(n5669), .A2(n5668), .ZN(n5672) );
  INV_X1 U7191 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8018) );
  INV_X1 U7192 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7625) );
  MUX2_X1 U7193 ( .A(n8018), .B(n7625), .S(n7795), .Z(n5675) );
  INV_X1 U7194 ( .A(SI_27_), .ZN(n5674) );
  NAND2_X1 U7195 ( .A1(n5675), .A2(n5674), .ZN(n6135) );
  INV_X1 U7196 ( .A(n5675), .ZN(n5676) );
  NAND2_X1 U7197 ( .A1(n5676), .A2(SI_27_), .ZN(n5677) );
  NAND2_X1 U7198 ( .A1(n7624), .A2(n7782), .ZN(n5679) );
  OR2_X1 U7199 ( .A1(n4341), .A2(n7625), .ZN(n5678) );
  NAND2_X1 U7200 ( .A1(n9352), .A2(n5150), .ZN(n5686) );
  XNOR2_X1 U7201 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n5680), .ZN(n9160) );
  NAND2_X1 U7202 ( .A1(n6478), .A2(n9160), .ZN(n5684) );
  NAND2_X1 U7203 ( .A1(n4345), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7204 ( .A1(n5520), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7205 ( .A1(n4335), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5681) );
  NAND4_X1 U7206 ( .A1(n5684), .A2(n5683), .A3(n5682), .A4(n5681), .ZN(n9039)
         );
  NAND2_X1 U7207 ( .A1(n9039), .A2(n5159), .ZN(n5685) );
  NAND2_X1 U7208 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  XNOR2_X1 U7209 ( .A(n5687), .B(n8894), .ZN(n5691) );
  NAND2_X1 U7210 ( .A1(n9352), .A2(n5159), .ZN(n5689) );
  NAND2_X1 U7211 ( .A1(n9039), .A2(n8896), .ZN(n5688) );
  NAND2_X1 U7212 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  NOR2_X1 U7213 ( .A1(n5691), .A2(n5690), .ZN(n8907) );
  AOI21_X1 U7214 ( .B1(n5691), .B2(n5690), .A(n8907), .ZN(n5696) );
  INV_X1 U7215 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U7216 ( .A1(n5694), .A2(n5693), .ZN(n5697) );
  AOI21_X1 U7217 ( .B1(n9003), .B2(n5697), .A(n5696), .ZN(n5721) );
  NAND2_X1 U7218 ( .A1(n7565), .A2(P1_B_REG_SCAN_IN), .ZN(n5699) );
  INV_X1 U7219 ( .A(P1_B_REG_SCAN_IN), .ZN(n10211) );
  NAND2_X1 U7220 ( .A1(n5711), .A2(n10211), .ZN(n5698) );
  OAI211_X1 U7221 ( .C1(n7576), .C2(n5699), .A(n7615), .B(n5698), .ZN(n9421)
         );
  NOR4_X1 U7222 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5703) );
  NOR4_X1 U7223 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5702) );
  NOR4_X1 U7224 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5701) );
  NOR4_X1 U7225 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5700) );
  NAND4_X1 U7226 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .ZN(n5709)
         );
  NOR2_X1 U7227 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .ZN(
        n5707) );
  NOR4_X1 U7228 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5706) );
  NOR4_X1 U7229 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5705) );
  NOR4_X1 U7230 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5704) );
  NAND4_X1 U7231 ( .A1(n5707), .A2(n5706), .A3(n5705), .A4(n5704), .ZN(n5708)
         );
  NOR2_X1 U7232 ( .A1(n5709), .A2(n5708), .ZN(n7257) );
  AND2_X1 U7233 ( .A1(n7257), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5710) );
  OR2_X1 U7234 ( .A1(n7615), .A2(n7576), .ZN(n9424) );
  OAI21_X1 U7235 ( .B1(n9421), .B2(n5710), .A(n9424), .ZN(n6486) );
  OR2_X1 U7236 ( .A1(n9421), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5712) );
  OR2_X1 U7237 ( .A1(n5711), .A2(n7615), .ZN(n9425) );
  NAND2_X1 U7238 ( .A1(n5712), .A2(n9425), .ZN(n9333) );
  NOR2_X1 U7239 ( .A1(n6486), .A2(n9333), .ZN(n5730) );
  NAND2_X1 U7240 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  NAND2_X1 U7241 ( .A1(n5715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5717) );
  INV_X1 U7242 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5716) );
  INV_X1 U7243 ( .A(n9423), .ZN(n5719) );
  AND2_X1 U7244 ( .A1(n5730), .A2(n5719), .ZN(n5746) );
  NAND2_X1 U7245 ( .A1(n5096), .A2(n7739), .ZN(n7980) );
  INV_X1 U7246 ( .A(n7980), .ZN(n6570) );
  NOR2_X1 U7247 ( .A1(n9787), .A2(n6570), .ZN(n5722) );
  OAI21_X1 U7248 ( .B1(n4757), .B2(n5721), .A(n9021), .ZN(n5755) );
  INV_X1 U7249 ( .A(n5722), .ZN(n5725) );
  INV_X1 U7250 ( .A(n8008), .ZN(n6490) );
  NOR2_X1 U7251 ( .A1(n7980), .A2(n6490), .ZN(n6485) );
  NOR2_X1 U7252 ( .A1(n6485), .A2(n5723), .ZN(n5724) );
  OAI21_X1 U7253 ( .B1(n5725), .B2(n5730), .A(n5724), .ZN(n5726) );
  NAND2_X1 U7254 ( .A1(n5726), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5736) );
  INV_X1 U7255 ( .A(n5727), .ZN(n6491) );
  NAND2_X1 U7256 ( .A1(n6491), .A2(n5728), .ZN(n9743) );
  AND2_X1 U7257 ( .A1(n9763), .A2(n8000), .ZN(n6522) );
  NAND2_X1 U7258 ( .A1(n6522), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5729) );
  OAI21_X1 U7259 ( .B1(n9743), .B2(n9423), .A(n5729), .ZN(n5734) );
  INV_X1 U7260 ( .A(n5730), .ZN(n5733) );
  INV_X1 U7261 ( .A(n6569), .ZN(n5731) );
  NAND2_X1 U7262 ( .A1(n5731), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8015) );
  INV_X1 U7263 ( .A(n8015), .ZN(n5732) );
  AOI21_X1 U7264 ( .B1(n5734), .B2(n5733), .A(n5732), .ZN(n5735) );
  INV_X1 U7265 ( .A(n5737), .ZN(n6647) );
  NAND3_X1 U7266 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .A3(n5738), .ZN(n6477) );
  INV_X1 U7267 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7268 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5738), .ZN(n5739) );
  NAND2_X1 U7269 ( .A1(n5740), .A2(n5739), .ZN(n5741) );
  NAND2_X1 U7270 ( .A1(n6478), .A2(n8902), .ZN(n5745) );
  NAND2_X1 U7271 ( .A1(n4345), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7272 ( .A1(n5520), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7273 ( .A1(n5521), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5742) );
  NAND4_X1 U7274 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n9038)
         );
  AOI22_X1 U7275 ( .A1(n9311), .A2(n9038), .B1(n9040), .B2(n9309), .ZN(n9167)
         );
  INV_X1 U7276 ( .A(n5746), .ZN(n5750) );
  OR2_X1 U7277 ( .A1(n5750), .A2(n8008), .ZN(n8959) );
  INV_X1 U7278 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5747) );
  OAI22_X1 U7279 ( .A1(n9167), .A2(n8959), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5747), .ZN(n5748) );
  AOI21_X1 U7280 ( .B1(n9160), .B2(n9030), .A(n5748), .ZN(n5754) );
  INV_X1 U7281 ( .A(n9352), .ZN(n6473) );
  NAND2_X1 U7282 ( .A1(n9734), .A2(n9747), .ZN(n7261) );
  INV_X1 U7283 ( .A(n6522), .ZN(n9745) );
  OR2_X1 U7284 ( .A1(n5750), .A2(n9745), .ZN(n5751) );
  NAND2_X1 U7285 ( .A1(n9352), .A2(n5752), .ZN(n5753) );
  NAND3_X1 U7286 ( .A1(n5755), .A2(n5754), .A3(n5753), .ZN(P1_U3214) );
  NOR2_X1 U7287 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5762) );
  NAND4_X1 U7288 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n5764)
         );
  NAND3_X1 U7289 ( .A1(n6016), .A2(n6021), .A3(n6037), .ZN(n5763) );
  INV_X1 U7290 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8861) );
  INV_X1 U7291 ( .A(n7666), .ZN(n5771) );
  INV_X1 U7292 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6955) );
  NAND2_X1 U7293 ( .A1(n5771), .A2(n5770), .ZN(n5790) );
  INV_X1 U7294 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6689) );
  OR2_X1 U7295 ( .A1(n5790), .A2(n6689), .ZN(n5773) );
  AND2_X4 U7296 ( .A1(n7666), .A2(n7654), .ZN(n6095) );
  NAND2_X1 U7297 ( .A1(n6095), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5772) );
  INV_X1 U7298 ( .A(n6303), .ZN(n6809) );
  NAND2_X2 U7299 ( .A1(n5827), .A2(n7795), .ZN(n5824) );
  INV_X1 U7300 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5780) );
  OAI22_X1 U7301 ( .A1(n5824), .A2(n6550), .B1(n5827), .B2(n6714), .ZN(n5781)
         );
  INV_X1 U7302 ( .A(n5781), .ZN(n5783) );
  OR2_X1 U7303 ( .A1(n5842), .A2(n6549), .ZN(n5782) );
  NAND2_X1 U7304 ( .A1(n6809), .A2(n4339), .ZN(n8077) );
  NAND2_X2 U7305 ( .A1(n8077), .A2(n8081), .ZN(n6213) );
  INV_X1 U7306 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6606) );
  OR2_X1 U7307 ( .A1(n5828), .A2(n6606), .ZN(n5787) );
  INV_X1 U7308 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6662) );
  OR2_X1 U7309 ( .A1(n5790), .A2(n6662), .ZN(n5786) );
  NAND2_X1 U7310 ( .A1(n5885), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7311 ( .A1(n6095), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5784) );
  INV_X1 U7312 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U7313 ( .A1(n4992), .A2(SI_0_), .ZN(n5789) );
  INV_X1 U7314 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5788) );
  XNOR2_X1 U7315 ( .A(n5789), .B(n5788), .ZN(n8867) );
  MUX2_X1 U7316 ( .A(n6712), .B(n8867), .S(n5827), .Z(n6848) );
  NAND2_X1 U7317 ( .A1(n6946), .A2(n6214), .ZN(n6948) );
  NAND2_X1 U7318 ( .A1(n6303), .A2(n4339), .ZN(n8721) );
  NAND2_X1 U7319 ( .A1(n6947), .A2(n8721), .ZN(n5802) );
  INV_X1 U7320 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5791) );
  INV_X1 U7321 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5792) );
  OR2_X1 U7322 ( .A1(n5832), .A2(n5792), .ZN(n5797) );
  INV_X1 U7323 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5793) );
  INV_X1 U7324 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5794) );
  OR2_X1 U7325 ( .A1(n5842), .A2(n6553), .ZN(n5801) );
  NAND2_X1 U7326 ( .A1(n8357), .A2(n6733), .ZN(n8087) );
  NAND2_X2 U7327 ( .A1(n8086), .A2(n8087), .ZN(n8082) );
  NAND2_X1 U7328 ( .A1(n5802), .A2(n8082), .ZN(n8724) );
  OR2_X1 U7329 ( .A1(n8357), .A2(n9948), .ZN(n5803) );
  NAND2_X1 U7330 ( .A1(n6095), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5807) );
  OR2_X1 U7331 ( .A1(n4344), .A2(n10000), .ZN(n5805) );
  INV_X1 U7332 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6984) );
  NAND2_X1 U7333 ( .A1(n5808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U7334 ( .A(n5809), .B(n5756), .ZN(n6762) );
  INV_X1 U7335 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6551) );
  OR2_X1 U7336 ( .A1(n5824), .A2(n6551), .ZN(n5811) );
  OR2_X1 U7337 ( .A1(n5842), .A2(n6552), .ZN(n5810) );
  OAI211_X1 U7338 ( .C1(n5827), .C2(n6762), .A(n5811), .B(n5810), .ZN(n6986)
         );
  INV_X1 U7339 ( .A(n6986), .ZN(n9954) );
  OR2_X1 U7340 ( .A1(n8719), .A2(n9954), .ZN(n5812) );
  NAND2_X1 U7341 ( .A1(n8719), .A2(n9954), .ZN(n6960) );
  NAND2_X1 U7342 ( .A1(n5885), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7343 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5814) );
  AND2_X1 U7344 ( .A1(n5830), .A2(n5814), .ZN(n7104) );
  OR2_X1 U7345 ( .A1(n5790), .A2(n7104), .ZN(n5818) );
  INV_X1 U7346 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5815) );
  OR2_X1 U7347 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  INV_X1 U7348 ( .A(n5839), .ZN(n5823) );
  NAND2_X1 U7349 ( .A1(n5820), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5821) );
  MUX2_X1 U7350 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5821), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5822) );
  OR2_X1 U7351 ( .A1(n5824), .A2(n4977), .ZN(n5826) );
  OR2_X1 U7352 ( .A1(n5842), .A2(n6554), .ZN(n5825) );
  OAI211_X1 U7353 ( .C1(n5827), .C2(n6799), .A(n5826), .B(n5825), .ZN(n8100)
         );
  INV_X1 U7354 ( .A(n8100), .ZN(n7105) );
  AND2_X1 U7355 ( .A1(n6960), .A2(n4967), .ZN(n7091) );
  INV_X1 U7356 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6794) );
  NAND2_X1 U7357 ( .A1(n5830), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5831) );
  AND2_X1 U7358 ( .A1(n5850), .A2(n5831), .ZN(n7100) );
  OR2_X1 U7359 ( .A1(n5790), .A2(n7100), .ZN(n5835) );
  INV_X1 U7360 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6793) );
  OR2_X1 U7361 ( .A1(n4344), .A2(n6793), .ZN(n5834) );
  NAND2_X1 U7362 ( .A1(n6095), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5833) );
  NOR2_X1 U7363 ( .A1(n5839), .A2(n4603), .ZN(n5837) );
  MUX2_X1 U7364 ( .A(n4603), .B(n5837), .S(P2_IR_REG_5__SCAN_IN), .Z(n5841) );
  NAND2_X1 U7365 ( .A1(n5839), .A2(n5838), .ZN(n5858) );
  INV_X1 U7366 ( .A(n5858), .ZN(n5840) );
  OR2_X1 U7367 ( .A1(n5842), .A2(n6544), .ZN(n5844) );
  INV_X1 U7368 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6545) );
  OR2_X1 U7369 ( .A1(n5824), .A2(n6545), .ZN(n5843) );
  OAI211_X1 U7370 ( .C1(n5827), .C2(n6869), .A(n5844), .B(n5843), .ZN(n6914)
         );
  OR2_X1 U7371 ( .A1(n9932), .A2(n6914), .ZN(n7088) );
  AND2_X1 U7372 ( .A1(n7091), .A2(n7088), .ZN(n5845) );
  INV_X1 U7373 ( .A(n7088), .ZN(n5846) );
  OR2_X1 U7374 ( .A1(n6312), .A2(n7105), .ZN(n7093) );
  OR2_X1 U7375 ( .A1(n5846), .A2(n7093), .ZN(n5847) );
  NAND2_X1 U7376 ( .A1(n9932), .A2(n6914), .ZN(n7087) );
  NAND2_X1 U7377 ( .A1(n5848), .A2(n7087), .ZN(n9927) );
  NAND2_X1 U7378 ( .A1(n6095), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5856) );
  INV_X1 U7379 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5849) );
  OR2_X1 U7380 ( .A1(n4344), .A2(n5849), .ZN(n5855) );
  NAND2_X1 U7381 ( .A1(n5850), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5851) );
  AND2_X1 U7382 ( .A1(n5867), .A2(n5851), .ZN(n9937) );
  OR2_X1 U7383 ( .A1(n6028), .A2(n9937), .ZN(n5854) );
  INV_X1 U7384 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5852) );
  OR2_X1 U7385 ( .A1(n5816), .A2(n5852), .ZN(n5853) );
  NAND2_X1 U7386 ( .A1(n5858), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5857) );
  MUX2_X1 U7387 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5857), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5859) );
  OR2_X1 U7388 ( .A1(n5842), .A2(n6542), .ZN(n5861) );
  INV_X1 U7389 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6543) );
  OR2_X1 U7390 ( .A1(n5824), .A2(n6543), .ZN(n5860) );
  OAI211_X1 U7391 ( .C1(n5827), .C2(n7043), .A(n5861), .B(n5860), .ZN(n9967)
         );
  INV_X1 U7392 ( .A(n9967), .ZN(n9938) );
  NAND2_X1 U7393 ( .A1(n9924), .A2(n9938), .ZN(n5862) );
  OR2_X1 U7394 ( .A1(n9924), .A2(n9938), .ZN(n5863) );
  NAND2_X1 U7395 ( .A1(n6095), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5873) );
  INV_X1 U7396 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5864) );
  OR2_X1 U7397 ( .A1(n4344), .A2(n5864), .ZN(n5872) );
  NAND2_X1 U7398 ( .A1(n5867), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5868) );
  AND2_X1 U7399 ( .A1(n5888), .A2(n5868), .ZN(n7214) );
  OR2_X1 U7400 ( .A1(n6028), .A2(n7214), .ZN(n5871) );
  INV_X1 U7401 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5869) );
  OR2_X1 U7402 ( .A1(n5816), .A2(n5869), .ZN(n5870) );
  NAND4_X1 U7403 ( .A1(n5873), .A2(n5872), .A3(n5871), .A4(n5870), .ZN(n9931)
         );
  NAND2_X1 U7404 ( .A1(n5880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5875) );
  XNOR2_X1 U7405 ( .A(n5875), .B(n5874), .ZN(n7116) );
  OR2_X1 U7406 ( .A1(n6547), .A2(n5842), .ZN(n5877) );
  INV_X1 U7407 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6548) );
  OR2_X1 U7408 ( .A1(n5824), .A2(n6548), .ZN(n5876) );
  OAI211_X1 U7409 ( .C1(n5827), .C2(n7116), .A(n5877), .B(n5876), .ZN(n7216)
         );
  OR2_X1 U7410 ( .A1(n9931), .A2(n7216), .ZN(n5878) );
  NAND2_X1 U7411 ( .A1(n6555), .A2(n8025), .ZN(n5884) );
  OAI21_X1 U7412 ( .B1(n5880), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5882) );
  INV_X1 U7413 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U7414 ( .A(n5882), .B(n5881), .ZN(n7299) );
  INV_X1 U7415 ( .A(n7299), .ZN(n7131) );
  AOI22_X1 U7416 ( .A1(n6039), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6535), .B2(
        n7131), .ZN(n5883) );
  INV_X2 U7417 ( .A(n5832), .ZN(n5885) );
  NAND2_X1 U7418 ( .A1(n5885), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5893) );
  INV_X1 U7419 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5887) );
  OR2_X1 U7420 ( .A1(n5886), .A2(n5887), .ZN(n5892) );
  NAND2_X1 U7421 ( .A1(n5888), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5889) );
  AND2_X1 U7422 ( .A1(n5905), .A2(n5889), .ZN(n7309) );
  OR2_X1 U7423 ( .A1(n6028), .A2(n7309), .ZN(n5891) );
  INV_X1 U7424 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7310) );
  OR2_X1 U7425 ( .A1(n5816), .A2(n7310), .ZN(n5890) );
  NAND4_X1 U7426 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n8353)
         );
  INV_X1 U7427 ( .A(n8353), .ZN(n7136) );
  AND2_X1 U7428 ( .A1(n7244), .A2(n7136), .ZN(n5895) );
  OR2_X1 U7429 ( .A1(n7136), .A2(n7244), .ZN(n5894) );
  NAND2_X1 U7430 ( .A1(n6564), .A2(n8025), .ZN(n5901) );
  NOR2_X1 U7431 ( .A1(n5896), .A2(n4603), .ZN(n5897) );
  MUX2_X1 U7432 ( .A(n4603), .B(n5897), .S(P2_IR_REG_9__SCAN_IN), .Z(n5899) );
  OR2_X1 U7433 ( .A1(n5899), .A2(n5898), .ZN(n7373) );
  AOI22_X1 U7434 ( .A1(n6039), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6535), .B2(
        n7374), .ZN(n5900) );
  NAND2_X1 U7435 ( .A1(n6095), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5911) );
  INV_X1 U7436 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5902) );
  OR2_X1 U7437 ( .A1(n4344), .A2(n5902), .ZN(n5910) );
  NAND2_X1 U7438 ( .A1(n5905), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5906) );
  AND2_X1 U7439 ( .A1(n5916), .A2(n5906), .ZN(n7270) );
  OR2_X1 U7440 ( .A1(n6028), .A2(n7270), .ZN(n5909) );
  INV_X1 U7441 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5907) );
  AND2_X1 U7442 ( .A1(n9980), .A2(n8352), .ZN(n5912) );
  OR2_X1 U7443 ( .A1(n6566), .A2(n5842), .ZN(n5915) );
  OR2_X1 U7444 ( .A1(n5898), .A2(n4603), .ZN(n5913) );
  XNOR2_X1 U7445 ( .A(n5913), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7447) );
  AOI22_X1 U7446 ( .A1(n6039), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6535), .B2(
        n7447), .ZN(n5914) );
  NAND2_X1 U7447 ( .A1(n6095), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5921) );
  INV_X1 U7448 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7361) );
  OR2_X1 U7449 ( .A1(n4344), .A2(n7361), .ZN(n5920) );
  NAND2_X1 U7450 ( .A1(n5916), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5917) );
  AND2_X1 U7451 ( .A1(n5928), .A2(n5917), .ZN(n7458) );
  OR2_X1 U7452 ( .A1(n6028), .A2(n7458), .ZN(n5919) );
  INV_X1 U7453 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7459) );
  OR2_X1 U7454 ( .A1(n5816), .A2(n7459), .ZN(n5918) );
  NAND4_X1 U7455 ( .A1(n5921), .A2(n5920), .A3(n5919), .A4(n5918), .ZN(n8351)
         );
  NOR2_X1 U7456 ( .A1(n9986), .A2(n8351), .ZN(n5923) );
  NAND2_X1 U7457 ( .A1(n9986), .A2(n8351), .ZN(n5922) );
  NAND2_X1 U7458 ( .A1(n6577), .A2(n8025), .ZN(n5926) );
  NAND2_X1 U7459 ( .A1(n5937), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5924) );
  XNOR2_X1 U7460 ( .A(n5924), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7386) );
  AOI22_X1 U7461 ( .A1(n6039), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6535), .B2(
        n7386), .ZN(n5925) );
  NAND2_X1 U7462 ( .A1(n5926), .A2(n5925), .ZN(n7342) );
  NAND2_X1 U7463 ( .A1(n6095), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5934) );
  INV_X1 U7464 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5927) );
  OR2_X1 U7465 ( .A1(n4344), .A2(n5927), .ZN(n5933) );
  NAND2_X1 U7466 ( .A1(n5928), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5929) );
  AND2_X1 U7467 ( .A1(n5942), .A2(n5929), .ZN(n7404) );
  OR2_X1 U7468 ( .A1(n6028), .A2(n7404), .ZN(n5932) );
  INV_X1 U7469 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5930) );
  OR2_X1 U7470 ( .A1(n5816), .A2(n5930), .ZN(n5931) );
  OR2_X1 U7471 ( .A1(n7342), .A2(n7510), .ZN(n8126) );
  NAND2_X1 U7472 ( .A1(n7342), .A2(n7510), .ZN(n8128) );
  NAND2_X1 U7473 ( .A1(n8126), .A2(n8128), .ZN(n7337) );
  NAND2_X1 U7474 ( .A1(n7336), .A2(n7337), .ZN(n5936) );
  INV_X1 U7475 ( .A(n7510), .ZN(n8350) );
  NAND2_X1 U7476 ( .A1(n7342), .A2(n8350), .ZN(n5935) );
  OR2_X1 U7477 ( .A1(n6592), .A2(n5842), .ZN(n5940) );
  NAND2_X1 U7478 ( .A1(n5949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5938) );
  XNOR2_X1 U7479 ( .A(n5938), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8377) );
  AOI22_X1 U7480 ( .A1(n6039), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6535), .B2(
        n8377), .ZN(n5939) );
  NAND2_X1 U7481 ( .A1(n6095), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5947) );
  INV_X1 U7482 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8376) );
  OR2_X1 U7483 ( .A1(n4344), .A2(n8376), .ZN(n5946) );
  INV_X1 U7484 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7485 ( .A1(n5942), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5943) );
  AND2_X1 U7486 ( .A1(n5955), .A2(n5943), .ZN(n7507) );
  OR2_X1 U7487 ( .A1(n6028), .A2(n7507), .ZN(n5945) );
  INV_X1 U7488 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8367) );
  OR2_X1 U7489 ( .A1(n5816), .A2(n8367), .ZN(n5944) );
  NAND4_X1 U7490 ( .A1(n5947), .A2(n5946), .A3(n5945), .A4(n5944), .ZN(n8349)
         );
  AND2_X1 U7491 ( .A1(n7547), .A2(n8349), .ZN(n5948) );
  OR2_X1 U7492 ( .A1(n6613), .A2(n5842), .ZN(n5952) );
  OR2_X1 U7493 ( .A1(n6024), .A2(n4603), .ZN(n5950) );
  XNOR2_X1 U7494 ( .A(n5950), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8387) );
  AOI22_X1 U7495 ( .A1(n6039), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6535), .B2(
        n8387), .ZN(n5951) );
  INV_X1 U7496 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7600) );
  OR2_X1 U7497 ( .A1(n5886), .A2(n7600), .ZN(n5960) );
  INV_X1 U7498 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8382) );
  OR2_X1 U7499 ( .A1(n4344), .A2(n8382), .ZN(n5959) );
  INV_X1 U7500 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7501 ( .A1(n5955), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5956) );
  AND2_X1 U7502 ( .A1(n5964), .A2(n5956), .ZN(n7607) );
  OR2_X1 U7503 ( .A1(n6028), .A2(n7607), .ZN(n5958) );
  INV_X1 U7504 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8362) );
  OR2_X1 U7505 ( .A1(n5816), .A2(n8362), .ZN(n5957) );
  NAND2_X1 U7506 ( .A1(n7606), .A2(n8348), .ZN(n7595) );
  NAND2_X1 U7507 ( .A1(n7598), .A2(n7595), .ZN(n5961) );
  NAND2_X1 U7508 ( .A1(n5961), .A2(n7596), .ZN(n7618) );
  NAND2_X1 U7509 ( .A1(n6680), .A2(n8025), .ZN(n5963) );
  NAND2_X1 U7510 ( .A1(n6024), .A2(n6021), .ZN(n6013) );
  NAND2_X1 U7511 ( .A1(n6013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U7512 ( .A(n5988), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8413) );
  AOI22_X1 U7513 ( .A1(n6039), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6535), .B2(
        n8413), .ZN(n5962) );
  INV_X1 U7514 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8853) );
  OR2_X1 U7515 ( .A1(n5886), .A2(n8853), .ZN(n5969) );
  INV_X1 U7516 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8395) );
  OR2_X1 U7517 ( .A1(n4344), .A2(n8395), .ZN(n5968) );
  NAND2_X1 U7518 ( .A1(n5964), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5965) );
  AND2_X1 U7519 ( .A1(n5977), .A2(n5965), .ZN(n8708) );
  OR2_X1 U7520 ( .A1(n6028), .A2(n8708), .ZN(n5967) );
  INV_X1 U7521 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8407) );
  OR2_X1 U7522 ( .A1(n5816), .A2(n8407), .ZN(n5966) );
  NAND4_X1 U7523 ( .A1(n5969), .A2(n5968), .A3(n5967), .A4(n5966), .ZN(n8347)
         );
  NAND2_X1 U7524 ( .A1(n8855), .A2(n8347), .ZN(n5970) );
  NAND2_X1 U7525 ( .A1(n7618), .A2(n5970), .ZN(n5972) );
  OR2_X1 U7526 ( .A1(n8855), .A2(n8347), .ZN(n5971) );
  NAND2_X1 U7527 ( .A1(n6775), .A2(n8025), .ZN(n5976) );
  INV_X1 U7528 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7529 ( .A1(n5988), .A2(n5986), .ZN(n5973) );
  NAND2_X1 U7530 ( .A1(n5973), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5974) );
  XNOR2_X1 U7531 ( .A(n5974), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8455) );
  AOI22_X1 U7532 ( .A1(n6039), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6535), .B2(
        n8455), .ZN(n5975) );
  NAND2_X1 U7533 ( .A1(n6095), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5982) );
  INV_X1 U7534 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8418) );
  OR2_X1 U7535 ( .A1(n5832), .A2(n8418), .ZN(n5981) );
  NAND2_X1 U7536 ( .A1(n5977), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5978) );
  AND2_X1 U7537 ( .A1(n5993), .A2(n5978), .ZN(n8332) );
  OR2_X1 U7538 ( .A1(n6028), .A2(n8332), .ZN(n5980) );
  INV_X1 U7539 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8419) );
  OR2_X1 U7540 ( .A1(n5828), .A2(n8419), .ZN(n5979) );
  NAND4_X1 U7541 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n8699)
         );
  NOR2_X1 U7542 ( .A1(n8326), .A2(n8699), .ZN(n5984) );
  NAND2_X1 U7543 ( .A1(n8326), .A2(n8699), .ZN(n5983) );
  NAND2_X1 U7544 ( .A1(n6855), .A2(n8025), .ZN(n5992) );
  INV_X1 U7545 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7546 ( .A1(n5986), .A2(n5985), .ZN(n6014) );
  NAND2_X1 U7547 ( .A1(n6014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7548 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  OR2_X1 U7549 ( .A1(n5989), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7550 ( .A1(n5989), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5990) );
  AOI22_X1 U7551 ( .A1(n6039), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6535), .B2(
        n8450), .ZN(n5991) );
  NAND2_X1 U7552 ( .A1(n6095), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5998) );
  INV_X1 U7553 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8779) );
  OR2_X1 U7554 ( .A1(n4344), .A2(n8779), .ZN(n5997) );
  NAND2_X1 U7555 ( .A1(n5993), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5994) );
  AND2_X1 U7556 ( .A1(n6005), .A2(n5994), .ZN(n8703) );
  OR2_X1 U7557 ( .A1(n6028), .A2(n8703), .ZN(n5996) );
  INV_X1 U7558 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8702) );
  OR2_X1 U7559 ( .A1(n5828), .A2(n8702), .ZN(n5995) );
  NAND4_X1 U7560 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n8686)
         );
  INV_X1 U7561 ( .A(n8686), .ZN(n8334) );
  NAND2_X1 U7562 ( .A1(n8848), .A2(n8334), .ZN(n8148) );
  NAND2_X1 U7563 ( .A1(n8153), .A2(n8148), .ZN(n8697) );
  NAND2_X1 U7564 ( .A1(n6940), .A2(n8025), .ZN(n6002) );
  NAND2_X1 U7565 ( .A1(n5999), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6000) );
  XNOR2_X1 U7566 ( .A(n6000), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8501) );
  AOI22_X1 U7567 ( .A1(n6039), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6535), .B2(
        n8501), .ZN(n6001) );
  INV_X1 U7568 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7569 ( .A1(n6005), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6006) );
  AND2_X1 U7570 ( .A1(n6029), .A2(n6006), .ZN(n8690) );
  OR2_X1 U7571 ( .A1(n6028), .A2(n8690), .ZN(n6010) );
  INV_X1 U7572 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10071) );
  OR2_X1 U7573 ( .A1(n5832), .A2(n10071), .ZN(n6009) );
  INV_X1 U7574 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8689) );
  OR2_X1 U7575 ( .A1(n5828), .A2(n8689), .ZN(n6008) );
  INV_X1 U7576 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8841) );
  OR2_X1 U7577 ( .A1(n5886), .A2(n8841), .ZN(n6007) );
  NAND4_X1 U7578 ( .A1(n6010), .A2(n6009), .A3(n6008), .A4(n6007), .ZN(n8700)
         );
  INV_X1 U7579 ( .A(n8700), .ZN(n8321) );
  NAND2_X1 U7580 ( .A1(n8842), .A2(n8321), .ZN(n8677) );
  NAND2_X1 U7581 ( .A1(n8165), .A2(n8677), .ZN(n8150) );
  NAND2_X1 U7582 ( .A1(n8685), .A2(n8150), .ZN(n6012) );
  NAND2_X1 U7583 ( .A1(n8842), .A2(n8700), .ZN(n6011) );
  NAND2_X1 U7584 ( .A1(n7012), .A2(n8025), .ZN(n6027) );
  INV_X1 U7585 ( .A(n6013), .ZN(n6017) );
  INV_X1 U7586 ( .A(n6014), .ZN(n6015) );
  AND2_X1 U7587 ( .A1(n6016), .A2(n6015), .ZN(n6019) );
  NAND2_X1 U7588 ( .A1(n4431), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6018) );
  MUX2_X1 U7589 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6018), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n6025) );
  INV_X1 U7590 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7591 ( .A1(n6025), .A2(n6150), .ZN(n8511) );
  INV_X1 U7592 ( .A(n8511), .ZN(n8528) );
  AOI22_X1 U7593 ( .A1(n6039), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6535), .B2(
        n8528), .ZN(n6026) );
  NAND2_X1 U7594 ( .A1(n6029), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7595 ( .A1(n6044), .A2(n6030), .ZN(n8669) );
  NAND2_X1 U7596 ( .A1(n6046), .A2(n8669), .ZN(n6036) );
  INV_X1 U7597 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6031) );
  OR2_X1 U7598 ( .A1(n5886), .A2(n6031), .ZN(n6035) );
  INV_X1 U7599 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7600 ( .A1(n4344), .A2(n6032), .ZN(n6034) );
  INV_X1 U7601 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8671) );
  OR2_X1 U7602 ( .A1(n5828), .A2(n8671), .ZN(n6033) );
  INV_X1 U7603 ( .A(n8658), .ZN(n8687) );
  AND2_X1 U7604 ( .A1(n8673), .A2(n8687), .ZN(n8650) );
  NAND2_X1 U7605 ( .A1(n7159), .A2(n8025), .ZN(n6041) );
  NAND2_X1 U7606 ( .A1(n6150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6038) );
  AOI22_X1 U7607 ( .A1(n6039), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6535), .B2(
        n8062), .ZN(n6040) );
  INV_X1 U7608 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8768) );
  OR2_X1 U7609 ( .A1(n5832), .A2(n8768), .ZN(n6043) );
  INV_X1 U7610 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8663) );
  OR2_X1 U7611 ( .A1(n5828), .A2(n8663), .ZN(n6042) );
  AND2_X1 U7612 ( .A1(n6043), .A2(n6042), .ZN(n6049) );
  NAND2_X1 U7613 ( .A1(n6044), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7614 ( .A1(n6052), .A2(n6045), .ZN(n8664) );
  NAND2_X1 U7615 ( .A1(n8664), .A2(n6046), .ZN(n6048) );
  NAND2_X1 U7616 ( .A1(n6095), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6047) );
  INV_X1 U7617 ( .A(n8636), .ZN(n8667) );
  AND2_X1 U7618 ( .A1(n8769), .A2(n8667), .ZN(n6058) );
  OR2_X1 U7619 ( .A1(n8650), .A2(n6058), .ZN(n8631) );
  NAND2_X1 U7620 ( .A1(n7188), .A2(n8025), .ZN(n6051) );
  INV_X1 U7621 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7203) );
  OR2_X1 U7622 ( .A1(n5824), .A2(n7203), .ZN(n6050) );
  NAND2_X1 U7623 ( .A1(n6052), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7624 ( .A1(n6062), .A2(n6053), .ZN(n8643) );
  NAND2_X1 U7625 ( .A1(n8643), .A2(n6046), .ZN(n6056) );
  AOI22_X1 U7626 ( .A1(n6095), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n5885), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7627 ( .A1(n6160), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7628 ( .A1(n8831), .A2(n8659), .ZN(n8173) );
  NAND2_X1 U7629 ( .A1(n8769), .A2(n8636), .ZN(n8170) );
  INV_X1 U7630 ( .A(n8654), .ZN(n6057) );
  OR2_X1 U7631 ( .A1(n8673), .A2(n8687), .ZN(n8652) );
  AND2_X1 U7632 ( .A1(n6057), .A2(n8652), .ZN(n8651) );
  OR2_X1 U7633 ( .A1(n6058), .A2(n8651), .ZN(n8632) );
  INV_X1 U7634 ( .A(n8659), .ZN(n8624) );
  NAND2_X1 U7635 ( .A1(n7204), .A2(n8025), .ZN(n6060) );
  OR2_X1 U7636 ( .A1(n5824), .A2(n7235), .ZN(n6059) );
  INV_X1 U7637 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U7638 ( .A1(n6062), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7639 ( .A1(n6071), .A2(n6063), .ZN(n8627) );
  NAND2_X1 U7640 ( .A1(n8627), .A2(n6046), .ZN(n6066) );
  AOI22_X1 U7641 ( .A1(n6095), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n5885), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7642 ( .A1(n6160), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7643 ( .A1(n8825), .A2(n8637), .ZN(n8179) );
  NAND2_X1 U7644 ( .A1(n8178), .A2(n8179), .ZN(n8621) );
  NAND2_X1 U7645 ( .A1(n8622), .A2(n8621), .ZN(n6068) );
  INV_X1 U7646 ( .A(n8637), .ZN(n8346) );
  OR2_X1 U7647 ( .A1(n8825), .A2(n8346), .ZN(n6067) );
  NAND2_X1 U7648 ( .A1(n6068), .A2(n6067), .ZN(n8611) );
  NAND2_X1 U7649 ( .A1(n7317), .A2(n8025), .ZN(n6070) );
  OR2_X1 U7650 ( .A1(n5824), .A2(n10086), .ZN(n6069) );
  NAND2_X1 U7651 ( .A1(n6071), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7652 ( .A1(n6081), .A2(n6072), .ZN(n8615) );
  INV_X1 U7653 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U7654 ( .A1(n6160), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7655 ( .A1(n5885), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6073) );
  OAI211_X1 U7656 ( .C1(n5886), .C2(n8820), .A(n6074), .B(n6073), .ZN(n6075)
         );
  AOI21_X1 U7657 ( .B1(n8615), .B2(n6046), .A(n6075), .ZN(n8263) );
  OR2_X1 U7658 ( .A1(n8756), .A2(n8263), .ZN(n8065) );
  NAND2_X1 U7659 ( .A1(n8756), .A2(n8263), .ZN(n8064) );
  NAND2_X1 U7660 ( .A1(n8065), .A2(n8064), .ZN(n8177) );
  NAND2_X1 U7661 ( .A1(n8611), .A2(n8177), .ZN(n6077) );
  INV_X1 U7662 ( .A(n8263), .ZN(n8623) );
  OR2_X1 U7663 ( .A1(n8756), .A2(n8623), .ZN(n6076) );
  NAND2_X1 U7664 ( .A1(n6077), .A2(n6076), .ZN(n8604) );
  NAND2_X1 U7665 ( .A1(n6078), .A2(n8025), .ZN(n6080) );
  OR2_X1 U7666 ( .A1(n5824), .A2(n7413), .ZN(n6079) );
  NAND2_X1 U7667 ( .A1(n6081), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7668 ( .A1(n6093), .A2(n6082), .ZN(n8608) );
  NAND2_X1 U7669 ( .A1(n8608), .A2(n6046), .ZN(n6087) );
  INV_X1 U7670 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U7671 ( .A1(n5885), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7672 ( .A1(n6160), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6083) );
  OAI211_X1 U7673 ( .C1(n8814), .C2(n5886), .A(n6084), .B(n6083), .ZN(n6085)
         );
  INV_X1 U7674 ( .A(n6085), .ZN(n6086) );
  NOR2_X1 U7675 ( .A1(n8815), .A2(n8591), .ZN(n6088) );
  NAND2_X1 U7676 ( .A1(n8815), .A2(n8591), .ZN(n6089) );
  NAND2_X1 U7677 ( .A1(n7563), .A2(n8025), .ZN(n6091) );
  OR2_X1 U7678 ( .A1(n5824), .A2(n10055), .ZN(n6090) );
  INV_X1 U7679 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7680 ( .A1(n6093), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7681 ( .A1(n6106), .A2(n6094), .ZN(n8593) );
  NAND2_X1 U7682 ( .A1(n8593), .A2(n6046), .ZN(n6100) );
  INV_X1 U7683 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U7684 ( .A1(n5885), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7685 ( .A1(n6095), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6096) );
  OAI211_X1 U7686 ( .C1(n5828), .C2(n8599), .A(n6097), .B(n6096), .ZN(n6098)
         );
  INV_X1 U7687 ( .A(n6098), .ZN(n6099) );
  AND2_X1 U7688 ( .A1(n8809), .A2(n8605), .ZN(n6101) );
  NAND2_X1 U7689 ( .A1(n7575), .A2(n8025), .ZN(n6103) );
  OR2_X1 U7690 ( .A1(n5824), .A2(n7594), .ZN(n6102) );
  INV_X1 U7691 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7692 ( .A1(n6106), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7693 ( .A1(n6117), .A2(n6107), .ZN(n8583) );
  NAND2_X1 U7694 ( .A1(n8583), .A2(n6046), .ZN(n6112) );
  INV_X1 U7695 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10193) );
  NAND2_X1 U7696 ( .A1(n6160), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7697 ( .A1(n5885), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6108) );
  OAI211_X1 U7698 ( .C1(n5886), .C2(n10193), .A(n6109), .B(n6108), .ZN(n6110)
         );
  INV_X1 U7699 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7700 ( .A1(n8803), .A2(n8285), .ZN(n8194) );
  NAND2_X1 U7701 ( .A1(n6232), .A2(n8194), .ZN(n8585) );
  OR2_X1 U7702 ( .A1(n8803), .A2(n8590), .ZN(n6113) );
  NAND2_X1 U7703 ( .A1(n6114), .A2(n6113), .ZN(n8570) );
  INV_X1 U7704 ( .A(n8570), .ZN(n6122) );
  NAND2_X1 U7705 ( .A1(n7614), .A2(n8025), .ZN(n6116) );
  OR2_X1 U7706 ( .A1(n5824), .A2(n10218), .ZN(n6115) );
  NAND2_X1 U7707 ( .A1(n6117), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6118) );
  INV_X1 U7708 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U7709 ( .A1(n6160), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7710 ( .A1(n5885), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6119) );
  OAI211_X1 U7711 ( .C1(n5886), .C2(n8797), .A(n6120), .B(n6119), .ZN(n6121)
         );
  NAND2_X1 U7712 ( .A1(n7624), .A2(n8025), .ZN(n6124) );
  OR2_X1 U7713 ( .A1(n5824), .A2(n8018), .ZN(n6123) );
  INV_X1 U7714 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7715 ( .A1(n4571), .A2(n6125), .ZN(n6139) );
  NAND2_X1 U7716 ( .A1(n6126), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7717 ( .A1(n6139), .A2(n6127), .ZN(n8562) );
  NAND2_X1 U7718 ( .A1(n8562), .A2(n6046), .ZN(n6132) );
  INV_X1 U7719 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U7720 ( .A1(n5885), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7721 ( .A1(n6160), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6128) );
  OAI211_X1 U7722 ( .C1(n8793), .C2(n5886), .A(n6129), .B(n6128), .ZN(n6130)
         );
  INV_X1 U7723 ( .A(n6130), .ZN(n6131) );
  NAND2_X1 U7724 ( .A1(n8738), .A2(n7713), .ZN(n8204) );
  NAND2_X1 U7725 ( .A1(n8203), .A2(n8204), .ZN(n8560) );
  NAND2_X1 U7726 ( .A1(n8554), .A2(n8560), .ZN(n6149) );
  OR2_X1 U7727 ( .A1(n8738), .A2(n8571), .ZN(n6147) );
  NAND2_X1 U7728 ( .A1(n6149), .A2(n6147), .ZN(n6146) );
  NAND2_X1 U7729 ( .A1(n6134), .A2(n6133), .ZN(n6136) );
  NAND2_X1 U7730 ( .A1(n6136), .A2(n6135), .ZN(n6257) );
  MUX2_X1 U7731 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7795), .Z(n6258) );
  INV_X1 U7732 ( .A(SI_28_), .ZN(n10056) );
  XNOR2_X1 U7733 ( .A(n6258), .B(n10056), .ZN(n6256) );
  NAND2_X1 U7734 ( .A1(n8020), .A2(n8025), .ZN(n6138) );
  INV_X1 U7735 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7652) );
  OR2_X1 U7736 ( .A1(n5824), .A2(n7652), .ZN(n6137) );
  NAND2_X1 U7737 ( .A1(n6139), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7738 ( .A1(n7678), .A2(n6140), .ZN(n8546) );
  NAND2_X1 U7739 ( .A1(n8546), .A2(n6046), .ZN(n6145) );
  INV_X1 U7740 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7741 ( .A1(n6160), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7742 ( .A1(n5885), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6141) );
  OAI211_X1 U7743 ( .C1(n5886), .C2(n6212), .A(n6142), .B(n6141), .ZN(n6143)
         );
  INV_X1 U7744 ( .A(n6143), .ZN(n6144) );
  XNOR2_X1 U7745 ( .A(n8547), .B(n6266), .ZN(n6234) );
  INV_X1 U7746 ( .A(n6234), .ZN(n8055) );
  NAND2_X1 U7747 ( .A1(n6146), .A2(n8055), .ZN(n6169) );
  AND2_X1 U7748 ( .A1(n6234), .A2(n6147), .ZN(n6148) );
  NAND2_X1 U7749 ( .A1(n6149), .A2(n6148), .ZN(n6265) );
  INV_X1 U7750 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7751 ( .A1(n4401), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6153) );
  INV_X1 U7752 ( .A(n7201), .ZN(n8224) );
  NAND2_X1 U7753 ( .A1(n6296), .A2(n8224), .ZN(n6156) );
  NAND2_X1 U7754 ( .A1(n4355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7755 ( .A1(n8062), .A2(n8229), .ZN(n6206) );
  NAND2_X2 U7756 ( .A1(n6156), .A2(n6206), .ZN(n9928) );
  INV_X1 U7757 ( .A(n7678), .ZN(n6159) );
  NAND2_X1 U7758 ( .A1(n6159), .A2(n6046), .ZN(n7675) );
  INV_X1 U7759 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7760 ( .A1(n6160), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7761 ( .A1(n5885), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6161) );
  OAI211_X1 U7762 ( .C1(n5886), .C2(n6288), .A(n6162), .B(n6161), .ZN(n6163)
         );
  INV_X1 U7763 ( .A(n6163), .ZN(n6164) );
  NAND2_X1 U7764 ( .A1(n7675), .A2(n6164), .ZN(n8345) );
  INV_X1 U7765 ( .A(n6165), .ZN(n8226) );
  XNOR2_X1 U7766 ( .A(n8226), .B(n8530), .ZN(n6390) );
  INV_X1 U7767 ( .A(n6390), .ZN(n6167) );
  AOI22_X1 U7768 ( .A1(n8345), .A2(n9930), .B1(n9933), .B2(n8571), .ZN(n6168)
         );
  NAND2_X1 U7769 ( .A1(n8547), .A2(n9987), .ZN(n6170) );
  INV_X1 U7770 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7771 ( .A1(n6205), .A2(n6204), .ZN(n6172) );
  AND2_X1 U7772 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6171) );
  NAND2_X1 U7773 ( .A1(n6172), .A2(n6171), .ZN(n6176) );
  INV_X1 U7774 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6173) );
  AND2_X1 U7775 ( .A1(n6204), .A2(n6173), .ZN(n6175) );
  NOR2_X1 U7776 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6174) );
  AOI21_X1 U7777 ( .B1(n6205), .B2(n6175), .A(n6174), .ZN(n6177) );
  NAND2_X1 U7778 ( .A1(n6176), .A2(n6177), .ZN(n6186) );
  XNOR2_X1 U7779 ( .A(n6186), .B(P2_B_REG_SCAN_IN), .ZN(n6180) );
  INV_X1 U7780 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7781 ( .A1(n6180), .A2(n6189), .ZN(n6185) );
  NAND2_X1 U7782 ( .A1(n6181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6182) );
  MUX2_X1 U7783 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6182), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6184) );
  NAND2_X1 U7784 ( .A1(n6185), .A2(n6187), .ZN(n6188) );
  NAND2_X1 U7785 ( .A1(n6186), .A2(n7622), .ZN(n6583) );
  OR2_X1 U7786 ( .A1(n6188), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7787 ( .A1(n6189), .A2(n7622), .ZN(n6580) );
  NAND2_X1 U7788 ( .A1(n6295), .A2(n6244), .ZN(n6239) );
  NOR2_X1 U7789 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .ZN(
        n6194) );
  NOR4_X1 U7790 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6193) );
  NOR4_X1 U7791 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6192) );
  NOR4_X1 U7792 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6191) );
  NAND4_X1 U7793 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(n6200)
         );
  NOR4_X1 U7794 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6198) );
  NOR4_X1 U7795 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6197) );
  NOR4_X1 U7796 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6196) );
  NOR4_X1 U7797 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6195) );
  NAND4_X1 U7798 ( .A1(n6198), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n6199)
         );
  NOR2_X1 U7799 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  NOR2_X1 U7800 ( .A1(n6188), .A2(n6201), .ZN(n6241) );
  NOR2_X1 U7801 ( .A1(n6239), .A2(n6241), .ZN(n6392) );
  INV_X1 U7802 ( .A(n6189), .ZN(n6203) );
  NOR2_X1 U7803 ( .A1(n6186), .A2(n7622), .ZN(n6202) );
  NAND2_X1 U7804 ( .A1(n6203), .A2(n6202), .ZN(n6537) );
  XNOR2_X1 U7805 ( .A(n6205), .B(n6204), .ZN(n6533) );
  NAND2_X1 U7806 ( .A1(n6392), .A2(n6559), .ZN(n6385) );
  INV_X1 U7807 ( .A(n6297), .ZN(n8221) );
  NOR2_X1 U7808 ( .A1(n6206), .A2(n7201), .ZN(n6207) );
  NAND2_X1 U7809 ( .A1(n8072), .A2(n6207), .ZN(n6398) );
  INV_X1 U7810 ( .A(n6398), .ZN(n6377) );
  NOR2_X1 U7811 ( .A1(n6840), .A2(n6377), .ZN(n6208) );
  OR2_X1 U7812 ( .A1(n6385), .A2(n6208), .ZN(n6211) );
  INV_X1 U7813 ( .A(n6244), .ZN(n6833) );
  INV_X1 U7814 ( .A(n6241), .ZN(n6209) );
  NAND3_X1 U7815 ( .A1(n6293), .A2(n6833), .A3(n6209), .ZN(n6403) );
  NOR2_X1 U7816 ( .A1(n6403), .A2(n6401), .ZN(n6388) );
  NAND3_X1 U7817 ( .A1(n6398), .A2(n9989), .A3(n8206), .ZN(n6376) );
  NAND2_X1 U7818 ( .A1(n6376), .A2(n8709), .ZN(n6393) );
  NAND2_X1 U7819 ( .A1(n6388), .A2(n6393), .ZN(n6210) );
  INV_X1 U7820 ( .A(n6213), .ZN(n6216) );
  NAND2_X1 U7821 ( .A1(n4376), .A2(n6214), .ZN(n6305) );
  INV_X1 U7822 ( .A(n6305), .ZN(n6215) );
  NAND2_X1 U7823 ( .A1(n6944), .A2(n8081), .ZN(n8716) );
  NAND2_X1 U7824 ( .A1(n8716), .A2(n8722), .ZN(n6978) );
  NAND2_X1 U7825 ( .A1(n6978), .A2(n8086), .ZN(n6217) );
  NAND2_X1 U7826 ( .A1(n6217), .A2(n8038), .ZN(n6957) );
  NAND2_X1 U7827 ( .A1(n6957), .A2(n8097), .ZN(n6218) );
  NAND2_X1 U7828 ( .A1(n7093), .A2(n4967), .ZN(n8037) );
  NAND2_X1 U7829 ( .A1(n6312), .A2(n8100), .ZN(n8092) );
  INV_X1 U7830 ( .A(n6914), .ZN(n9959) );
  OR2_X1 U7831 ( .A1(n9924), .A2(n9967), .ZN(n8101) );
  NAND2_X1 U7832 ( .A1(n9932), .A2(n9959), .ZN(n9922) );
  NAND2_X1 U7833 ( .A1(n9923), .A2(n8096), .ZN(n6219) );
  NAND2_X1 U7834 ( .A1(n9924), .A2(n9967), .ZN(n8071) );
  INV_X1 U7835 ( .A(n7216), .ZN(n9972) );
  OR2_X1 U7836 ( .A1(n9931), .A2(n9972), .ZN(n8115) );
  NAND2_X1 U7837 ( .A1(n9931), .A2(n9972), .ZN(n7237) );
  NAND2_X1 U7838 ( .A1(n8115), .A2(n7237), .ZN(n8040) );
  NAND2_X1 U7839 ( .A1(n7244), .A2(n8353), .ZN(n8107) );
  AND2_X1 U7840 ( .A1(n8107), .A2(n7237), .ZN(n8114) );
  NOR2_X1 U7841 ( .A1(n7244), .A2(n8353), .ZN(n8117) );
  NAND2_X1 U7842 ( .A1(n9980), .A2(n6220), .ZN(n8118) );
  NAND2_X1 U7843 ( .A1(n7265), .A2(n8045), .ZN(n7450) );
  OR2_X1 U7844 ( .A1(n9986), .A2(n7339), .ZN(n8125) );
  NAND2_X1 U7845 ( .A1(n9986), .A2(n7339), .ZN(n8123) );
  NAND2_X1 U7846 ( .A1(n8125), .A2(n8123), .ZN(n8042) );
  INV_X1 U7847 ( .A(n8042), .ZN(n6221) );
  AND2_X1 U7848 ( .A1(n8113), .A2(n6221), .ZN(n6222) );
  NAND2_X1 U7849 ( .A1(n7450), .A2(n6222), .ZN(n7451) );
  NAND2_X1 U7850 ( .A1(n7451), .A2(n8123), .ZN(n7341) );
  INV_X1 U7851 ( .A(n7337), .ZN(n8046) );
  NAND2_X1 U7852 ( .A1(n7341), .A2(n8046), .ZN(n7340) );
  NAND2_X1 U7853 ( .A1(n7340), .A2(n8128), .ZN(n7535) );
  NAND2_X1 U7854 ( .A1(n7547), .A2(n7569), .ZN(n8132) );
  NAND2_X1 U7855 ( .A1(n8133), .A2(n8132), .ZN(n8136) );
  NOR2_X1 U7856 ( .A1(n7606), .A2(n8238), .ZN(n8139) );
  NAND2_X1 U7857 ( .A1(n7606), .A2(n8238), .ZN(n8138) );
  INV_X1 U7858 ( .A(n8347), .ZN(n6223) );
  OR2_X1 U7859 ( .A1(n8855), .A2(n6223), .ZN(n8143) );
  NAND2_X1 U7860 ( .A1(n8855), .A2(n6223), .ZN(n8144) );
  NAND2_X1 U7861 ( .A1(n6224), .A2(n8144), .ZN(n7695) );
  INV_X1 U7862 ( .A(n8699), .ZN(n6345) );
  OR2_X1 U7863 ( .A1(n8326), .A2(n6345), .ZN(n8147) );
  NAND2_X1 U7864 ( .A1(n7695), .A2(n8147), .ZN(n8695) );
  NAND2_X1 U7865 ( .A1(n8326), .A2(n6345), .ZN(n8694) );
  AND2_X1 U7866 ( .A1(n8148), .A2(n8694), .ZN(n8155) );
  NAND2_X1 U7867 ( .A1(n8695), .A2(n8155), .ZN(n6225) );
  NAND2_X1 U7868 ( .A1(n6225), .A2(n8153), .ZN(n8674) );
  INV_X1 U7869 ( .A(n8165), .ZN(n8675) );
  INV_X1 U7870 ( .A(n8166), .ZN(n6227) );
  NAND2_X1 U7871 ( .A1(n8673), .A2(n8658), .ZN(n8160) );
  NAND2_X1 U7872 ( .A1(n8166), .A2(n8160), .ZN(n8679) );
  INV_X1 U7873 ( .A(n8679), .ZN(n6226) );
  AND2_X1 U7874 ( .A1(n6226), .A2(n8677), .ZN(n8676) );
  INV_X1 U7875 ( .A(n8169), .ZN(n6228) );
  OAI21_X1 U7876 ( .B1(n8642), .B2(n6228), .A(n8173), .ZN(n8620) );
  INV_X1 U7877 ( .A(n8179), .ZN(n6229) );
  OAI21_X1 U7878 ( .B1(n8620), .B2(n6229), .A(n8178), .ZN(n8614) );
  INV_X1 U7879 ( .A(n8065), .ZN(n6230) );
  AOI21_X1 U7880 ( .B1(n8614), .B2(n8064), .A(n6230), .ZN(n8602) );
  NAND2_X1 U7881 ( .A1(n8602), .A2(n8183), .ZN(n8595) );
  NAND2_X1 U7882 ( .A1(n8809), .A2(n8248), .ZN(n8185) );
  NAND2_X1 U7883 ( .A1(n8815), .A2(n6368), .ZN(n8596) );
  AND2_X1 U7884 ( .A1(n8185), .A2(n8596), .ZN(n8187) );
  NAND2_X1 U7885 ( .A1(n8595), .A2(n8187), .ZN(n6231) );
  INV_X1 U7886 ( .A(n6232), .ZN(n8198) );
  NAND2_X1 U7887 ( .A1(n8798), .A2(n8557), .ZN(n8197) );
  NAND2_X1 U7888 ( .A1(n8561), .A2(n8203), .ZN(n6233) );
  NAND2_X1 U7889 ( .A1(n6233), .A2(n8204), .ZN(n6255) );
  XNOR2_X1 U7890 ( .A(n6255), .B(n6234), .ZN(n8550) );
  OAI21_X1 U7891 ( .B1(n8062), .B2(n7318), .A(n6297), .ZN(n6235) );
  NAND2_X1 U7892 ( .A1(n9989), .A2(n6235), .ZN(n6236) );
  INV_X1 U7893 ( .A(n9994), .ZN(n9965) );
  NAND2_X1 U7894 ( .A1(n6238), .A2(n6237), .ZN(P2_U3455) );
  INV_X1 U7895 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6250) );
  INV_X1 U7896 ( .A(n6239), .ZN(n6240) );
  NOR2_X1 U7897 ( .A1(n9982), .A2(n6296), .ZN(n6386) );
  NOR2_X1 U7898 ( .A1(n6240), .A2(n6386), .ZN(n6248) );
  OR2_X1 U7899 ( .A1(n8206), .A2(n8221), .ZN(n6395) );
  NOR2_X1 U7900 ( .A1(n6241), .A2(n6401), .ZN(n6242) );
  NAND3_X1 U7901 ( .A1(n8224), .A2(n8229), .A3(n8539), .ZN(n6243) );
  NAND2_X1 U7902 ( .A1(n8206), .A2(n6243), .ZN(n6245) );
  OR2_X1 U7903 ( .A1(n6293), .A2(n6245), .ZN(n6247) );
  NAND2_X1 U7904 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  NAND2_X1 U7905 ( .A1(n6247), .A2(n6246), .ZN(n6836) );
  MUX2_X1 U7906 ( .A(n6250), .B(n6249), .S(n10008), .Z(n6252) );
  NAND2_X1 U7907 ( .A1(n6252), .A2(n6251), .ZN(P2_U3487) );
  INV_X1 U7908 ( .A(n9982), .ZN(n9949) );
  AND2_X1 U7909 ( .A1(n8547), .A2(n6266), .ZN(n6254) );
  OR2_X1 U7910 ( .A1(n8547), .A2(n6266), .ZN(n6253) );
  NAND2_X1 U7911 ( .A1(n6257), .A2(n6256), .ZN(n6261) );
  INV_X1 U7912 ( .A(n6258), .ZN(n6259) );
  NAND2_X1 U7913 ( .A1(n6259), .A2(n10056), .ZN(n6260) );
  NAND2_X1 U7914 ( .A1(n6261), .A2(n6260), .ZN(n7659) );
  INV_X1 U7915 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7653) );
  INV_X1 U7916 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7655) );
  MUX2_X1 U7917 ( .A(n7653), .B(n7655), .S(n7795), .Z(n7658) );
  NAND2_X1 U7918 ( .A1(n6474), .A2(n8025), .ZN(n6263) );
  OR2_X1 U7919 ( .A1(n5824), .A2(n7653), .ZN(n6262) );
  INV_X1 U7920 ( .A(n8345), .ZN(n6264) );
  NAND2_X1 U7921 ( .A1(n6283), .A2(n6264), .ZN(n8029) );
  INV_X1 U7922 ( .A(n6278), .ZN(n6282) );
  INV_X1 U7923 ( .A(n8547), .ZN(n6267) );
  OAI21_X1 U7924 ( .B1(n6267), .B2(n6266), .A(n6265), .ZN(n6268) );
  XNOR2_X1 U7925 ( .A(n6268), .B(n4406), .ZN(n6269) );
  NAND2_X1 U7926 ( .A1(n6269), .A2(n9928), .ZN(n6281) );
  INV_X1 U7927 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7928 ( .A1(n6095), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6272) );
  INV_X1 U7929 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6270) );
  OR2_X1 U7930 ( .A1(n5828), .A2(n6270), .ZN(n6271) );
  OAI211_X1 U7931 ( .C1(n4344), .C2(n6273), .A(n6272), .B(n6271), .ZN(n6274)
         );
  INV_X1 U7932 ( .A(n6274), .ZN(n6275) );
  NAND2_X1 U7933 ( .A1(n7675), .A2(n6275), .ZN(n8344) );
  AND2_X1 U7934 ( .A1(n5827), .A2(P2_B_REG_SCAN_IN), .ZN(n6276) );
  NOR2_X1 U7935 ( .A1(n8718), .A2(n6276), .ZN(n7676) );
  AOI22_X1 U7936 ( .A1(n9933), .A2(n8555), .B1(n8344), .B2(n7676), .ZN(n6277)
         );
  NAND2_X1 U7937 ( .A1(n10008), .A2(n9987), .ZN(n8737) );
  INV_X1 U7938 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7939 ( .B1(n6292), .B2(n6287), .A(n6286), .ZN(P2_U3488) );
  OR2_X1 U7940 ( .A1(n9995), .A2(n6288), .ZN(n6289) );
  OAI21_X1 U7941 ( .B1(n6292), .B2(n9997), .A(n6291), .ZN(P2_U3456) );
  INV_X1 U7942 ( .A(n6293), .ZN(n6295) );
  NAND2_X1 U7943 ( .A1(n6296), .A2(n7201), .ZN(n6298) );
  XNOR2_X1 U7944 ( .A(n7547), .B(n6375), .ZN(n6337) );
  INV_X1 U7945 ( .A(n6337), .ZN(n6338) );
  NAND2_X1 U7946 ( .A1(n6809), .A2(n6301), .ZN(n6304) );
  NAND2_X1 U7947 ( .A1(n6303), .A2(n6302), .ZN(n6306) );
  AND2_X1 U7948 ( .A1(n6304), .A2(n6306), .ZN(n6684) );
  OAI21_X1 U7949 ( .B1(n6412), .B2(n6214), .A(n6305), .ZN(n6683) );
  NAND2_X1 U7950 ( .A1(n6684), .A2(n6683), .ZN(n6682) );
  NAND2_X1 U7951 ( .A1(n6682), .A2(n6306), .ZN(n6730) );
  XNOR2_X1 U7952 ( .A(n6307), .B(n8357), .ZN(n6731) );
  NAND2_X1 U7953 ( .A1(n6730), .A2(n6731), .ZN(n6729) );
  NAND2_X1 U7954 ( .A1(n6307), .A2(n4615), .ZN(n6308) );
  NAND2_X1 U7955 ( .A1(n6729), .A2(n6308), .ZN(n6822) );
  XNOR2_X1 U7956 ( .A(n6310), .B(n8719), .ZN(n6823) );
  XNOR2_X1 U7957 ( .A(n6412), .B(n8100), .ZN(n6313) );
  NAND2_X1 U7958 ( .A1(n6313), .A2(n6312), .ZN(n6315) );
  INV_X1 U7959 ( .A(n6315), .ZN(n6309) );
  OR2_X1 U7960 ( .A1(n6823), .A2(n6309), .ZN(n6318) );
  INV_X1 U7961 ( .A(n6310), .ZN(n6311) );
  INV_X1 U7962 ( .A(n6312), .ZN(n8355) );
  INV_X1 U7963 ( .A(n6313), .ZN(n6314) );
  NAND2_X1 U7964 ( .A1(n8355), .A2(n6314), .ZN(n6882) );
  NAND3_X1 U7965 ( .A1(n6881), .A2(n6882), .A3(n6315), .ZN(n6883) );
  NAND2_X1 U7966 ( .A1(n6883), .A2(n6315), .ZN(n6316) );
  XNOR2_X1 U7967 ( .A(n6412), .B(n6914), .ZN(n6319) );
  XNOR2_X1 U7968 ( .A(n6319), .B(n9932), .ZN(n6906) );
  AND2_X1 U7969 ( .A1(n6316), .A2(n6906), .ZN(n6317) );
  INV_X1 U7970 ( .A(n9932), .ZN(n6963) );
  XNOR2_X1 U7971 ( .A(n6412), .B(n9967), .ZN(n6322) );
  XNOR2_X1 U7972 ( .A(n6322), .B(n9924), .ZN(n6932) );
  INV_X1 U7973 ( .A(n6322), .ZN(n6323) );
  INV_X1 U7974 ( .A(n9924), .ZN(n8354) );
  NAND2_X1 U7975 ( .A1(n6323), .A2(n8354), .ZN(n6324) );
  XNOR2_X1 U7976 ( .A(n6412), .B(n7216), .ZN(n6325) );
  XNOR2_X1 U7977 ( .A(n6325), .B(n9931), .ZN(n7055) );
  INV_X1 U7978 ( .A(n9931), .ZN(n7141) );
  XNOR2_X1 U7979 ( .A(n7244), .B(n6412), .ZN(n7137) );
  NAND2_X1 U7980 ( .A1(n7137), .A2(n8353), .ZN(n6326) );
  NAND2_X1 U7981 ( .A1(n7135), .A2(n6326), .ZN(n6329) );
  INV_X1 U7982 ( .A(n7137), .ZN(n6327) );
  NAND2_X1 U7983 ( .A1(n6327), .A2(n7136), .ZN(n6328) );
  XNOR2_X1 U7984 ( .A(n9980), .B(n6375), .ZN(n6331) );
  XNOR2_X1 U7985 ( .A(n6331), .B(n8352), .ZN(n7193) );
  INV_X1 U7986 ( .A(n7193), .ZN(n6330) );
  NAND2_X1 U7987 ( .A1(n6331), .A2(n8352), .ZN(n6332) );
  XNOR2_X1 U7988 ( .A(n6333), .B(n7339), .ZN(n7347) );
  XOR2_X1 U7989 ( .A(n6375), .B(n9986), .Z(n7348) );
  INV_X1 U7990 ( .A(n6333), .ZN(n6334) );
  XNOR2_X1 U7991 ( .A(n7337), .B(n6375), .ZN(n7403) );
  XOR2_X1 U7992 ( .A(n8349), .B(n6337), .Z(n7505) );
  XNOR2_X1 U7993 ( .A(n7606), .B(n6412), .ZN(n7566) );
  NAND2_X1 U7994 ( .A1(n7566), .A2(n8238), .ZN(n6340) );
  INV_X1 U7995 ( .A(n7566), .ZN(n6339) );
  XNOR2_X1 U7996 ( .A(n8855), .B(n6375), .ZN(n6341) );
  XOR2_X1 U7997 ( .A(n8347), .B(n6341), .Z(n8234) );
  OR2_X1 U7998 ( .A1(n6341), .A2(n8347), .ZN(n6342) );
  XNOR2_X1 U7999 ( .A(n8326), .B(n6375), .ZN(n6344) );
  XNOR2_X1 U8000 ( .A(n6344), .B(n8699), .ZN(n8328) );
  INV_X1 U8001 ( .A(n8328), .ZN(n6343) );
  INV_X1 U8002 ( .A(n6344), .ZN(n6346) );
  XNOR2_X1 U8003 ( .A(n8848), .B(n6375), .ZN(n6347) );
  XOR2_X1 U8004 ( .A(n8686), .B(n6347), .Z(n7681) );
  XNOR2_X1 U8005 ( .A(n8842), .B(n6375), .ZN(n6348) );
  NOR2_X1 U8006 ( .A1(n6348), .A2(n8700), .ZN(n8313) );
  AOI21_X1 U8007 ( .B1(n6348), .B2(n8700), .A(n8313), .ZN(n8269) );
  XNOR2_X1 U8008 ( .A(n8673), .B(n6412), .ZN(n6349) );
  NAND2_X1 U8009 ( .A1(n6349), .A2(n8658), .ZN(n8254) );
  INV_X1 U8010 ( .A(n6349), .ZN(n6350) );
  NAND2_X1 U8011 ( .A1(n6350), .A2(n8687), .ZN(n6351) );
  AND2_X1 U8012 ( .A1(n8254), .A2(n6351), .ZN(n8312) );
  XNOR2_X1 U8013 ( .A(n8769), .B(n6412), .ZN(n6352) );
  NAND2_X1 U8014 ( .A1(n6352), .A2(n8636), .ZN(n6355) );
  INV_X1 U8015 ( .A(n6352), .ZN(n6353) );
  NAND2_X1 U8016 ( .A1(n6353), .A2(n8667), .ZN(n6354) );
  NAND2_X1 U8017 ( .A1(n6355), .A2(n6354), .ZN(n8253) );
  INV_X1 U8018 ( .A(n6355), .ZN(n8292) );
  XNOR2_X1 U8019 ( .A(n8831), .B(n6412), .ZN(n6356) );
  NAND2_X1 U8020 ( .A1(n6356), .A2(n8659), .ZN(n8261) );
  INV_X1 U8021 ( .A(n6356), .ZN(n6357) );
  NAND2_X1 U8022 ( .A1(n6357), .A2(n8624), .ZN(n6358) );
  OAI21_X2 U8023 ( .B1(n8293), .B2(n8292), .A(n8291), .ZN(n8290) );
  XNOR2_X1 U8024 ( .A(n8825), .B(n6412), .ZN(n6359) );
  NAND2_X1 U8025 ( .A1(n6359), .A2(n8637), .ZN(n6362) );
  INV_X1 U8026 ( .A(n6359), .ZN(n6360) );
  NAND2_X1 U8027 ( .A1(n6360), .A2(n8346), .ZN(n6361) );
  NAND2_X1 U8028 ( .A1(n6362), .A2(n6361), .ZN(n8260) );
  AOI21_X2 U8029 ( .B1(n8290), .B2(n8261), .A(n8260), .ZN(n8303) );
  INV_X1 U8030 ( .A(n6362), .ZN(n8302) );
  XNOR2_X1 U8031 ( .A(n8756), .B(n6375), .ZN(n6363) );
  XNOR2_X1 U8032 ( .A(n6363), .B(n8263), .ZN(n8301) );
  OAI21_X2 U8033 ( .B1(n8303), .B2(n8302), .A(n8301), .ZN(n8300) );
  NAND2_X1 U8034 ( .A1(n8300), .A2(n6364), .ZN(n6366) );
  XOR2_X1 U8035 ( .A(n6375), .B(n8815), .Z(n6365) );
  XNOR2_X1 U8036 ( .A(n8809), .B(n6412), .ZN(n6369) );
  NAND2_X1 U8037 ( .A1(n6369), .A2(n8248), .ZN(n7721) );
  INV_X1 U8038 ( .A(n6369), .ZN(n6370) );
  NAND2_X1 U8039 ( .A1(n6370), .A2(n8605), .ZN(n6371) );
  XNOR2_X1 U8040 ( .A(n8803), .B(n6412), .ZN(n6373) );
  XNOR2_X1 U8041 ( .A(n6373), .B(n8590), .ZN(n6372) );
  INV_X1 U8042 ( .A(n6372), .ZN(n7722) );
  XOR2_X1 U8043 ( .A(n6375), .B(n8798), .Z(n7708) );
  XNOR2_X1 U8044 ( .A(n8738), .B(n6375), .ZN(n6417) );
  NAND2_X1 U8045 ( .A1(n6417), .A2(n8571), .ZN(n6421) );
  OAI21_X1 U8046 ( .B1(n6417), .B2(n8571), .A(n6421), .ZN(n6381) );
  OR2_X1 U8047 ( .A1(n6385), .A2(n6376), .ZN(n6379) );
  NAND2_X1 U8048 ( .A1(n6388), .A2(n6377), .ZN(n6378) );
  AOI21_X1 U8049 ( .B1(n6380), .B2(n6381), .A(n8327), .ZN(n6384) );
  INV_X1 U8050 ( .A(n6381), .ZN(n6382) );
  NAND2_X1 U8051 ( .A1(n6383), .A2(n6382), .ZN(n6426) );
  NAND2_X1 U8052 ( .A1(n6384), .A2(n6426), .ZN(n6411) );
  INV_X1 U8053 ( .A(n8738), .ZN(n8564) );
  OR2_X1 U8054 ( .A1(n6385), .A2(n9989), .ZN(n6387) );
  INV_X1 U8055 ( .A(n8250), .ZN(n8341) );
  AND2_X1 U8056 ( .A1(n6388), .A2(n6840), .ZN(n6389) );
  INV_X1 U8057 ( .A(n6389), .ZN(n6391) );
  INV_X1 U8058 ( .A(n6403), .ZN(n6399) );
  INV_X1 U8059 ( .A(n6392), .ZN(n6394) );
  NAND2_X1 U8060 ( .A1(n6394), .A2(n6393), .ZN(n6397) );
  AND3_X1 U8061 ( .A1(n6395), .A2(n6537), .A3(n6533), .ZN(n6396) );
  OAI211_X1 U8062 ( .C1(n6399), .C2(n6398), .A(n6397), .B(n6396), .ZN(n6400)
         );
  NAND2_X1 U8063 ( .A1(n6400), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6405) );
  INV_X1 U8064 ( .A(n6840), .ZN(n6402) );
  NOR2_X1 U8065 ( .A1(n6402), .A2(n6401), .ZN(n8227) );
  NAND2_X1 U8066 ( .A1(n8227), .A2(n6403), .ZN(n6404) );
  AOI22_X1 U8067 ( .A1(n8562), .A2(n8323), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6406) );
  OAI21_X1 U8068 ( .B1(n8557), .B2(n8320), .A(n6406), .ZN(n6407) );
  AOI21_X1 U8069 ( .B1(n8318), .B2(n8555), .A(n6407), .ZN(n6408) );
  OAI21_X1 U8070 ( .B1(n8564), .B2(n8341), .A(n6408), .ZN(n6409) );
  INV_X1 U8071 ( .A(n6409), .ZN(n6410) );
  NAND2_X1 U8072 ( .A1(n6411), .A2(n6410), .ZN(P2_U3154) );
  XNOR2_X1 U8073 ( .A(n8555), .B(n6412), .ZN(n6413) );
  XNOR2_X1 U8074 ( .A(n8547), .B(n6413), .ZN(n6422) );
  INV_X1 U8075 ( .A(n6422), .ZN(n6414) );
  NAND2_X1 U8076 ( .A1(n6414), .A2(n8315), .ZN(n6425) );
  NAND2_X1 U8077 ( .A1(n8345), .A2(n8318), .ZN(n6416) );
  AOI22_X1 U8078 ( .A1(n8546), .A2(n8323), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n6415) );
  OAI211_X1 U8079 ( .C1(n7713), .C2(n8320), .A(n6416), .B(n6415), .ZN(n6420)
         );
  INV_X1 U8080 ( .A(n6417), .ZN(n6418) );
  NOR4_X1 U8081 ( .A1(n6422), .A2(n6418), .A3(n7713), .A4(n8327), .ZN(n6419)
         );
  AOI211_X1 U8082 ( .C1(n8547), .C2(n8250), .A(n6420), .B(n6419), .ZN(n6424)
         );
  NAND2_X1 U8083 ( .A1(n6426), .A2(n4957), .ZN(n6423) );
  OAI211_X1 U8084 ( .C1(n6426), .C2(n6425), .A(n6424), .B(n6423), .ZN(P2_U3160) );
  NAND2_X1 U8085 ( .A1(n8020), .A2(n7782), .ZN(n6428) );
  INV_X1 U8086 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8021) );
  OR2_X1 U8087 ( .A1(n4342), .A2(n8021), .ZN(n6427) );
  INV_X1 U8088 ( .A(n9038), .ZN(n6516) );
  INV_X1 U8089 ( .A(n9040), .ZN(n7776) );
  INV_X1 U8090 ( .A(n9356), .ZN(n9017) );
  INV_X1 U8091 ( .A(n8928), .ZN(n9042) );
  INV_X1 U8092 ( .A(n9367), .ZN(n9207) );
  INV_X1 U8093 ( .A(n8980), .ZN(n9043) );
  INV_X1 U8094 ( .A(n9371), .ZN(n9215) );
  XNOR2_X2 U8095 ( .A(n6493), .B(n6429), .ZN(n9727) );
  AND2_X1 U8096 ( .A1(n7737), .A2(n9762), .ZN(n9726) );
  NAND2_X1 U8097 ( .A1(n6780), .A2(n7949), .ZN(n6431) );
  NAND2_X1 U8098 ( .A1(n6851), .A2(n9774), .ZN(n6430) );
  NAND2_X1 U8099 ( .A1(n6431), .A2(n6430), .ZN(n6921) );
  NAND2_X1 U8100 ( .A1(n9058), .A2(n9780), .ZN(n7823) );
  AND2_X1 U8101 ( .A1(n4387), .A2(n7823), .ZN(n7947) );
  INV_X1 U8102 ( .A(n7947), .ZN(n6922) );
  NAND2_X1 U8103 ( .A1(n6921), .A2(n6922), .ZN(n6433) );
  INV_X1 U8104 ( .A(n9058), .ZN(n6816) );
  NAND2_X1 U8105 ( .A1(n6816), .A2(n9780), .ZN(n6432) );
  NAND2_X1 U8106 ( .A1(n6433), .A2(n6432), .ZN(n7065) );
  INV_X1 U8107 ( .A(n9057), .ZN(n7081) );
  NAND2_X1 U8108 ( .A1(n7081), .A2(n9786), .ZN(n7825) );
  AND2_X1 U8109 ( .A1(n9057), .A2(n7073), .ZN(n7812) );
  NAND2_X1 U8110 ( .A1(n7825), .A2(n7827), .ZN(n7950) );
  NAND2_X1 U8111 ( .A1(n7065), .A2(n7950), .ZN(n6435) );
  NAND2_X1 U8112 ( .A1(n7081), .A2(n7073), .ZN(n6434) );
  NAND2_X1 U8113 ( .A1(n6435), .A2(n6434), .ZN(n6969) );
  INV_X1 U8114 ( .A(n9056), .ZN(n7154) );
  INV_X1 U8115 ( .A(n6971), .ZN(n9795) );
  NAND2_X1 U8116 ( .A1(n9056), .A2(n9795), .ZN(n7814) );
  NAND2_X1 U8117 ( .A1(n7154), .A2(n9795), .ZN(n6436) );
  NAND2_X1 U8118 ( .A1(n7165), .A2(n6519), .ZN(n7819) );
  NAND2_X1 U8119 ( .A1(n9055), .A2(n9721), .ZN(n7815) );
  NAND2_X1 U8120 ( .A1(n7330), .A2(n7182), .ZN(n7219) );
  INV_X1 U8121 ( .A(n7330), .ZN(n9054) );
  NAND2_X1 U8122 ( .A1(n9802), .A2(n9054), .ZN(n7834) );
  INV_X1 U8123 ( .A(n7832), .ZN(n7179) );
  NAND2_X1 U8124 ( .A1(n7178), .A2(n7179), .ZN(n6438) );
  NAND2_X1 U8125 ( .A1(n7330), .A2(n9802), .ZN(n6437) );
  NAND2_X1 U8126 ( .A1(n6438), .A2(n6437), .ZN(n7225) );
  OR2_X1 U8127 ( .A1(n7228), .A2(n7426), .ZN(n7835) );
  NAND2_X1 U8128 ( .A1(n7228), .A2(n7426), .ZN(n7839) );
  NAND2_X1 U8129 ( .A1(n7835), .A2(n7839), .ZN(n7226) );
  INV_X1 U8130 ( .A(n7426), .ZN(n9053) );
  OR2_X1 U8131 ( .A1(n7228), .A2(n9053), .ZN(n6439) );
  INV_X1 U8132 ( .A(n9052), .ZN(n6440) );
  OR2_X1 U8133 ( .A1(n9706), .A2(n6440), .ZN(n7850) );
  NAND2_X1 U8134 ( .A1(n4343), .A2(n6440), .ZN(n7840) );
  NAND2_X1 U8135 ( .A1(n7850), .A2(n7840), .ZN(n7278) );
  INV_X1 U8136 ( .A(n9051), .ZN(n6441) );
  OR2_X1 U8137 ( .A1(n9818), .A2(n6441), .ZN(n7852) );
  AND2_X1 U8138 ( .A1(n9818), .A2(n6441), .ZN(n7849) );
  INV_X1 U8139 ( .A(n7849), .ZN(n7748) );
  INV_X1 U8140 ( .A(n9699), .ZN(n9705) );
  OR2_X1 U8141 ( .A1(n9691), .A2(n9050), .ZN(n6446) );
  INV_X1 U8142 ( .A(n6446), .ZN(n6443) );
  INV_X1 U8143 ( .A(n9050), .ZN(n6442) );
  OR2_X1 U8144 ( .A1(n9691), .A2(n6442), .ZN(n9682) );
  NAND2_X1 U8145 ( .A1(n9691), .A2(n6442), .ZN(n7853) );
  NAND2_X1 U8146 ( .A1(n9682), .A2(n7853), .ZN(n9678) );
  OR2_X1 U8147 ( .A1(n6443), .A2(n9678), .ZN(n6445) );
  AND2_X1 U8148 ( .A1(n9705), .A2(n6445), .ZN(n6444) );
  NAND2_X1 U8149 ( .A1(n9673), .A2(n6444), .ZN(n6450) );
  INV_X1 U8150 ( .A(n6445), .ZN(n6448) );
  OR2_X1 U8151 ( .A1(n9818), .A2(n9051), .ZN(n9674) );
  AND2_X1 U8152 ( .A1(n9674), .A2(n6446), .ZN(n6447) );
  OR2_X1 U8153 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  NAND2_X1 U8154 ( .A1(n6450), .A2(n6449), .ZN(n9666) );
  OR2_X1 U8155 ( .A1(n9665), .A2(n7585), .ZN(n7857) );
  NAND2_X1 U8156 ( .A1(n9665), .A2(n7585), .ZN(n7854) );
  NAND2_X1 U8157 ( .A1(n7857), .A2(n7854), .ZN(n9667) );
  INV_X1 U8158 ( .A(n7585), .ZN(n9049) );
  OR2_X1 U8159 ( .A1(n9665), .A2(n9049), .ZN(n6451) );
  NAND2_X1 U8160 ( .A1(n9839), .A2(n9048), .ZN(n7861) );
  NAND2_X1 U8161 ( .A1(n7560), .A2(n9047), .ZN(n6452) );
  NAND2_X1 U8162 ( .A1(n7524), .A2(n6452), .ZN(n6454) );
  OR2_X1 U8163 ( .A1(n7560), .A2(n9047), .ZN(n6453) );
  NOR2_X1 U8164 ( .A1(n9402), .A2(n9046), .ZN(n6455) );
  NAND2_X1 U8165 ( .A1(n9402), .A2(n9046), .ZN(n6456) );
  OR2_X1 U8166 ( .A1(n9512), .A2(n9026), .ZN(n7871) );
  NAND2_X1 U8167 ( .A1(n9512), .A2(n9026), .ZN(n7872) );
  NAND2_X1 U8168 ( .A1(n7871), .A2(n7872), .ZN(n9324) );
  OR2_X1 U8169 ( .A1(n9323), .A2(n9301), .ZN(n7878) );
  AND2_X1 U8170 ( .A1(n9324), .A2(n7878), .ZN(n6457) );
  INV_X1 U8171 ( .A(n7878), .ZN(n6459) );
  NAND2_X1 U8172 ( .A1(n9323), .A2(n9301), .ZN(n7879) );
  INV_X1 U8173 ( .A(n9026), .ZN(n9310) );
  NAND2_X1 U8174 ( .A1(n9512), .A2(n9310), .ZN(n9325) );
  AND2_X1 U8175 ( .A1(n7879), .A2(n9325), .ZN(n6458) );
  OR2_X1 U8176 ( .A1(n6459), .A2(n6458), .ZN(n6460) );
  NAND2_X1 U8177 ( .A1(n6461), .A2(n6460), .ZN(n9291) );
  NAND2_X1 U8178 ( .A1(n9297), .A2(n8886), .ZN(n6463) );
  NOR2_X1 U8179 ( .A1(n9297), .A2(n8886), .ZN(n6462) );
  NAND2_X1 U8180 ( .A1(n9286), .A2(n9302), .ZN(n6464) );
  INV_X1 U8181 ( .A(n9257), .ZN(n6466) );
  NAND2_X1 U8182 ( .A1(n9381), .A2(n8982), .ZN(n7901) );
  NAND2_X1 U8183 ( .A1(n7903), .A2(n7901), .ZN(n9242) );
  INV_X1 U8184 ( .A(n9225), .ZN(n6469) );
  OAI21_X1 U8185 ( .B1(n9367), .B2(n9042), .A(n6470), .ZN(n9183) );
  INV_X1 U8186 ( .A(n9183), .ZN(n6472) );
  INV_X1 U8187 ( .A(n9041), .ZN(n9009) );
  NAND2_X1 U8188 ( .A1(n9352), .A2(n9007), .ZN(n7917) );
  NAND2_X1 U8189 ( .A1(n9346), .A2(n6516), .ZN(n7927) );
  NAND2_X1 U8190 ( .A1(n9138), .A2(n9145), .ZN(n9137) );
  NAND2_X1 U8191 ( .A1(n6474), .A2(n7782), .ZN(n6476) );
  OR2_X1 U8192 ( .A1(n4342), .A2(n7655), .ZN(n6475) );
  INV_X1 U8193 ( .A(n6477), .ZN(n6523) );
  NAND2_X1 U8194 ( .A1(n6478), .A2(n6523), .ZN(n6482) );
  NAND2_X1 U8195 ( .A1(n4340), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U8196 ( .A1(n4335), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8197 ( .A1(n5520), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6479) );
  NAND4_X1 U8198 ( .A1(n6482), .A2(n6481), .A3(n6480), .A4(n6479), .ZN(n9037)
         );
  INV_X1 U8199 ( .A(n9037), .ZN(n6483) );
  NAND2_X1 U8200 ( .A1(n9341), .A2(n6483), .ZN(n7929) );
  INV_X1 U8201 ( .A(n9334), .ZN(n6488) );
  INV_X1 U8202 ( .A(n9333), .ZN(n7262) );
  NOR2_X1 U8203 ( .A1(n7262), .A2(n6486), .ZN(n6487) );
  NAND2_X1 U8204 ( .A1(n6488), .A2(n6487), .ZN(n6521) );
  NAND2_X1 U8205 ( .A1(n9752), .A2(n6489), .ZN(n9686) );
  INV_X1 U8206 ( .A(n9763), .ZN(n9746) );
  OAI211_X1 U8207 ( .C1(n6491), .C2(n6490), .A(n9746), .B(n9743), .ZN(n7529)
         );
  INV_X1 U8208 ( .A(n7529), .ZN(n9732) );
  NAND2_X1 U8209 ( .A1(n9752), .A2(n9732), .ZN(n6492) );
  NAND2_X1 U8210 ( .A1(n9727), .A2(n7945), .ZN(n6495) );
  INV_X1 U8211 ( .A(n6493), .ZN(n6815) );
  NAND2_X1 U8212 ( .A1(n6815), .A2(n9740), .ZN(n6494) );
  NAND2_X1 U8213 ( .A1(n6495), .A2(n6494), .ZN(n6778) );
  NAND2_X1 U8214 ( .A1(n7813), .A2(n7825), .ZN(n7066) );
  NAND2_X1 U8215 ( .A1(n7066), .A2(n7827), .ZN(n6965) );
  OR2_X1 U8216 ( .A1(n6965), .A2(n6970), .ZN(n6496) );
  AND2_X1 U8217 ( .A1(n6496), .A2(n7816), .ZN(n7173) );
  AND2_X1 U8218 ( .A1(n7850), .A2(n7835), .ZN(n7841) );
  INV_X1 U8219 ( .A(n7841), .ZN(n6502) );
  NAND2_X1 U8220 ( .A1(n7839), .A2(n7219), .ZN(n7836) );
  INV_X1 U8221 ( .A(n7836), .ZN(n6497) );
  OR2_X1 U8222 ( .A1(n6502), .A2(n6497), .ZN(n6498) );
  NAND2_X1 U8223 ( .A1(n6498), .A2(n7840), .ZN(n6499) );
  INV_X1 U8224 ( .A(n7815), .ZN(n6504) );
  INV_X1 U8225 ( .A(n7834), .ZN(n6501) );
  NOR2_X1 U8226 ( .A1(n6502), .A2(n6501), .ZN(n7957) );
  INV_X1 U8227 ( .A(n7957), .ZN(n6503) );
  OAI21_X1 U8228 ( .B1(n6504), .B2(n6503), .A(n7744), .ZN(n7747) );
  AOI21_X1 U8229 ( .B1(n7173), .B2(n6506), .A(n6505), .ZN(n9698) );
  NAND2_X1 U8230 ( .A1(n9698), .A2(n9699), .ZN(n9697) );
  NAND2_X1 U8231 ( .A1(n9680), .A2(n7853), .ZN(n9660) );
  NAND2_X1 U8232 ( .A1(n7857), .A2(n9682), .ZN(n7736) );
  INV_X1 U8233 ( .A(n7736), .ZN(n7751) );
  NAND2_X1 U8234 ( .A1(n7390), .A2(n7854), .ZN(n6507) );
  OR2_X1 U8235 ( .A1(n7560), .A2(n9024), .ZN(n7865) );
  AND2_X1 U8236 ( .A1(n7560), .A2(n9024), .ZN(n7876) );
  INV_X1 U8237 ( .A(n7876), .ZN(n7862) );
  NAND2_X1 U8238 ( .A1(n7865), .A2(n7862), .ZN(n7963) );
  INV_X1 U8239 ( .A(n9046), .ZN(n8944) );
  OR2_X1 U8240 ( .A1(n9402), .A2(n8944), .ZN(n7755) );
  NAND2_X1 U8241 ( .A1(n9402), .A2(n8944), .ZN(n7754) );
  NAND2_X1 U8242 ( .A1(n7755), .A2(n7754), .ZN(n7962) );
  NAND2_X1 U8243 ( .A1(n7645), .A2(n7644), .ZN(n7643) );
  NAND2_X1 U8244 ( .A1(n7643), .A2(n7754), .ZN(n7629) );
  INV_X1 U8245 ( .A(n9301), .ZN(n8996) );
  OR2_X1 U8246 ( .A1(n9323), .A2(n8996), .ZN(n7757) );
  NAND2_X1 U8247 ( .A1(n9323), .A2(n8996), .ZN(n7760) );
  OR2_X1 U8248 ( .A1(n9397), .A2(n8886), .ZN(n7763) );
  NAND2_X1 U8249 ( .A1(n9397), .A2(n8886), .ZN(n7761) );
  NAND2_X1 U8250 ( .A1(n9300), .A2(n9299), .ZN(n9298) );
  NAND2_X1 U8251 ( .A1(n9298), .A2(n7761), .ZN(n9275) );
  AND2_X1 U8252 ( .A1(n9392), .A2(n9302), .ZN(n7894) );
  INV_X1 U8253 ( .A(n7894), .ZN(n7764) );
  AND2_X1 U8254 ( .A1(n9265), .A2(n9278), .ZN(n7810) );
  INV_X1 U8255 ( .A(n7810), .ZN(n9241) );
  AND2_X1 U8256 ( .A1(n9386), .A2(n8917), .ZN(n7808) );
  INV_X1 U8257 ( .A(n7808), .ZN(n6508) );
  NAND2_X1 U8258 ( .A1(n7901), .A2(n6508), .ZN(n6509) );
  NAND2_X1 U8259 ( .A1(n6509), .A2(n7903), .ZN(n7904) );
  NAND2_X1 U8260 ( .A1(n9376), .A2(n8918), .ZN(n7770) );
  NAND2_X1 U8261 ( .A1(n9371), .A2(n8980), .ZN(n7908) );
  OR2_X1 U8262 ( .A1(n9367), .A2(n8928), .ZN(n7911) );
  NAND2_X1 U8263 ( .A1(n9367), .A2(n8928), .ZN(n7910) );
  INV_X1 U8264 ( .A(n9199), .ZN(n7969) );
  INV_X1 U8265 ( .A(n7911), .ZN(n6510) );
  INV_X1 U8266 ( .A(n7921), .ZN(n7734) );
  NAND2_X1 U8267 ( .A1(n9361), .A2(n9009), .ZN(n7923) );
  NAND2_X1 U8268 ( .A1(n7734), .A2(n7923), .ZN(n9190) );
  XNOR2_X1 U8269 ( .A(n9356), .B(n7776), .ZN(n7971) );
  AND2_X1 U8270 ( .A1(n9356), .A2(n7776), .ZN(n7926) );
  NAND2_X1 U8271 ( .A1(n9166), .A2(n9165), .ZN(n9149) );
  AOI21_X1 U8272 ( .B1(n9149), .B2(n7925), .A(n9145), .ZN(n9148) );
  NOR2_X1 U8273 ( .A1(n9148), .A2(n7919), .ZN(n6511) );
  XOR2_X1 U8274 ( .A(n6511), .B(n7972), .Z(n6518) );
  AND2_X1 U8275 ( .A1(n5096), .A2(n9747), .ZN(n7944) );
  INV_X1 U8276 ( .A(n7944), .ZN(n6512) );
  NAND2_X1 U8277 ( .A1(n7739), .A2(n8000), .ZN(n8005) );
  INV_X1 U8278 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U8279 ( .A1(n5520), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8280 ( .A1(n4335), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6513) );
  OAI211_X1 U8281 ( .C1(n4337), .C2(n9132), .A(n6514), .B(n6513), .ZN(n9036)
         );
  INV_X1 U8282 ( .A(n9036), .ZN(n7786) );
  OR2_X1 U8283 ( .A1(n7626), .A2(n10211), .ZN(n6515) );
  NAND2_X1 U8284 ( .A1(n9311), .A2(n6515), .ZN(n9124) );
  OAI22_X1 U8285 ( .A1(n6516), .A2(n9008), .B1(n7786), .B2(n9124), .ZN(n6517)
         );
  NAND2_X1 U8286 ( .A1(n9767), .A2(n9735), .ZN(n9733) );
  INV_X1 U8287 ( .A(n7228), .ZN(n9809) );
  NAND2_X1 U8288 ( .A1(n9265), .A2(n9282), .ZN(n9267) );
  INV_X1 U8289 ( .A(n9734), .ZN(n9246) );
  AOI211_X1 U8290 ( .C1(n9341), .C2(n9141), .A(n9246), .B(n9131), .ZN(n9340)
         );
  INV_X1 U8291 ( .A(n9341), .ZN(n6525) );
  NAND2_X1 U8292 ( .A1(n9752), .A2(n6522), .ZN(n9720) );
  AOI22_X1 U8293 ( .A1(n9754), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n6523), .B2(
        n9749), .ZN(n6524) );
  OAI21_X1 U8294 ( .B1(n6525), .B2(n9720), .A(n6524), .ZN(n6526) );
  AOI21_X1 U8295 ( .B1(n9340), .B2(n9738), .A(n6526), .ZN(n6527) );
  INV_X1 U8296 ( .A(n6527), .ZN(n6528) );
  NOR2_X1 U8297 ( .A1(n6531), .A2(P1_U3086), .ZN(n6532) );
  INV_X1 U8298 ( .A(n6533), .ZN(n7411) );
  OR2_X1 U8299 ( .A1(n8206), .A2(n7411), .ZN(n6534) );
  OR2_X1 U8300 ( .A1(n6537), .A2(n7411), .ZN(n6601) );
  NAND2_X1 U8301 ( .A1(n6534), .A2(n6601), .ZN(n6605) );
  OAI21_X1 U8302 ( .B1(n6605), .B2(n6535), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  INV_X1 U8303 ( .A(n6584), .ZN(n6536) );
  NOR2_X1 U8304 ( .A1(n7795), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9431) );
  INV_X1 U8305 ( .A(n9431), .ZN(n9438) );
  NAND2_X1 U8306 ( .A1(n7795), .A2(P1_U3086), .ZN(n9436) );
  OAI222_X1 U8307 ( .A1(n9438), .A2(n4476), .B1(n6745), .B2(P1_U3086), .C1(
        n9436), .C2(n6553), .ZN(P1_U3353) );
  OAI222_X1 U8308 ( .A1(n9438), .A2(n6587), .B1(n9537), .B2(P1_U3086), .C1(
        n9436), .C2(n6549), .ZN(P1_U3354) );
  OAI222_X1 U8309 ( .A1(n9438), .A2(n6538), .B1(n6678), .B2(P1_U3086), .C1(
        n9436), .C2(n6554), .ZN(P1_U3351) );
  INV_X1 U8310 ( .A(n9436), .ZN(n7414) );
  INV_X1 U8311 ( .A(n7414), .ZN(n8023) );
  OAI222_X1 U8312 ( .A1(n8023), .A2(n6544), .B1(n9551), .B2(P1_U3086), .C1(
        n6539), .C2(n9438), .ZN(P1_U3350) );
  OAI222_X1 U8313 ( .A1(n8023), .A2(n6542), .B1(n9565), .B2(P1_U3086), .C1(
        n6540), .C2(n9438), .ZN(P1_U3349) );
  OAI222_X1 U8314 ( .A1(n9438), .A2(n6541), .B1(n9484), .B2(P1_U3086), .C1(
        n8023), .C2(n6552), .ZN(P1_U3352) );
  NOR2_X1 U8315 ( .A1(n7795), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8865) );
  INV_X2 U8316 ( .A(n8865), .ZN(n8017) );
  OAI222_X1 U8317 ( .A1(n8019), .A2(n6543), .B1(n8017), .B2(n6542), .C1(n7043), 
        .C2(P2_U3151), .ZN(P2_U3289) );
  OAI222_X1 U8318 ( .A1(n8019), .A2(n6545), .B1(n8017), .B2(n6544), .C1(n6869), 
        .C2(P2_U3151), .ZN(P2_U3290) );
  INV_X1 U8319 ( .A(n6641), .ZN(n9467) );
  INV_X1 U8320 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6546) );
  OAI222_X1 U8321 ( .A1(n8023), .A2(n6547), .B1(n9467), .B2(P1_U3086), .C1(
        n6546), .C2(n9438), .ZN(P1_U3348) );
  OAI222_X1 U8322 ( .A1(n8019), .A2(n6548), .B1(n8017), .B2(n6547), .C1(n7116), 
        .C2(P2_U3151), .ZN(P2_U3288) );
  OAI222_X1 U8323 ( .A1(P2_U3151), .A2(n6714), .B1(n8019), .B2(n6550), .C1(
        n8017), .C2(n6549), .ZN(P2_U3294) );
  OAI222_X1 U8324 ( .A1(P2_U3151), .A2(n6762), .B1(n8017), .B2(n6552), .C1(
        n6551), .C2(n8019), .ZN(P2_U3292) );
  OAI222_X1 U8325 ( .A1(P2_U3151), .A2(n9912), .B1(n8017), .B2(n6553), .C1(
        n4982), .C2(n8019), .ZN(P2_U3293) );
  OAI222_X1 U8326 ( .A1(P2_U3151), .A2(n6799), .B1(n8017), .B2(n6554), .C1(
        n4977), .C2(n8019), .ZN(P2_U3291) );
  INV_X1 U8327 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6556) );
  INV_X1 U8328 ( .A(n6555), .ZN(n6557) );
  INV_X1 U8329 ( .A(n6644), .ZN(n9503) );
  OAI222_X1 U8330 ( .A1(n9438), .A2(n6556), .B1(n9436), .B2(n6557), .C1(
        P1_U3086), .C2(n9503), .ZN(P1_U3347) );
  INV_X1 U8331 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6558) );
  OAI222_X1 U8332 ( .A1(n8019), .A2(n6558), .B1(n8017), .B2(n6557), .C1(
        P2_U3151), .C2(n7299), .ZN(P2_U3287) );
  INV_X1 U8333 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6560) );
  NOR2_X1 U8334 ( .A1(n6579), .A2(n6560), .ZN(P2_U3256) );
  INV_X1 U8335 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10199) );
  NOR2_X1 U8336 ( .A1(n6579), .A2(n10199), .ZN(P2_U3238) );
  INV_X1 U8337 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10195) );
  NOR2_X1 U8338 ( .A1(n6579), .A2(n10195), .ZN(P2_U3260) );
  INV_X1 U8339 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6561) );
  NOR2_X1 U8340 ( .A1(n6579), .A2(n6561), .ZN(P2_U3253) );
  INV_X1 U8341 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6562) );
  NOR2_X1 U8342 ( .A1(n6579), .A2(n6562), .ZN(P2_U3242) );
  INV_X1 U8343 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10172) );
  NOR2_X1 U8344 ( .A1(n6579), .A2(n10172), .ZN(P2_U3237) );
  INV_X1 U8345 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U8346 ( .A1(n6579), .A2(n10208), .ZN(P2_U3258) );
  AOI22_X1 U8347 ( .A1(n9449), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9431), .ZN(n6563) );
  OAI21_X1 U8348 ( .B1(n6566), .B2(n9436), .A(n6563), .ZN(P1_U3345) );
  INV_X1 U8349 ( .A(n6564), .ZN(n6572) );
  INV_X1 U8350 ( .A(n7000), .ZN(n6650) );
  OAI222_X1 U8351 ( .A1(n8023), .A2(n6572), .B1(n6650), .B2(P1_U3086), .C1(
        n6565), .C2(n9438), .ZN(P1_U3346) );
  INV_X1 U8352 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6567) );
  INV_X1 U8353 ( .A(n7447), .ZN(n7378) );
  OAI222_X1 U8354 ( .A1(n8019), .A2(n6567), .B1(n8017), .B2(n6566), .C1(n7378), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  AOI21_X1 U8355 ( .B1(n6570), .B2(n6569), .A(n6568), .ZN(n6597) );
  INV_X1 U8356 ( .A(n6597), .ZN(n6571) );
  NAND2_X1 U8357 ( .A1(n9423), .A2(n8015), .ZN(n6596) );
  AND2_X1 U8358 ( .A1(n6571), .A2(n6596), .ZN(n9522) );
  NOR2_X1 U8359 ( .A1(n9522), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI222_X1 U8360 ( .A1(n8019), .A2(n6573), .B1(n8017), .B2(n6572), .C1(n7373), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8361 ( .A(n6579), .ZN(n6574) );
  AND2_X1 U8362 ( .A1(n6574), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8363 ( .A1(n6574), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8364 ( .A1(n6574), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8365 ( .A1(n6574), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8366 ( .A1(n6574), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8367 ( .A1(n6574), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8368 ( .A1(n6574), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8369 ( .A1(n6574), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  NAND2_X1 U8370 ( .A1(n7737), .A2(P1_U3973), .ZN(n6575) );
  OAI21_X1 U8371 ( .B1(P1_U3973), .B2(n5788), .A(n6575), .ZN(P1_U3554) );
  NAND2_X1 U8372 ( .A1(n6946), .A2(P2_U3893), .ZN(n6576) );
  OAI21_X1 U8373 ( .B1(P2_U3893), .B2(n5148), .A(n6576), .ZN(P2_U3491) );
  INV_X1 U8374 ( .A(n6577), .ZN(n6589) );
  AOI22_X1 U8375 ( .A1(n9570), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9431), .ZN(n6578) );
  OAI21_X1 U8376 ( .B1(n6589), .B2(n8023), .A(n6578), .ZN(P1_U3344) );
  AND2_X1 U8377 ( .A1(n6574), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8378 ( .A1(n6574), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8379 ( .A1(n6574), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8380 ( .A1(n6574), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8381 ( .A1(n6574), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8382 ( .A1(n6574), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8383 ( .A1(n6574), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8384 ( .A1(n6574), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8385 ( .A1(n6574), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8386 ( .A1(n6574), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8387 ( .A1(n6574), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8388 ( .A1(n6574), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8389 ( .A1(n6574), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8390 ( .A1(n6574), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8391 ( .A1(n6574), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  INV_X1 U8392 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6582) );
  INV_X1 U8393 ( .A(n6580), .ZN(n6581) );
  AOI22_X1 U8394 ( .A1(n6574), .A2(n6582), .B1(n6584), .B2(n6581), .ZN(
        P2_U3377) );
  INV_X1 U8395 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6586) );
  INV_X1 U8396 ( .A(n6583), .ZN(n6585) );
  AOI22_X1 U8397 ( .A1(n6574), .A2(n6586), .B1(n6585), .B2(n6584), .ZN(
        P2_U3376) );
  MUX2_X1 U8398 ( .A(n6587), .B(n6303), .S(P2_U3893), .Z(n6588) );
  INV_X1 U8399 ( .A(n6588), .ZN(P2_U3492) );
  INV_X1 U8400 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6590) );
  INV_X1 U8401 ( .A(n7386), .ZN(n7486) );
  OAI222_X1 U8402 ( .A1(n8019), .A2(n6590), .B1(n8017), .B2(n6589), .C1(
        P2_U3151), .C2(n7486), .ZN(P2_U3284) );
  INV_X1 U8403 ( .A(n9077), .ZN(n7011) );
  INV_X1 U8404 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6591) );
  OAI222_X1 U8405 ( .A1(n8023), .A2(n6592), .B1(n7011), .B2(P1_U3086), .C1(
        n6591), .C2(n9438), .ZN(P1_U3343) );
  INV_X1 U8406 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6593) );
  INV_X1 U8407 ( .A(n8377), .ZN(n7475) );
  OAI222_X1 U8408 ( .A1(n8019), .A2(n6593), .B1(n8017), .B2(n6592), .C1(n7475), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8409 ( .A(n7626), .ZN(n6663) );
  INV_X1 U8410 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6594) );
  AOI21_X1 U8411 ( .B1(n6663), .B2(n6594), .A(n5737), .ZN(n6664) );
  OAI21_X1 U8412 ( .B1(n6663), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6664), .ZN(
        n6595) );
  MUX2_X1 U8413 ( .A(n6664), .B(n6595), .S(n6625), .Z(n6600) );
  NAND2_X1 U8414 ( .A1(n6597), .A2(n6596), .ZN(n6648) );
  AOI22_X1 U8415 ( .A1(n9522), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6599) );
  INV_X1 U8416 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9855) );
  NAND3_X1 U8417 ( .A1(n9112), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9855), .ZN(
        n6598) );
  OAI211_X1 U8418 ( .C1(n6600), .C2(n6648), .A(n6599), .B(n6598), .ZN(P1_U3243) );
  NOR2_X1 U8419 ( .A1(n6605), .A2(n8503), .ZN(n6602) );
  INV_X1 U8420 ( .A(n6601), .ZN(n6604) );
  MUX2_X1 U8421 ( .A(n6602), .B(n6604), .S(n8226), .Z(n6603) );
  NAND2_X1 U8422 ( .A1(n6603), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9913) );
  OR2_X1 U8423 ( .A1(n6165), .A2(P2_U3151), .ZN(n7650) );
  NOR2_X1 U8424 ( .A1(n6605), .A2(n7650), .ZN(n6723) );
  OR2_X1 U8425 ( .A1(n8507), .A2(n8226), .ZN(n8509) );
  INV_X1 U8426 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6832) );
  MUX2_X1 U8427 ( .A(n6606), .B(n6832), .S(n8503), .Z(n6607) );
  NAND2_X1 U8428 ( .A1(n6607), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9884) );
  OAI21_X1 U8429 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6607), .A(n9884), .ZN(n6608) );
  OAI21_X1 U8430 ( .B1(n6723), .B2(n9906), .A(n6608), .ZN(n6609) );
  OAI21_X1 U8431 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6662), .A(n6609), .ZN(n6610) );
  AOI21_X1 U8432 ( .B1(n9905), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6610), .ZN(
        n6611) );
  OAI21_X1 U8433 ( .B1(n6712), .B2(n9913), .A(n6611), .ZN(P2_U3182) );
  AOI22_X1 U8434 ( .A1(n9589), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9431), .ZN(n6612) );
  OAI21_X1 U8435 ( .B1(n6613), .B2(n9436), .A(n6612), .ZN(P1_U3342) );
  INV_X1 U8436 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6614) );
  INV_X1 U8437 ( .A(n8387), .ZN(n8380) );
  OAI222_X1 U8438 ( .A1(n8019), .A2(n6614), .B1(n8017), .B2(n6613), .C1(n8380), 
        .C2(P2_U3151), .ZN(P2_U3282) );
  INV_X1 U8439 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6615) );
  AOI22_X1 U8440 ( .A1(n7000), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6615), .B2(
        n6650), .ZN(n6622) );
  INV_X1 U8441 ( .A(n9565), .ZN(n6638) );
  INV_X1 U8442 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7071) );
  MUX2_X1 U8443 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7071), .S(n6678), .Z(n6669)
         );
  NAND2_X1 U8444 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9523) );
  NOR2_X1 U8445 ( .A1(n9524), .A2(n9523), .ZN(n9525) );
  AOI21_X1 U8446 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n6626), .A(n9525), .ZN(
        n6740) );
  INV_X1 U8447 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10058) );
  AOI22_X1 U8448 ( .A1(n6628), .A2(n10058), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n6745), .ZN(n6739) );
  NOR2_X1 U8449 ( .A1(n6740), .A2(n6739), .ZN(n6738) );
  AOI21_X1 U8450 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6628), .A(n6738), .ZN(
        n9473) );
  NAND2_X1 U8451 ( .A1(n6629), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6616) );
  OAI21_X1 U8452 ( .B1(n6629), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6616), .ZN(
        n9472) );
  NOR2_X1 U8453 ( .A1(n6669), .A2(n6670), .ZN(n6668) );
  NOR2_X1 U8454 ( .A1(n6678), .A2(n7071), .ZN(n6617) );
  NOR2_X1 U8455 ( .A1(n6668), .A2(n6617), .ZN(n9542) );
  NAND2_X1 U8456 ( .A1(n6634), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6618) );
  OAI21_X1 U8457 ( .B1(n6634), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6618), .ZN(
        n9541) );
  INV_X1 U8458 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U8459 ( .A1(n6638), .A2(n10200), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n9565), .ZN(n9555) );
  NAND2_X1 U8460 ( .A1(n6641), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6619) );
  OAI21_X1 U8461 ( .B1(n6641), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6619), .ZN(
        n9454) );
  NOR2_X1 U8462 ( .A1(n9453), .A2(n9454), .ZN(n9455) );
  NAND2_X1 U8463 ( .A1(n6644), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6620) );
  OAI21_X1 U8464 ( .B1(n6644), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6620), .ZN(
        n9490) );
  OAI21_X1 U8465 ( .B1(n6622), .B2(n6621), .A(n6995), .ZN(n6623) );
  NAND2_X1 U8466 ( .A1(n6647), .A2(n6663), .ZN(n8012) );
  INV_X1 U8467 ( .A(n9649), .ZN(n9116) );
  NAND2_X1 U8468 ( .A1(n6623), .A2(n9116), .ZN(n6654) );
  INV_X1 U8469 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9870) );
  AOI22_X1 U8470 ( .A1(n7000), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n9870), .B2(
        n6650), .ZN(n6646) );
  INV_X1 U8471 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9862) );
  MUX2_X1 U8472 ( .A(n9862), .B(P1_REG1_REG_4__SCAN_IN), .S(n6678), .Z(n6675)
         );
  NAND2_X1 U8473 ( .A1(n6629), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6631) );
  INV_X1 U8474 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6624) );
  AOI21_X1 U8475 ( .B1(n6626), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9531), .ZN(
        n6743) );
  NAND2_X1 U8476 ( .A1(n6628), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6627) );
  OAI21_X1 U8477 ( .B1(n6628), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6627), .ZN(
        n6742) );
  NOR2_X1 U8478 ( .A1(n6743), .A2(n6742), .ZN(n6741) );
  OR2_X1 U8479 ( .A1(n6629), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U8480 ( .A1(n6630), .A2(n6631), .ZN(n9477) );
  INV_X1 U8481 ( .A(n6678), .ZN(n6632) );
  NAND2_X1 U8482 ( .A1(n6632), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U8483 ( .A1(n6673), .A2(n6633), .ZN(n9546) );
  OR2_X1 U8484 ( .A1(n6634), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U8485 ( .A1(n6634), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6636) );
  AND2_X1 U8486 ( .A1(n6635), .A2(n6636), .ZN(n9547) );
  NAND2_X1 U8487 ( .A1(n9546), .A2(n9547), .ZN(n9545) );
  INV_X1 U8488 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6637) );
  MUX2_X1 U8489 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6637), .S(n9565), .Z(n9560)
         );
  OR2_X1 U8490 ( .A1(n6641), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U8491 ( .A1(n6641), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U8492 ( .A1(n6640), .A2(n6639), .ZN(n9459) );
  AOI21_X1 U8493 ( .B1(n6641), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9461), .ZN(
        n9495) );
  OR2_X1 U8494 ( .A1(n6644), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U8495 ( .A1(n6644), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U8496 ( .A1(n6643), .A2(n6642), .ZN(n9496) );
  OAI21_X1 U8497 ( .B1(n6646), .B2(n6645), .A(n6999), .ZN(n6652) );
  NAND2_X1 U8498 ( .A1(n9522), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U8499 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7424) );
  OAI211_X1 U8500 ( .C1(n9625), .C2(n6650), .A(n6649), .B(n7424), .ZN(n6651)
         );
  AOI21_X1 U8501 ( .B1(n6652), .B2(n9112), .A(n6651), .ZN(n6653) );
  NAND2_X1 U8502 ( .A1(n6654), .A2(n6653), .ZN(P1_U3252) );
  OAI21_X1 U8503 ( .B1(n6657), .B2(n6656), .A(n6655), .ZN(n6667) );
  NAND2_X1 U8504 ( .A1(n9012), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6819) );
  NAND2_X1 U8505 ( .A1(n6493), .A2(n9311), .ZN(n9757) );
  OAI22_X1 U8506 ( .A1(n9034), .A2(n9735), .B1(n9757), .B2(n8959), .ZN(n6658)
         );
  AOI21_X1 U8507 ( .B1(n6819), .B2(P1_REG3_REG_0__SCAN_IN), .A(n6658), .ZN(
        n6659) );
  OAI21_X1 U8508 ( .B1(n6667), .B2(n8999), .A(n6659), .ZN(P1_U3232) );
  NOR2_X1 U8509 ( .A1(n8323), .A2(P2_U3151), .ZN(n6737) );
  NAND2_X1 U8510 ( .A1(n6946), .A2(n6848), .ZN(n8076) );
  NAND2_X1 U8511 ( .A1(n6305), .A2(n8076), .ZN(n8035) );
  AOI22_X1 U8512 ( .A1(n6214), .A2(n8250), .B1(n8315), .B2(n8035), .ZN(n6661)
         );
  NAND2_X1 U8513 ( .A1(n8318), .A2(n6809), .ZN(n6660) );
  OAI211_X1 U8514 ( .C1(n6737), .C2(n6662), .A(n6661), .B(n6660), .ZN(P2_U3172) );
  NOR2_X1 U8515 ( .A1(n6663), .A2(n5737), .ZN(n6666) );
  INV_X2 U8516 ( .A(P1_U3973), .ZN(n9060) );
  OAI22_X1 U8517 ( .A1(n6664), .A2(P1_IR_REG_0__SCAN_IN), .B1(n9523), .B2(
        n8012), .ZN(n6665) );
  AOI211_X1 U8518 ( .C1(n6667), .C2(n6666), .A(n9060), .B(n6665), .ZN(n6748)
         );
  NAND2_X1 U8519 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6901) );
  INV_X1 U8520 ( .A(n6901), .ZN(n6672) );
  AOI211_X1 U8521 ( .C1(n6670), .C2(n6669), .A(n6668), .B(n9649), .ZN(n6671)
         );
  AOI211_X1 U8522 ( .C1(n9522), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n6672), .B(
        n6671), .ZN(n6677) );
  OAI211_X1 U8523 ( .C1(n6675), .C2(n6674), .A(n9112), .B(n6673), .ZN(n6676)
         );
  OAI211_X1 U8524 ( .C1(n9625), .C2(n6678), .A(n6677), .B(n6676), .ZN(n6679)
         );
  OR2_X1 U8525 ( .A1(n6748), .A2(n6679), .ZN(P1_U3247) );
  INV_X1 U8526 ( .A(n6680), .ZN(n6690) );
  AOI22_X1 U8527 ( .A1(n9609), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9431), .ZN(n6681) );
  OAI21_X1 U8528 ( .B1(n6690), .B2(n9436), .A(n6681), .ZN(P1_U3341) );
  OAI21_X1 U8529 ( .B1(n6684), .B2(n6683), .A(n6682), .ZN(n6685) );
  NAND2_X1 U8530 ( .A1(n6685), .A2(n8315), .ZN(n6688) );
  OAI22_X1 U8531 ( .A1(n8341), .A2(n4339), .B1(n4376), .B2(n8320), .ZN(n6686)
         );
  AOI21_X1 U8532 ( .B1(n8318), .B2(n8357), .A(n6686), .ZN(n6687) );
  OAI211_X1 U8533 ( .C1(n6737), .C2(n6689), .A(n6688), .B(n6687), .ZN(P2_U3162) );
  INV_X1 U8534 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6691) );
  INV_X1 U8535 ( .A(n8413), .ZN(n8431) );
  OAI222_X1 U8536 ( .A1(n8019), .A2(n6691), .B1(n8017), .B2(n6690), .C1(
        P2_U3151), .C2(n8431), .ZN(P2_U3281) );
  INV_X1 U8537 ( .A(n6762), .ZN(n6699) );
  MUX2_X1 U8538 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8503), .Z(n6697) );
  INV_X1 U8539 ( .A(n6697), .ZN(n6698) );
  INV_X1 U8540 ( .A(n9912), .ZN(n6696) );
  MUX2_X1 U8541 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8503), .Z(n6694) );
  INV_X1 U8542 ( .A(n6694), .ZN(n6695) );
  INV_X1 U8543 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6692) );
  OAI21_X1 U8544 ( .B1(n4592), .B2(n6693), .A(n9883), .ZN(n9909) );
  XOR2_X1 U8545 ( .A(n9912), .B(n6694), .Z(n9908) );
  NAND2_X1 U8546 ( .A1(n9909), .A2(n9908), .ZN(n9907) );
  OAI21_X1 U8547 ( .B1(n6696), .B2(n6695), .A(n9907), .ZN(n6751) );
  XNOR2_X1 U8548 ( .A(n6697), .B(n6762), .ZN(n6752) );
  NOR2_X1 U8549 ( .A1(n6751), .A2(n6752), .ZN(n6750) );
  MUX2_X1 U8550 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8503), .Z(n6789) );
  XOR2_X1 U8551 ( .A(n6799), .B(n6789), .Z(n6700) );
  NAND2_X1 U8552 ( .A1(n6701), .A2(n6700), .ZN(n6790) );
  OAI211_X1 U8553 ( .C1(n6701), .C2(n6700), .A(n6790), .B(n9906), .ZN(n6728)
         );
  NAND2_X1 U8554 ( .A1(n5799), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8555 ( .A1(n9917), .A2(n9916), .ZN(n9915) );
  NAND2_X1 U8556 ( .A1(n9912), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6704) );
  NAND2_X1 U8557 ( .A1(n9915), .A2(n6704), .ZN(n6705) );
  NAND2_X1 U8558 ( .A1(n6705), .A2(n6762), .ZN(n6707) );
  XNOR2_X1 U8559 ( .A(n6799), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6708) );
  AND3_X1 U8560 ( .A1(n6758), .A2(n6708), .A3(n6707), .ZN(n6709) );
  AND2_X1 U8561 ( .A1(n6723), .A2(n8530), .ZN(n9919) );
  OAI21_X1 U8562 ( .B1(n6797), .B2(n6709), .A(n9919), .ZN(n6710) );
  NAND2_X1 U8563 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U8564 ( .A1(n6710), .A2(n6889), .ZN(n6726) );
  AND2_X1 U8565 ( .A1(n6712), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U8566 ( .A1(n5799), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6715) );
  OAI21_X1 U8567 ( .B1(n6714), .B2(n6713), .A(n6715), .ZN(n9882) );
  OR2_X1 U8568 ( .A1(n9882), .A2(n6692), .ZN(n9880) );
  NAND2_X1 U8569 ( .A1(n9880), .A2(n6715), .ZN(n9901) );
  NAND2_X1 U8570 ( .A1(n9912), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U8571 ( .A1(n6717), .A2(n6762), .ZN(n6721) );
  OAI21_X1 U8572 ( .B1(n6717), .B2(n6762), .A(n6721), .ZN(n6753) );
  INV_X1 U8573 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10000) );
  NAND2_X1 U8574 ( .A1(n6755), .A2(n6721), .ZN(n6719) );
  INV_X1 U8575 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6718) );
  XNOR2_X1 U8576 ( .A(n6799), .B(n6718), .ZN(n6720) );
  NAND2_X1 U8577 ( .A1(n6719), .A2(n6720), .ZN(n6801) );
  INV_X1 U8578 ( .A(n6720), .ZN(n6722) );
  NAND3_X1 U8579 ( .A1(n6755), .A2(n6722), .A3(n6721), .ZN(n6724) );
  NAND2_X1 U8580 ( .A1(n6723), .A2(n8503), .ZN(n9889) );
  AOI21_X1 U8581 ( .B1(n6801), .B2(n6724), .A(n9889), .ZN(n6725) );
  AOI211_X1 U8582 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9905), .A(n6726), .B(
        n6725), .ZN(n6727) );
  OAI211_X1 U8583 ( .C1(n9913), .C2(n6799), .A(n6728), .B(n6727), .ZN(P2_U3186) );
  OAI21_X1 U8584 ( .B1(n6731), .B2(n6730), .A(n6729), .ZN(n6732) );
  NAND2_X1 U8585 ( .A1(n6732), .A2(n8315), .ZN(n6736) );
  OAI22_X1 U8586 ( .A1(n8341), .A2(n6733), .B1(n6303), .B2(n8320), .ZN(n6734)
         );
  AOI21_X1 U8587 ( .B1(n8318), .B2(n8356), .A(n6734), .ZN(n6735) );
  OAI211_X1 U8588 ( .C1(n6737), .C2(n5791), .A(n6736), .B(n6735), .ZN(P2_U3177) );
  AOI211_X1 U8589 ( .C1(n6740), .C2(n6739), .A(n6738), .B(n9649), .ZN(n6749)
         );
  AOI211_X1 U8590 ( .C1(n6743), .C2(n6742), .A(n6741), .B(n9644), .ZN(n6747)
         );
  AOI22_X1 U8591 ( .A1(n9522), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6744) );
  OAI21_X1 U8592 ( .B1(n6745), .B2(n9625), .A(n6744), .ZN(n6746) );
  OR4_X1 U8593 ( .A1(n6749), .A2(n6748), .A3(n6747), .A4(n6746), .ZN(P1_U3245)
         );
  AOI21_X1 U8594 ( .B1(n6752), .B2(n6751), .A(n6750), .ZN(n6766) );
  NAND2_X1 U8595 ( .A1(n6753), .A2(n10000), .ZN(n6754) );
  AND2_X1 U8596 ( .A1(n6755), .A2(n6754), .ZN(n6761) );
  NAND2_X1 U8597 ( .A1(n6756), .A2(n6984), .ZN(n6757) );
  NAND2_X1 U8598 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  NAND2_X1 U8599 ( .A1(n9919), .A2(n6759), .ZN(n6760) );
  NAND2_X1 U8600 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6825) );
  OAI211_X1 U8601 ( .C1(n6761), .C2(n9889), .A(n6760), .B(n6825), .ZN(n6764)
         );
  NOR2_X1 U8602 ( .A1(n9913), .A2(n6762), .ZN(n6763) );
  AOI211_X1 U8603 ( .C1(n9905), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6764), .B(
        n6763), .ZN(n6765) );
  OAI21_X1 U8604 ( .B1(n6766), .B2(n8509), .A(n6765), .ZN(P2_U3185) );
  INV_X1 U8605 ( .A(n6819), .ZN(n6774) );
  OAI21_X1 U8606 ( .B1(n6769), .B2(n6768), .A(n6767), .ZN(n6770) );
  NAND2_X1 U8607 ( .A1(n6770), .A2(n9021), .ZN(n6773) );
  INV_X1 U8608 ( .A(n7737), .ZN(n6771) );
  OAI22_X1 U8609 ( .A1(n6771), .A2(n9008), .B1(n6851), .B2(n9006), .ZN(n9731)
         );
  AOI22_X1 U8610 ( .A1(n9731), .A2(n9014), .B1(n9740), .B2(n5752), .ZN(n6772)
         );
  OAI211_X1 U8611 ( .C1(n6774), .C2(n5125), .A(n6773), .B(n6772), .ZN(P1_U3222) );
  INV_X1 U8612 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10170) );
  INV_X1 U8613 ( .A(n6775), .ZN(n6776) );
  INV_X1 U8614 ( .A(n9638), .ZN(n9079) );
  OAI222_X1 U8615 ( .A1(n9438), .A2(n10170), .B1(n9436), .B2(n6776), .C1(
        P1_U3086), .C2(n9079), .ZN(P1_U3340) );
  INV_X1 U8616 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6777) );
  INV_X1 U8617 ( .A(n8455), .ZN(n8432) );
  OAI222_X1 U8618 ( .A1(n8019), .A2(n6777), .B1(n8017), .B2(n6776), .C1(
        P2_U3151), .C2(n8432), .ZN(P2_U3280) );
  XNOR2_X1 U8619 ( .A(n6778), .B(n7949), .ZN(n6779) );
  OAI222_X1 U8620 ( .A1(n9006), .A2(n6816), .B1(n9008), .B2(n6815), .C1(n6779), 
        .C2(n9759), .ZN(n9775) );
  INV_X1 U8621 ( .A(n9775), .ZN(n6788) );
  XNOR2_X1 U8622 ( .A(n7949), .B(n6780), .ZN(n9777) );
  INV_X1 U8623 ( .A(n9733), .ZN(n6781) );
  OAI211_X1 U8624 ( .C1(n6781), .C2(n9774), .A(n9734), .B(n6923), .ZN(n9773)
         );
  INV_X1 U8625 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6782) );
  OAI22_X1 U8626 ( .A1(n9752), .A2(n10058), .B1(n6782), .B2(n9315), .ZN(n6783)
         );
  AOI21_X1 U8627 ( .B1(n9739), .B2(n6784), .A(n6783), .ZN(n6785) );
  OAI21_X1 U8628 ( .B1(n9694), .B2(n9773), .A(n6785), .ZN(n6786) );
  AOI21_X1 U8629 ( .B1(n9777), .B2(n9715), .A(n6786), .ZN(n6787) );
  OAI21_X1 U8630 ( .B1(n6788), .B2(n9754), .A(n6787), .ZN(P1_U3291) );
  INV_X1 U8631 ( .A(n6799), .ZN(n6792) );
  INV_X1 U8632 ( .A(n6789), .ZN(n6791) );
  OAI21_X1 U8633 ( .B1(n6792), .B2(n6791), .A(n6790), .ZN(n6796) );
  MUX2_X1 U8634 ( .A(n6794), .B(n6793), .S(n8503), .Z(n6860) );
  XNOR2_X1 U8635 ( .A(n6860), .B(n6869), .ZN(n6795) );
  NAND2_X1 U8636 ( .A1(n6796), .A2(n6795), .ZN(n6859) );
  OAI211_X1 U8637 ( .C1(n6796), .C2(n6795), .A(n6859), .B(n9906), .ZN(n6808)
         );
  AOI21_X1 U8638 ( .B1(n6794), .B2(n6798), .A(n6866), .ZN(n6805) );
  NAND2_X1 U8639 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U8640 ( .A1(n6799), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U8641 ( .A1(n6801), .A2(n6800), .ZN(n6870) );
  NOR2_X1 U8642 ( .A1(n6802), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6803) );
  INV_X1 U8643 ( .A(n9889), .ZN(n9904) );
  OAI21_X1 U8644 ( .B1(n6872), .B2(n6803), .A(n9904), .ZN(n6804) );
  OAI211_X1 U8645 ( .C1(n9896), .C2(n6805), .A(n6911), .B(n6804), .ZN(n6806)
         );
  AOI21_X1 U8646 ( .B1(n9905), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6806), .ZN(
        n6807) );
  OAI211_X1 U8647 ( .C1(n9913), .C2(n6869), .A(n6808), .B(n6807), .ZN(P2_U3187) );
  INV_X1 U8648 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6812) );
  OAI21_X1 U8649 ( .B1(n9994), .B2(n9928), .A(n8035), .ZN(n6810) );
  NAND2_X1 U8650 ( .A1(n6809), .A2(n9930), .ZN(n6842) );
  OAI211_X1 U8651 ( .C1(n9989), .C2(n6848), .A(n6810), .B(n6842), .ZN(n6830)
         );
  NAND2_X1 U8652 ( .A1(n9995), .A2(n6830), .ZN(n6811) );
  OAI21_X1 U8653 ( .B1(n9995), .B2(n6812), .A(n6811), .ZN(P2_U3390) );
  XOR2_X1 U8654 ( .A(n6813), .B(n6814), .Z(n6821) );
  NAND2_X1 U8655 ( .A1(n9014), .A2(n9309), .ZN(n9025) );
  OAI22_X1 U8656 ( .A1(n9025), .A2(n6815), .B1(n9034), .B2(n9774), .ZN(n6818)
         );
  NOR2_X1 U8657 ( .A1(n8959), .A2(n9006), .ZN(n8993) );
  INV_X1 U8658 ( .A(n8993), .ZN(n9027) );
  NOR2_X1 U8659 ( .A1(n9027), .A2(n6816), .ZN(n6817) );
  AOI211_X1 U8660 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n6819), .A(n6818), .B(
        n6817), .ZN(n6820) );
  OAI21_X1 U8661 ( .B1(n6821), .B2(n8999), .A(n6820), .ZN(P1_U3237) );
  AOI21_X1 U8662 ( .B1(n6822), .B2(n6823), .A(n8327), .ZN(n6824) );
  OR2_X1 U8663 ( .A1(n6822), .A2(n6823), .ZN(n6885) );
  NAND2_X1 U8664 ( .A1(n6824), .A2(n6885), .ZN(n6829) );
  INV_X1 U8665 ( .A(n6825), .ZN(n6827) );
  OAI22_X1 U8666 ( .A1(n8335), .A2(n6312), .B1(n4615), .B2(n8320), .ZN(n6826)
         );
  AOI211_X1 U8667 ( .C1(n6986), .C2(n8250), .A(n6827), .B(n6826), .ZN(n6828)
         );
  OAI211_X1 U8668 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8333), .A(n6829), .B(
        n6828), .ZN(P2_U3158) );
  NAND2_X1 U8669 ( .A1(n6830), .A2(n10008), .ZN(n6831) );
  OAI21_X1 U8670 ( .B1(n10008), .B2(n6832), .A(n6831), .ZN(P2_U3459) );
  NAND2_X1 U8671 ( .A1(n6833), .A2(n6293), .ZN(n6834) );
  AND2_X1 U8672 ( .A1(n6835), .A2(n6834), .ZN(n6838) );
  INV_X1 U8673 ( .A(n6836), .ZN(n6837) );
  NAND2_X1 U8674 ( .A1(n6838), .A2(n6837), .ZN(n6843) );
  INV_X1 U8675 ( .A(n6843), .ZN(n6839) );
  INV_X1 U8676 ( .A(n8709), .ZN(n8728) );
  INV_X1 U8677 ( .A(n8035), .ZN(n6841) );
  NOR3_X1 U8678 ( .A1(n6841), .A2(n9987), .A3(n6840), .ZN(n6845) );
  INV_X1 U8679 ( .A(n6842), .ZN(n6844) );
  NAND2_X2 U8680 ( .A1(n6843), .A2(n9936), .ZN(n8733) );
  OAI21_X1 U8681 ( .B1(n6845), .B2(n6844), .A(n8733), .ZN(n6847) );
  AOI22_X1 U8682 ( .A1(n8713), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n8729), .ZN(n6846) );
  OAI211_X1 U8683 ( .C1(n9939), .C2(n6848), .A(n6847), .B(n6846), .ZN(P2_U3233) );
  XOR2_X1 U8684 ( .A(n6849), .B(n6850), .Z(n6854) );
  OAI22_X1 U8685 ( .A1(n7081), .A2(n9006), .B1(n6851), .B2(n9008), .ZN(n6918)
         );
  AOI22_X1 U8686 ( .A1(n6918), .A2(n9014), .B1(n6926), .B2(n5752), .ZN(n6853)
         );
  MUX2_X1 U8687 ( .A(P1_STATE_REG_SCAN_IN), .B(n9012), .S(n6925), .Z(n6852) );
  OAI211_X1 U8688 ( .C1(n6854), .C2(n8999), .A(n6853), .B(n6852), .ZN(P1_U3218) );
  INV_X1 U8689 ( .A(n6855), .ZN(n6857) );
  INV_X1 U8690 ( .A(n8450), .ZN(n8471) );
  OAI222_X1 U8691 ( .A1(n8019), .A2(n6856), .B1(n8017), .B2(n6857), .C1(n8471), 
        .C2(P2_U3151), .ZN(P2_U3279) );
  INV_X1 U8692 ( .A(n9095), .ZN(n9074) );
  OAI222_X1 U8693 ( .A1(n9438), .A2(n6858), .B1(n9074), .B2(P1_U3086), .C1(
        n9436), .C2(n6857), .ZN(P1_U3339) );
  MUX2_X1 U8694 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8503), .Z(n7033) );
  XNOR2_X1 U8695 ( .A(n7033), .B(n7043), .ZN(n6863) );
  OAI21_X1 U8696 ( .B1(n6861), .B2(n6860), .A(n6859), .ZN(n6862) );
  NOR2_X1 U8697 ( .A1(n6862), .A2(n6863), .ZN(n7034) );
  AOI21_X1 U8698 ( .B1(n6863), .B2(n6862), .A(n7034), .ZN(n6880) );
  INV_X1 U8699 ( .A(n7043), .ZN(n7036) );
  INV_X1 U8700 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6865) );
  NOR2_X1 U8701 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4581), .ZN(n6937) );
  INV_X1 U8702 ( .A(n6937), .ZN(n6864) );
  OAI21_X1 U8703 ( .B1(n9899), .B2(n6865), .A(n6864), .ZN(n6878) );
  NAND2_X1 U8704 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n7043), .ZN(n6867) );
  OAI21_X1 U8705 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7043), .A(n6867), .ZN(
        n6868) );
  AOI21_X1 U8706 ( .B1(n4445), .B2(n6868), .A(n7042), .ZN(n6876) );
  NAND2_X1 U8707 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n7043), .ZN(n6873) );
  OAI21_X1 U8708 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n7043), .A(n6873), .ZN(
        n6874) );
  AOI21_X1 U8709 ( .B1(n4441), .B2(n6874), .A(n7038), .ZN(n6875) );
  OAI22_X1 U8710 ( .A1(n9896), .A2(n6876), .B1(n6875), .B2(n9889), .ZN(n6877)
         );
  AOI211_X1 U8711 ( .C1(n7036), .C2(n9891), .A(n6878), .B(n6877), .ZN(n6879)
         );
  OAI21_X1 U8712 ( .B1(n6880), .B2(n8509), .A(n6879), .ZN(P2_U3188) );
  AND2_X1 U8713 ( .A1(n6881), .A2(n6885), .ZN(n6887) );
  AND2_X1 U8714 ( .A1(n6315), .A2(n6882), .ZN(n6886) );
  INV_X1 U8715 ( .A(n6883), .ZN(n6884) );
  NAND2_X1 U8716 ( .A1(n6885), .A2(n6884), .ZN(n6905) );
  OAI21_X1 U8717 ( .B1(n6887), .B2(n6886), .A(n6905), .ZN(n6888) );
  NAND2_X1 U8718 ( .A1(n6888), .A2(n8315), .ZN(n6893) );
  INV_X1 U8719 ( .A(n6889), .ZN(n6891) );
  OAI22_X1 U8720 ( .A1(n8335), .A2(n6963), .B1(n8719), .B2(n8320), .ZN(n6890)
         );
  AOI211_X1 U8721 ( .C1(n8100), .C2(n8250), .A(n6891), .B(n6890), .ZN(n6892)
         );
  OAI211_X1 U8722 ( .C1(n7104), .C2(n8333), .A(n6893), .B(n6892), .ZN(P2_U3170) );
  INV_X1 U8723 ( .A(n6894), .ZN(n7072) );
  AOI21_X1 U8724 ( .B1(n6896), .B2(n6895), .A(n8999), .ZN(n6898) );
  NAND2_X1 U8725 ( .A1(n6898), .A2(n6897), .ZN(n6904) );
  NAND2_X1 U8726 ( .A1(n9058), .A2(n9309), .ZN(n6900) );
  NAND2_X1 U8727 ( .A1(n9056), .A2(n9311), .ZN(n6899) );
  NAND2_X1 U8728 ( .A1(n6900), .A2(n6899), .ZN(n7069) );
  OAI21_X1 U8729 ( .B1(n9034), .B2(n7073), .A(n6901), .ZN(n6902) );
  AOI21_X1 U8730 ( .B1(n9014), .B2(n7069), .A(n6902), .ZN(n6903) );
  OAI211_X1 U8731 ( .C1(n9012), .C2(n7072), .A(n6904), .B(n6903), .ZN(P1_U3230) );
  INV_X1 U8732 ( .A(n6905), .ZN(n6907) );
  NOR3_X1 U8733 ( .A1(n6907), .A2(n6309), .A3(n6906), .ZN(n6910) );
  INV_X1 U8734 ( .A(n6908), .ZN(n6909) );
  OAI21_X1 U8735 ( .B1(n6910), .B2(n6909), .A(n8315), .ZN(n6916) );
  INV_X1 U8736 ( .A(n6911), .ZN(n6913) );
  OAI22_X1 U8737 ( .A1(n8335), .A2(n9924), .B1(n6312), .B2(n8320), .ZN(n6912)
         );
  AOI211_X1 U8738 ( .C1(n6914), .C2(n8250), .A(n6913), .B(n6912), .ZN(n6915)
         );
  OAI211_X1 U8739 ( .C1(n7100), .C2(n8333), .A(n6916), .B(n6915), .ZN(P2_U3167) );
  XNOR2_X1 U8740 ( .A(n6917), .B(n6922), .ZN(n6920) );
  INV_X1 U8741 ( .A(n6918), .ZN(n6919) );
  OAI21_X1 U8742 ( .B1(n6920), .B2(n9759), .A(n6919), .ZN(n9781) );
  INV_X1 U8743 ( .A(n9781), .ZN(n6931) );
  XNOR2_X1 U8744 ( .A(n6921), .B(n6922), .ZN(n9783) );
  INV_X1 U8745 ( .A(n6923), .ZN(n6924) );
  OAI211_X1 U8746 ( .C1(n9780), .C2(n6924), .A(n4439), .B(n9734), .ZN(n9779)
         );
  AOI22_X1 U8747 ( .A1(n9754), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9749), .B2(
        n6925), .ZN(n6928) );
  NAND2_X1 U8748 ( .A1(n9739), .A2(n6926), .ZN(n6927) );
  OAI211_X1 U8749 ( .C1(n9779), .C2(n9694), .A(n6928), .B(n6927), .ZN(n6929)
         );
  AOI21_X1 U8750 ( .B1(n9783), .B2(n9715), .A(n6929), .ZN(n6930) );
  OAI21_X1 U8751 ( .B1(n6931), .B2(n9754), .A(n6930), .ZN(P1_U3290) );
  AOI21_X1 U8752 ( .B1(n6933), .B2(n6932), .A(n8327), .ZN(n6935) );
  NAND2_X1 U8753 ( .A1(n6935), .A2(n6934), .ZN(n6939) );
  OAI22_X1 U8754 ( .A1(n8335), .A2(n7141), .B1(n6963), .B2(n8320), .ZN(n6936)
         );
  AOI211_X1 U8755 ( .C1(n9967), .C2(n8250), .A(n6937), .B(n6936), .ZN(n6938)
         );
  OAI211_X1 U8756 ( .C1(n9937), .C2(n8333), .A(n6939), .B(n6938), .ZN(P2_U3179) );
  INV_X1 U8757 ( .A(n6940), .ZN(n6942) );
  INV_X1 U8758 ( .A(n9110), .ZN(n9104) );
  OAI222_X1 U8759 ( .A1(n9438), .A2(n6941), .B1(n9436), .B2(n6942), .C1(
        P1_U3086), .C2(n9104), .ZN(P1_U3338) );
  INV_X1 U8760 ( .A(n8501), .ZN(n8480) );
  OAI222_X1 U8761 ( .A1(n8019), .A2(n6943), .B1(n8017), .B2(n6942), .C1(
        P2_U3151), .C2(n8480), .ZN(P2_U3278) );
  AND2_X1 U8762 ( .A1(n6296), .A2(n8222), .ZN(n7090) );
  INV_X1 U8763 ( .A(n6944), .ZN(n6945) );
  AOI21_X1 U8764 ( .B1(n6305), .B2(n6213), .A(n6945), .ZN(n9944) );
  INV_X1 U8765 ( .A(n9944), .ZN(n6953) );
  NOR2_X1 U8766 ( .A1(n9936), .A2(n6689), .ZN(n6952) );
  AOI22_X1 U8767 ( .A1(n9933), .A2(n6946), .B1(n8357), .B2(n9930), .ZN(n6951)
         );
  OAI21_X1 U8768 ( .B1(n6948), .B2(n6213), .A(n6947), .ZN(n6949) );
  NAND2_X1 U8769 ( .A1(n6949), .A2(n9928), .ZN(n6950) );
  OAI211_X1 U8770 ( .C1(n9944), .C2(n8717), .A(n6951), .B(n6950), .ZN(n9946)
         );
  AOI211_X1 U8771 ( .C1(n7090), .C2(n6953), .A(n6952), .B(n9946), .ZN(n6954)
         );
  MUX2_X1 U8772 ( .A(n6955), .B(n6954), .S(n8733), .Z(n6956) );
  OAI21_X1 U8773 ( .B1(n4339), .B2(n9939), .A(n6956), .ZN(P2_U3232) );
  INV_X1 U8774 ( .A(n8037), .ZN(n8088) );
  NAND3_X1 U8775 ( .A1(n6957), .A2(n8088), .A3(n8097), .ZN(n6958) );
  NAND2_X1 U8776 ( .A1(n6959), .A2(n6958), .ZN(n7109) );
  NAND2_X1 U8777 ( .A1(n7092), .A2(n6960), .ZN(n6961) );
  XNOR2_X1 U8778 ( .A(n6961), .B(n8037), .ZN(n6962) );
  OAI222_X1 U8779 ( .A1(n8718), .A2(n6963), .B1(n8720), .B2(n8719), .C1(n6962), 
        .C2(n6157), .ZN(n7106) );
  AOI21_X1 U8780 ( .B1(n9994), .B2(n7109), .A(n7106), .ZN(n6991) );
  AOI22_X1 U8781 ( .A1(n8854), .A2(n8100), .B1(n9997), .B2(
        P2_REG0_REG_4__SCAN_IN), .ZN(n6964) );
  OAI21_X1 U8782 ( .B1(n6991), .B2(n9997), .A(n6964), .ZN(P2_U3402) );
  XNOR2_X1 U8783 ( .A(n6965), .B(n6970), .ZN(n6966) );
  NAND2_X1 U8784 ( .A1(n6966), .A2(n9702), .ZN(n6968) );
  AOI22_X1 U8785 ( .A1(n9309), .A2(n9057), .B1(n9055), .B2(n9311), .ZN(n6967)
         );
  NAND2_X1 U8786 ( .A1(n6968), .A2(n6967), .ZN(n9796) );
  INV_X1 U8787 ( .A(n9796), .ZN(n6976) );
  XNOR2_X1 U8788 ( .A(n6970), .B(n6969), .ZN(n9798) );
  OAI211_X1 U8789 ( .C1(n4365), .C2(n9795), .A(n9734), .B(n7252), .ZN(n9794)
         );
  AOI22_X1 U8790 ( .A1(n9754), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7084), .B2(
        n9749), .ZN(n6973) );
  NAND2_X1 U8791 ( .A1(n9739), .A2(n6971), .ZN(n6972) );
  OAI211_X1 U8792 ( .C1(n9794), .C2(n9694), .A(n6973), .B(n6972), .ZN(n6974)
         );
  AOI21_X1 U8793 ( .B1(n9798), .B2(n9715), .A(n6974), .ZN(n6975) );
  OAI21_X1 U8794 ( .B1(n6976), .B2(n9754), .A(n6975), .ZN(P1_U3288) );
  INV_X1 U8795 ( .A(n8086), .ZN(n6977) );
  NOR2_X1 U8796 ( .A1(n8038), .A2(n6977), .ZN(n6980) );
  INV_X1 U8797 ( .A(n6957), .ZN(n6979) );
  AOI21_X1 U8798 ( .B1(n6980), .B2(n6978), .A(n6979), .ZN(n9955) );
  INV_X1 U8799 ( .A(n7090), .ZN(n8731) );
  NAND2_X1 U8800 ( .A1(n8717), .A2(n8731), .ZN(n6981) );
  XOR2_X1 U8801 ( .A(n8038), .B(n6982), .Z(n6983) );
  AOI222_X1 U8802 ( .A1(n9928), .A2(n6983), .B1(n8355), .B2(n9930), .C1(n8357), 
        .C2(n9933), .ZN(n9953) );
  MUX2_X1 U8803 ( .A(n6984), .B(n9953), .S(n8733), .Z(n6988) );
  AOI22_X1 U8804 ( .A1(n8705), .A2(n6986), .B1(n8729), .B2(n6985), .ZN(n6987)
         );
  OAI211_X1 U8805 ( .C1(n9955), .C2(n9943), .A(n6988), .B(n6987), .ZN(P2_U3230) );
  OAI22_X1 U8806 ( .A1(n8737), .A2(n7105), .B1(n10008), .B2(n6718), .ZN(n6989)
         );
  INV_X1 U8807 ( .A(n6989), .ZN(n6990) );
  OAI21_X1 U8808 ( .B1(n6991), .B2(n6287), .A(n6990), .ZN(P2_U3463) );
  NOR2_X1 U8809 ( .A1(n9077), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6992) );
  AOI21_X1 U8810 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9077), .A(n6992), .ZN(
        n6997) );
  INV_X1 U8811 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6993) );
  NAND2_X1 U8812 ( .A1(n9449), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6994) );
  OAI21_X1 U8813 ( .B1(n9449), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6994), .ZN(
        n9445) );
  OAI21_X1 U8814 ( .B1(n7000), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6995), .ZN(
        n9446) );
  NOR2_X1 U8815 ( .A1(n9445), .A2(n9446), .ZN(n9444) );
  AOI21_X1 U8816 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9449), .A(n9444), .ZN(
        n9571) );
  NAND2_X1 U8817 ( .A1(n6997), .A2(n6996), .ZN(n9076) );
  OAI21_X1 U8818 ( .B1(n6997), .B2(n6996), .A(n9076), .ZN(n7007) );
  INV_X1 U8819 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9873) );
  MUX2_X1 U8820 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9873), .S(n9570), .Z(n9575)
         );
  NAND2_X1 U8821 ( .A1(n9449), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7002) );
  INV_X1 U8822 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6998) );
  MUX2_X1 U8823 ( .A(n6998), .B(P1_REG1_REG_10__SCAN_IN), .S(n9449), .Z(n9442)
         );
  NOR2_X1 U8824 ( .A1(n9442), .A2(n9443), .ZN(n9441) );
  INV_X1 U8825 ( .A(n9441), .ZN(n7001) );
  NAND2_X1 U8826 ( .A1(n7002), .A2(n7001), .ZN(n9576) );
  NAND2_X1 U8827 ( .A1(n9575), .A2(n9576), .ZN(n9580) );
  INV_X1 U8828 ( .A(n9580), .ZN(n7003) );
  AOI21_X1 U8829 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9570), .A(n7003), .ZN(
        n7005) );
  INV_X1 U8830 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9875) );
  AOI22_X1 U8831 ( .A1(n9077), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9875), .B2(
        n7011), .ZN(n7004) );
  OAI21_X1 U8832 ( .B1(n7005), .B2(n7004), .A(n9062), .ZN(n7006) );
  AOI22_X1 U8833 ( .A1(n9116), .A2(n7007), .B1(n9112), .B2(n7006), .ZN(n7010)
         );
  NAND2_X1 U8834 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7466) );
  INV_X1 U8835 ( .A(n7466), .ZN(n7008) );
  AOI21_X1 U8836 ( .B1(n9522), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7008), .ZN(
        n7009) );
  OAI211_X1 U8837 ( .C1(n7011), .C2(n9625), .A(n7010), .B(n7009), .ZN(P1_U3255) );
  INV_X1 U8838 ( .A(n7012), .ZN(n7064) );
  AOI22_X1 U8839 ( .A1(n9654), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9431), .ZN(n7013) );
  OAI21_X1 U8840 ( .B1(n7064), .B2(n9436), .A(n7013), .ZN(P1_U3337) );
  INV_X1 U8841 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10015) );
  NOR2_X1 U8842 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7014) );
  AOI21_X1 U8843 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7014), .ZN(n10021) );
  NOR2_X1 U8844 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7015) );
  AOI21_X1 U8845 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7015), .ZN(n10024) );
  NOR2_X1 U8846 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7016) );
  AOI21_X1 U8847 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7016), .ZN(n10027) );
  NOR2_X1 U8848 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7017) );
  AOI21_X1 U8849 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7017), .ZN(n10030) );
  NOR2_X1 U8850 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7018) );
  AOI21_X1 U8851 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7018), .ZN(n10033) );
  INV_X1 U8852 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10196) );
  INV_X1 U8853 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7482) );
  AOI22_X1 U8854 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .B1(n10196), .B2(n7482), .ZN(n10036) );
  NOR2_X1 U8855 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7019) );
  AOI21_X1 U8856 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7019), .ZN(n10039) );
  NOR2_X1 U8857 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7020) );
  AOI21_X1 U8858 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7020), .ZN(n10042) );
  NOR2_X1 U8859 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7021) );
  AOI21_X1 U8860 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7021), .ZN(n10241) );
  NOR2_X1 U8861 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P2_ADDR_REG_8__SCAN_IN), 
        .ZN(n7022) );
  AOI21_X1 U8862 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n7022), .ZN(n10250) );
  NOR2_X1 U8863 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7023) );
  AOI21_X1 U8864 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7023), .ZN(n10247) );
  NOR2_X1 U8865 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n7024) );
  AOI21_X1 U8866 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n7024), .ZN(n10244) );
  NOR2_X1 U8867 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n7025) );
  AOI21_X1 U8868 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n7025), .ZN(n10238) );
  AND2_X1 U8869 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7026) );
  NOR2_X1 U8870 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7026), .ZN(n10010) );
  INV_X1 U8871 ( .A(n10010), .ZN(n10011) );
  INV_X1 U8872 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10013) );
  NAND3_X1 U8873 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U8874 ( .A1(n10013), .A2(n10012), .ZN(n10009) );
  NAND2_X1 U8875 ( .A1(n10011), .A2(n10009), .ZN(n10253) );
  NAND2_X1 U8876 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7027) );
  OAI21_X1 U8877 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7027), .ZN(n10252) );
  NOR2_X1 U8878 ( .A1(n10253), .A2(n10252), .ZN(n10251) );
  AOI21_X1 U8879 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10251), .ZN(n10256) );
  NAND2_X1 U8880 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7028) );
  OAI21_X1 U8881 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7028), .ZN(n10255) );
  NOR2_X1 U8882 ( .A1(n10256), .A2(n10255), .ZN(n10254) );
  AOI21_X1 U8883 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10254), .ZN(n10259) );
  NOR2_X1 U8884 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7029) );
  AOI21_X1 U8885 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7029), .ZN(n10258) );
  NAND2_X1 U8886 ( .A1(n10259), .A2(n10258), .ZN(n10257) );
  OAI21_X1 U8887 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10257), .ZN(n10237) );
  NAND2_X1 U8888 ( .A1(n10238), .A2(n10237), .ZN(n10236) );
  OAI21_X1 U8889 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10236), .ZN(n10243) );
  NAND2_X1 U8890 ( .A1(n10244), .A2(n10243), .ZN(n10242) );
  OAI21_X1 U8891 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10242), .ZN(n10246) );
  NAND2_X1 U8892 ( .A1(n10247), .A2(n10246), .ZN(n10245) );
  OAI21_X1 U8893 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10245), .ZN(n10249) );
  NAND2_X1 U8894 ( .A1(n10250), .A2(n10249), .ZN(n10248) );
  OAI21_X1 U8895 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10248), .ZN(n10240) );
  NAND2_X1 U8896 ( .A1(n10241), .A2(n10240), .ZN(n10239) );
  OAI21_X1 U8897 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10239), .ZN(n10041) );
  NAND2_X1 U8898 ( .A1(n10042), .A2(n10041), .ZN(n10040) );
  OAI21_X1 U8899 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10040), .ZN(n10038) );
  NAND2_X1 U8900 ( .A1(n10039), .A2(n10038), .ZN(n10037) );
  OAI21_X1 U8901 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10037), .ZN(n10035) );
  NAND2_X1 U8902 ( .A1(n10036), .A2(n10035), .ZN(n10034) );
  OAI21_X1 U8903 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10034), .ZN(n10032) );
  NAND2_X1 U8904 ( .A1(n10033), .A2(n10032), .ZN(n10031) );
  OAI21_X1 U8905 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10031), .ZN(n10029) );
  NAND2_X1 U8906 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  OAI21_X1 U8907 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10028), .ZN(n10026) );
  NAND2_X1 U8908 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  OAI21_X1 U8909 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10025), .ZN(n10023) );
  NAND2_X1 U8910 ( .A1(n10024), .A2(n10023), .ZN(n10022) );
  OAI21_X1 U8911 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10022), .ZN(n10020) );
  NAND2_X1 U8912 ( .A1(n10021), .A2(n10020), .ZN(n10019) );
  OAI21_X1 U8913 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10019), .ZN(n10016) );
  NAND2_X1 U8914 ( .A1(n10015), .A2(n10016), .ZN(n7030) );
  NOR2_X1 U8915 ( .A1(n10015), .A2(n10016), .ZN(n10014) );
  AOI21_X1 U8916 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7030), .A(n10014), .ZN(
        n7032) );
  XNOR2_X1 U8917 ( .A(n9122), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7031) );
  XNOR2_X1 U8918 ( .A(n7032), .B(n7031), .ZN(ADD_1068_U4) );
  INV_X1 U8919 ( .A(n7033), .ZN(n7035) );
  MUX2_X1 U8920 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8503), .Z(n7117) );
  XNOR2_X1 U8921 ( .A(n7117), .B(n7116), .ZN(n7118) );
  XNOR2_X1 U8922 ( .A(n7119), .B(n7118), .ZN(n7037) );
  NAND2_X1 U8923 ( .A1(n7037), .A2(n9906), .ZN(n7053) );
  AOI21_X1 U8924 ( .B1(n7043), .B2(P2_REG1_REG_6__SCAN_IN), .A(n7038), .ZN(
        n7039) );
  INV_X1 U8925 ( .A(n7116), .ZN(n7044) );
  AOI21_X1 U8926 ( .B1(n4975), .B2(n5864), .A(n4438), .ZN(n7041) );
  NOR2_X1 U8927 ( .A1(n9889), .A2(n7041), .ZN(n7051) );
  NOR2_X1 U8928 ( .A1(n7045), .A2(n7044), .ZN(n7112) );
  INV_X1 U8929 ( .A(n7112), .ZN(n7047) );
  NOR2_X1 U8930 ( .A1(n5869), .A2(n7048), .ZN(n7111) );
  AOI21_X1 U8931 ( .B1(n7048), .B2(n5869), .A(n7111), .ZN(n7049) );
  NAND2_X1 U8932 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7058) );
  OAI21_X1 U8933 ( .B1(n9896), .B2(n7049), .A(n7058), .ZN(n7050) );
  AOI211_X1 U8934 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9905), .A(n7051), .B(
        n7050), .ZN(n7052) );
  OAI211_X1 U8935 ( .C1(n9913), .C2(n7116), .A(n7053), .B(n7052), .ZN(P2_U3189) );
  OAI21_X1 U8936 ( .B1(n7056), .B2(n7055), .A(n7054), .ZN(n7057) );
  NAND2_X1 U8937 ( .A1(n7057), .A2(n8315), .ZN(n7062) );
  INV_X1 U8938 ( .A(n7058), .ZN(n7060) );
  OAI22_X1 U8939 ( .A1(n8335), .A2(n7136), .B1(n9924), .B2(n8320), .ZN(n7059)
         );
  AOI211_X1 U8940 ( .C1(n7216), .C2(n8250), .A(n7060), .B(n7059), .ZN(n7061)
         );
  OAI211_X1 U8941 ( .C1(n7214), .C2(n8333), .A(n7062), .B(n7061), .ZN(P2_U3153) );
  OAI222_X1 U8942 ( .A1(P2_U3151), .A2(n8511), .B1(n8017), .B2(n7064), .C1(
        n7063), .C2(n8019), .ZN(P2_U3277) );
  XOR2_X1 U8943 ( .A(n7065), .B(n7950), .Z(n9790) );
  INV_X1 U8944 ( .A(n7813), .ZN(n7068) );
  NOR2_X1 U8945 ( .A1(n7066), .A2(n7812), .ZN(n7067) );
  AOI211_X1 U8946 ( .C1(n7068), .C2(n7950), .A(n9759), .B(n7067), .ZN(n7070)
         );
  NOR2_X1 U8947 ( .A1(n7070), .A2(n7069), .ZN(n9789) );
  MUX2_X1 U8948 ( .A(n7071), .B(n9789), .S(n9752), .Z(n7076) );
  AOI211_X1 U8949 ( .C1(n9786), .C2(n4439), .A(n9246), .B(n4365), .ZN(n9785)
         );
  OAI22_X1 U8950 ( .A1(n9720), .A2(n7073), .B1(n7072), .B2(n9315), .ZN(n7074)
         );
  AOI21_X1 U8951 ( .B1(n9785), .B2(n9738), .A(n7074), .ZN(n7075) );
  OAI211_X1 U8952 ( .C1(n9307), .C2(n9790), .A(n7076), .B(n7075), .ZN(P1_U3289) );
  NAND2_X1 U8953 ( .A1(n7078), .A2(n7077), .ZN(n7079) );
  XOR2_X1 U8954 ( .A(n7080), .B(n7079), .Z(n7086) );
  INV_X1 U8955 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10059) );
  OAI22_X1 U8956 ( .A1(n9034), .A2(n9795), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10059), .ZN(n7083) );
  OAI22_X1 U8957 ( .A1(n9027), .A2(n7165), .B1(n7081), .B2(n9025), .ZN(n7082)
         );
  AOI211_X1 U8958 ( .C1(n7084), .C2(n9030), .A(n7083), .B(n7082), .ZN(n7085)
         );
  OAI21_X1 U8959 ( .B1(n7086), .B2(n8999), .A(n7085), .ZN(P1_U3227) );
  NAND2_X1 U8960 ( .A1(n7088), .A2(n7087), .ZN(n7095) );
  XOR2_X1 U8961 ( .A(n7095), .B(n7089), .Z(n9960) );
  NAND2_X1 U8962 ( .A1(n8733), .A2(n7090), .ZN(n7694) );
  NAND2_X1 U8963 ( .A1(n7092), .A2(n7091), .ZN(n7094) );
  NAND2_X1 U8964 ( .A1(n7094), .A2(n7093), .ZN(n7096) );
  XNOR2_X1 U8965 ( .A(n7096), .B(n7095), .ZN(n7098) );
  OAI22_X1 U8966 ( .A1(n6312), .A2(n8720), .B1(n9924), .B2(n8718), .ZN(n7097)
         );
  AOI21_X1 U8967 ( .B1(n7098), .B2(n9928), .A(n7097), .ZN(n7099) );
  OAI21_X1 U8968 ( .B1(n9960), .B2(n8717), .A(n7099), .ZN(n9962) );
  NAND2_X1 U8969 ( .A1(n9962), .A2(n8733), .ZN(n7103) );
  OAI22_X1 U8970 ( .A1(n9939), .A2(n9959), .B1(n7100), .B2(n9936), .ZN(n7101)
         );
  AOI21_X1 U8971 ( .B1(n8713), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7101), .ZN(
        n7102) );
  OAI211_X1 U8972 ( .C1(n9960), .C2(n7694), .A(n7103), .B(n7102), .ZN(P2_U3228) );
  INV_X1 U8973 ( .A(n9943), .ZN(n8681) );
  OAI22_X1 U8974 ( .A1(n9939), .A2(n7105), .B1(n7104), .B2(n9936), .ZN(n7108)
         );
  MUX2_X1 U8975 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7106), .S(n8733), .Z(n7107)
         );
  AOI211_X1 U8976 ( .C1(n8681), .C2(n7109), .A(n7108), .B(n7107), .ZN(n7110)
         );
  INV_X1 U8977 ( .A(n7110), .ZN(P2_U3229) );
  NOR2_X1 U8978 ( .A1(n7112), .A2(n7111), .ZN(n7115) );
  NAND2_X1 U8979 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7299), .ZN(n7113) );
  OAI21_X1 U8980 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7299), .A(n7113), .ZN(
        n7114) );
  NOR2_X1 U8981 ( .A1(n7115), .A2(n7114), .ZN(n7287) );
  AOI21_X1 U8982 ( .B1(n7115), .B2(n7114), .A(n7287), .ZN(n7134) );
  OAI22_X1 U8983 ( .A1(n7119), .A2(n7118), .B1(n7117), .B2(n7116), .ZN(n7121)
         );
  MUX2_X1 U8984 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8503), .Z(n7289) );
  XNOR2_X1 U8985 ( .A(n7289), .B(n7131), .ZN(n7120) );
  NAND2_X1 U8986 ( .A1(n7121), .A2(n7120), .ZN(n7290) );
  OAI21_X1 U8987 ( .B1(n7121), .B2(n7120), .A(n7290), .ZN(n7122) );
  NAND2_X1 U8988 ( .A1(n7122), .A2(n9906), .ZN(n7133) );
  INV_X1 U8989 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7125) );
  INV_X1 U8990 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7123) );
  NOR2_X1 U8991 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7123), .ZN(n7139) );
  INV_X1 U8992 ( .A(n7139), .ZN(n7124) );
  OAI21_X1 U8993 ( .B1(n9899), .B2(n7125), .A(n7124), .ZN(n7130) );
  NAND2_X1 U8994 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7299), .ZN(n7126) );
  OAI21_X1 U8995 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7299), .A(n7126), .ZN(
        n7127) );
  AOI21_X1 U8996 ( .B1(n4443), .B2(n7127), .A(n7301), .ZN(n7128) );
  NOR2_X1 U8997 ( .A1(n7128), .A2(n9889), .ZN(n7129) );
  AOI211_X1 U8998 ( .C1(n9891), .C2(n7131), .A(n7130), .B(n7129), .ZN(n7132)
         );
  OAI211_X1 U8999 ( .C1(n7134), .C2(n9896), .A(n7133), .B(n7132), .ZN(P2_U3190) );
  XNOR2_X1 U9000 ( .A(n7137), .B(n7136), .ZN(n7138) );
  XNOR2_X1 U9001 ( .A(n7135), .B(n7138), .ZN(n7147) );
  AOI21_X1 U9002 ( .B1(n8318), .B2(n8352), .A(n7139), .ZN(n7145) );
  INV_X1 U9003 ( .A(n7244), .ZN(n7314) );
  NAND2_X1 U9004 ( .A1(n8250), .A2(n7314), .ZN(n7144) );
  INV_X1 U9005 ( .A(n7309), .ZN(n7140) );
  NAND2_X1 U9006 ( .A1(n8323), .A2(n7140), .ZN(n7143) );
  OR2_X1 U9007 ( .A1(n8320), .A2(n7141), .ZN(n7142) );
  NAND4_X1 U9008 ( .A1(n7145), .A2(n7144), .A3(n7143), .A4(n7142), .ZN(n7146)
         );
  AOI21_X1 U9009 ( .B1(n7147), .B2(n8315), .A(n7146), .ZN(n7148) );
  INV_X1 U9010 ( .A(n7148), .ZN(P2_U3161) );
  INV_X1 U9011 ( .A(n7149), .ZN(n7150) );
  AOI21_X1 U9012 ( .B1(n7152), .B2(n7151), .A(n7150), .ZN(n7158) );
  INV_X1 U9013 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7153) );
  OAI22_X1 U9014 ( .A1(n9025), .A2(n7154), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7153), .ZN(n7156) );
  OAI22_X1 U9015 ( .A1(n9027), .A2(n7330), .B1(n9721), .B2(n9034), .ZN(n7155)
         );
  AOI211_X1 U9016 ( .C1(n9718), .C2(n9030), .A(n7156), .B(n7155), .ZN(n7157)
         );
  OAI21_X1 U9017 ( .B1(n7158), .B2(n8999), .A(n7157), .ZN(P1_U3239) );
  INV_X1 U9018 ( .A(n7159), .ZN(n7727) );
  OAI222_X1 U9019 ( .A1(n8019), .A2(n7160), .B1(n8017), .B2(n7727), .C1(
        P2_U3151), .C2(n8539), .ZN(P2_U3276) );
  XNOR2_X1 U9020 ( .A(n7163), .B(n7162), .ZN(n7164) );
  XNOR2_X1 U9021 ( .A(n7161), .B(n7164), .ZN(n7171) );
  AOI22_X1 U9022 ( .A1(n8993), .A2(n9053), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7169) );
  NAND2_X1 U9023 ( .A1(n5752), .A2(n7182), .ZN(n7168) );
  NAND2_X1 U9024 ( .A1(n9030), .A2(n7181), .ZN(n7167) );
  OR2_X1 U9025 ( .A1(n9025), .A2(n7165), .ZN(n7166) );
  NAND4_X1 U9026 ( .A1(n7169), .A2(n7168), .A3(n7167), .A4(n7166), .ZN(n7170)
         );
  AOI21_X1 U9027 ( .B1(n7171), .B2(n9021), .A(n7170), .ZN(n7172) );
  INV_X1 U9028 ( .A(n7172), .ZN(P1_U3213) );
  INV_X1 U9029 ( .A(n7173), .ZN(n7250) );
  NAND2_X1 U9030 ( .A1(n7250), .A2(n4911), .ZN(n7249) );
  NAND2_X1 U9031 ( .A1(n7249), .A2(n7819), .ZN(n7174) );
  NAND2_X1 U9032 ( .A1(n7174), .A2(n7832), .ZN(n7220) );
  OAI21_X1 U9033 ( .B1(n7832), .B2(n7174), .A(n7220), .ZN(n7175) );
  NAND2_X1 U9034 ( .A1(n7175), .A2(n9702), .ZN(n7177) );
  AOI22_X1 U9035 ( .A1(n9053), .A2(n9311), .B1(n9309), .B2(n9055), .ZN(n7176)
         );
  NAND2_X1 U9036 ( .A1(n7177), .A2(n7176), .ZN(n9805) );
  INV_X1 U9037 ( .A(n9805), .ZN(n7187) );
  XNOR2_X1 U9038 ( .A(n7178), .B(n7179), .ZN(n9800) );
  OAI21_X1 U9039 ( .B1(n7253), .B2(n9802), .A(n9734), .ZN(n7180) );
  OR2_X1 U9040 ( .A1(n7180), .A2(n7227), .ZN(n9801) );
  AOI22_X1 U9041 ( .A1(n9754), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7181), .B2(
        n9749), .ZN(n7184) );
  NAND2_X1 U9042 ( .A1(n9739), .A2(n7182), .ZN(n7183) );
  OAI211_X1 U9043 ( .C1(n9801), .C2(n9694), .A(n7184), .B(n7183), .ZN(n7185)
         );
  AOI21_X1 U9044 ( .B1(n9800), .B2(n9715), .A(n7185), .ZN(n7186) );
  OAI21_X1 U9045 ( .B1(n7187), .B2(n9754), .A(n7186), .ZN(P1_U3286) );
  INV_X1 U9046 ( .A(n7188), .ZN(n7202) );
  OAI222_X1 U9047 ( .A1(n8023), .A2(n7202), .B1(n5749), .B2(P1_U3086), .C1(
        n7189), .C2(n9438), .ZN(P1_U3335) );
  INV_X1 U9048 ( .A(n7190), .ZN(n7191) );
  AOI211_X1 U9049 ( .C1(n7193), .C2(n7192), .A(n8327), .B(n7191), .ZN(n7200)
         );
  AND2_X1 U9050 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7295) );
  AOI21_X1 U9051 ( .B1(n8338), .B2(n8353), .A(n7295), .ZN(n7198) );
  NAND2_X1 U9052 ( .A1(n8250), .A2(n9980), .ZN(n7197) );
  INV_X1 U9053 ( .A(n7270), .ZN(n7194) );
  NAND2_X1 U9054 ( .A1(n8323), .A2(n7194), .ZN(n7196) );
  NAND2_X1 U9055 ( .A1(n8318), .A2(n8351), .ZN(n7195) );
  NAND4_X1 U9056 ( .A1(n7198), .A2(n7197), .A3(n7196), .A4(n7195), .ZN(n7199)
         );
  OR2_X1 U9057 ( .A1(n7200), .A2(n7199), .ZN(P2_U3171) );
  OAI222_X1 U9058 ( .A1(n8019), .A2(n7203), .B1(n8017), .B2(n7202), .C1(n7201), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  INV_X1 U9059 ( .A(n7204), .ZN(n7234) );
  OAI222_X1 U9060 ( .A1(n8023), .A2(n7234), .B1(n5720), .B2(P1_U3086), .C1(
        n7205), .C2(n9438), .ZN(P1_U3334) );
  NAND2_X1 U9061 ( .A1(n7207), .A2(n8040), .ZN(n7208) );
  NAND2_X1 U9062 ( .A1(n7206), .A2(n7208), .ZN(n9973) );
  AOI22_X1 U9063 ( .A1(n8354), .A2(n9933), .B1(n9930), .B2(n8353), .ZN(n7212)
         );
  INV_X1 U9064 ( .A(n8040), .ZN(n8111) );
  XNOR2_X1 U9065 ( .A(n7209), .B(n8111), .ZN(n7210) );
  NAND2_X1 U9066 ( .A1(n7210), .A2(n9928), .ZN(n7211) );
  OAI211_X1 U9067 ( .C1(n9973), .C2(n8717), .A(n7212), .B(n7211), .ZN(n9975)
         );
  MUX2_X1 U9068 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9975), .S(n8733), .Z(n7213)
         );
  INV_X1 U9069 ( .A(n7213), .ZN(n7218) );
  INV_X1 U9070 ( .A(n7214), .ZN(n7215) );
  AOI22_X1 U9071 ( .A1(n8705), .A2(n7216), .B1(n8729), .B2(n7215), .ZN(n7217)
         );
  OAI211_X1 U9072 ( .C1(n9973), .C2(n7694), .A(n7218), .B(n7217), .ZN(P2_U3226) );
  NAND2_X1 U9073 ( .A1(n7220), .A2(n7219), .ZN(n7221) );
  NAND2_X1 U9074 ( .A1(n7221), .A2(n4899), .ZN(n7274) );
  OAI21_X1 U9075 ( .B1(n4899), .B2(n7221), .A(n7274), .ZN(n7222) );
  NAND2_X1 U9076 ( .A1(n7222), .A2(n9702), .ZN(n7224) );
  AOI22_X1 U9077 ( .A1(n9054), .A2(n9309), .B1(n9311), .B2(n9052), .ZN(n7223)
         );
  NAND2_X1 U9078 ( .A1(n7224), .A2(n7223), .ZN(n9812) );
  INV_X1 U9079 ( .A(n9812), .ZN(n7233) );
  XNOR2_X1 U9080 ( .A(n7225), .B(n7226), .ZN(n9807) );
  OAI211_X1 U9081 ( .C1(n7227), .C2(n9809), .A(n9707), .B(n9734), .ZN(n9808)
         );
  AOI22_X1 U9082 ( .A1(n9754), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7333), .B2(
        n9749), .ZN(n7230) );
  NAND2_X1 U9083 ( .A1(n9739), .A2(n7228), .ZN(n7229) );
  OAI211_X1 U9084 ( .C1(n9808), .C2(n9694), .A(n7230), .B(n7229), .ZN(n7231)
         );
  AOI21_X1 U9085 ( .B1(n9807), .B2(n9715), .A(n7231), .ZN(n7232) );
  OAI21_X1 U9086 ( .B1(n7233), .B2(n9754), .A(n7232), .ZN(P1_U3285) );
  OAI222_X1 U9087 ( .A1(n8019), .A2(n7235), .B1(n8017), .B2(n7234), .C1(n8072), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  INV_X1 U9088 ( .A(n8107), .ZN(n7236) );
  OR2_X1 U9089 ( .A1(n8117), .A2(n7236), .ZN(n8041) );
  NAND2_X1 U9090 ( .A1(n7206), .A2(n7237), .ZN(n7238) );
  XOR2_X1 U9091 ( .A(n8041), .B(n7238), .Z(n7311) );
  XNOR2_X1 U9092 ( .A(n7239), .B(n8041), .ZN(n7240) );
  AOI222_X1 U9093 ( .A1(n9928), .A2(n7240), .B1(n8352), .B2(n9930), .C1(n9931), 
        .C2(n9933), .ZN(n7316) );
  OAI21_X1 U9094 ( .B1(n9965), .B2(n7311), .A(n7316), .ZN(n7246) );
  OAI22_X1 U9095 ( .A1(n7244), .A2(n8834), .B1(n9995), .B2(n5887), .ZN(n7241)
         );
  AOI21_X1 U9096 ( .B1(n7246), .B2(n9995), .A(n7241), .ZN(n7242) );
  INV_X1 U9097 ( .A(n7242), .ZN(P2_U3414) );
  INV_X1 U9098 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7243) );
  OAI22_X1 U9099 ( .A1(n8737), .A2(n7244), .B1(n10008), .B2(n7243), .ZN(n7245)
         );
  AOI21_X1 U9100 ( .B1(n7246), .B2(n10008), .A(n7245), .ZN(n7247) );
  INV_X1 U9101 ( .A(n7247), .ZN(P2_U3467) );
  NAND2_X1 U9102 ( .A1(n7319), .A2(n9747), .ZN(n7932) );
  OR2_X1 U9103 ( .A1(n7932), .A2(n8000), .ZN(n9765) );
  XNOR2_X1 U9104 ( .A(n7248), .B(n7954), .ZN(n9716) );
  OAI21_X1 U9105 ( .B1(n4911), .B2(n7250), .A(n7249), .ZN(n7251) );
  AOI222_X1 U9106 ( .A1(n9702), .A2(n7251), .B1(n9054), .B2(n9311), .C1(n9056), 
        .C2(n9309), .ZN(n9717) );
  INV_X1 U9107 ( .A(n7252), .ZN(n7255) );
  INV_X1 U9108 ( .A(n7253), .ZN(n7254) );
  OAI211_X1 U9109 ( .C1(n9721), .C2(n7255), .A(n7254), .B(n9734), .ZN(n9713)
         );
  OAI211_X1 U9110 ( .C1(n9721), .C2(n9846), .A(n9717), .B(n9713), .ZN(n7256)
         );
  AOI21_X1 U9111 ( .B1(n9842), .B2(n9716), .A(n7256), .ZN(n10231) );
  OR2_X1 U9112 ( .A1(n9421), .A2(n7257), .ZN(n7259) );
  OAI21_X1 U9113 ( .B1(n9421), .B2(P1_D_REG_1__SCAN_IN), .A(n9424), .ZN(n7258)
         );
  AND2_X1 U9114 ( .A1(n7259), .A2(n7258), .ZN(n7260) );
  NOR2_X1 U9115 ( .A1(n9334), .A2(n7262), .ZN(n7263) );
  NAND2_X1 U9116 ( .A1(n9852), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7264) );
  OAI21_X1 U9117 ( .B1(n10231), .B2(n9852), .A(n7264), .ZN(P1_U3471) );
  XNOR2_X1 U9118 ( .A(n7265), .B(n8045), .ZN(n9977) );
  AOI22_X1 U9119 ( .A1(n9933), .A2(n8353), .B1(n8351), .B2(n9930), .ZN(n7269)
         );
  XNOR2_X1 U9120 ( .A(n7266), .B(n8045), .ZN(n7267) );
  NAND2_X1 U9121 ( .A1(n7267), .A2(n9928), .ZN(n7268) );
  OAI211_X1 U9122 ( .C1(n9977), .C2(n8717), .A(n7269), .B(n7268), .ZN(n9978)
         );
  NAND2_X1 U9123 ( .A1(n9978), .A2(n8733), .ZN(n7273) );
  OAI22_X1 U9124 ( .A1(n8733), .A2(n5907), .B1(n7270), .B2(n9936), .ZN(n7271)
         );
  AOI21_X1 U9125 ( .B1(n8705), .B2(n9980), .A(n7271), .ZN(n7272) );
  OAI211_X1 U9126 ( .C1(n9977), .C2(n7694), .A(n7273), .B(n7272), .ZN(P2_U3224) );
  NAND2_X1 U9127 ( .A1(n7274), .A2(n7839), .ZN(n7275) );
  XNOR2_X1 U9128 ( .A(n7275), .B(n7278), .ZN(n7276) );
  OAI22_X1 U9129 ( .A1(n7276), .A2(n9759), .B1(n7426), .B2(n9008), .ZN(n9814)
         );
  INV_X1 U9130 ( .A(n9814), .ZN(n7285) );
  XNOR2_X1 U9131 ( .A(n7277), .B(n7278), .ZN(n9816) );
  XNOR2_X1 U9132 ( .A(n9707), .B(n4569), .ZN(n7280) );
  AND2_X1 U9133 ( .A1(n9051), .A2(n9311), .ZN(n7279) );
  AOI21_X1 U9134 ( .B1(n7280), .B2(n9734), .A(n7279), .ZN(n9813) );
  AOI22_X1 U9135 ( .A1(n9754), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7428), .B2(
        n9749), .ZN(n7282) );
  NAND2_X1 U9136 ( .A1(n4343), .A2(n9739), .ZN(n7281) );
  OAI211_X1 U9137 ( .C1(n9813), .C2(n9694), .A(n7282), .B(n7281), .ZN(n7283)
         );
  AOI21_X1 U9138 ( .B1(n9816), .B2(n9715), .A(n7283), .ZN(n7284) );
  OAI21_X1 U9139 ( .B1(n7285), .B2(n9754), .A(n7284), .ZN(P1_U3284) );
  XNOR2_X1 U9140 ( .A(n7372), .B(n7374), .ZN(n7288) );
  NOR2_X1 U9141 ( .A1(n7288), .A2(n5907), .ZN(n7376) );
  AOI21_X1 U9142 ( .B1(n5907), .B2(n7288), .A(n7376), .ZN(n7308) );
  INV_X1 U9143 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7298) );
  MUX2_X1 U9144 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8503), .Z(n7365) );
  XNOR2_X1 U9145 ( .A(n7365), .B(n7374), .ZN(n7293) );
  OR2_X1 U9146 ( .A1(n7289), .A2(n7299), .ZN(n7291) );
  NAND2_X1 U9147 ( .A1(n7291), .A2(n7290), .ZN(n7292) );
  NAND2_X1 U9148 ( .A1(n7293), .A2(n7292), .ZN(n7366) );
  OAI21_X1 U9149 ( .B1(n7293), .B2(n7292), .A(n7366), .ZN(n7294) );
  NAND2_X1 U9150 ( .A1(n7294), .A2(n9906), .ZN(n7297) );
  INV_X1 U9151 ( .A(n7295), .ZN(n7296) );
  OAI211_X1 U9152 ( .C1(n9899), .C2(n7298), .A(n7297), .B(n7296), .ZN(n7306)
         );
  AND2_X1 U9153 ( .A1(n7299), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7300) );
  NAND2_X1 U9154 ( .A1(n7302), .A2(n7373), .ZN(n7358) );
  AOI21_X1 U9155 ( .B1(n7303), .B2(n5902), .A(n7359), .ZN(n7304) );
  NOR2_X1 U9156 ( .A1(n7304), .A2(n9889), .ZN(n7305) );
  AOI211_X1 U9157 ( .C1(n9891), .C2(n7374), .A(n7306), .B(n7305), .ZN(n7307)
         );
  OAI21_X1 U9158 ( .B1(n7308), .B2(n9896), .A(n7307), .ZN(P2_U3191) );
  OAI22_X1 U9159 ( .A1(n8733), .A2(n7310), .B1(n7309), .B2(n9936), .ZN(n7313)
         );
  NOR2_X1 U9160 ( .A1(n7311), .A2(n9943), .ZN(n7312) );
  AOI211_X1 U9161 ( .C1(n8705), .C2(n7314), .A(n7313), .B(n7312), .ZN(n7315)
         );
  OAI21_X1 U9162 ( .B1(n8713), .B2(n7316), .A(n7315), .ZN(P2_U3225) );
  INV_X1 U9163 ( .A(n7317), .ZN(n7320) );
  OAI222_X1 U9164 ( .A1(n8019), .A2(n10086), .B1(n8017), .B2(n7320), .C1(n7318), .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9165 ( .A1(n9438), .A2(n7321), .B1(n9436), .B2(n7320), .C1(
        P1_U3086), .C2(n7319), .ZN(P1_U3333) );
  INV_X1 U9166 ( .A(n7322), .ZN(n7325) );
  INV_X1 U9167 ( .A(n7323), .ZN(n7324) );
  AND2_X1 U9168 ( .A1(n7323), .A2(n7322), .ZN(n7419) );
  AOI21_X1 U9169 ( .B1(n7325), .B2(n7324), .A(n7419), .ZN(n7326) );
  NAND2_X1 U9170 ( .A1(n7326), .A2(n7327), .ZN(n7421) );
  OAI21_X1 U9171 ( .B1(n7327), .B2(n7326), .A(n7421), .ZN(n7328) );
  NAND2_X1 U9172 ( .A1(n7328), .A2(n9021), .ZN(n7335) );
  NAND2_X1 U9173 ( .A1(n8993), .A2(n9052), .ZN(n7329) );
  NAND2_X1 U9174 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9505) );
  OAI211_X1 U9175 ( .C1(n9025), .C2(n7330), .A(n7329), .B(n9505), .ZN(n7332)
         );
  NOR2_X1 U9176 ( .A1(n9809), .A2(n9034), .ZN(n7331) );
  AOI211_X1 U9177 ( .C1(n7333), .C2(n9030), .A(n7332), .B(n7331), .ZN(n7334)
         );
  NAND2_X1 U9178 ( .A1(n7335), .A2(n7334), .ZN(P1_U3221) );
  XNOR2_X1 U9179 ( .A(n7336), .B(n7337), .ZN(n7338) );
  OAI222_X1 U9180 ( .A1(n8720), .A2(n7339), .B1(n8718), .B2(n7569), .C1(n7338), 
        .C2(n6157), .ZN(n9991) );
  INV_X1 U9181 ( .A(n9991), .ZN(n7346) );
  OAI21_X1 U9182 ( .B1(n7341), .B2(n8046), .A(n7340), .ZN(n9993) );
  INV_X1 U9183 ( .A(n7342), .ZN(n9990) );
  NOR2_X1 U9184 ( .A1(n9990), .A2(n9939), .ZN(n7344) );
  OAI22_X1 U9185 ( .A1(n8733), .A2(n5930), .B1(n7404), .B2(n9936), .ZN(n7343)
         );
  AOI211_X1 U9186 ( .C1(n9993), .C2(n8681), .A(n7344), .B(n7343), .ZN(n7345)
         );
  OAI21_X1 U9187 ( .B1(n7346), .B2(n8713), .A(n7345), .ZN(P2_U3222) );
  XNOR2_X1 U9188 ( .A(n7347), .B(n7348), .ZN(n7356) );
  NAND2_X1 U9189 ( .A1(n9986), .A2(n8250), .ZN(n7354) );
  INV_X1 U9190 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7349) );
  NOR2_X1 U9191 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7349), .ZN(n7438) );
  AOI21_X1 U9192 ( .B1(n8338), .B2(n8352), .A(n7438), .ZN(n7353) );
  INV_X1 U9193 ( .A(n7458), .ZN(n7350) );
  NAND2_X1 U9194 ( .A1(n8323), .A2(n7350), .ZN(n7352) );
  NAND2_X1 U9195 ( .A1(n8318), .A2(n8350), .ZN(n7351) );
  NAND4_X1 U9196 ( .A1(n7354), .A2(n7353), .A3(n7352), .A4(n7351), .ZN(n7355)
         );
  AOI21_X1 U9197 ( .B1(n7356), .B2(n8315), .A(n7355), .ZN(n7357) );
  INV_X1 U9198 ( .A(n7357), .ZN(P2_U3157) );
  INV_X1 U9199 ( .A(n7358), .ZN(n7360) );
  AOI22_X1 U9200 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7447), .B1(n7378), .B2(
        n7361), .ZN(n7443) );
  NAND2_X1 U9201 ( .A1(n7362), .A2(n7486), .ZN(n7470) );
  OAI21_X1 U9202 ( .B1(n7362), .B2(n7486), .A(n7470), .ZN(n7363) );
  NOR2_X1 U9203 ( .A1(n7363), .A2(n5927), .ZN(n7471) );
  AOI21_X1 U9204 ( .B1(n7363), .B2(n5927), .A(n7471), .ZN(n7389) );
  MUX2_X1 U9205 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8503), .Z(n7477) );
  XNOR2_X1 U9206 ( .A(n7477), .B(n7386), .ZN(n7370) );
  MUX2_X1 U9207 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8503), .Z(n7364) );
  OR2_X1 U9208 ( .A1(n7364), .A2(n7378), .ZN(n7368) );
  XNOR2_X1 U9209 ( .A(n7364), .B(n7447), .ZN(n7436) );
  OR2_X1 U9210 ( .A1(n7365), .A2(n7373), .ZN(n7367) );
  NAND2_X1 U9211 ( .A1(n7367), .A2(n7366), .ZN(n7435) );
  NAND2_X1 U9212 ( .A1(n7436), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U9213 ( .A1(n7368), .A2(n7434), .ZN(n7369) );
  NAND2_X1 U9214 ( .A1(n7370), .A2(n7369), .ZN(n7478) );
  OAI21_X1 U9215 ( .B1(n7370), .B2(n7369), .A(n7478), .ZN(n7385) );
  INV_X1 U9216 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7371) );
  NOR2_X1 U9217 ( .A1(n9899), .A2(n7371), .ZN(n7384) );
  MUX2_X1 U9218 ( .A(n7459), .B(P2_REG2_REG_10__SCAN_IN), .S(n7447), .Z(n7377)
         );
  INV_X1 U9219 ( .A(n7377), .ZN(n7432) );
  AOI21_X1 U9220 ( .B1(n5930), .B2(n7380), .A(n7484), .ZN(n7382) );
  NOR2_X1 U9221 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4573), .ZN(n7405) );
  INV_X1 U9222 ( .A(n7405), .ZN(n7381) );
  OAI21_X1 U9223 ( .B1(n9896), .B2(n7382), .A(n7381), .ZN(n7383) );
  AOI211_X1 U9224 ( .C1(n9906), .C2(n7385), .A(n7384), .B(n7383), .ZN(n7388)
         );
  NAND2_X1 U9225 ( .A1(n9891), .A2(n7386), .ZN(n7387) );
  OAI211_X1 U9226 ( .C1(n7389), .C2(n9889), .A(n7388), .B(n7387), .ZN(P2_U3193) );
  NAND3_X1 U9227 ( .A1(n7390), .A2(n7854), .A3(n7398), .ZN(n7391) );
  NAND2_X1 U9228 ( .A1(n7392), .A2(n7391), .ZN(n7393) );
  AOI222_X1 U9229 ( .A1(n9702), .A2(n7393), .B1(n9047), .B2(n9311), .C1(n9049), 
        .C2(n9309), .ZN(n9838) );
  OAI211_X1 U9230 ( .C1(n9839), .C2(n9669), .A(n4770), .B(n9734), .ZN(n9837)
         );
  INV_X1 U9231 ( .A(n9837), .ZN(n7396) );
  AOI22_X1 U9232 ( .A1(n9754), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7517), .B2(
        n9749), .ZN(n7394) );
  OAI21_X1 U9233 ( .B1(n9839), .B2(n9720), .A(n7394), .ZN(n7395) );
  AOI21_X1 U9234 ( .B1(n7396), .B2(n9738), .A(n7395), .ZN(n7400) );
  XNOR2_X1 U9235 ( .A(n7397), .B(n7398), .ZN(n9841) );
  NAND2_X1 U9236 ( .A1(n9841), .A2(n9715), .ZN(n7399) );
  OAI211_X1 U9237 ( .C1(n9838), .C2(n9754), .A(n7400), .B(n7399), .ZN(P1_U3280) );
  OAI211_X1 U9238 ( .C1(n7401), .C2(n7403), .A(n7402), .B(n8315), .ZN(n7410)
         );
  INV_X1 U9239 ( .A(n7404), .ZN(n7408) );
  AOI21_X1 U9240 ( .B1(n8338), .B2(n8351), .A(n7405), .ZN(n7406) );
  OAI21_X1 U9241 ( .B1(n8335), .B2(n7569), .A(n7406), .ZN(n7407) );
  AOI21_X1 U9242 ( .B1(n7408), .B2(n8323), .A(n7407), .ZN(n7409) );
  OAI211_X1 U9243 ( .C1(n9990), .C2(n8341), .A(n7410), .B(n7409), .ZN(P2_U3176) );
  NAND2_X1 U9244 ( .A1(n6078), .A2(n8865), .ZN(n7412) );
  NAND2_X1 U9245 ( .A1(n7411), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8231) );
  OAI211_X1 U9246 ( .C1(n7413), .C2(n8019), .A(n7412), .B(n8231), .ZN(P2_U3272) );
  NAND2_X1 U9247 ( .A1(n6078), .A2(n7414), .ZN(n7415) );
  OAI211_X1 U9248 ( .C1(n7416), .C2(n9438), .A(n7415), .B(n8015), .ZN(P1_U3332) );
  NOR2_X1 U9249 ( .A1(n7418), .A2(n7417), .ZN(n7423) );
  INV_X1 U9250 ( .A(n7419), .ZN(n7420) );
  NAND2_X1 U9251 ( .A1(n7421), .A2(n7420), .ZN(n7422) );
  XOR2_X1 U9252 ( .A(n7423), .B(n7422), .Z(n7431) );
  NAND2_X1 U9253 ( .A1(n8993), .A2(n9051), .ZN(n7425) );
  OAI211_X1 U9254 ( .C1(n9025), .C2(n7426), .A(n7425), .B(n7424), .ZN(n7427)
         );
  AOI21_X1 U9255 ( .B1(n7428), .B2(n9030), .A(n7427), .ZN(n7430) );
  NAND2_X1 U9256 ( .A1(n4343), .A2(n5752), .ZN(n7429) );
  OAI211_X1 U9257 ( .C1(n7431), .C2(n8999), .A(n7430), .B(n7429), .ZN(P1_U3231) );
  AOI21_X1 U9258 ( .B1(n7433), .B2(n7432), .A(n4436), .ZN(n7449) );
  INV_X1 U9259 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7441) );
  OAI21_X1 U9260 ( .B1(n7436), .B2(n7435), .A(n7434), .ZN(n7437) );
  NAND2_X1 U9261 ( .A1(n7437), .A2(n9906), .ZN(n7440) );
  INV_X1 U9262 ( .A(n7438), .ZN(n7439) );
  OAI211_X1 U9263 ( .C1(n9899), .C2(n7441), .A(n7440), .B(n7439), .ZN(n7446)
         );
  AOI21_X1 U9264 ( .B1(n4437), .B2(n7443), .A(n7442), .ZN(n7444) );
  NOR2_X1 U9265 ( .A1(n7444), .A2(n9889), .ZN(n7445) );
  AOI211_X1 U9266 ( .C1(n9891), .C2(n7447), .A(n7446), .B(n7445), .ZN(n7448)
         );
  OAI21_X1 U9267 ( .B1(n7449), .B2(n9896), .A(n7448), .ZN(P2_U3192) );
  NAND2_X1 U9268 ( .A1(n7450), .A2(n8113), .ZN(n7453) );
  INV_X1 U9269 ( .A(n7451), .ZN(n7452) );
  AOI21_X1 U9270 ( .B1(n8042), .B2(n7453), .A(n7452), .ZN(n9983) );
  AOI22_X1 U9271 ( .A1(n8350), .A2(n9930), .B1(n9933), .B2(n8352), .ZN(n7457)
         );
  XNOR2_X1 U9272 ( .A(n7454), .B(n8042), .ZN(n7455) );
  NAND2_X1 U9273 ( .A1(n7455), .A2(n9928), .ZN(n7456) );
  OAI211_X1 U9274 ( .C1(n9983), .C2(n8717), .A(n7457), .B(n7456), .ZN(n9984)
         );
  NAND2_X1 U9275 ( .A1(n9984), .A2(n8733), .ZN(n7462) );
  OAI22_X1 U9276 ( .A1(n8733), .A2(n7459), .B1(n7458), .B2(n9936), .ZN(n7460)
         );
  AOI21_X1 U9277 ( .B1(n8705), .B2(n9986), .A(n7460), .ZN(n7461) );
  OAI211_X1 U9278 ( .C1(n9983), .C2(n7694), .A(n7462), .B(n7461), .ZN(P2_U3223) );
  XOR2_X1 U9279 ( .A(n7464), .B(n7463), .Z(n7469) );
  AOI22_X1 U9280 ( .A1(n9311), .A2(n9048), .B1(n9050), .B2(n9309), .ZN(n9662)
         );
  NAND2_X1 U9281 ( .A1(n9030), .A2(n4962), .ZN(n7465) );
  OAI211_X1 U9282 ( .C1(n9662), .C2(n8959), .A(n7466), .B(n7465), .ZN(n7467)
         );
  AOI21_X1 U9283 ( .B1(n9665), .B2(n5752), .A(n7467), .ZN(n7468) );
  OAI21_X1 U9284 ( .B1(n7469), .B2(n8999), .A(n7468), .ZN(P1_U3224) );
  INV_X1 U9285 ( .A(n7470), .ZN(n7472) );
  NOR2_X1 U9286 ( .A1(n7472), .A2(n7471), .ZN(n7474) );
  AOI22_X1 U9287 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8377), .B1(n7475), .B2(
        n8376), .ZN(n7473) );
  NOR2_X1 U9288 ( .A1(n7474), .A2(n7473), .ZN(n8379) );
  AOI21_X1 U9289 ( .B1(n7474), .B2(n7473), .A(n8379), .ZN(n7495) );
  MUX2_X1 U9290 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8503), .Z(n7476) );
  AND2_X1 U9291 ( .A1(n7476), .A2(n7475), .ZN(n8358) );
  NOR2_X1 U9292 ( .A1(n7476), .A2(n7475), .ZN(n8361) );
  NOR2_X1 U9293 ( .A1(n8358), .A2(n8361), .ZN(n7480) );
  OR2_X1 U9294 ( .A1(n7477), .A2(n7486), .ZN(n7479) );
  NAND2_X1 U9295 ( .A1(n7479), .A2(n7478), .ZN(n8360) );
  XNOR2_X1 U9296 ( .A(n7480), .B(n8360), .ZN(n7481) );
  NAND2_X1 U9297 ( .A1(n7481), .A2(n9906), .ZN(n7494) );
  NOR2_X1 U9298 ( .A1(n9899), .A2(n7482), .ZN(n7492) );
  INV_X1 U9299 ( .A(n7483), .ZN(n7485) );
  MUX2_X1 U9300 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8367), .S(n8377), .Z(n7487)
         );
  NOR2_X1 U9301 ( .A1(n7488), .A2(n7487), .ZN(n8368) );
  AOI21_X1 U9302 ( .B1(n7488), .B2(n7487), .A(n8368), .ZN(n7490) );
  AND2_X1 U9303 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7508) );
  INV_X1 U9304 ( .A(n7508), .ZN(n7489) );
  OAI21_X1 U9305 ( .B1(n9896), .B2(n7490), .A(n7489), .ZN(n7491) );
  AOI211_X1 U9306 ( .C1(n9891), .C2(n8377), .A(n7492), .B(n7491), .ZN(n7493)
         );
  OAI211_X1 U9307 ( .C1(n7495), .C2(n9889), .A(n7494), .B(n7493), .ZN(P2_U3194) );
  XNOR2_X1 U9308 ( .A(n7496), .B(n7580), .ZN(n7497) );
  NOR2_X1 U9309 ( .A1(n7497), .A2(n7498), .ZN(n7579) );
  AOI21_X1 U9310 ( .B1(n7498), .B2(n7497), .A(n7579), .ZN(n7503) );
  AOI22_X1 U9311 ( .A1(n9309), .A2(n9052), .B1(n9050), .B2(n9311), .ZN(n9700)
         );
  OAI22_X1 U9312 ( .A1(n9700), .A2(n8959), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7499), .ZN(n7500) );
  AOI21_X1 U9313 ( .B1(n9704), .B2(n9030), .A(n7500), .ZN(n7502) );
  NAND2_X1 U9314 ( .A1(n9818), .A2(n5752), .ZN(n7501) );
  OAI211_X1 U9315 ( .C1(n7503), .C2(n8999), .A(n7502), .B(n7501), .ZN(P1_U3217) );
  INV_X1 U9316 ( .A(n7547), .ZN(n7514) );
  OAI211_X1 U9317 ( .C1(n7506), .C2(n7505), .A(n7504), .B(n8315), .ZN(n7513)
         );
  INV_X1 U9318 ( .A(n7507), .ZN(n7540) );
  AOI21_X1 U9319 ( .B1(n8318), .B2(n8348), .A(n7508), .ZN(n7509) );
  OAI21_X1 U9320 ( .B1(n7510), .B2(n8320), .A(n7509), .ZN(n7511) );
  AOI21_X1 U9321 ( .B1(n7540), .B2(n8323), .A(n7511), .ZN(n7512) );
  OAI211_X1 U9322 ( .C1(n7514), .C2(n8341), .A(n7513), .B(n7512), .ZN(P2_U3164) );
  XOR2_X1 U9323 ( .A(n7516), .B(n7515), .Z(n7523) );
  AOI22_X1 U9324 ( .A1(n8993), .A2(n9047), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n7519) );
  NAND2_X1 U9325 ( .A1(n9030), .A2(n7517), .ZN(n7518) );
  OAI211_X1 U9326 ( .C1(n7585), .C2(n9025), .A(n7519), .B(n7518), .ZN(n7520)
         );
  AOI21_X1 U9327 ( .B1(n7521), .B2(n5752), .A(n7520), .ZN(n7522) );
  OAI21_X1 U9328 ( .B1(n7523), .B2(n8999), .A(n7522), .ZN(P1_U3234) );
  XOR2_X1 U9329 ( .A(n7524), .B(n7963), .Z(n9844) );
  XOR2_X1 U9330 ( .A(n7963), .B(n7525), .Z(n7527) );
  OAI22_X1 U9331 ( .A1(n7558), .A2(n9008), .B1(n8944), .B2(n9006), .ZN(n7526)
         );
  AOI21_X1 U9332 ( .B1(n7527), .B2(n9702), .A(n7526), .ZN(n7528) );
  OAI21_X1 U9333 ( .B1(n9844), .B2(n7529), .A(n7528), .ZN(n9848) );
  NAND2_X1 U9334 ( .A1(n9848), .A2(n9752), .ZN(n7534) );
  OAI211_X1 U9335 ( .C1(n4767), .C2(n9847), .A(n9734), .B(n4347), .ZN(n9845)
         );
  INV_X1 U9336 ( .A(n9845), .ZN(n7532) );
  AOI22_X1 U9337 ( .A1(n9754), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7555), .B2(
        n9749), .ZN(n7530) );
  OAI21_X1 U9338 ( .B1(n9847), .B2(n9720), .A(n7530), .ZN(n7531) );
  AOI21_X1 U9339 ( .B1(n7532), .B2(n9738), .A(n7531), .ZN(n7533) );
  OAI211_X1 U9340 ( .C1(n9844), .C2(n9686), .A(n7534), .B(n7533), .ZN(P1_U3279) );
  INV_X1 U9341 ( .A(n7535), .ZN(n7537) );
  INV_X1 U9342 ( .A(n8136), .ZN(n8047) );
  OAI21_X1 U9343 ( .B1(n7537), .B2(n8047), .A(n7536), .ZN(n7550) );
  XNOR2_X1 U9344 ( .A(n7538), .B(n8047), .ZN(n7539) );
  AOI222_X1 U9345 ( .A1(n9928), .A2(n7539), .B1(n8350), .B2(n9933), .C1(n8348), 
        .C2(n9930), .ZN(n7546) );
  MUX2_X1 U9346 ( .A(n8367), .B(n7546), .S(n8733), .Z(n7542) );
  AOI22_X1 U9347 ( .A1(n7547), .A2(n8705), .B1(n8729), .B2(n7540), .ZN(n7541)
         );
  OAI211_X1 U9348 ( .C1(n9943), .C2(n7550), .A(n7542), .B(n7541), .ZN(P2_U3221) );
  INV_X1 U9349 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7543) );
  MUX2_X1 U9350 ( .A(n7543), .B(n7546), .S(n9995), .Z(n7545) );
  NAND2_X1 U9351 ( .A1(n7547), .A2(n8854), .ZN(n7544) );
  OAI211_X1 U9352 ( .C1(n7550), .C2(n8858), .A(n7545), .B(n7544), .ZN(P2_U3426) );
  MUX2_X1 U9353 ( .A(n8376), .B(n7546), .S(n10008), .Z(n7549) );
  NAND2_X1 U9354 ( .A1(n7547), .A2(n8780), .ZN(n7548) );
  OAI211_X1 U9355 ( .C1(n7550), .C2(n8783), .A(n7549), .B(n7548), .ZN(P2_U3471) );
  XNOR2_X1 U9356 ( .A(n7552), .B(n7551), .ZN(n7553) );
  XNOR2_X1 U9357 ( .A(n7554), .B(n7553), .ZN(n7562) );
  AOI22_X1 U9358 ( .A1(n8993), .A2(n9046), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n7557) );
  NAND2_X1 U9359 ( .A1(n9030), .A2(n7555), .ZN(n7556) );
  OAI211_X1 U9360 ( .C1(n7558), .C2(n9025), .A(n7557), .B(n7556), .ZN(n7559)
         );
  AOI21_X1 U9361 ( .B1(n7560), .B2(n5752), .A(n7559), .ZN(n7561) );
  OAI21_X1 U9362 ( .B1(n7562), .B2(n8999), .A(n7561), .ZN(P1_U3215) );
  INV_X1 U9363 ( .A(n7563), .ZN(n7657) );
  OAI222_X1 U9364 ( .A1(n8023), .A2(n7657), .B1(n7565), .B2(P1_U3086), .C1(
        n7564), .C2(n9438), .ZN(P1_U3331) );
  XNOR2_X1 U9365 ( .A(n7566), .B(n8348), .ZN(n7567) );
  XNOR2_X1 U9366 ( .A(n7568), .B(n7567), .ZN(n7574) );
  AND2_X1 U9367 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8372) );
  NOR2_X1 U9368 ( .A1(n8320), .A2(n7569), .ZN(n7570) );
  AOI211_X1 U9369 ( .C1(n8318), .C2(n8347), .A(n8372), .B(n7570), .ZN(n7571)
         );
  OAI21_X1 U9370 ( .B1(n7607), .B2(n8333), .A(n7571), .ZN(n7572) );
  AOI21_X1 U9371 ( .B1(n7606), .B2(n8250), .A(n7572), .ZN(n7573) );
  OAI21_X1 U9372 ( .B1(n7574), .B2(n8327), .A(n7573), .ZN(P2_U3174) );
  INV_X1 U9373 ( .A(n7575), .ZN(n7593) );
  INV_X1 U9374 ( .A(n7576), .ZN(n7578) );
  OAI222_X1 U9375 ( .A1(n8023), .A2(n7593), .B1(n7578), .B2(P1_U3086), .C1(
        n7577), .C2(n9438), .ZN(P1_U3330) );
  AOI21_X1 U9376 ( .B1(n7580), .B2(n7496), .A(n7579), .ZN(n7584) );
  XOR2_X1 U9377 ( .A(n7582), .B(n7581), .Z(n7583) );
  XNOR2_X1 U9378 ( .A(n7584), .B(n7583), .ZN(n7592) );
  OR2_X1 U9379 ( .A1(n7585), .A2(n9006), .ZN(n7587) );
  NAND2_X1 U9380 ( .A1(n9051), .A2(n9309), .ZN(n7586) );
  AND2_X1 U9381 ( .A1(n7587), .A2(n7586), .ZN(n9677) );
  OAI22_X1 U9382 ( .A1(n9677), .A2(n8959), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7588), .ZN(n7589) );
  AOI21_X1 U9383 ( .B1(n9690), .B2(n9030), .A(n7589), .ZN(n7591) );
  NAND2_X1 U9384 ( .A1(n9691), .A2(n5752), .ZN(n7590) );
  OAI211_X1 U9385 ( .C1(n7592), .C2(n8999), .A(n7591), .B(n7590), .ZN(P1_U3236) );
  OAI222_X1 U9386 ( .A1(n8019), .A2(n7594), .B1(n8017), .B2(n7593), .C1(n6189), 
        .C2(P2_U3151), .ZN(P2_U3270) );
  NAND2_X1 U9387 ( .A1(n7596), .A2(n7595), .ZN(n8135) );
  XNOR2_X1 U9388 ( .A(n7597), .B(n8135), .ZN(n7613) );
  XOR2_X1 U9389 ( .A(n7598), .B(n8135), .Z(n7599) );
  AOI222_X1 U9390 ( .A1(n9928), .A2(n7599), .B1(n8347), .B2(n9930), .C1(n8349), 
        .C2(n9933), .ZN(n7605) );
  MUX2_X1 U9391 ( .A(n7600), .B(n7605), .S(n9995), .Z(n7602) );
  NAND2_X1 U9392 ( .A1(n7606), .A2(n8854), .ZN(n7601) );
  OAI211_X1 U9393 ( .C1(n7613), .C2(n8858), .A(n7602), .B(n7601), .ZN(P2_U3429) );
  MUX2_X1 U9394 ( .A(n8382), .B(n7605), .S(n10008), .Z(n7604) );
  NAND2_X1 U9395 ( .A1(n7606), .A2(n8780), .ZN(n7603) );
  OAI211_X1 U9396 ( .C1(n8783), .C2(n7613), .A(n7604), .B(n7603), .ZN(P2_U3472) );
  INV_X1 U9397 ( .A(n7605), .ZN(n7610) );
  INV_X1 U9398 ( .A(n7606), .ZN(n7608) );
  OAI22_X1 U9399 ( .A1(n7608), .A2(n8709), .B1(n7607), .B2(n9936), .ZN(n7609)
         );
  OAI21_X1 U9400 ( .B1(n7610), .B2(n7609), .A(n8733), .ZN(n7612) );
  NAND2_X1 U9401 ( .A1(n8713), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7611) );
  OAI211_X1 U9402 ( .C1(n7613), .C2(n9943), .A(n7612), .B(n7611), .ZN(P2_U3220) );
  INV_X1 U9403 ( .A(n7614), .ZN(n7623) );
  INV_X1 U9404 ( .A(n7615), .ZN(n7616) );
  OAI222_X1 U9405 ( .A1(n8023), .A2(n7623), .B1(n7616), .B2(P1_U3086), .C1(
        n10169), .C2(n9438), .ZN(P1_U3329) );
  AND2_X1 U9406 ( .A1(n8143), .A2(n8144), .ZN(n8049) );
  XNOR2_X1 U9407 ( .A(n7617), .B(n8142), .ZN(n8859) );
  XNOR2_X1 U9408 ( .A(n7618), .B(n8142), .ZN(n7619) );
  AOI222_X1 U9409 ( .A1(n9928), .A2(n7619), .B1(n8699), .B2(n9930), .C1(n8348), 
        .C2(n9933), .ZN(n8852) );
  MUX2_X1 U9410 ( .A(n8395), .B(n8852), .S(n10008), .Z(n7621) );
  NAND2_X1 U9411 ( .A1(n8855), .A2(n8780), .ZN(n7620) );
  OAI211_X1 U9412 ( .C1(n8783), .C2(n8859), .A(n7621), .B(n7620), .ZN(P2_U3473) );
  OAI222_X1 U9413 ( .A1(n8019), .A2(n10218), .B1(n8017), .B2(n7623), .C1(n7622), .C2(P2_U3151), .ZN(P2_U3269) );
  INV_X1 U9414 ( .A(n7624), .ZN(n8016) );
  OAI222_X1 U9415 ( .A1(n8023), .A2(n8016), .B1(P1_U3086), .B2(n7626), .C1(
        n7625), .C2(n9438), .ZN(P1_U3328) );
  XNOR2_X1 U9416 ( .A(n7627), .B(n7630), .ZN(n9517) );
  INV_X1 U9417 ( .A(n9517), .ZN(n7638) );
  INV_X1 U9418 ( .A(n8946), .ZN(n7632) );
  OAI21_X1 U9419 ( .B1(n7630), .B2(n7629), .A(n7628), .ZN(n7631) );
  AOI222_X1 U9420 ( .A1(n9702), .A2(n7631), .B1(n9301), .B2(n9311), .C1(n9046), 
        .C2(n9309), .ZN(n9514) );
  OAI21_X1 U9421 ( .B1(n7632), .B2(n9315), .A(n9514), .ZN(n7636) );
  AOI21_X1 U9422 ( .B1(n9512), .B2(n7640), .A(n9246), .ZN(n7633) );
  NAND2_X1 U9423 ( .A1(n7633), .A2(n9318), .ZN(n9513) );
  AOI22_X1 U9424 ( .A1(n9512), .A2(n9739), .B1(n9754), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n7634) );
  OAI21_X1 U9425 ( .B1(n9513), .B2(n9694), .A(n7634), .ZN(n7635) );
  AOI21_X1 U9426 ( .B1(n7636), .B2(n9752), .A(n7635), .ZN(n7637) );
  OAI21_X1 U9427 ( .B1(n9307), .B2(n7638), .A(n7637), .ZN(P1_U3277) );
  XNOR2_X1 U9428 ( .A(n7639), .B(n7644), .ZN(n9405) );
  INV_X1 U9429 ( .A(n7640), .ZN(n7641) );
  AOI211_X1 U9430 ( .C1(n9402), .C2(n4347), .A(n9246), .B(n7641), .ZN(n9401)
         );
  INV_X1 U9431 ( .A(n9402), .ZN(n9035) );
  AOI22_X1 U9432 ( .A1(n9754), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9031), .B2(
        n9749), .ZN(n7642) );
  OAI21_X1 U9433 ( .B1(n9035), .B2(n9720), .A(n7642), .ZN(n7648) );
  OAI21_X1 U9434 ( .B1(n7645), .B2(n7644), .A(n7643), .ZN(n7646) );
  AOI222_X1 U9435 ( .A1(n9702), .A2(n7646), .B1(n9310), .B2(n9311), .C1(n9047), 
        .C2(n9309), .ZN(n9404) );
  NOR2_X1 U9436 ( .A1(n9404), .A2(n9754), .ZN(n7647) );
  AOI211_X1 U9437 ( .C1(n9401), .C2(n9738), .A(n7648), .B(n7647), .ZN(n7649)
         );
  OAI21_X1 U9438 ( .B1(n9307), .B2(n9405), .A(n7649), .ZN(P1_U3278) );
  NAND2_X1 U9439 ( .A1(n8020), .A2(n8865), .ZN(n7651) );
  OAI211_X1 U9440 ( .C1(n8019), .C2(n7652), .A(n7651), .B(n7650), .ZN(P2_U3267) );
  INV_X1 U9441 ( .A(n6474), .ZN(n7656) );
  OAI222_X1 U9442 ( .A1(n7654), .A2(P2_U3151), .B1(n8017), .B2(n7656), .C1(
        n7653), .C2(n8019), .ZN(P2_U3266) );
  OAI222_X1 U9443 ( .A1(n8023), .A2(n7656), .B1(P1_U3086), .B2(n5109), .C1(
        n7655), .C2(n9438), .ZN(P1_U3326) );
  OAI222_X1 U9444 ( .A1(n8019), .A2(n10055), .B1(n8017), .B2(n7657), .C1(n6186), .C2(P2_U3151), .ZN(P2_U3271) );
  INV_X1 U9445 ( .A(SI_29_), .ZN(n7661) );
  INV_X1 U9446 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7667) );
  INV_X1 U9447 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9437) );
  MUX2_X1 U9448 ( .A(n7667), .B(n9437), .S(n7795), .Z(n7663) );
  INV_X1 U9449 ( .A(SI_30_), .ZN(n10212) );
  NAND2_X1 U9450 ( .A1(n7663), .A2(n10212), .ZN(n7788) );
  INV_X1 U9451 ( .A(n7663), .ZN(n7664) );
  NAND2_X1 U9452 ( .A1(n7664), .A2(SI_30_), .ZN(n7665) );
  NAND2_X1 U9453 ( .A1(n7788), .A2(n7665), .ZN(n7789) );
  INV_X1 U9454 ( .A(n7783), .ZN(n9435) );
  NOR2_X1 U9455 ( .A1(n5824), .A2(n7667), .ZN(n7668) );
  INV_X1 U9456 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U9457 ( .A1(n6095), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7671) );
  INV_X1 U9458 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7669) );
  OR2_X1 U9459 ( .A1(n5828), .A2(n7669), .ZN(n7670) );
  OAI211_X1 U9460 ( .C1(n5832), .C2(n7672), .A(n7671), .B(n7670), .ZN(n7673)
         );
  INV_X1 U9461 ( .A(n7673), .ZN(n7674) );
  NAND2_X1 U9462 ( .A1(n7675), .A2(n7674), .ZN(n8343) );
  NAND2_X1 U9463 ( .A1(n8343), .A2(n7676), .ZN(n8784) );
  NOR2_X1 U9464 ( .A1(n8784), .A2(n6287), .ZN(n8735) );
  AOI21_X1 U9465 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n6287), .A(n8735), .ZN(
        n7677) );
  OAI21_X1 U9466 ( .B1(n8027), .B2(n8737), .A(n7677), .ZN(P2_U3489) );
  INV_X1 U9467 ( .A(n8784), .ZN(n7679) );
  NOR2_X1 U9468 ( .A1(n7678), .A2(n9936), .ZN(n7691) );
  AOI21_X1 U9469 ( .B1(n7679), .B2(n8733), .A(n7691), .ZN(n8545) );
  NAND2_X1 U9470 ( .A1(n8713), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7680) );
  OAI211_X1 U9471 ( .C1(n8027), .C2(n9939), .A(n8545), .B(n7680), .ZN(P2_U3203) );
  XNOR2_X1 U9472 ( .A(n7682), .B(n7681), .ZN(n7687) );
  NAND2_X1 U9473 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8451) );
  OAI21_X1 U9474 ( .B1(n8335), .B2(n8321), .A(n8451), .ZN(n7683) );
  AOI21_X1 U9475 ( .B1(n8338), .B2(n8699), .A(n7683), .ZN(n7684) );
  OAI21_X1 U9476 ( .B1(n8703), .B2(n8333), .A(n7684), .ZN(n7685) );
  AOI21_X1 U9477 ( .B1(n8848), .B2(n8250), .A(n7685), .ZN(n7686) );
  OAI21_X1 U9478 ( .B1(n7687), .B2(n8327), .A(n7686), .ZN(P2_U3166) );
  NAND2_X1 U9479 ( .A1(n7688), .A2(n8733), .ZN(n7693) );
  NOR2_X1 U9480 ( .A1(n7689), .A2(n9939), .ZN(n7690) );
  AOI211_X1 U9481 ( .C1(n8713), .C2(P2_REG2_REG_29__SCAN_IN), .A(n7691), .B(
        n7690), .ZN(n7692) );
  OAI211_X1 U9482 ( .C1(n6278), .C2(n7694), .A(n7693), .B(n7692), .ZN(P2_U3204) );
  XOR2_X1 U9483 ( .A(n7695), .B(n8146), .Z(n7707) );
  INV_X1 U9484 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7698) );
  XOR2_X1 U9485 ( .A(n8146), .B(n7696), .Z(n7697) );
  AOI222_X1 U9486 ( .A1(n9928), .A2(n7697), .B1(n8347), .B2(n9933), .C1(n8686), 
        .C2(n9930), .ZN(n7703) );
  MUX2_X1 U9487 ( .A(n7698), .B(n7703), .S(n9995), .Z(n7700) );
  NAND2_X1 U9488 ( .A1(n8326), .A2(n8854), .ZN(n7699) );
  OAI211_X1 U9489 ( .C1(n7707), .C2(n8858), .A(n7700), .B(n7699), .ZN(P2_U3435) );
  MUX2_X1 U9490 ( .A(n8418), .B(n7703), .S(n10008), .Z(n7702) );
  NAND2_X1 U9491 ( .A1(n8326), .A2(n8780), .ZN(n7701) );
  OAI211_X1 U9492 ( .C1(n8783), .C2(n7707), .A(n7702), .B(n7701), .ZN(P2_U3474) );
  MUX2_X1 U9493 ( .A(n8419), .B(n7703), .S(n8733), .Z(n7706) );
  INV_X1 U9494 ( .A(n8332), .ZN(n7704) );
  AOI22_X1 U9495 ( .A1(n8326), .A2(n8705), .B1(n8729), .B2(n7704), .ZN(n7705)
         );
  OAI211_X1 U9496 ( .C1(n7707), .C2(n9943), .A(n7706), .B(n7705), .ZN(P2_U3218) );
  XNOR2_X1 U9497 ( .A(n7708), .B(n8557), .ZN(n7709) );
  XNOR2_X1 U9498 ( .A(n7710), .B(n7709), .ZN(n7716) );
  AOI22_X1 U9499 ( .A1(n8590), .A2(n8338), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7712) );
  NAND2_X1 U9500 ( .A1(n8574), .A2(n8323), .ZN(n7711) );
  OAI211_X1 U9501 ( .C1(n7713), .C2(n8335), .A(n7712), .B(n7711), .ZN(n7714)
         );
  AOI21_X1 U9502 ( .B1(n8798), .B2(n8250), .A(n7714), .ZN(n7715) );
  OAI21_X1 U9503 ( .B1(n7716), .B2(n8327), .A(n7715), .ZN(P2_U3180) );
  AOI22_X1 U9504 ( .A1(n8605), .A2(n8338), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7718) );
  NAND2_X1 U9505 ( .A1(n8583), .A2(n8323), .ZN(n7717) );
  OAI211_X1 U9506 ( .C1(n8557), .C2(n8335), .A(n7718), .B(n7717), .ZN(n7725)
         );
  NAND2_X1 U9507 ( .A1(n7720), .A2(n8278), .ZN(n8281) );
  NAND3_X1 U9508 ( .A1(n8281), .A2(n7722), .A3(n7721), .ZN(n7723) );
  AOI21_X1 U9509 ( .B1(n7719), .B2(n7723), .A(n8327), .ZN(n7724) );
  AOI211_X1 U9510 ( .C1(n8803), .C2(n8250), .A(n7725), .B(n7724), .ZN(n7726)
         );
  INV_X1 U9511 ( .A(n7726), .ZN(P2_U3165) );
  OAI222_X1 U9512 ( .A1(n9438), .A2(n7728), .B1(n9436), .B2(n7727), .C1(
        P1_U3086), .C2(n8003), .ZN(P1_U3336) );
  NAND2_X1 U9513 ( .A1(n7931), .A2(n7729), .ZN(n7989) );
  NAND2_X1 U9514 ( .A1(n7927), .A2(n7917), .ZN(n7985) );
  INV_X1 U9515 ( .A(n7985), .ZN(n7780) );
  NAND2_X1 U9516 ( .A1(n7902), .A2(n7730), .ZN(n7804) );
  NAND2_X1 U9517 ( .A1(n7804), .A2(n7908), .ZN(n7731) );
  NAND2_X1 U9518 ( .A1(n7911), .A2(n7731), .ZN(n7732) );
  NAND2_X1 U9519 ( .A1(n7732), .A2(n7910), .ZN(n7733) );
  AND2_X1 U9520 ( .A1(n7734), .A2(n7733), .ZN(n7773) );
  INV_X1 U9521 ( .A(n7773), .ZN(n7984) );
  INV_X1 U9522 ( .A(n7852), .ZN(n7735) );
  NOR2_X1 U9523 ( .A1(n7736), .A2(n7735), .ZN(n7844) );
  NAND2_X1 U9524 ( .A1(n7737), .A2(n9735), .ZN(n7946) );
  NAND2_X1 U9525 ( .A1(n6493), .A2(n9767), .ZN(n7738) );
  AND4_X1 U9526 ( .A1(n7822), .A2(n7946), .A3(n7739), .A4(n7738), .ZN(n7740)
         );
  OAI211_X1 U9527 ( .C1(n7741), .C2(n7740), .A(n7823), .B(n7827), .ZN(n7742)
         );
  NAND3_X1 U9528 ( .A1(n7742), .A2(n7816), .A3(n7825), .ZN(n7743) );
  NAND2_X1 U9529 ( .A1(n7743), .A2(n7814), .ZN(n7745) );
  NAND3_X1 U9530 ( .A1(n7745), .A2(n7744), .A3(n7819), .ZN(n7746) );
  NAND3_X1 U9531 ( .A1(n7844), .A2(n7747), .A3(n7746), .ZN(n7752) );
  NAND2_X1 U9532 ( .A1(n7853), .A2(n7748), .ZN(n7750) );
  INV_X1 U9533 ( .A(n7854), .ZN(n7749) );
  AOI21_X1 U9534 ( .B1(n7751), .B2(n7750), .A(n7749), .ZN(n7847) );
  AND3_X1 U9535 ( .A1(n7752), .A2(n7847), .A3(n7874), .ZN(n7753) );
  NAND2_X1 U9536 ( .A1(n7865), .A2(n7861), .ZN(n7873) );
  OAI21_X1 U9537 ( .B1(n7753), .B2(n7873), .A(n7862), .ZN(n7758) );
  NAND2_X1 U9538 ( .A1(n7872), .A2(n7754), .ZN(n7877) );
  NAND2_X1 U9539 ( .A1(n7871), .A2(n7755), .ZN(n7868) );
  NAND2_X1 U9540 ( .A1(n7868), .A2(n7872), .ZN(n7756) );
  OAI211_X1 U9541 ( .C1(n7758), .C2(n7877), .A(n7757), .B(n7756), .ZN(n7759)
         );
  NAND3_X1 U9542 ( .A1(n7761), .A2(n7760), .A3(n7759), .ZN(n7762) );
  NAND3_X1 U9543 ( .A1(n7764), .A2(n7763), .A3(n7762), .ZN(n7766) );
  NAND2_X1 U9544 ( .A1(n7766), .A2(n7765), .ZN(n7767) );
  NAND3_X1 U9545 ( .A1(n7903), .A2(n9241), .A3(n7767), .ZN(n7768) );
  NOR2_X1 U9546 ( .A1(n7984), .A2(n7768), .ZN(n7778) );
  INV_X1 U9547 ( .A(n7926), .ZN(n7769) );
  NAND2_X1 U9548 ( .A1(n7769), .A2(n7923), .ZN(n7915) );
  INV_X1 U9549 ( .A(n7915), .ZN(n7775) );
  NAND2_X1 U9550 ( .A1(n7908), .A2(n7770), .ZN(n7805) );
  INV_X1 U9551 ( .A(n7805), .ZN(n7771) );
  NAND3_X1 U9552 ( .A1(n7910), .A2(n7771), .A3(n7904), .ZN(n7772) );
  NAND2_X1 U9553 ( .A1(n7773), .A2(n7772), .ZN(n7774) );
  AND2_X1 U9554 ( .A1(n7775), .A2(n7774), .ZN(n7982) );
  INV_X1 U9555 ( .A(n7982), .ZN(n7777) );
  OR2_X1 U9556 ( .A1(n9356), .A2(n7776), .ZN(n7914) );
  NAND2_X1 U9557 ( .A1(n7925), .A2(n7914), .ZN(n7920) );
  INV_X1 U9558 ( .A(n7920), .ZN(n7987) );
  OAI21_X1 U9559 ( .B1(n7778), .B2(n7777), .A(n7987), .ZN(n7779) );
  AND2_X1 U9560 ( .A1(n7780), .A2(n7779), .ZN(n7781) );
  NOR2_X1 U9561 ( .A1(n7989), .A2(n7781), .ZN(n7787) );
  NAND2_X1 U9562 ( .A1(n7783), .A2(n7782), .ZN(n7785) );
  OR2_X1 U9563 ( .A1(n4341), .A2(n9437), .ZN(n7784) );
  NAND2_X1 U9564 ( .A1(n9135), .A2(n7786), .ZN(n7975) );
  NAND2_X1 U9565 ( .A1(n7975), .A2(n7929), .ZN(n7991) );
  OR2_X1 U9566 ( .A1(n9135), .A2(n7786), .ZN(n7976) );
  OAI21_X1 U9567 ( .B1(n7787), .B2(n7991), .A(n7976), .ZN(n7801) );
  INV_X1 U9568 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8862) );
  INV_X1 U9569 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7791) );
  MUX2_X1 U9570 ( .A(n8862), .B(n7791), .S(n7795), .Z(n7792) );
  XNOR2_X1 U9571 ( .A(n7792), .B(SI_31_), .ZN(n7793) );
  MUX2_X1 U9572 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9426), .S(n7795), .Z(n7797) );
  INV_X1 U9573 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U9574 ( .A1(n5520), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U9575 ( .A1(n5521), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7798) );
  OAI211_X1 U9576 ( .C1(n4336), .C2(n9127), .A(n7799), .B(n7798), .ZN(n9125)
         );
  NAND2_X1 U9577 ( .A1(n9332), .A2(n9125), .ZN(n7993) );
  NAND2_X1 U9578 ( .A1(n7801), .A2(n7993), .ZN(n7802) );
  NOR2_X1 U9579 ( .A1(n8007), .A2(n8003), .ZN(n8001) );
  INV_X1 U9580 ( .A(n7932), .ZN(n7937) );
  INV_X1 U9581 ( .A(n7902), .ZN(n7803) );
  NOR2_X1 U9582 ( .A1(n7803), .A2(n7937), .ZN(n7806) );
  AOI22_X1 U9583 ( .A1(n7806), .A2(n7805), .B1(n7937), .B2(n7804), .ZN(n7907)
         );
  NOR3_X1 U9584 ( .A1(n7810), .A2(n7894), .A3(n9286), .ZN(n7807) );
  AOI21_X1 U9585 ( .B1(n9302), .B2(n7932), .A(n7807), .ZN(n7809) );
  NOR2_X1 U9586 ( .A1(n7809), .A2(n7808), .ZN(n7900) );
  NOR3_X1 U9587 ( .A1(n7810), .A2(n7894), .A3(n7932), .ZN(n7899) );
  INV_X1 U9588 ( .A(n7871), .ZN(n7870) );
  INV_X1 U9589 ( .A(n7840), .ZN(n7846) );
  AND4_X1 U9590 ( .A1(n7819), .A2(n7816), .A3(n7825), .A4(n7932), .ZN(n7811)
         );
  OAI21_X1 U9591 ( .B1(n7813), .B2(n7812), .A(n7811), .ZN(n7833) );
  INV_X1 U9592 ( .A(n7816), .ZN(n7817) );
  NAND3_X1 U9593 ( .A1(n7828), .A2(n7817), .A3(n7937), .ZN(n7818) );
  INV_X1 U9594 ( .A(n7820), .ZN(n7831) );
  INV_X1 U9595 ( .A(n7821), .ZN(n7824) );
  OAI211_X1 U9596 ( .C1(n6778), .C2(n7824), .A(n7823), .B(n7822), .ZN(n7826)
         );
  NAND3_X1 U9597 ( .A1(n7826), .A2(n4387), .A3(n7825), .ZN(n7829) );
  NAND4_X1 U9598 ( .A1(n7829), .A2(n7937), .A3(n7828), .A4(n7827), .ZN(n7830)
         );
  NAND2_X1 U9599 ( .A1(n7835), .A2(n7834), .ZN(n7837) );
  MUX2_X1 U9600 ( .A(n7837), .B(n7836), .S(n7932), .Z(n7838) );
  AND2_X1 U9601 ( .A1(n7840), .A2(n7839), .ZN(n7842) );
  MUX2_X1 U9602 ( .A(n7842), .B(n7841), .S(n7932), .Z(n7843) );
  INV_X1 U9603 ( .A(n7851), .ZN(n7845) );
  OAI21_X1 U9604 ( .B1(n7846), .B2(n7845), .A(n7844), .ZN(n7848) );
  NAND2_X1 U9605 ( .A1(n7848), .A2(n7847), .ZN(n7860) );
  NAND2_X1 U9606 ( .A1(n9682), .A2(n7852), .ZN(n7855) );
  OAI211_X1 U9607 ( .C1(n7856), .C2(n7855), .A(n7854), .B(n7853), .ZN(n7858)
         );
  NAND2_X1 U9608 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  INV_X1 U9609 ( .A(n7875), .ZN(n7864) );
  INV_X1 U9610 ( .A(n7861), .ZN(n7863) );
  OAI211_X1 U9611 ( .C1(n7864), .C2(n7863), .A(n7862), .B(n7874), .ZN(n7866)
         );
  NAND2_X1 U9612 ( .A1(n7866), .A2(n7865), .ZN(n7867) );
  NOR2_X1 U9613 ( .A1(n7868), .A2(n7867), .ZN(n7869) );
  MUX2_X1 U9614 ( .A(n7870), .B(n7869), .S(n7932), .Z(n7897) );
  AOI22_X1 U9615 ( .A1(n7877), .A2(n7871), .B1(n9035), .B2(n7937), .ZN(n7882)
         );
  AOI21_X1 U9616 ( .B1(n7872), .B2(n9046), .A(n7932), .ZN(n7881) );
  OAI211_X1 U9617 ( .C1(n7882), .C2(n7881), .A(n7880), .B(n9299), .ZN(n7896)
         );
  NOR2_X1 U9618 ( .A1(n9301), .A2(n7932), .ZN(n7885) );
  AOI22_X1 U9619 ( .A1(n9323), .A2(n7885), .B1(n8886), .B2(n7937), .ZN(n7891)
         );
  NAND2_X1 U9620 ( .A1(n9301), .A2(n7932), .ZN(n7884) );
  OAI22_X1 U9621 ( .A1(n9323), .A2(n7884), .B1(n8886), .B2(n7937), .ZN(n7883)
         );
  NAND2_X1 U9622 ( .A1(n9297), .A2(n7883), .ZN(n7890) );
  NOR2_X1 U9623 ( .A1(n7884), .A2(n8886), .ZN(n7888) );
  NAND2_X1 U9624 ( .A1(n7885), .A2(n8886), .ZN(n7886) );
  NAND2_X1 U9625 ( .A1(n9323), .A2(n7886), .ZN(n7887) );
  OAI21_X1 U9626 ( .B1(n9323), .B2(n7888), .A(n7887), .ZN(n7889) );
  OAI211_X1 U9627 ( .C1(n9297), .C2(n7891), .A(n7890), .B(n7889), .ZN(n7892)
         );
  NOR3_X1 U9628 ( .A1(n7894), .A2(n7893), .A3(n7892), .ZN(n7895) );
  OAI21_X1 U9629 ( .B1(n7897), .B2(n7896), .A(n7895), .ZN(n7898) );
  OAI21_X1 U9630 ( .B1(n7900), .B2(n7899), .A(n7898), .ZN(n7906) );
  INV_X1 U9631 ( .A(n7903), .ZN(n7905) );
  NAND3_X1 U9632 ( .A1(n7909), .A2(n9199), .A3(n4970), .ZN(n7913) );
  MUX2_X1 U9633 ( .A(n7911), .B(n7910), .S(n7932), .Z(n7912) );
  NAND2_X1 U9634 ( .A1(n7913), .A2(n7912), .ZN(n7922) );
  OAI21_X1 U9635 ( .B1(n7916), .B2(n7915), .A(n7914), .ZN(n7918) );
  INV_X1 U9636 ( .A(n7925), .ZN(n9146) );
  INV_X1 U9637 ( .A(n7927), .ZN(n7928) );
  INV_X1 U9638 ( .A(n7929), .ZN(n7930) );
  MUX2_X1 U9639 ( .A(n7937), .B(n7939), .S(n9135), .Z(n7943) );
  NAND2_X1 U9640 ( .A1(n4790), .A2(n9036), .ZN(n7942) );
  NAND2_X1 U9641 ( .A1(n7937), .A2(n9135), .ZN(n7938) );
  OAI21_X1 U9642 ( .B1(n7939), .B2(n9135), .A(n7938), .ZN(n7940) );
  NAND2_X1 U9643 ( .A1(n9125), .A2(n9036), .ZN(n7990) );
  NAND3_X1 U9644 ( .A1(n7940), .A2(n7990), .A3(n7993), .ZN(n7941) );
  AOI22_X1 U9645 ( .A1(n8002), .A2(n7944), .B1(n9747), .B2(n5720), .ZN(n7999)
         );
  INV_X1 U9646 ( .A(n8004), .ZN(n7981) );
  XNOR2_X1 U9647 ( .A(n9386), .B(n9278), .ZN(n9258) );
  INV_X1 U9648 ( .A(n7945), .ZN(n9728) );
  AND2_X1 U9649 ( .A1(n9728), .A2(n7946), .ZN(n9758) );
  NAND4_X1 U9650 ( .A1(n7948), .A2(n7947), .A3(n9758), .A4(n5720), .ZN(n7952)
         );
  OR2_X1 U9651 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  NOR2_X1 U9652 ( .A1(n7952), .A2(n7951), .ZN(n7956) );
  INV_X1 U9653 ( .A(n9727), .ZN(n7953) );
  NOR2_X1 U9654 ( .A1(n7954), .A2(n7953), .ZN(n7955) );
  NAND4_X1 U9655 ( .A1(n9699), .A2(n7957), .A3(n7956), .A4(n7955), .ZN(n7958)
         );
  NOR4_X1 U9656 ( .A1(n9667), .A2(n9678), .A3(n7958), .A4(n6499), .ZN(n7959)
         );
  NAND2_X1 U9657 ( .A1(n7960), .A2(n7959), .ZN(n7961) );
  OR4_X1 U9658 ( .A1(n9324), .A2(n7963), .A3(n7962), .A4(n7961), .ZN(n7964) );
  NOR2_X1 U9659 ( .A1(n9328), .A2(n7964), .ZN(n7965) );
  NAND4_X1 U9660 ( .A1(n9258), .A2(n9276), .A3(n9299), .A4(n7965), .ZN(n7966)
         );
  NOR2_X1 U9661 ( .A1(n9242), .A2(n7966), .ZN(n7967) );
  NAND3_X1 U9662 ( .A1(n9218), .A2(n9224), .A3(n7967), .ZN(n7968) );
  OR4_X1 U9663 ( .A1(n7970), .A2(n9190), .A3(n7969), .A4(n7968), .ZN(n7973) );
  OR4_X1 U9664 ( .A1(n7973), .A2(n7972), .A3(n7971), .A4(n9145), .ZN(n7974) );
  NOR2_X1 U9665 ( .A1(n7981), .A2(n7974), .ZN(n7979) );
  INV_X1 U9666 ( .A(n7993), .ZN(n8006) );
  NAND2_X1 U9667 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  NOR2_X1 U9668 ( .A1(n8006), .A2(n7977), .ZN(n7978) );
  NOR2_X1 U9669 ( .A1(n7981), .A2(n7980), .ZN(n7996) );
  OAI21_X1 U9670 ( .B1(n7984), .B2(n7983), .A(n7982), .ZN(n7986) );
  AOI21_X1 U9671 ( .B1(n7987), .B2(n7986), .A(n7985), .ZN(n7988) );
  NOR2_X1 U9672 ( .A1(n7989), .A2(n7988), .ZN(n7992) );
  OAI22_X1 U9673 ( .A1(n7992), .A2(n7991), .B1(n9135), .B2(n7990), .ZN(n7994)
         );
  OAI211_X1 U9674 ( .C1(n9339), .C2(n9125), .A(n7994), .B(n7993), .ZN(n7995)
         );
  AOI21_X1 U9675 ( .B1(n7996), .B2(n7995), .A(n7998), .ZN(n7997) );
  OAI21_X1 U9676 ( .B1(n8004), .B2(n8003), .A(n8002), .ZN(n8011) );
  AOI211_X1 U9677 ( .C1(n8006), .C2(n9747), .A(n5096), .B(n8005), .ZN(n8010)
         );
  INV_X1 U9678 ( .A(n8007), .ZN(n8009) );
  NOR3_X1 U9679 ( .A1(n9743), .A2(n9423), .A3(n8012), .ZN(n8014) );
  OAI21_X1 U9680 ( .B1(n8015), .B2(n5096), .A(P1_B_REG_SCAN_IN), .ZN(n8013) );
  OAI222_X1 U9681 ( .A1(n8019), .A2(n8018), .B1(n8017), .B2(n8016), .C1(n8503), 
        .C2(P2_U3151), .ZN(P2_U3268) );
  INV_X1 U9682 ( .A(n8020), .ZN(n8022) );
  OAI222_X1 U9683 ( .A1(n8023), .A2(n8022), .B1(n5737), .B2(P1_U3086), .C1(
        n8021), .C2(n9438), .ZN(P1_U3327) );
  AND2_X1 U9684 ( .A1(n8027), .A2(n8344), .ZN(n8215) );
  NOR2_X1 U9685 ( .A1(n5824), .A2(n8862), .ZN(n8024) );
  INV_X1 U9686 ( .A(n8786), .ZN(n8032) );
  NAND2_X1 U9687 ( .A1(n8786), .A2(n8343), .ZN(n8220) );
  OAI21_X1 U9688 ( .B1(n8027), .B2(n8032), .A(n8220), .ZN(n8030) );
  INV_X1 U9689 ( .A(n8027), .ZN(n8787) );
  INV_X1 U9690 ( .A(n8344), .ZN(n8028) );
  NAND2_X1 U9691 ( .A1(n8787), .A2(n8028), .ZN(n8216) );
  NAND2_X1 U9692 ( .A1(n8216), .A2(n8029), .ZN(n8212) );
  INV_X1 U9693 ( .A(n8343), .ZN(n8031) );
  NAND2_X1 U9694 ( .A1(n8032), .A2(n8031), .ZN(n8217) );
  AND2_X1 U9695 ( .A1(n6296), .A2(n8217), .ZN(n8061) );
  INV_X1 U9696 ( .A(n8217), .ZN(n8060) );
  INV_X1 U9697 ( .A(n8220), .ZN(n8057) );
  INV_X1 U9698 ( .A(n8215), .ZN(n8034) );
  NAND2_X1 U9699 ( .A1(n8034), .A2(n8033), .ZN(n8211) );
  INV_X1 U9700 ( .A(n8560), .ZN(n8201) );
  NAND2_X1 U9701 ( .A1(n8195), .A2(n8197), .ZN(n8569) );
  NOR2_X1 U9702 ( .A1(n8569), .A2(n8585), .ZN(n8193) );
  NAND2_X1 U9703 ( .A1(n8189), .A2(n8185), .ZN(n8597) );
  NAND2_X1 U9704 ( .A1(n8183), .A2(n8596), .ZN(n8603) );
  INV_X1 U9705 ( .A(n8621), .ZN(n8052) );
  INV_X1 U9706 ( .A(n8096), .ZN(n8036) );
  NOR4_X1 U9707 ( .A1(n8036), .A2(n8035), .A3(n6213), .A4(n8082), .ZN(n8039)
         );
  AND2_X1 U9708 ( .A1(n4959), .A2(n8071), .ZN(n8103) );
  NAND4_X1 U9709 ( .A1(n8039), .A2(n8103), .A3(n8038), .A4(n8037), .ZN(n8043)
         );
  NOR4_X1 U9710 ( .A1(n8043), .A2(n8042), .A3(n8041), .A4(n8040), .ZN(n8044)
         );
  AND4_X1 U9711 ( .A1(n8047), .A2(n8046), .A3(n8045), .A4(n8044), .ZN(n8048)
         );
  NAND4_X1 U9712 ( .A1(n8146), .A2(n8135), .A3(n8049), .A4(n8048), .ZN(n8050)
         );
  NOR4_X1 U9713 ( .A1(n8679), .A2(n8150), .A3(n8697), .A4(n8050), .ZN(n8051)
         );
  NAND4_X1 U9714 ( .A1(n8640), .A2(n8052), .A3(n8654), .A4(n8051), .ZN(n8053)
         );
  NOR4_X1 U9715 ( .A1(n8597), .A2(n8603), .A3(n8177), .A4(n8053), .ZN(n8054)
         );
  NAND4_X1 U9716 ( .A1(n8055), .A2(n8201), .A3(n8193), .A4(n8054), .ZN(n8056)
         );
  NOR4_X1 U9717 ( .A1(n8057), .A2(n8211), .A3(n8212), .A4(n8056), .ZN(n8058)
         );
  NAND2_X1 U9718 ( .A1(n8058), .A2(n8072), .ZN(n8059) );
  XNOR2_X1 U9719 ( .A(n8063), .B(n8062), .ZN(n8225) );
  INV_X1 U9720 ( .A(n8064), .ZN(n8067) );
  NAND2_X1 U9721 ( .A1(n8183), .A2(n8065), .ZN(n8066) );
  MUX2_X1 U9722 ( .A(n8067), .B(n8066), .S(n8219), .Z(n8068) );
  INV_X1 U9723 ( .A(n8068), .ZN(n8182) );
  NAND2_X1 U9724 ( .A1(n8179), .A2(n8173), .ZN(n8070) );
  NAND2_X1 U9725 ( .A1(n8178), .A2(n8169), .ZN(n8069) );
  MUX2_X1 U9726 ( .A(n8070), .B(n8069), .S(n8219), .Z(n8181) );
  NAND2_X1 U9727 ( .A1(n6305), .A2(n8072), .ZN(n8073) );
  NAND2_X1 U9728 ( .A1(n8073), .A2(n8076), .ZN(n8074) );
  NAND2_X1 U9729 ( .A1(n8074), .A2(n8081), .ZN(n8075) );
  NAND3_X1 U9730 ( .A1(n8075), .A2(n8206), .A3(n8077), .ZN(n8080) );
  NAND2_X1 U9731 ( .A1(n8077), .A2(n8076), .ZN(n8078) );
  NAND2_X1 U9732 ( .A1(n8078), .A2(n8219), .ZN(n8079) );
  NAND2_X1 U9733 ( .A1(n8080), .A2(n8079), .ZN(n8085) );
  INV_X1 U9734 ( .A(n8081), .ZN(n8083) );
  AOI21_X1 U9735 ( .B1(n8083), .B2(n8219), .A(n8082), .ZN(n8084) );
  NAND2_X1 U9736 ( .A1(n8085), .A2(n8084), .ZN(n8090) );
  AOI21_X1 U9737 ( .B1(n8090), .B2(n8089), .A(n8088), .ZN(n8098) );
  INV_X1 U9738 ( .A(n8098), .ZN(n8094) );
  INV_X1 U9739 ( .A(n8091), .ZN(n8093) );
  OAI211_X1 U9740 ( .C1(n8094), .C2(n8093), .A(n8103), .B(n8092), .ZN(n8095)
         );
  OAI21_X1 U9741 ( .B1(n4685), .B2(n8096), .A(n8095), .ZN(n8106) );
  NAND2_X1 U9742 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  OAI211_X1 U9743 ( .C1(n6312), .C2(n8100), .A(n8099), .B(n9922), .ZN(n8104)
         );
  INV_X1 U9744 ( .A(n8101), .ZN(n8102) );
  AOI21_X1 U9745 ( .B1(n8104), .B2(n8103), .A(n8102), .ZN(n8105) );
  AND2_X1 U9746 ( .A1(n8113), .A2(n8107), .ZN(n8110) );
  INV_X1 U9747 ( .A(n8117), .ZN(n8108) );
  AND2_X1 U9748 ( .A1(n8108), .A2(n8118), .ZN(n8109) );
  MUX2_X1 U9749 ( .A(n8110), .B(n8109), .S(n8206), .Z(n8112) );
  INV_X1 U9750 ( .A(n8112), .ZN(n8120) );
  OAI211_X1 U9751 ( .C1(n8120), .C2(n8114), .A(n8113), .B(n8125), .ZN(n8122)
         );
  INV_X1 U9752 ( .A(n8115), .ZN(n8116) );
  NOR2_X1 U9753 ( .A1(n8117), .A2(n8116), .ZN(n8119) );
  OAI211_X1 U9754 ( .C1(n8120), .C2(n8119), .A(n8118), .B(n8123), .ZN(n8121)
         );
  NAND2_X1 U9755 ( .A1(n8124), .A2(n8126), .ZN(n8131) );
  NAND3_X1 U9756 ( .A1(n8127), .A2(n8126), .A3(n8125), .ZN(n8129) );
  NAND2_X1 U9757 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  MUX2_X1 U9758 ( .A(n8131), .B(n8130), .S(n8219), .Z(n8137) );
  MUX2_X1 U9759 ( .A(n8133), .B(n8132), .S(n8206), .Z(n8134) );
  INV_X1 U9760 ( .A(n8138), .ZN(n8140) );
  MUX2_X1 U9761 ( .A(n8140), .B(n8139), .S(n8206), .Z(n8141) );
  MUX2_X1 U9762 ( .A(n8144), .B(n8143), .S(n8219), .Z(n8145) );
  NAND3_X1 U9763 ( .A1(n8156), .A2(n8153), .A3(n8147), .ZN(n8149) );
  NAND3_X1 U9764 ( .A1(n8149), .A2(n8219), .A3(n8148), .ZN(n8151) );
  NAND2_X1 U9765 ( .A1(n8151), .A2(n8684), .ZN(n8159) );
  NAND2_X1 U9766 ( .A1(n8160), .A2(n8677), .ZN(n8152) );
  NAND2_X1 U9767 ( .A1(n8152), .A2(n8219), .ZN(n8158) );
  NAND2_X1 U9768 ( .A1(n8153), .A2(n8206), .ZN(n8154) );
  AOI21_X1 U9769 ( .B1(n8156), .B2(n8155), .A(n8154), .ZN(n8157) );
  AOI21_X1 U9770 ( .B1(n8159), .B2(n8158), .A(n8157), .ZN(n8164) );
  NAND3_X1 U9771 ( .A1(n8164), .A2(n8654), .A3(n8166), .ZN(n8162) );
  NAND2_X1 U9772 ( .A1(n8170), .A2(n8160), .ZN(n8161) );
  MUX2_X1 U9773 ( .A(n8162), .B(n8161), .S(n8206), .Z(n8163) );
  INV_X1 U9774 ( .A(n8164), .ZN(n8167) );
  NAND2_X1 U9775 ( .A1(n8169), .A2(n8168), .ZN(n8172) );
  INV_X1 U9776 ( .A(n8170), .ZN(n8171) );
  MUX2_X1 U9777 ( .A(n8172), .B(n8171), .S(n8219), .Z(n8175) );
  INV_X1 U9778 ( .A(n8173), .ZN(n8174) );
  NOR2_X1 U9779 ( .A1(n8175), .A2(n8174), .ZN(n8176) );
  MUX2_X1 U9780 ( .A(n8179), .B(n8178), .S(n8206), .Z(n8180) );
  INV_X1 U9781 ( .A(n8596), .ZN(n8184) );
  OAI211_X1 U9782 ( .C1(n8188), .C2(n8184), .A(n8189), .B(n8183), .ZN(n8186)
         );
  NAND2_X1 U9783 ( .A1(n8186), .A2(n8185), .ZN(n8192) );
  NAND2_X1 U9784 ( .A1(n8188), .A2(n8187), .ZN(n8190) );
  NAND2_X1 U9785 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  INV_X1 U9786 ( .A(n8194), .ZN(n8196) );
  OAI21_X1 U9787 ( .B1(n8569), .B2(n8196), .A(n8195), .ZN(n8200) );
  OAI21_X1 U9788 ( .B1(n8569), .B2(n8198), .A(n8197), .ZN(n8199) );
  MUX2_X1 U9789 ( .A(n8200), .B(n8199), .S(n8219), .Z(n8202) );
  MUX2_X1 U9790 ( .A(n8204), .B(n8203), .S(n8206), .Z(n8205) );
  MUX2_X1 U9791 ( .A(n8555), .B(n8547), .S(n8206), .Z(n8210) );
  INV_X1 U9792 ( .A(n8210), .ZN(n8208) );
  MUX2_X1 U9793 ( .A(n8555), .B(n8547), .S(n8219), .Z(n8207) );
  AOI21_X1 U9794 ( .B1(n8219), .B2(n8216), .A(n8215), .ZN(n8218) );
  AOI21_X1 U9795 ( .B1(n8225), .B2(n8224), .A(n8223), .ZN(n8232) );
  NAND3_X1 U9796 ( .A1(n8227), .A2(n8226), .A3(n8503), .ZN(n8228) );
  OAI211_X1 U9797 ( .C1(n8229), .C2(n8231), .A(n8228), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8230) );
  OAI21_X1 U9798 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(P2_U3296) );
  INV_X1 U9799 ( .A(n8855), .ZN(n8710) );
  OAI21_X1 U9800 ( .B1(n8235), .B2(n8234), .A(n8233), .ZN(n8236) );
  NAND2_X1 U9801 ( .A1(n8236), .A2(n8315), .ZN(n8242) );
  INV_X1 U9802 ( .A(n8708), .ZN(n8240) );
  NOR2_X1 U9803 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4577), .ZN(n8401) );
  AOI21_X1 U9804 ( .B1(n8318), .B2(n8699), .A(n8401), .ZN(n8237) );
  OAI21_X1 U9805 ( .B1(n8238), .B2(n8320), .A(n8237), .ZN(n8239) );
  AOI21_X1 U9806 ( .B1(n8240), .B2(n8323), .A(n8239), .ZN(n8241) );
  OAI211_X1 U9807 ( .C1(n8710), .C2(n8341), .A(n8242), .B(n8241), .ZN(P2_U3155) );
  INV_X1 U9809 ( .A(n8245), .ZN(n8280) );
  AOI21_X1 U9810 ( .B1(n8591), .B2(n8243), .A(n8280), .ZN(n8252) );
  AOI22_X1 U9811 ( .A1(n8623), .A2(n8338), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8247) );
  NAND2_X1 U9812 ( .A1(n8608), .A2(n8323), .ZN(n8246) );
  OAI211_X1 U9813 ( .C1(n8248), .C2(n8335), .A(n8247), .B(n8246), .ZN(n8249)
         );
  AOI21_X1 U9814 ( .B1(n8815), .B2(n8250), .A(n8249), .ZN(n8251) );
  OAI21_X1 U9815 ( .B1(n8252), .B2(n8327), .A(n8251), .ZN(P2_U3156) );
  INV_X1 U9816 ( .A(n8769), .ZN(n8835) );
  AND3_X1 U9817 ( .A1(n8311), .A2(n8254), .A3(n8253), .ZN(n8255) );
  OAI21_X1 U9818 ( .B1(n8293), .B2(n8255), .A(n8315), .ZN(n8259) );
  NAND2_X1 U9819 ( .A1(n8624), .A2(n8318), .ZN(n8256) );
  NAND2_X1 U9820 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8535) );
  OAI211_X1 U9821 ( .C1(n8658), .C2(n8320), .A(n8256), .B(n8535), .ZN(n8257)
         );
  AOI21_X1 U9822 ( .B1(n8664), .B2(n8323), .A(n8257), .ZN(n8258) );
  OAI211_X1 U9823 ( .C1(n8835), .C2(n8341), .A(n8259), .B(n8258), .ZN(P2_U3159) );
  INV_X1 U9824 ( .A(n8825), .ZN(n8268) );
  AND3_X1 U9825 ( .A1(n8290), .A2(n8261), .A3(n8260), .ZN(n8262) );
  OAI21_X1 U9826 ( .B1(n8303), .B2(n8262), .A(n8315), .ZN(n8267) );
  NOR2_X1 U9827 ( .A1(n8320), .A2(n8659), .ZN(n8265) );
  OAI22_X1 U9828 ( .A1(n8263), .A2(n8335), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10077), .ZN(n8264) );
  AOI211_X1 U9829 ( .C1(n8627), .C2(n8323), .A(n8265), .B(n8264), .ZN(n8266)
         );
  OAI211_X1 U9830 ( .C1(n8268), .C2(n8341), .A(n8267), .B(n8266), .ZN(P2_U3163) );
  INV_X1 U9831 ( .A(n8842), .ZN(n8276) );
  NOR2_X1 U9832 ( .A1(n8270), .A2(n8269), .ZN(n8271) );
  OAI21_X1 U9833 ( .B1(n8271), .B2(n8314), .A(n8315), .ZN(n8275) );
  NOR2_X1 U9834 ( .A1(n8333), .A2(n8690), .ZN(n8273) );
  NAND2_X1 U9835 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8473) );
  OAI21_X1 U9836 ( .B1(n8335), .B2(n8658), .A(n8473), .ZN(n8272) );
  AOI211_X1 U9837 ( .C1(n8338), .C2(n8686), .A(n8273), .B(n8272), .ZN(n8274)
         );
  OAI211_X1 U9838 ( .C1(n8276), .C2(n8341), .A(n8275), .B(n8274), .ZN(P2_U3168) );
  INV_X1 U9839 ( .A(n8809), .ZN(n8289) );
  INV_X1 U9840 ( .A(n8277), .ZN(n8279) );
  NOR3_X1 U9841 ( .A1(n8280), .A2(n8279), .A3(n8278), .ZN(n8283) );
  INV_X1 U9842 ( .A(n8281), .ZN(n8282) );
  OAI21_X1 U9843 ( .B1(n8283), .B2(n8282), .A(n8315), .ZN(n8288) );
  AOI22_X1 U9844 ( .A1(n8591), .A2(n8338), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8284) );
  OAI21_X1 U9845 ( .B1(n8285), .B2(n8335), .A(n8284), .ZN(n8286) );
  AOI21_X1 U9846 ( .B1(n8593), .B2(n8323), .A(n8286), .ZN(n8287) );
  OAI211_X1 U9847 ( .C1(n8289), .C2(n8341), .A(n8288), .B(n8287), .ZN(P2_U3169) );
  INV_X1 U9848 ( .A(n8831), .ZN(n8645) );
  INV_X1 U9849 ( .A(n8290), .ZN(n8295) );
  NOR3_X1 U9850 ( .A1(n8293), .A2(n8292), .A3(n8291), .ZN(n8294) );
  OAI21_X1 U9851 ( .B1(n8295), .B2(n8294), .A(n8315), .ZN(n8299) );
  AOI22_X1 U9852 ( .A1(n8346), .A2(n8318), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8296) );
  OAI21_X1 U9853 ( .B1(n8636), .B2(n8320), .A(n8296), .ZN(n8297) );
  AOI21_X1 U9854 ( .B1(n8643), .B2(n8323), .A(n8297), .ZN(n8298) );
  OAI211_X1 U9855 ( .C1(n8645), .C2(n8341), .A(n8299), .B(n8298), .ZN(P2_U3173) );
  INV_X1 U9856 ( .A(n8756), .ZN(n8310) );
  INV_X1 U9857 ( .A(n8300), .ZN(n8305) );
  NOR3_X1 U9858 ( .A1(n8303), .A2(n8302), .A3(n8301), .ZN(n8304) );
  OAI21_X1 U9859 ( .B1(n8305), .B2(n8304), .A(n8315), .ZN(n8309) );
  AOI22_X1 U9860 ( .A1(n8346), .A2(n8338), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8306) );
  OAI21_X1 U9861 ( .B1(n6368), .B2(n8335), .A(n8306), .ZN(n8307) );
  AOI21_X1 U9862 ( .B1(n8615), .B2(n8323), .A(n8307), .ZN(n8308) );
  OAI211_X1 U9863 ( .C1(n8310), .C2(n8341), .A(n8309), .B(n8308), .ZN(P2_U3175) );
  INV_X1 U9864 ( .A(n8673), .ZN(n8776) );
  INV_X1 U9865 ( .A(n8311), .ZN(n8317) );
  NOR3_X1 U9866 ( .A1(n8314), .A2(n8313), .A3(n8312), .ZN(n8316) );
  OAI21_X1 U9867 ( .B1(n8317), .B2(n8316), .A(n8315), .ZN(n8325) );
  NAND2_X1 U9868 ( .A1(n8318), .A2(n8667), .ZN(n8319) );
  NAND2_X1 U9869 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8513) );
  OAI211_X1 U9870 ( .C1(n8321), .C2(n8320), .A(n8319), .B(n8513), .ZN(n8322)
         );
  AOI21_X1 U9871 ( .B1(n8669), .B2(n8323), .A(n8322), .ZN(n8324) );
  OAI211_X1 U9872 ( .C1(n8776), .C2(n8341), .A(n8325), .B(n8324), .ZN(P2_U3178) );
  INV_X1 U9873 ( .A(n8326), .ZN(n8342) );
  AOI21_X1 U9874 ( .B1(n8329), .B2(n8328), .A(n8327), .ZN(n8331) );
  NAND2_X1 U9875 ( .A1(n8331), .A2(n8330), .ZN(n8340) );
  NOR2_X1 U9876 ( .A1(n8333), .A2(n8332), .ZN(n8337) );
  NAND2_X1 U9877 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8428) );
  OAI21_X1 U9878 ( .B1(n8335), .B2(n8334), .A(n8428), .ZN(n8336) );
  AOI211_X1 U9879 ( .C1(n8338), .C2(n8347), .A(n8337), .B(n8336), .ZN(n8339)
         );
  OAI211_X1 U9880 ( .C1(n8342), .C2(n8341), .A(n8340), .B(n8339), .ZN(P2_U3181) );
  MUX2_X1 U9881 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8343), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9882 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8344), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9883 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8345), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9884 ( .A(n8555), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8507), .Z(
        P2_U3519) );
  MUX2_X1 U9885 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8571), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9886 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8579), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9887 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8590), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9888 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8605), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9889 ( .A(n8591), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8507), .Z(
        P2_U3514) );
  MUX2_X1 U9890 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8623), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9891 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8346), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9892 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8624), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9893 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8667), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9894 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8687), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9895 ( .A(n8700), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8507), .Z(
        P2_U3508) );
  MUX2_X1 U9896 ( .A(n8686), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8507), .Z(
        P2_U3507) );
  MUX2_X1 U9897 ( .A(n8699), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8507), .Z(
        P2_U3506) );
  MUX2_X1 U9898 ( .A(n8347), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8507), .Z(
        P2_U3505) );
  MUX2_X1 U9899 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8348), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9900 ( .A(n8349), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8507), .Z(
        P2_U3503) );
  MUX2_X1 U9901 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8350), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9902 ( .A(n8351), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8507), .Z(
        P2_U3501) );
  MUX2_X1 U9903 ( .A(n8352), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8507), .Z(
        P2_U3500) );
  MUX2_X1 U9904 ( .A(n8353), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8507), .Z(
        P2_U3499) );
  MUX2_X1 U9905 ( .A(n9931), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8507), .Z(
        P2_U3498) );
  MUX2_X1 U9906 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8354), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9907 ( .A(n9932), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8507), .Z(
        P2_U3496) );
  MUX2_X1 U9908 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8355), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9909 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8356), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9910 ( .A(n8357), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8507), .Z(
        P2_U3493) );
  INV_X1 U9911 ( .A(n8358), .ZN(n8359) );
  MUX2_X1 U9912 ( .A(n8362), .B(n8382), .S(n8503), .Z(n8364) );
  AND2_X1 U9913 ( .A1(n8364), .A2(n8387), .ZN(n8398) );
  INV_X1 U9914 ( .A(n8398), .ZN(n8363) );
  OAI21_X1 U9915 ( .B1(n8387), .B2(n8364), .A(n8363), .ZN(n8365) );
  AOI21_X1 U9916 ( .B1(n8366), .B2(n8365), .A(n4430), .ZN(n8389) );
  AOI21_X1 U9917 ( .B1(n8370), .B2(n8362), .A(n8405), .ZN(n8375) );
  INV_X1 U9918 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8371) );
  OR2_X1 U9919 ( .A1(n9899), .A2(n8371), .ZN(n8374) );
  INV_X1 U9920 ( .A(n8372), .ZN(n8373) );
  OAI211_X1 U9921 ( .C1(n9896), .C2(n8375), .A(n8374), .B(n8373), .ZN(n8386)
         );
  NOR2_X1 U9922 ( .A1(n8377), .A2(n8376), .ZN(n8378) );
  NAND2_X1 U9923 ( .A1(n8381), .A2(n8380), .ZN(n8390) );
  OAI21_X1 U9924 ( .B1(n8381), .B2(n8380), .A(n8390), .ZN(n8383) );
  NOR2_X1 U9925 ( .A1(n8382), .A2(n8383), .ZN(n8391) );
  AOI21_X1 U9926 ( .B1(n8383), .B2(n8382), .A(n8391), .ZN(n8384) );
  NOR2_X1 U9927 ( .A1(n8384), .A2(n9889), .ZN(n8385) );
  AOI211_X1 U9928 ( .C1(n9891), .C2(n8387), .A(n8386), .B(n8385), .ZN(n8388)
         );
  OAI21_X1 U9929 ( .B1(n8389), .B2(n8509), .A(n8388), .ZN(P2_U3195) );
  INV_X1 U9930 ( .A(n8390), .ZN(n8392) );
  AOI22_X1 U9931 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8413), .B1(n8431), .B2(
        n8395), .ZN(n8393) );
  AOI21_X1 U9932 ( .B1(n8394), .B2(n8393), .A(n8416), .ZN(n8415) );
  MUX2_X1 U9933 ( .A(n8407), .B(n8395), .S(n8503), .Z(n8397) );
  AND2_X1 U9934 ( .A1(n8397), .A2(n8413), .ZN(n8423) );
  INV_X1 U9935 ( .A(n8423), .ZN(n8396) );
  OAI21_X1 U9936 ( .B1(n8413), .B2(n8397), .A(n8396), .ZN(n8400) );
  AOI21_X1 U9937 ( .B1(n8400), .B2(n8399), .A(n8422), .ZN(n8404) );
  NAND2_X1 U9938 ( .A1(n9905), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8403) );
  INV_X1 U9939 ( .A(n8401), .ZN(n8402) );
  OAI211_X1 U9940 ( .C1(n8404), .C2(n8509), .A(n8403), .B(n8402), .ZN(n8412)
         );
  AOI22_X1 U9941 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8413), .B1(n8431), .B2(
        n8407), .ZN(n8408) );
  NOR2_X1 U9942 ( .A1(n8409), .A2(n8408), .ZN(n8430) );
  AOI21_X1 U9943 ( .B1(n8409), .B2(n8408), .A(n8430), .ZN(n8410) );
  NOR2_X1 U9944 ( .A1(n8410), .A2(n9896), .ZN(n8411) );
  AOI211_X1 U9945 ( .C1(n9891), .C2(n8413), .A(n8412), .B(n8411), .ZN(n8414)
         );
  OAI21_X1 U9946 ( .B1(n8415), .B2(n9889), .A(n8414), .ZN(P2_U3196) );
  NOR2_X1 U9947 ( .A1(n8418), .A2(n8417), .ZN(n8440) );
  AOI21_X1 U9948 ( .B1(n8418), .B2(n8417), .A(n8440), .ZN(n8438) );
  INV_X1 U9949 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8429) );
  MUX2_X1 U9950 ( .A(n8419), .B(n8418), .S(n8503), .Z(n8421) );
  AND2_X1 U9951 ( .A1(n8421), .A2(n8455), .ZN(n8445) );
  INV_X1 U9952 ( .A(n8445), .ZN(n8420) );
  OAI21_X1 U9953 ( .B1(n8455), .B2(n8421), .A(n8420), .ZN(n8425) );
  NOR2_X1 U9954 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  NOR2_X1 U9955 ( .A1(n8424), .A2(n8425), .ZN(n8444) );
  AOI21_X1 U9956 ( .B1(n8425), .B2(n8424), .A(n8444), .ZN(n8426) );
  OR2_X1 U9957 ( .A1(n8426), .A2(n8509), .ZN(n8427) );
  OAI211_X1 U9958 ( .C1(n9899), .C2(n8429), .A(n8428), .B(n8427), .ZN(n8436)
         );
  AOI21_X1 U9959 ( .B1(n8419), .B2(n8433), .A(n8456), .ZN(n8434) );
  NOR2_X1 U9960 ( .A1(n8434), .A2(n9896), .ZN(n8435) );
  AOI211_X1 U9961 ( .C1(n9891), .C2(n8455), .A(n8436), .B(n8435), .ZN(n8437)
         );
  OAI21_X1 U9962 ( .B1(n8438), .B2(n9889), .A(n8437), .ZN(P2_U3197) );
  NOR2_X1 U9963 ( .A1(n8455), .A2(n8439), .ZN(n8441) );
  NOR2_X1 U9964 ( .A1(n8441), .A2(n8440), .ZN(n8443) );
  AOI22_X1 U9965 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8450), .B1(n8471), .B2(
        n8779), .ZN(n8442) );
  AOI21_X1 U9966 ( .B1(n8443), .B2(n8442), .A(n8467), .ZN(n8466) );
  MUX2_X1 U9967 ( .A(n8702), .B(n8779), .S(n8503), .Z(n8446) );
  NAND2_X1 U9968 ( .A1(n8446), .A2(n8450), .ZN(n8477) );
  MUX2_X1 U9969 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8503), .Z(n8447) );
  AND2_X1 U9970 ( .A1(n8447), .A2(n8471), .ZN(n8479) );
  INV_X1 U9971 ( .A(n8479), .ZN(n8448) );
  NAND2_X1 U9972 ( .A1(n8477), .A2(n8448), .ZN(n8449) );
  XNOR2_X1 U9973 ( .A(n8478), .B(n8449), .ZN(n8464) );
  INV_X1 U9974 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U9975 ( .A1(n9891), .A2(n8450), .ZN(n8452) );
  OAI211_X1 U9976 ( .C1(n8453), .C2(n9899), .A(n8452), .B(n8451), .ZN(n8463)
         );
  NOR2_X1 U9977 ( .A1(n8455), .A2(n8454), .ZN(n8457) );
  NAND2_X1 U9978 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8471), .ZN(n8458) );
  OAI21_X1 U9979 ( .B1(n8471), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8458), .ZN(
        n8459) );
  AOI21_X1 U9980 ( .B1(n8460), .B2(n8459), .A(n8470), .ZN(n8461) );
  NOR2_X1 U9981 ( .A1(n8461), .A2(n9896), .ZN(n8462) );
  AOI211_X1 U9982 ( .C1(n9906), .C2(n8464), .A(n8463), .B(n8462), .ZN(n8465)
         );
  OAI21_X1 U9983 ( .B1(n8466), .B2(n9889), .A(n8465), .ZN(P2_U3198) );
  AOI21_X1 U9984 ( .B1(n10071), .B2(n8468), .A(n8488), .ZN(n8486) );
  INV_X1 U9985 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8469) );
  NOR2_X1 U9986 ( .A1(n9899), .A2(n8469), .ZN(n8476) );
  AOI21_X1 U9987 ( .B1(n8472), .B2(n8689), .A(n8493), .ZN(n8474) );
  OAI21_X1 U9988 ( .B1(n9896), .B2(n8474), .A(n8473), .ZN(n8475) );
  AOI211_X1 U9989 ( .C1(n9891), .C2(n8501), .A(n8476), .B(n8475), .ZN(n8485)
         );
  OAI21_X1 U9990 ( .B1(n8479), .B2(n8478), .A(n8477), .ZN(n8482) );
  MUX2_X1 U9991 ( .A(n8689), .B(n10071), .S(n8503), .Z(n8502) );
  XNOR2_X1 U9992 ( .A(n8480), .B(n8502), .ZN(n8481) );
  OAI21_X1 U9993 ( .B1(n8482), .B2(n8481), .A(n8500), .ZN(n8483) );
  NAND2_X1 U9994 ( .A1(n8483), .A2(n9906), .ZN(n8484) );
  OAI211_X1 U9995 ( .C1(n8486), .C2(n9889), .A(n8485), .B(n8484), .ZN(P2_U3199) );
  NOR2_X1 U9996 ( .A1(n8501), .A2(n8487), .ZN(n8489) );
  NAND2_X1 U9997 ( .A1(n8511), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8518) );
  OAI21_X1 U9998 ( .B1(n8511), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8518), .ZN(
        n8490) );
  NOR2_X1 U9999 ( .A1(n8491), .A2(n8490), .ZN(n8520) );
  AOI21_X1 U10000 ( .B1(n8491), .B2(n8490), .A(n8520), .ZN(n8517) );
  NOR2_X1 U10001 ( .A1(n8501), .A2(n8492), .ZN(n8494) );
  NOR2_X1 U10002 ( .A1(n8494), .A2(n8493), .ZN(n8496) );
  INV_X1 U10003 ( .A(n8496), .ZN(n8499) );
  NAND2_X1 U10004 ( .A1(n8511), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8523) );
  OAI21_X1 U10005 ( .B1(n8511), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8523), .ZN(
        n8495) );
  INV_X1 U10006 ( .A(n8495), .ZN(n8498) );
  NOR2_X1 U10007 ( .A1(n8496), .A2(n8495), .ZN(n8525) );
  INV_X1 U10008 ( .A(n8525), .ZN(n8497) );
  MUX2_X1 U10009 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8503), .Z(n8504) );
  INV_X1 U10010 ( .A(n8529), .ZN(n8506) );
  NAND2_X1 U10011 ( .A1(n8505), .A2(n8504), .ZN(n8527) );
  INV_X1 U10012 ( .A(n8508), .ZN(n8510) );
  NOR2_X1 U10013 ( .A1(n8510), .A2(n8509), .ZN(n8512) );
  INV_X1 U10014 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10017) );
  OAI21_X1 U10015 ( .B1(n9899), .B2(n10017), .A(n8513), .ZN(n8514) );
  OAI21_X1 U10016 ( .B1(n8517), .B2(n9889), .A(n8516), .ZN(P2_U3200) );
  INV_X1 U10017 ( .A(n8518), .ZN(n8519) );
  NOR2_X1 U10018 ( .A1(n8520), .A2(n8519), .ZN(n8522) );
  XNOR2_X1 U10019 ( .A(n8539), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8532) );
  INV_X1 U10020 ( .A(n8532), .ZN(n8521) );
  XNOR2_X1 U10021 ( .A(n8522), .B(n8521), .ZN(n8543) );
  INV_X1 U10022 ( .A(n8523), .ZN(n8524) );
  XNOR2_X1 U10023 ( .A(n8539), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8531) );
  XNOR2_X1 U10024 ( .A(n8526), .B(n8531), .ZN(n8541) );
  OAI21_X1 U10025 ( .B1(n8529), .B2(n8528), .A(n8527), .ZN(n8534) );
  MUX2_X1 U10026 ( .A(n8532), .B(n8531), .S(n8530), .Z(n8533) );
  XNOR2_X1 U10027 ( .A(n8534), .B(n8533), .ZN(n8537) );
  OAI21_X1 U10028 ( .B1(n9899), .B2(n4837), .A(n8535), .ZN(n8536) );
  AOI21_X1 U10029 ( .B1(n8537), .B2(n9906), .A(n8536), .ZN(n8538) );
  OAI21_X1 U10030 ( .B1(n8539), .B2(n9913), .A(n8538), .ZN(n8540) );
  AOI21_X1 U10031 ( .B1(n8541), .B2(n9919), .A(n8540), .ZN(n8542) );
  OAI21_X1 U10032 ( .B1(n8543), .B2(n9889), .A(n8542), .ZN(P2_U3201) );
  NAND2_X1 U10033 ( .A1(n8713), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8544) );
  OAI211_X1 U10034 ( .C1(n8786), .C2(n9939), .A(n8545), .B(n8544), .ZN(
        P2_U3202) );
  AOI22_X1 U10035 ( .A1(n8546), .A2(n8729), .B1(n8713), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10036 ( .A1(n8547), .A2(n8705), .ZN(n8548) );
  OAI211_X1 U10037 ( .C1(n8550), .C2(n9943), .A(n8549), .B(n8548), .ZN(n8551)
         );
  INV_X1 U10038 ( .A(n8551), .ZN(n8552) );
  OAI21_X1 U10039 ( .B1(n8553), .B2(n8713), .A(n8552), .ZN(P2_U3205) );
  OAI21_X1 U10040 ( .B1(n8554), .B2(n8560), .A(n6149), .ZN(n8559) );
  NAND2_X1 U10041 ( .A1(n8555), .A2(n9930), .ZN(n8556) );
  OAI21_X1 U10042 ( .B1(n8557), .B2(n8720), .A(n8556), .ZN(n8558) );
  AOI21_X1 U10043 ( .B1(n8559), .B2(n9928), .A(n8558), .ZN(n8740) );
  XNOR2_X1 U10044 ( .A(n8561), .B(n8560), .ZN(n8795) );
  INV_X1 U10045 ( .A(n8795), .ZN(n8566) );
  AOI22_X1 U10046 ( .A1(n8562), .A2(n8729), .B1(n8713), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8563) );
  OAI21_X1 U10047 ( .B1(n8564), .B2(n9939), .A(n8563), .ZN(n8565) );
  AOI21_X1 U10048 ( .B1(n8566), .B2(n8681), .A(n8565), .ZN(n8567) );
  OAI21_X1 U10049 ( .B1(n8740), .B2(n8713), .A(n8567), .ZN(P2_U3206) );
  XNOR2_X1 U10050 ( .A(n8568), .B(n8569), .ZN(n8801) );
  INV_X1 U10051 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8573) );
  XNOR2_X1 U10052 ( .A(n8570), .B(n8569), .ZN(n8572) );
  AOI222_X1 U10053 ( .A1(n9928), .A2(n8572), .B1(n8571), .B2(n9930), .C1(n8590), .C2(n9933), .ZN(n8796) );
  MUX2_X1 U10054 ( .A(n8573), .B(n8796), .S(n8733), .Z(n8576) );
  AOI22_X1 U10055 ( .A1(n8798), .A2(n8705), .B1(n8729), .B2(n8574), .ZN(n8575)
         );
  OAI211_X1 U10056 ( .C1(n8801), .C2(n9943), .A(n8576), .B(n8575), .ZN(
        P2_U3207) );
  INV_X1 U10057 ( .A(n8803), .ZN(n8577) );
  NOR2_X1 U10058 ( .A1(n8577), .A2(n8709), .ZN(n8582) );
  XNOR2_X1 U10059 ( .A(n8578), .B(n8585), .ZN(n8580) );
  AOI222_X1 U10060 ( .A1(n9928), .A2(n8580), .B1(n8579), .B2(n9930), .C1(n8605), .C2(n9933), .ZN(n8802) );
  INV_X1 U10061 ( .A(n8802), .ZN(n8581) );
  AOI211_X1 U10062 ( .C1(n8729), .C2(n8583), .A(n8582), .B(n8581), .ZN(n8588)
         );
  XOR2_X1 U10063 ( .A(n8585), .B(n8584), .Z(n8806) );
  INV_X1 U10064 ( .A(n8806), .ZN(n8586) );
  AOI22_X1 U10065 ( .A1(n8586), .A2(n8681), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8713), .ZN(n8587) );
  OAI21_X1 U10066 ( .B1(n8588), .B2(n8713), .A(n8587), .ZN(P2_U3208) );
  XOR2_X1 U10067 ( .A(n8589), .B(n8597), .Z(n8592) );
  AOI222_X1 U10068 ( .A1(n9928), .A2(n8592), .B1(n8591), .B2(n9933), .C1(n8590), .C2(n9930), .ZN(n8807) );
  AOI22_X1 U10069 ( .A1(n8809), .A2(n8728), .B1(n8729), .B2(n8593), .ZN(n8594)
         );
  AOI21_X1 U10070 ( .B1(n8807), .B2(n8594), .A(n8713), .ZN(n8601) );
  NAND2_X1 U10071 ( .A1(n8595), .A2(n8596), .ZN(n8598) );
  XNOR2_X1 U10072 ( .A(n8598), .B(n8597), .ZN(n8812) );
  OAI22_X1 U10073 ( .A1(n8812), .A2(n9943), .B1(n8599), .B2(n8733), .ZN(n8600)
         );
  OR2_X1 U10074 ( .A1(n8601), .A2(n8600), .ZN(P2_U3209) );
  XNOR2_X1 U10075 ( .A(n8602), .B(n8603), .ZN(n8818) );
  INV_X1 U10076 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U10077 ( .A(n8604), .B(n8603), .ZN(n8606) );
  AOI222_X1 U10078 ( .A1(n9928), .A2(n8606), .B1(n8605), .B2(n9930), .C1(n8623), .C2(n9933), .ZN(n8813) );
  MUX2_X1 U10079 ( .A(n8607), .B(n8813), .S(n8733), .Z(n8610) );
  AOI22_X1 U10080 ( .A1(n8815), .A2(n8705), .B1(n8729), .B2(n8608), .ZN(n8609)
         );
  OAI211_X1 U10081 ( .C1(n8818), .C2(n9943), .A(n8610), .B(n8609), .ZN(
        P2_U3210) );
  XNOR2_X1 U10082 ( .A(n8611), .B(n8613), .ZN(n8612) );
  OAI222_X1 U10083 ( .A1(n8720), .A2(n8637), .B1(n8718), .B2(n6368), .C1(n6157), .C2(n8612), .ZN(n8755) );
  XNOR2_X1 U10084 ( .A(n8614), .B(n8613), .ZN(n8822) );
  AOI22_X1 U10085 ( .A1(n8713), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8729), .B2(
        n8615), .ZN(n8617) );
  NAND2_X1 U10086 ( .A1(n8756), .A2(n8705), .ZN(n8616) );
  OAI211_X1 U10087 ( .C1(n8822), .C2(n9943), .A(n8617), .B(n8616), .ZN(n8618)
         );
  AOI21_X1 U10088 ( .B1(n8755), .B2(n8733), .A(n8618), .ZN(n8619) );
  INV_X1 U10089 ( .A(n8619), .ZN(P2_U3211) );
  XNOR2_X1 U10090 ( .A(n8620), .B(n8621), .ZN(n8828) );
  INV_X1 U10091 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8626) );
  XNOR2_X1 U10092 ( .A(n8622), .B(n8621), .ZN(n8625) );
  AOI222_X1 U10093 ( .A1(n9928), .A2(n8625), .B1(n8624), .B2(n9933), .C1(n8623), .C2(n9930), .ZN(n8823) );
  MUX2_X1 U10094 ( .A(n8626), .B(n8823), .S(n8733), .Z(n8629) );
  AOI22_X1 U10095 ( .A1(n8825), .A2(n8705), .B1(n8729), .B2(n8627), .ZN(n8628)
         );
  OAI211_X1 U10096 ( .C1(n8828), .C2(n9943), .A(n8629), .B(n8628), .ZN(
        P2_U3212) );
  OR2_X1 U10097 ( .A1(n8630), .A2(n8631), .ZN(n8633) );
  AND2_X1 U10098 ( .A1(n8633), .A2(n8632), .ZN(n8634) );
  NAND2_X1 U10099 ( .A1(n8634), .A2(n8640), .ZN(n8635) );
  NAND2_X1 U10100 ( .A1(n4434), .A2(n8635), .ZN(n8639) );
  OAI22_X1 U10101 ( .A1(n8637), .A2(n8718), .B1(n8636), .B2(n8720), .ZN(n8638)
         );
  AOI21_X1 U10102 ( .B1(n8639), .B2(n9928), .A(n8638), .ZN(n8764) );
  INV_X1 U10103 ( .A(n8640), .ZN(n8641) );
  XNOR2_X1 U10104 ( .A(n8642), .B(n8641), .ZN(n8762) );
  AOI22_X1 U10105 ( .A1(n8713), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8729), .B2(
        n8643), .ZN(n8644) );
  OAI21_X1 U10106 ( .B1(n8645), .B2(n9939), .A(n8644), .ZN(n8646) );
  AOI21_X1 U10107 ( .B1(n8762), .B2(n8681), .A(n8646), .ZN(n8647) );
  OAI21_X1 U10108 ( .B1(n8764), .B2(n8713), .A(n8647), .ZN(P2_U3213) );
  OAI21_X1 U10109 ( .B1(n8649), .B2(n8654), .A(n8648), .ZN(n8836) );
  OR2_X1 U10110 ( .A1(n8630), .A2(n8650), .ZN(n8653) );
  NAND2_X1 U10111 ( .A1(n8653), .A2(n8651), .ZN(n8657) );
  NAND2_X1 U10112 ( .A1(n8653), .A2(n8652), .ZN(n8655) );
  NAND2_X1 U10113 ( .A1(n8655), .A2(n8654), .ZN(n8656) );
  NAND3_X1 U10114 ( .A1(n8657), .A2(n9928), .A3(n8656), .ZN(n8662) );
  OAI22_X1 U10115 ( .A1(n8659), .A2(n8718), .B1(n8658), .B2(n8720), .ZN(n8660)
         );
  INV_X1 U10116 ( .A(n8660), .ZN(n8661) );
  NAND2_X1 U10117 ( .A1(n8662), .A2(n8661), .ZN(n8833) );
  INV_X1 U10118 ( .A(n8833), .ZN(n8767) );
  MUX2_X1 U10119 ( .A(n8663), .B(n8767), .S(n8733), .Z(n8666) );
  AOI22_X1 U10120 ( .A1(n8769), .A2(n8705), .B1(n8729), .B2(n8664), .ZN(n8665)
         );
  OAI211_X1 U10121 ( .C1(n8836), .C2(n9943), .A(n8666), .B(n8665), .ZN(
        P2_U3214) );
  XOR2_X1 U10122 ( .A(n8630), .B(n8679), .Z(n8668) );
  AOI222_X1 U10123 ( .A1(n9928), .A2(n8668), .B1(n8667), .B2(n9930), .C1(n8700), .C2(n9933), .ZN(n8775) );
  INV_X1 U10124 ( .A(n8669), .ZN(n8670) );
  OAI22_X1 U10125 ( .A1(n8733), .A2(n8671), .B1(n8670), .B2(n9936), .ZN(n8672)
         );
  AOI21_X1 U10126 ( .B1(n8673), .B2(n8705), .A(n8672), .ZN(n8683) );
  OR2_X1 U10127 ( .A1(n8674), .A2(n8675), .ZN(n8678) );
  NAND2_X1 U10128 ( .A1(n8678), .A2(n8676), .ZN(n8773) );
  NAND2_X1 U10129 ( .A1(n8678), .A2(n8677), .ZN(n8680) );
  NAND2_X1 U10130 ( .A1(n8680), .A2(n8679), .ZN(n8772) );
  NAND3_X1 U10131 ( .A1(n8773), .A2(n8772), .A3(n8681), .ZN(n8682) );
  OAI211_X1 U10132 ( .C1(n8775), .C2(n8713), .A(n8683), .B(n8682), .ZN(
        P2_U3215) );
  XNOR2_X1 U10133 ( .A(n8674), .B(n8684), .ZN(n8845) );
  XNOR2_X1 U10134 ( .A(n8685), .B(n8684), .ZN(n8688) );
  AOI222_X1 U10135 ( .A1(n9928), .A2(n8688), .B1(n8687), .B2(n9930), .C1(n8686), .C2(n9933), .ZN(n8840) );
  MUX2_X1 U10136 ( .A(n8689), .B(n8840), .S(n8733), .Z(n8693) );
  INV_X1 U10137 ( .A(n8690), .ZN(n8691) );
  AOI22_X1 U10138 ( .A1(n8842), .A2(n8705), .B1(n8729), .B2(n8691), .ZN(n8692)
         );
  OAI211_X1 U10139 ( .C1(n8845), .C2(n9943), .A(n8693), .B(n8692), .ZN(
        P2_U3216) );
  NAND2_X1 U10140 ( .A1(n8695), .A2(n8694), .ZN(n8696) );
  XNOR2_X1 U10141 ( .A(n8696), .B(n8697), .ZN(n8851) );
  XOR2_X1 U10142 ( .A(n8698), .B(n8697), .Z(n8701) );
  AOI222_X1 U10143 ( .A1(n9928), .A2(n8701), .B1(n8700), .B2(n9930), .C1(n8699), .C2(n9933), .ZN(n8846) );
  MUX2_X1 U10144 ( .A(n8702), .B(n8846), .S(n8733), .Z(n8707) );
  INV_X1 U10145 ( .A(n8703), .ZN(n8704) );
  AOI22_X1 U10146 ( .A1(n8848), .A2(n8705), .B1(n8729), .B2(n8704), .ZN(n8706)
         );
  OAI211_X1 U10147 ( .C1(n8851), .C2(n9943), .A(n8707), .B(n8706), .ZN(
        P2_U3217) );
  INV_X1 U10148 ( .A(n8852), .ZN(n8712) );
  OAI22_X1 U10149 ( .A1(n8710), .A2(n8709), .B1(n8708), .B2(n9936), .ZN(n8711)
         );
  OAI21_X1 U10150 ( .B1(n8712), .B2(n8711), .A(n8733), .ZN(n8715) );
  NAND2_X1 U10151 ( .A1(n8713), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8714) );
  OAI211_X1 U10152 ( .C1(n8859), .C2(n9943), .A(n8715), .B(n8714), .ZN(
        P2_U3219) );
  OAI21_X1 U10153 ( .B1(n8716), .B2(n8722), .A(n6978), .ZN(n9950) );
  INV_X1 U10154 ( .A(n9950), .ZN(n8732) );
  INV_X1 U10155 ( .A(n8717), .ZN(n8727) );
  OAI22_X1 U10156 ( .A1(n6303), .A2(n8720), .B1(n8719), .B2(n8718), .ZN(n8726)
         );
  NAND3_X1 U10157 ( .A1(n6947), .A2(n8722), .A3(n8721), .ZN(n8723) );
  AOI21_X1 U10158 ( .B1(n8724), .B2(n8723), .A(n6157), .ZN(n8725) );
  AOI211_X1 U10159 ( .C1(n8727), .C2(n9950), .A(n8726), .B(n8725), .ZN(n9952)
         );
  AOI22_X1 U10160 ( .A1(n8729), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8728), .B2(
        n9948), .ZN(n8730) );
  OAI211_X1 U10161 ( .C1(n8732), .C2(n8731), .A(n9952), .B(n8730), .ZN(n8734)
         );
  MUX2_X1 U10162 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8734), .S(n8733), .Z(
        P2_U3231) );
  AOI21_X1 U10163 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n6287), .A(n8735), .ZN(
        n8736) );
  OAI21_X1 U10164 ( .B1(n8786), .B2(n8737), .A(n8736), .ZN(P2_U3490) );
  INV_X1 U10165 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U10166 ( .A1(n8738), .A2(n9987), .ZN(n8739) );
  AND2_X1 U10167 ( .A1(n8740), .A2(n8739), .ZN(n8792) );
  MUX2_X1 U10168 ( .A(n8741), .B(n8792), .S(n10008), .Z(n8742) );
  OAI21_X1 U10169 ( .B1(n8783), .B2(n8795), .A(n8742), .ZN(P2_U3486) );
  INV_X1 U10170 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8743) );
  MUX2_X1 U10171 ( .A(n8743), .B(n8796), .S(n10008), .Z(n8745) );
  NAND2_X1 U10172 ( .A1(n8798), .A2(n8780), .ZN(n8744) );
  OAI211_X1 U10173 ( .C1(n8783), .C2(n8801), .A(n8745), .B(n8744), .ZN(
        P2_U3485) );
  INV_X1 U10174 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8746) );
  MUX2_X1 U10175 ( .A(n8746), .B(n8802), .S(n10008), .Z(n8748) );
  NAND2_X1 U10176 ( .A1(n8803), .A2(n8780), .ZN(n8747) );
  OAI211_X1 U10177 ( .C1(n8806), .C2(n8783), .A(n8748), .B(n8747), .ZN(
        P2_U3484) );
  INV_X1 U10178 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8749) );
  MUX2_X1 U10179 ( .A(n8749), .B(n8807), .S(n10008), .Z(n8751) );
  NAND2_X1 U10180 ( .A1(n8809), .A2(n8780), .ZN(n8750) );
  OAI211_X1 U10181 ( .C1(n8783), .C2(n8812), .A(n8751), .B(n8750), .ZN(
        P2_U3483) );
  INV_X1 U10182 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8752) );
  MUX2_X1 U10183 ( .A(n8752), .B(n8813), .S(n10008), .Z(n8754) );
  NAND2_X1 U10184 ( .A1(n8815), .A2(n8780), .ZN(n8753) );
  OAI211_X1 U10185 ( .C1(n8818), .C2(n8783), .A(n8754), .B(n8753), .ZN(
        P2_U3482) );
  INV_X1 U10186 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8757) );
  AOI21_X1 U10187 ( .B1(n9987), .B2(n8756), .A(n8755), .ZN(n8819) );
  MUX2_X1 U10188 ( .A(n8757), .B(n8819), .S(n10008), .Z(n8758) );
  OAI21_X1 U10189 ( .B1(n8822), .B2(n8783), .A(n8758), .ZN(P2_U3481) );
  INV_X1 U10190 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8759) );
  MUX2_X1 U10191 ( .A(n8759), .B(n8823), .S(n10008), .Z(n8761) );
  NAND2_X1 U10192 ( .A1(n8825), .A2(n8780), .ZN(n8760) );
  OAI211_X1 U10193 ( .C1(n8783), .C2(n8828), .A(n8761), .B(n8760), .ZN(
        P2_U3480) );
  NAND2_X1 U10194 ( .A1(n8762), .A2(n9994), .ZN(n8763) );
  NAND2_X1 U10195 ( .A1(n8764), .A2(n8763), .ZN(n8829) );
  MUX2_X1 U10196 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8829), .S(n10008), .Z(
        n8765) );
  AOI21_X1 U10197 ( .B1(n8780), .B2(n8831), .A(n8765), .ZN(n8766) );
  INV_X1 U10198 ( .A(n8766), .ZN(P2_U3479) );
  MUX2_X1 U10199 ( .A(n8768), .B(n8767), .S(n10008), .Z(n8771) );
  NAND2_X1 U10200 ( .A1(n8769), .A2(n8780), .ZN(n8770) );
  OAI211_X1 U10201 ( .C1(n8783), .C2(n8836), .A(n8771), .B(n8770), .ZN(
        P2_U3478) );
  NAND3_X1 U10202 ( .A1(n8773), .A2(n8772), .A3(n9994), .ZN(n8774) );
  OAI211_X1 U10203 ( .C1(n8776), .C2(n9989), .A(n8775), .B(n8774), .ZN(n8839)
         );
  MUX2_X1 U10204 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8839), .S(n10008), .Z(
        P2_U3477) );
  MUX2_X1 U10205 ( .A(n10071), .B(n8840), .S(n10008), .Z(n8778) );
  NAND2_X1 U10206 ( .A1(n8842), .A2(n8780), .ZN(n8777) );
  OAI211_X1 U10207 ( .C1(n8845), .C2(n8783), .A(n8778), .B(n8777), .ZN(
        P2_U3476) );
  MUX2_X1 U10208 ( .A(n8779), .B(n8846), .S(n10008), .Z(n8782) );
  NAND2_X1 U10209 ( .A1(n8848), .A2(n8780), .ZN(n8781) );
  OAI211_X1 U10210 ( .C1(n8783), .C2(n8851), .A(n8782), .B(n8781), .ZN(
        P2_U3475) );
  NOR2_X1 U10211 ( .A1(n8784), .A2(n9997), .ZN(n8788) );
  AOI21_X1 U10212 ( .B1(n9997), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8788), .ZN(
        n8785) );
  OAI21_X1 U10213 ( .B1(n8786), .B2(n8834), .A(n8785), .ZN(P2_U3458) );
  INV_X1 U10214 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U10215 ( .A1(n8787), .A2(n8854), .ZN(n8790) );
  INV_X1 U10216 ( .A(n8788), .ZN(n8789) );
  OAI211_X1 U10217 ( .C1(n8791), .C2(n9995), .A(n8790), .B(n8789), .ZN(
        P2_U3457) );
  MUX2_X1 U10218 ( .A(n8793), .B(n8792), .S(n9995), .Z(n8794) );
  OAI21_X1 U10219 ( .B1(n8795), .B2(n8858), .A(n8794), .ZN(P2_U3454) );
  MUX2_X1 U10220 ( .A(n8797), .B(n8796), .S(n9995), .Z(n8800) );
  NAND2_X1 U10221 ( .A1(n8798), .A2(n8854), .ZN(n8799) );
  OAI211_X1 U10222 ( .C1(n8801), .C2(n8858), .A(n8800), .B(n8799), .ZN(
        P2_U3453) );
  MUX2_X1 U10223 ( .A(n10193), .B(n8802), .S(n9995), .Z(n8805) );
  NAND2_X1 U10224 ( .A1(n8803), .A2(n8854), .ZN(n8804) );
  OAI211_X1 U10225 ( .C1(n8806), .C2(n8858), .A(n8805), .B(n8804), .ZN(
        P2_U3452) );
  INV_X1 U10226 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8808) );
  MUX2_X1 U10227 ( .A(n8808), .B(n8807), .S(n9995), .Z(n8811) );
  NAND2_X1 U10228 ( .A1(n8809), .A2(n8854), .ZN(n8810) );
  OAI211_X1 U10229 ( .C1(n8812), .C2(n8858), .A(n8811), .B(n8810), .ZN(
        P2_U3451) );
  MUX2_X1 U10230 ( .A(n8814), .B(n8813), .S(n9995), .Z(n8817) );
  NAND2_X1 U10231 ( .A1(n8815), .A2(n8854), .ZN(n8816) );
  OAI211_X1 U10232 ( .C1(n8818), .C2(n8858), .A(n8817), .B(n8816), .ZN(
        P2_U3450) );
  MUX2_X1 U10233 ( .A(n8820), .B(n8819), .S(n9995), .Z(n8821) );
  OAI21_X1 U10234 ( .B1(n8822), .B2(n8858), .A(n8821), .ZN(P2_U3449) );
  INV_X1 U10235 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8824) );
  MUX2_X1 U10236 ( .A(n8824), .B(n8823), .S(n9995), .Z(n8827) );
  NAND2_X1 U10237 ( .A1(n8825), .A2(n8854), .ZN(n8826) );
  OAI211_X1 U10238 ( .C1(n8828), .C2(n8858), .A(n8827), .B(n8826), .ZN(
        P2_U3448) );
  MUX2_X1 U10239 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8829), .S(n9995), .Z(n8830) );
  AOI21_X1 U10240 ( .B1(n8854), .B2(n8831), .A(n8830), .ZN(n8832) );
  INV_X1 U10241 ( .A(n8832), .ZN(P2_U3447) );
  MUX2_X1 U10242 ( .A(n8833), .B(P2_REG0_REG_19__SCAN_IN), .S(n9997), .Z(n8838) );
  OAI22_X1 U10243 ( .A1(n8836), .A2(n8858), .B1(n8835), .B2(n8834), .ZN(n8837)
         );
  OR2_X1 U10244 ( .A1(n8838), .A2(n8837), .ZN(P2_U3446) );
  MUX2_X1 U10245 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8839), .S(n9995), .Z(
        P2_U3444) );
  MUX2_X1 U10246 ( .A(n8841), .B(n8840), .S(n9995), .Z(n8844) );
  NAND2_X1 U10247 ( .A1(n8842), .A2(n8854), .ZN(n8843) );
  OAI211_X1 U10248 ( .C1(n8845), .C2(n8858), .A(n8844), .B(n8843), .ZN(
        P2_U3441) );
  INV_X1 U10249 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8847) );
  MUX2_X1 U10250 ( .A(n8847), .B(n8846), .S(n9995), .Z(n8850) );
  NAND2_X1 U10251 ( .A1(n8848), .A2(n8854), .ZN(n8849) );
  OAI211_X1 U10252 ( .C1(n8851), .C2(n8858), .A(n8850), .B(n8849), .ZN(
        P2_U3438) );
  MUX2_X1 U10253 ( .A(n8853), .B(n8852), .S(n9995), .Z(n8857) );
  NAND2_X1 U10254 ( .A1(n8855), .A2(n8854), .ZN(n8856) );
  OAI211_X1 U10255 ( .C1(n8859), .C2(n8858), .A(n8857), .B(n8856), .ZN(
        P2_U3432) );
  NAND3_X1 U10256 ( .A1(n8861), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8863) );
  OAI22_X1 U10257 ( .A1(n8860), .A2(n8863), .B1(n8862), .B2(n8019), .ZN(n8864)
         );
  AOI21_X1 U10258 ( .B1(n9426), .B2(n8865), .A(n8864), .ZN(n8866) );
  INV_X1 U10259 ( .A(n8866), .ZN(P2_U3264) );
  INV_X1 U10260 ( .A(n8867), .ZN(n8868) );
  MUX2_X1 U10261 ( .A(n8868), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10262 ( .A(n8869), .ZN(n8871) );
  INV_X1 U10263 ( .A(n8872), .ZN(n8873) );
  OAI21_X1 U10264 ( .B1(n8874), .B2(n8873), .A(n9021), .ZN(n8879) );
  OAI22_X1 U10265 ( .A1(n8928), .A2(n9006), .B1(n8918), .B2(n9008), .ZN(n9219)
         );
  INV_X1 U10266 ( .A(n9213), .ZN(n8876) );
  OAI22_X1 U10267 ( .A1(n8876), .A2(n9012), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8875), .ZN(n8877) );
  AOI21_X1 U10268 ( .B1(n9219), .B2(n9014), .A(n8877), .ZN(n8878) );
  OAI211_X1 U10269 ( .C1(n9215), .C2(n9034), .A(n8879), .B(n8878), .ZN(
        P1_U3216) );
  INV_X1 U10270 ( .A(n8880), .ZN(n8881) );
  NOR2_X1 U10271 ( .A1(n8882), .A2(n8881), .ZN(n8883) );
  XNOR2_X1 U10272 ( .A(n8884), .B(n8883), .ZN(n8891) );
  OAI22_X1 U10273 ( .A1(n9025), .A2(n8886), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8885), .ZN(n8887) );
  AOI21_X1 U10274 ( .B1(n8993), .B2(n9278), .A(n8887), .ZN(n8888) );
  OAI21_X1 U10275 ( .B1(n9012), .B2(n9283), .A(n8888), .ZN(n8889) );
  AOI21_X1 U10276 ( .B1(n9286), .B2(n5752), .A(n8889), .ZN(n8890) );
  OAI21_X1 U10277 ( .B1(n8891), .B2(n8999), .A(n8890), .ZN(P1_U3219) );
  NAND2_X1 U10278 ( .A1(n9346), .A2(n5150), .ZN(n8893) );
  NAND2_X1 U10279 ( .A1(n9038), .A2(n5159), .ZN(n8892) );
  NAND2_X1 U10280 ( .A1(n8893), .A2(n8892), .ZN(n8895) );
  XNOR2_X1 U10281 ( .A(n8895), .B(n8894), .ZN(n8898) );
  AOI22_X1 U10282 ( .A1(n9346), .A2(n5159), .B1(n8896), .B2(n9038), .ZN(n8897)
         );
  XNOR2_X1 U10283 ( .A(n8898), .B(n8897), .ZN(n8908) );
  NAND3_X1 U10284 ( .A1(n4757), .A2(n9021), .A3(n8908), .ZN(n8912) );
  INV_X1 U10285 ( .A(n8907), .ZN(n8900) );
  INV_X1 U10286 ( .A(n8908), .ZN(n8899) );
  NAND4_X1 U10287 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n9021), .ZN(n8911)
         );
  INV_X1 U10288 ( .A(n8902), .ZN(n9144) );
  NAND2_X1 U10289 ( .A1(n9037), .A2(n9311), .ZN(n8904) );
  NAND2_X1 U10290 ( .A1(n9039), .A2(n9309), .ZN(n8903) );
  NAND2_X1 U10291 ( .A1(n8904), .A2(n8903), .ZN(n9151) );
  AOI22_X1 U10292 ( .A1(n9151), .A2(n9014), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8905) );
  OAI21_X1 U10293 ( .B1(n9012), .B2(n9144), .A(n8905), .ZN(n8906) );
  AOI21_X1 U10294 ( .B1(n9346), .B2(n5752), .A(n8906), .ZN(n8910) );
  NAND3_X1 U10295 ( .A1(n8908), .A2(n9021), .A3(n8907), .ZN(n8909) );
  NAND4_X1 U10296 ( .A1(n8912), .A2(n8911), .A3(n8910), .A4(n8909), .ZN(
        P1_U3220) );
  INV_X1 U10297 ( .A(n9381), .ZN(n9252) );
  OAI21_X1 U10298 ( .B1(n8915), .B2(n8914), .A(n8913), .ZN(n8916) );
  NAND2_X1 U10299 ( .A1(n8916), .A2(n9021), .ZN(n8923) );
  OAI22_X1 U10300 ( .A1(n8918), .A2(n9006), .B1(n8917), .B2(n9008), .ZN(n9244)
         );
  INV_X1 U10301 ( .A(n9249), .ZN(n8920) );
  INV_X1 U10302 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8919) );
  OAI22_X1 U10303 ( .A1(n9012), .A2(n8920), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8919), .ZN(n8921) );
  AOI21_X1 U10304 ( .B1(n9244), .B2(n9014), .A(n8921), .ZN(n8922) );
  OAI211_X1 U10305 ( .C1(n9252), .C2(n9034), .A(n8923), .B(n8922), .ZN(
        P1_U3223) );
  NAND2_X1 U10306 ( .A1(n8924), .A2(n8960), .ZN(n8964) );
  NAND2_X1 U10307 ( .A1(n8964), .A2(n8925), .ZN(n8926) );
  OAI21_X1 U10308 ( .B1(n8927), .B2(n8926), .A(n9002), .ZN(n8934) );
  AOI22_X1 U10309 ( .A1(n9186), .A2(n9030), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8932) );
  OR2_X1 U10310 ( .A1(n8928), .A2(n9008), .ZN(n8930) );
  NAND2_X1 U10311 ( .A1(n9040), .A2(n9311), .ZN(n8929) );
  NAND2_X1 U10312 ( .A1(n8930), .A2(n8929), .ZN(n9192) );
  NAND2_X1 U10313 ( .A1(n9192), .A2(n9014), .ZN(n8931) );
  OAI211_X1 U10314 ( .C1(n9188), .C2(n9034), .A(n8932), .B(n8931), .ZN(n8933)
         );
  AOI21_X1 U10315 ( .B1(n8934), .B2(n9021), .A(n8933), .ZN(n8935) );
  INV_X1 U10316 ( .A(n8935), .ZN(P1_U3225) );
  XNOR2_X1 U10317 ( .A(n8936), .B(n8937), .ZN(n9019) );
  NAND2_X1 U10318 ( .A1(n9019), .A2(n9020), .ZN(n9018) );
  OAI21_X1 U10319 ( .B1(n8936), .B2(n8938), .A(n9018), .ZN(n8942) );
  XNOR2_X1 U10320 ( .A(n8940), .B(n8939), .ZN(n8941) );
  XNOR2_X1 U10321 ( .A(n8942), .B(n8941), .ZN(n8949) );
  NAND2_X1 U10322 ( .A1(n8993), .A2(n9301), .ZN(n8943) );
  NAND2_X1 U10323 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9072) );
  OAI211_X1 U10324 ( .C1(n9025), .C2(n8944), .A(n8943), .B(n9072), .ZN(n8945)
         );
  AOI21_X1 U10325 ( .B1(n8946), .B2(n9030), .A(n8945), .ZN(n8948) );
  NAND2_X1 U10326 ( .A1(n9512), .A2(n5752), .ZN(n8947) );
  OAI211_X1 U10327 ( .C1(n8949), .C2(n8999), .A(n8948), .B(n8947), .ZN(
        P1_U3226) );
  INV_X1 U10328 ( .A(n9323), .ZN(n9509) );
  OAI211_X1 U10329 ( .C1(n8952), .C2(n8951), .A(n8950), .B(n9021), .ZN(n8956)
         );
  NAND2_X1 U10330 ( .A1(n8993), .A2(n9312), .ZN(n8953) );
  NAND2_X1 U10331 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9098) );
  OAI211_X1 U10332 ( .C1(n9025), .C2(n9026), .A(n8953), .B(n9098), .ZN(n8954)
         );
  AOI21_X1 U10333 ( .B1(n9314), .B2(n9030), .A(n8954), .ZN(n8955) );
  OAI211_X1 U10334 ( .C1(n9509), .C2(n9034), .A(n8956), .B(n8955), .ZN(
        P1_U3228) );
  NOR2_X1 U10335 ( .A1(n8980), .A2(n9008), .ZN(n8957) );
  AOI21_X1 U10336 ( .B1(n9041), .B2(n9311), .A(n8957), .ZN(n9201) );
  AOI22_X1 U10337 ( .A1(n4968), .A2(n9030), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8958) );
  OAI21_X1 U10338 ( .B1(n9201), .B2(n8959), .A(n8958), .ZN(n8966) );
  INV_X1 U10339 ( .A(n8960), .ZN(n8961) );
  NAND3_X1 U10340 ( .A1(n8872), .A2(n8962), .A3(n8961), .ZN(n8963) );
  AOI21_X1 U10341 ( .B1(n8964), .B2(n8963), .A(n8999), .ZN(n8965) );
  AOI211_X1 U10342 ( .C1(n9367), .C2(n5752), .A(n8966), .B(n8965), .ZN(n8967)
         );
  INV_X1 U10343 ( .A(n8967), .ZN(P1_U3229) );
  OAI21_X1 U10344 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n8971) );
  NAND2_X1 U10345 ( .A1(n8971), .A2(n9021), .ZN(n8976) );
  OAI22_X1 U10346 ( .A1(n8982), .A2(n9006), .B1(n8972), .B2(n9008), .ZN(n9260)
         );
  INV_X1 U10347 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8973) );
  OAI22_X1 U10348 ( .A1(n9012), .A2(n9262), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8973), .ZN(n8974) );
  AOI21_X1 U10349 ( .B1(n9260), .B2(n9014), .A(n8974), .ZN(n8975) );
  OAI211_X1 U10350 ( .C1(n9265), .C2(n9034), .A(n8976), .B(n8975), .ZN(
        P1_U3233) );
  AOI21_X1 U10351 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(n8987) );
  OR2_X1 U10352 ( .A1(n8980), .A2(n9006), .ZN(n8981) );
  OAI21_X1 U10353 ( .B1(n8982), .B2(n9008), .A(n8981), .ZN(n9235) );
  OAI22_X1 U10354 ( .A1(n9012), .A2(n9229), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8983), .ZN(n8985) );
  NOR2_X1 U10355 ( .A1(n6520), .A2(n9034), .ZN(n8984) );
  AOI211_X1 U10356 ( .C1(n9014), .C2(n9235), .A(n8985), .B(n8984), .ZN(n8986)
         );
  OAI21_X1 U10357 ( .B1(n8987), .B2(n8999), .A(n8986), .ZN(P1_U3235) );
  INV_X1 U10358 ( .A(n8988), .ZN(n8990) );
  NAND2_X1 U10359 ( .A1(n8990), .A2(n8989), .ZN(n8992) );
  XNOR2_X1 U10360 ( .A(n8992), .B(n8991), .ZN(n9000) );
  AOI22_X1 U10361 ( .A1(n8993), .A2(n9302), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8995) );
  NAND2_X1 U10362 ( .A1(n9030), .A2(n9294), .ZN(n8994) );
  OAI211_X1 U10363 ( .C1(n8996), .C2(n9025), .A(n8995), .B(n8994), .ZN(n8997)
         );
  AOI21_X1 U10364 ( .B1(n9397), .B2(n5752), .A(n8997), .ZN(n8998) );
  OAI21_X1 U10365 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(P1_U3238) );
  AND2_X1 U10366 ( .A1(n9002), .A2(n9001), .ZN(n9005) );
  OAI211_X1 U10367 ( .C1(n9005), .C2(n9004), .A(n9021), .B(n9003), .ZN(n9016)
         );
  OAI22_X1 U10368 ( .A1(n9009), .A2(n9008), .B1(n9007), .B2(n9006), .ZN(n9178)
         );
  INV_X1 U10369 ( .A(n9010), .ZN(n9175) );
  OAI22_X1 U10370 ( .A1(n9012), .A2(n9175), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9011), .ZN(n9013) );
  AOI21_X1 U10371 ( .B1(n9178), .B2(n9014), .A(n9013), .ZN(n9015) );
  OAI211_X1 U10372 ( .C1(n9017), .C2(n9034), .A(n9016), .B(n9015), .ZN(
        P1_U3240) );
  OAI21_X1 U10373 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(n9022) );
  NAND2_X1 U10374 ( .A1(n9022), .A2(n9021), .ZN(n9033) );
  OAI22_X1 U10375 ( .A1(n9025), .A2(n9024), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9023), .ZN(n9029) );
  NOR2_X1 U10376 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  AOI211_X1 U10377 ( .C1(n9031), .C2(n9030), .A(n9029), .B(n9028), .ZN(n9032)
         );
  OAI211_X1 U10378 ( .C1(n9035), .C2(n9034), .A(n9033), .B(n9032), .ZN(
        P1_U3241) );
  MUX2_X1 U10379 ( .A(n9125), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9060), .Z(
        P1_U3585) );
  MUX2_X1 U10380 ( .A(n9036), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9060), .Z(
        P1_U3584) );
  MUX2_X1 U10381 ( .A(n9037), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9060), .Z(
        P1_U3583) );
  MUX2_X1 U10382 ( .A(n9038), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9060), .Z(
        P1_U3582) );
  MUX2_X1 U10383 ( .A(n9039), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9060), .Z(
        P1_U3581) );
  MUX2_X1 U10384 ( .A(n9040), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9060), .Z(
        P1_U3580) );
  MUX2_X1 U10385 ( .A(n9041), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9060), .Z(
        P1_U3579) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9042), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9043), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10388 ( .A(n9044), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9060), .Z(
        P1_U3576) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9045), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10390 ( .A(n9278), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9060), .Z(
        P1_U3574) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9302), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9312), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10393 ( .A(n9301), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9060), .Z(
        P1_U3571) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9310), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10395 ( .A(n9046), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9060), .Z(
        P1_U3569) );
  MUX2_X1 U10396 ( .A(n9047), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9060), .Z(
        P1_U3568) );
  MUX2_X1 U10397 ( .A(n9048), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9060), .Z(
        P1_U3567) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9049), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10399 ( .A(n9050), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9060), .Z(
        P1_U3565) );
  MUX2_X1 U10400 ( .A(n9051), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9060), .Z(
        P1_U3564) );
  MUX2_X1 U10401 ( .A(n9052), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9060), .Z(
        P1_U3563) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9053), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9054), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10404 ( .A(n9055), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9060), .Z(
        P1_U3560) );
  MUX2_X1 U10405 ( .A(n9056), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9060), .Z(
        P1_U3559) );
  MUX2_X1 U10406 ( .A(n9057), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9060), .Z(
        P1_U3558) );
  MUX2_X1 U10407 ( .A(n9058), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9060), .Z(
        P1_U3557) );
  MUX2_X1 U10408 ( .A(n9059), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9060), .Z(
        P1_U3556) );
  MUX2_X1 U10409 ( .A(n6493), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9060), .Z(
        P1_U3555) );
  INV_X1 U10410 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9061) );
  MUX2_X1 U10411 ( .A(n9061), .B(P1_REG1_REG_13__SCAN_IN), .S(n9589), .Z(n9597) );
  OR2_X1 U10412 ( .A1(n9077), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9063) );
  INV_X1 U10413 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9064) );
  OR2_X1 U10414 ( .A1(n9609), .A2(n9064), .ZN(n9066) );
  NAND2_X1 U10415 ( .A1(n9609), .A2(n9064), .ZN(n9065) );
  AND2_X1 U10416 ( .A1(n9066), .A2(n9065), .ZN(n9616) );
  NOR2_X1 U10417 ( .A1(n9617), .A2(n9616), .ZN(n9618) );
  AOI21_X1 U10418 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9609), .A(n9618), .ZN(
        n9067) );
  NOR2_X1 U10419 ( .A1(n9067), .A2(n9079), .ZN(n9068) );
  INV_X1 U10420 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9632) );
  INV_X1 U10421 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9069) );
  MUX2_X1 U10422 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9069), .S(n9095), .Z(n9070) );
  OAI21_X1 U10423 ( .B1(n9071), .B2(n9070), .A(n9094), .ZN(n9086) );
  NAND2_X1 U10424 ( .A1(n9522), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9073) );
  OAI211_X1 U10425 ( .C1(n9625), .C2(n9074), .A(n9073), .B(n9072), .ZN(n9085)
         );
  NAND2_X1 U10426 ( .A1(n9589), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9075) );
  OAI21_X1 U10427 ( .B1(n9589), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9075), .ZN(
        n9591) );
  NAND2_X1 U10428 ( .A1(n9609), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9078) );
  OAI21_X1 U10429 ( .B1(n9609), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9078), .ZN(
        n9611) );
  AOI21_X1 U10430 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9609), .A(n9612), .ZN(
        n9080) );
  INV_X1 U10431 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9634) );
  XNOR2_X1 U10432 ( .A(n9095), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9082) );
  INV_X1 U10433 ( .A(n9089), .ZN(n9081) );
  AOI211_X1 U10434 ( .C1(n9083), .C2(n9082), .A(n9649), .B(n9081), .ZN(n9084)
         );
  AOI211_X1 U10435 ( .C1(n9112), .C2(n9086), .A(n9085), .B(n9084), .ZN(n9087)
         );
  INV_X1 U10436 ( .A(n9087), .ZN(P1_U3259) );
  NAND2_X1 U10437 ( .A1(n9095), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9088) );
  INV_X1 U10438 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9317) );
  MUX2_X1 U10439 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n9317), .S(n9110), .Z(n9090) );
  NAND2_X1 U10440 ( .A1(n9091), .A2(n9090), .ZN(n9106) );
  OAI21_X1 U10441 ( .B1(n9091), .B2(n9090), .A(n9106), .ZN(n9092) );
  NAND2_X1 U10442 ( .A1(n9092), .A2(n9116), .ZN(n9103) );
  INV_X1 U10443 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9093) );
  MUX2_X1 U10444 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9093), .S(n9110), .Z(n9097) );
  OAI21_X1 U10445 ( .B1(n9095), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9094), .ZN(
        n9096) );
  NAND2_X1 U10446 ( .A1(n9096), .A2(n9097), .ZN(n9109) );
  OAI21_X1 U10447 ( .B1(n9097), .B2(n9096), .A(n9109), .ZN(n9101) );
  NAND2_X1 U10448 ( .A1(n9522), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9099) );
  OAI211_X1 U10449 ( .C1(n9625), .C2(n9104), .A(n9099), .B(n9098), .ZN(n9100)
         );
  AOI21_X1 U10450 ( .B1(n9101), .B2(n9112), .A(n9100), .ZN(n9102) );
  NAND2_X1 U10451 ( .A1(n9103), .A2(n9102), .ZN(P1_U3260) );
  NAND2_X1 U10452 ( .A1(n9104), .A2(n9317), .ZN(n9105) );
  NAND2_X1 U10453 ( .A1(n9106), .A2(n9105), .ZN(n9650) );
  NAND2_X1 U10454 ( .A1(n9654), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9107) );
  OAI21_X1 U10455 ( .B1(n9654), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9107), .ZN(
        n9651) );
  NAND2_X1 U10456 ( .A1(n9647), .A2(n9107), .ZN(n9108) );
  INV_X1 U10457 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9284) );
  XNOR2_X1 U10458 ( .A(n9108), .B(n9284), .ZN(n9113) );
  OAI21_X1 U10459 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9110), .A(n9109), .ZN(
        n9645) );
  NAND2_X1 U10460 ( .A1(n9654), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9111) );
  OAI21_X1 U10461 ( .B1(n9654), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9111), .ZN(
        n9646) );
  AOI22_X1 U10462 ( .A1(n9113), .A2(n9116), .B1(n9112), .B2(n9114), .ZN(n9119)
         );
  INV_X1 U10463 ( .A(n9113), .ZN(n9117) );
  AOI21_X1 U10464 ( .B1(n9117), .B2(n9116), .A(n9115), .ZN(n9118) );
  MUX2_X1 U10465 ( .A(n9119), .B(n9118), .S(n9747), .Z(n9121) );
  NAND2_X1 U10466 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9120) );
  OAI211_X1 U10467 ( .C1(n9122), .C2(n9659), .A(n9121), .B(n9120), .ZN(
        P1_U3262) );
  NAND2_X1 U10468 ( .A1(n9123), .A2(n9734), .ZN(n9331) );
  INV_X1 U10469 ( .A(n9124), .ZN(n9126) );
  NAND2_X1 U10470 ( .A1(n9126), .A2(n9125), .ZN(n9337) );
  NOR2_X1 U10471 ( .A1(n9754), .A2(n9337), .ZN(n9133) );
  NOR2_X1 U10472 ( .A1(n9752), .A2(n9127), .ZN(n9128) );
  AOI211_X1 U10473 ( .C1(n4790), .C2(n9739), .A(n9133), .B(n9128), .ZN(n9129)
         );
  OAI21_X1 U10474 ( .B1(n9331), .B2(n9694), .A(n9129), .ZN(P1_U3263) );
  OAI211_X1 U10475 ( .C1(n9339), .C2(n9131), .A(n9734), .B(n9130), .ZN(n9338)
         );
  NOR2_X1 U10476 ( .A1(n9752), .A2(n9132), .ZN(n9134) );
  AOI211_X1 U10477 ( .C1(n9135), .C2(n9739), .A(n9134), .B(n9133), .ZN(n9136)
         );
  OAI21_X1 U10478 ( .B1(n9338), .B2(n9694), .A(n9136), .ZN(P1_U3264) );
  OAI21_X1 U10479 ( .B1(n9138), .B2(n9145), .A(n9137), .ZN(n9349) );
  OR2_X1 U10480 ( .A1(n9139), .A2(n9159), .ZN(n9140) );
  AND3_X1 U10481 ( .A1(n9141), .A2(n9140), .A3(n9734), .ZN(n9345) );
  NAND2_X1 U10482 ( .A1(n9346), .A2(n9739), .ZN(n9143) );
  NAND2_X1 U10483 ( .A1(n9754), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9142) );
  OAI211_X1 U10484 ( .C1(n9315), .C2(n9144), .A(n9143), .B(n9142), .ZN(n9154)
         );
  INV_X1 U10485 ( .A(n9145), .ZN(n9147) );
  NOR2_X1 U10486 ( .A1(n9147), .A2(n9146), .ZN(n9150) );
  AOI211_X1 U10487 ( .C1(n9150), .C2(n9149), .A(n9759), .B(n9148), .ZN(n9152)
         );
  NOR2_X1 U10488 ( .A1(n9152), .A2(n9151), .ZN(n9348) );
  NOR2_X1 U10489 ( .A1(n9348), .A2(n9754), .ZN(n9153) );
  AOI211_X1 U10490 ( .C1(n9345), .C2(n9738), .A(n9154), .B(n9153), .ZN(n9155)
         );
  OAI21_X1 U10491 ( .B1(n9307), .B2(n9349), .A(n9155), .ZN(P1_U3265) );
  XNOR2_X1 U10492 ( .A(n9156), .B(n9165), .ZN(n9354) );
  NAND2_X1 U10493 ( .A1(n9352), .A2(n4973), .ZN(n9157) );
  NAND2_X1 U10494 ( .A1(n9157), .A2(n9734), .ZN(n9158) );
  NOR2_X1 U10495 ( .A1(n9159), .A2(n9158), .ZN(n9351) );
  INV_X1 U10496 ( .A(n9160), .ZN(n9163) );
  NAND2_X1 U10497 ( .A1(n9352), .A2(n9739), .ZN(n9162) );
  NAND2_X1 U10498 ( .A1(n9754), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9161) );
  OAI211_X1 U10499 ( .C1(n9163), .C2(n9315), .A(n9162), .B(n9161), .ZN(n9164)
         );
  AOI21_X1 U10500 ( .B1(n9351), .B2(n9738), .A(n9164), .ZN(n9170) );
  XNOR2_X1 U10501 ( .A(n9166), .B(n9165), .ZN(n9168) );
  OAI21_X1 U10502 ( .B1(n9168), .B2(n9759), .A(n9167), .ZN(n9350) );
  NAND2_X1 U10503 ( .A1(n9350), .A2(n9752), .ZN(n9169) );
  OAI211_X1 U10504 ( .C1(n9354), .C2(n9307), .A(n9170), .B(n9169), .ZN(
        P1_U3266) );
  XNOR2_X1 U10505 ( .A(n9171), .B(n9176), .ZN(n9359) );
  AOI21_X1 U10506 ( .B1(n9356), .B2(n9184), .A(n9246), .ZN(n9172) );
  AND2_X1 U10507 ( .A1(n9172), .A2(n4973), .ZN(n9355) );
  NAND2_X1 U10508 ( .A1(n9356), .A2(n9739), .ZN(n9174) );
  NAND2_X1 U10509 ( .A1(n9754), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9173) );
  OAI211_X1 U10510 ( .C1(n9315), .C2(n9175), .A(n9174), .B(n9173), .ZN(n9181)
         );
  XNOR2_X1 U10511 ( .A(n9177), .B(n9176), .ZN(n9179) );
  AOI21_X1 U10512 ( .B1(n9179), .B2(n9702), .A(n9178), .ZN(n9358) );
  NOR2_X1 U10513 ( .A1(n9358), .A2(n9754), .ZN(n9180) );
  AOI211_X1 U10514 ( .C1(n9355), .C2(n9738), .A(n9181), .B(n9180), .ZN(n9182)
         );
  OAI21_X1 U10515 ( .B1(n9307), .B2(n9359), .A(n9182), .ZN(P1_U3267) );
  XOR2_X1 U10516 ( .A(n9183), .B(n9190), .Z(n9364) );
  INV_X1 U10517 ( .A(n9184), .ZN(n9185) );
  AOI211_X1 U10518 ( .C1(n9361), .C2(n4812), .A(n9246), .B(n9185), .ZN(n9360)
         );
  AOI22_X1 U10519 ( .A1(n9186), .A2(n9749), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9754), .ZN(n9187) );
  OAI21_X1 U10520 ( .B1(n9188), .B2(n9720), .A(n9187), .ZN(n9195) );
  AOI211_X1 U10521 ( .C1(n9191), .C2(n9190), .A(n9759), .B(n9189), .ZN(n9193)
         );
  NOR2_X1 U10522 ( .A1(n9193), .A2(n9192), .ZN(n9363) );
  NOR2_X1 U10523 ( .A1(n9363), .A2(n9754), .ZN(n9194) );
  AOI211_X1 U10524 ( .C1(n9360), .C2(n9738), .A(n9195), .B(n9194), .ZN(n9196)
         );
  OAI21_X1 U10525 ( .B1(n9307), .B2(n9364), .A(n9196), .ZN(P1_U3268) );
  XNOR2_X1 U10526 ( .A(n9197), .B(n9199), .ZN(n9369) );
  INV_X1 U10527 ( .A(n9198), .ZN(n9200) );
  OAI21_X1 U10528 ( .B1(n9200), .B2(n9199), .A(n9702), .ZN(n9203) );
  OAI21_X1 U10529 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n9365) );
  AOI211_X1 U10530 ( .C1(n9367), .C2(n9211), .A(n9246), .B(n9204), .ZN(n9366)
         );
  NAND2_X1 U10531 ( .A1(n9366), .A2(n9738), .ZN(n9206) );
  AOI22_X1 U10532 ( .A1(n4968), .A2(n9749), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9754), .ZN(n9205) );
  OAI211_X1 U10533 ( .C1(n9207), .C2(n9720), .A(n9206), .B(n9205), .ZN(n9208)
         );
  AOI21_X1 U10534 ( .B1(n9365), .B2(n9752), .A(n9208), .ZN(n9209) );
  OAI21_X1 U10535 ( .B1(n9369), .B2(n9307), .A(n9209), .ZN(P1_U3269) );
  XNOR2_X1 U10536 ( .A(n9210), .B(n9218), .ZN(n9374) );
  INV_X1 U10537 ( .A(n9211), .ZN(n9212) );
  AOI211_X1 U10538 ( .C1(n9371), .C2(n9227), .A(n9246), .B(n9212), .ZN(n9370)
         );
  AOI22_X1 U10539 ( .A1(n9213), .A2(n9749), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9754), .ZN(n9214) );
  OAI21_X1 U10540 ( .B1(n9215), .B2(n9720), .A(n9214), .ZN(n9222) );
  OAI21_X1 U10541 ( .B1(n9218), .B2(n9217), .A(n9216), .ZN(n9220) );
  AOI21_X1 U10542 ( .B1(n9220), .B2(n9702), .A(n9219), .ZN(n9373) );
  NOR2_X1 U10543 ( .A1(n9373), .A2(n9754), .ZN(n9221) );
  AOI211_X1 U10544 ( .C1(n9370), .C2(n9738), .A(n9222), .B(n9221), .ZN(n9223)
         );
  OAI21_X1 U10545 ( .B1(n9307), .B2(n9374), .A(n9223), .ZN(P1_U3270) );
  XNOR2_X1 U10546 ( .A(n9225), .B(n9224), .ZN(n9379) );
  INV_X1 U10547 ( .A(n9227), .ZN(n9228) );
  AOI211_X1 U10548 ( .C1(n9376), .C2(n9247), .A(n9246), .B(n9228), .ZN(n9375)
         );
  INV_X1 U10549 ( .A(n9229), .ZN(n9230) );
  AOI22_X1 U10550 ( .A1(n9230), .A2(n9749), .B1(n9754), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9231) );
  OAI21_X1 U10551 ( .B1(n6520), .B2(n9720), .A(n9231), .ZN(n9238) );
  AOI211_X1 U10552 ( .C1(n9234), .C2(n9233), .A(n9759), .B(n9232), .ZN(n9236)
         );
  NOR2_X1 U10553 ( .A1(n9236), .A2(n9235), .ZN(n9378) );
  NOR2_X1 U10554 ( .A1(n9378), .A2(n9754), .ZN(n9237) );
  AOI211_X1 U10555 ( .C1(n9375), .C2(n9738), .A(n9238), .B(n9237), .ZN(n9239)
         );
  OAI21_X1 U10556 ( .B1(n9307), .B2(n9379), .A(n9239), .ZN(P1_U3271) );
  XNOR2_X1 U10557 ( .A(n9240), .B(n9242), .ZN(n9384) );
  INV_X1 U10558 ( .A(n9258), .ZN(n9256) );
  OAI21_X1 U10559 ( .B1(n9259), .B2(n9256), .A(n9241), .ZN(n9243) );
  XNOR2_X1 U10560 ( .A(n9243), .B(n9242), .ZN(n9245) );
  AOI21_X1 U10561 ( .B1(n9245), .B2(n9702), .A(n9244), .ZN(n9383) );
  INV_X1 U10562 ( .A(n9383), .ZN(n9254) );
  AOI21_X1 U10563 ( .B1(n9381), .B2(n9267), .A(n9246), .ZN(n9248) );
  AND2_X1 U10564 ( .A1(n9248), .A2(n9247), .ZN(n9380) );
  NAND2_X1 U10565 ( .A1(n9380), .A2(n9738), .ZN(n9251) );
  AOI22_X1 U10566 ( .A1(n9754), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9249), .B2(
        n9749), .ZN(n9250) );
  OAI211_X1 U10567 ( .C1(n9252), .C2(n9720), .A(n9251), .B(n9250), .ZN(n9253)
         );
  AOI21_X1 U10568 ( .B1(n9254), .B2(n9752), .A(n9253), .ZN(n9255) );
  OAI21_X1 U10569 ( .B1(n9384), .B2(n9307), .A(n9255), .ZN(P1_U3272) );
  XNOR2_X1 U10570 ( .A(n9257), .B(n9256), .ZN(n9389) );
  XNOR2_X1 U10571 ( .A(n9259), .B(n9258), .ZN(n9261) );
  AOI21_X1 U10572 ( .B1(n9261), .B2(n9702), .A(n9260), .ZN(n9388) );
  INV_X1 U10573 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9263) );
  OAI22_X1 U10574 ( .A1(n9752), .A2(n9263), .B1(n9262), .B2(n9315), .ZN(n9264)
         );
  AOI21_X1 U10575 ( .B1(n9386), .B2(n9739), .A(n9264), .ZN(n9269) );
  OR2_X1 U10576 ( .A1(n9265), .A2(n9282), .ZN(n9266) );
  AND3_X1 U10577 ( .A1(n9267), .A2(n9734), .A3(n9266), .ZN(n9385) );
  NAND2_X1 U10578 ( .A1(n9385), .A2(n9738), .ZN(n9268) );
  OAI211_X1 U10579 ( .C1(n9388), .C2(n9754), .A(n9269), .B(n9268), .ZN(n9270)
         );
  INV_X1 U10580 ( .A(n9270), .ZN(n9271) );
  OAI21_X1 U10581 ( .B1(n9307), .B2(n9389), .A(n9271), .ZN(P1_U3273) );
  INV_X1 U10582 ( .A(n9276), .ZN(n9273) );
  XNOR2_X1 U10583 ( .A(n9272), .B(n9273), .ZN(n9390) );
  INV_X1 U10584 ( .A(n9390), .ZN(n9290) );
  OAI21_X1 U10585 ( .B1(n9276), .B2(n9275), .A(n9274), .ZN(n9277) );
  NAND2_X1 U10586 ( .A1(n9277), .A2(n9702), .ZN(n9280) );
  AOI22_X1 U10587 ( .A1(n9278), .A2(n9311), .B1(n9309), .B2(n9312), .ZN(n9279)
         );
  NAND2_X1 U10588 ( .A1(n9280), .A2(n9279), .ZN(n9394) );
  OAI21_X1 U10589 ( .B1(n9392), .B2(n9293), .A(n9734), .ZN(n9281) );
  OR2_X1 U10590 ( .A1(n9282), .A2(n9281), .ZN(n9391) );
  OAI22_X1 U10591 ( .A1(n9752), .A2(n9284), .B1(n9283), .B2(n9315), .ZN(n9285)
         );
  AOI21_X1 U10592 ( .B1(n9286), .B2(n9739), .A(n9285), .ZN(n9287) );
  OAI21_X1 U10593 ( .B1(n9391), .B2(n9694), .A(n9287), .ZN(n9288) );
  AOI21_X1 U10594 ( .B1(n9394), .B2(n9752), .A(n9288), .ZN(n9289) );
  OAI21_X1 U10595 ( .B1(n9290), .B2(n9307), .A(n9289), .ZN(P1_U3274) );
  XOR2_X1 U10596 ( .A(n9291), .B(n9299), .Z(n9400) );
  OAI21_X1 U10597 ( .B1(n9297), .B2(n9319), .A(n9734), .ZN(n9292) );
  NAND2_X1 U10598 ( .A1(n9754), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U10599 ( .A1(n9749), .A2(n9294), .ZN(n9295) );
  OAI211_X1 U10600 ( .C1(n9297), .C2(n9720), .A(n9296), .B(n9295), .ZN(n9305)
         );
  OAI21_X1 U10601 ( .B1(n9300), .B2(n9299), .A(n9298), .ZN(n9303) );
  AOI222_X1 U10602 ( .A1(n9702), .A2(n9303), .B1(n9302), .B2(n9311), .C1(n9301), .C2(n9309), .ZN(n9399) );
  NOR2_X1 U10603 ( .A1(n9399), .A2(n9754), .ZN(n9304) );
  AOI211_X1 U10604 ( .C1(n4424), .C2(n9738), .A(n9305), .B(n9304), .ZN(n9306)
         );
  OAI21_X1 U10605 ( .B1(n9307), .B2(n9400), .A(n9306), .ZN(P1_U3275) );
  XOR2_X1 U10606 ( .A(n9308), .B(n9328), .Z(n9313) );
  AOI222_X1 U10607 ( .A1(n9702), .A2(n9313), .B1(n9312), .B2(n9311), .C1(n9310), .C2(n9309), .ZN(n9508) );
  INV_X1 U10608 ( .A(n9314), .ZN(n9316) );
  OAI22_X1 U10609 ( .A1(n9752), .A2(n9317), .B1(n9316), .B2(n9315), .ZN(n9322)
         );
  INV_X1 U10610 ( .A(n9319), .ZN(n9320) );
  OAI211_X1 U10611 ( .C1(n9509), .C2(n4817), .A(n9320), .B(n9734), .ZN(n9507)
         );
  NOR2_X1 U10612 ( .A1(n9507), .A2(n9694), .ZN(n9321) );
  AOI211_X1 U10613 ( .C1(n9739), .C2(n9323), .A(n9322), .B(n9321), .ZN(n9330)
         );
  NAND2_X1 U10614 ( .A1(n7627), .A2(n9324), .ZN(n9326) );
  NAND2_X1 U10615 ( .A1(n9326), .A2(n9325), .ZN(n9327) );
  XOR2_X1 U10616 ( .A(n9328), .B(n9327), .Z(n9511) );
  NAND2_X1 U10617 ( .A1(n9511), .A2(n9715), .ZN(n9329) );
  OAI211_X1 U10618 ( .C1(n9508), .C2(n9754), .A(n9330), .B(n9329), .ZN(
        P1_U3276) );
  OAI211_X1 U10619 ( .C1(n9332), .C2(n9846), .A(n9331), .B(n9337), .ZN(n9406)
         );
  NOR2_X1 U10620 ( .A1(n9334), .A2(n9333), .ZN(n9335) );
  MUX2_X1 U10621 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9406), .S(n10233), .Z(
        P1_U3553) );
  OAI211_X1 U10622 ( .C1(n9339), .C2(n9846), .A(n9338), .B(n9337), .ZN(n9407)
         );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9407), .S(n10233), .Z(
        P1_U3552) );
  AOI21_X1 U10624 ( .B1(n9787), .B2(n9341), .A(n9340), .ZN(n9342) );
  OAI211_X1 U10625 ( .C1(n9344), .C2(n9791), .A(n9343), .B(n9342), .ZN(n9408)
         );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9408), .S(n10233), .Z(
        P1_U3551) );
  AOI21_X1 U10627 ( .B1(n9787), .B2(n9346), .A(n9345), .ZN(n9347) );
  OAI211_X1 U10628 ( .C1(n9349), .C2(n9791), .A(n9348), .B(n9347), .ZN(n9409)
         );
  MUX2_X1 U10629 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9409), .S(n10233), .Z(
        P1_U3550) );
  AOI211_X1 U10630 ( .C1(n9787), .C2(n9352), .A(n9351), .B(n9350), .ZN(n9353)
         );
  OAI21_X1 U10631 ( .B1(n9354), .B2(n9791), .A(n9353), .ZN(n9410) );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9410), .S(n10233), .Z(
        P1_U3549) );
  AOI21_X1 U10633 ( .B1(n9787), .B2(n9356), .A(n9355), .ZN(n9357) );
  OAI211_X1 U10634 ( .C1(n9359), .C2(n9791), .A(n9358), .B(n9357), .ZN(n9411)
         );
  MUX2_X1 U10635 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9411), .S(n10233), .Z(
        P1_U3548) );
  AOI21_X1 U10636 ( .B1(n9787), .B2(n9361), .A(n9360), .ZN(n9362) );
  OAI211_X1 U10637 ( .C1(n9364), .C2(n9791), .A(n9363), .B(n9362), .ZN(n9412)
         );
  MUX2_X1 U10638 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9412), .S(n10233), .Z(
        P1_U3547) );
  AOI211_X1 U10639 ( .C1(n9787), .C2(n9367), .A(n9366), .B(n9365), .ZN(n9368)
         );
  OAI21_X1 U10640 ( .B1(n9369), .B2(n9791), .A(n9368), .ZN(n9413) );
  MUX2_X1 U10641 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9413), .S(n10233), .Z(
        P1_U3546) );
  AOI21_X1 U10642 ( .B1(n9787), .B2(n9371), .A(n9370), .ZN(n9372) );
  OAI211_X1 U10643 ( .C1(n9374), .C2(n9791), .A(n9373), .B(n9372), .ZN(n9414)
         );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9414), .S(n10233), .Z(
        P1_U3545) );
  AOI21_X1 U10645 ( .B1(n9787), .B2(n9376), .A(n9375), .ZN(n9377) );
  OAI211_X1 U10646 ( .C1(n9379), .C2(n9791), .A(n9378), .B(n9377), .ZN(n9415)
         );
  MUX2_X1 U10647 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9415), .S(n10233), .Z(
        P1_U3544) );
  AOI21_X1 U10648 ( .B1(n9787), .B2(n9381), .A(n9380), .ZN(n9382) );
  OAI211_X1 U10649 ( .C1(n9384), .C2(n9791), .A(n9383), .B(n9382), .ZN(n9416)
         );
  MUX2_X1 U10650 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9416), .S(n10233), .Z(
        P1_U3543) );
  AOI21_X1 U10651 ( .B1(n9787), .B2(n9386), .A(n9385), .ZN(n9387) );
  OAI211_X1 U10652 ( .C1(n9389), .C2(n9791), .A(n9388), .B(n9387), .ZN(n9417)
         );
  MUX2_X1 U10653 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9417), .S(n10233), .Z(
        P1_U3542) );
  NAND2_X1 U10654 ( .A1(n9390), .A2(n9842), .ZN(n9396) );
  OAI21_X1 U10655 ( .B1(n9392), .B2(n9846), .A(n9391), .ZN(n9393) );
  NOR2_X1 U10656 ( .A1(n9394), .A2(n9393), .ZN(n9395) );
  NAND2_X1 U10657 ( .A1(n9396), .A2(n9395), .ZN(n9418) );
  MUX2_X1 U10658 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9418), .S(n10233), .Z(
        P1_U3541) );
  AOI21_X1 U10659 ( .B1(n9787), .B2(n9397), .A(n4424), .ZN(n9398) );
  OAI211_X1 U10660 ( .C1(n9400), .C2(n9791), .A(n9399), .B(n9398), .ZN(n9419)
         );
  MUX2_X1 U10661 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9419), .S(n10233), .Z(
        P1_U3540) );
  AOI21_X1 U10662 ( .B1(n9787), .B2(n9402), .A(n9401), .ZN(n9403) );
  OAI211_X1 U10663 ( .C1(n9791), .C2(n9405), .A(n9404), .B(n9403), .ZN(n9420)
         );
  MUX2_X1 U10664 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9420), .S(n10233), .Z(
        P1_U3537) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9406), .S(n9854), .Z(
        P1_U3521) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9407), .S(n9854), .Z(
        P1_U3520) );
  MUX2_X1 U10667 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9408), .S(n9854), .Z(
        P1_U3519) );
  MUX2_X1 U10668 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9409), .S(n9854), .Z(
        P1_U3518) );
  MUX2_X1 U10669 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9410), .S(n9854), .Z(
        P1_U3517) );
  MUX2_X1 U10670 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9411), .S(n9854), .Z(
        P1_U3516) );
  MUX2_X1 U10671 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9412), .S(n9854), .Z(
        P1_U3515) );
  MUX2_X1 U10672 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9413), .S(n9854), .Z(
        P1_U3514) );
  MUX2_X1 U10673 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9414), .S(n9854), .Z(
        P1_U3513) );
  MUX2_X1 U10674 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9415), .S(n9854), .Z(
        P1_U3512) );
  MUX2_X1 U10675 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9416), .S(n9854), .Z(
        P1_U3511) );
  MUX2_X1 U10676 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9417), .S(n9854), .Z(
        P1_U3510) );
  MUX2_X1 U10677 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9418), .S(n9854), .Z(
        P1_U3509) );
  MUX2_X1 U10678 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9419), .S(n9854), .Z(
        P1_U3507) );
  MUX2_X1 U10679 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9420), .S(n9854), .Z(
        P1_U3498) );
  INV_X1 U10680 ( .A(n9421), .ZN(n9422) );
  MUX2_X1 U10681 ( .A(n9424), .B(P1_D_REG_1__SCAN_IN), .S(n9756), .Z(P1_U3440)
         );
  MUX2_X1 U10682 ( .A(n9425), .B(P1_D_REG_0__SCAN_IN), .S(n9756), .Z(P1_U3439)
         );
  INV_X1 U10683 ( .A(n9426), .ZN(n9433) );
  NAND3_X1 U10684 ( .A1(n9427), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9428) );
  NOR4_X1 U10685 ( .A1(n9429), .A2(P1_IR_REG_30__SCAN_IN), .A3(
        P1_IR_REG_28__SCAN_IN), .A4(n9428), .ZN(n9430) );
  AOI21_X1 U10686 ( .B1(n9431), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9430), .ZN(
        n9432) );
  OAI21_X1 U10687 ( .B1(n9433), .B2(n9436), .A(n9432), .ZN(P1_U3324) );
  OAI222_X1 U10688 ( .A1(n9438), .A2(n9437), .B1(n9436), .B2(n9435), .C1(
        P1_U3086), .C2(n9434), .ZN(P1_U3325) );
  INV_X1 U10689 ( .A(n9439), .ZN(n9440) );
  MUX2_X1 U10690 ( .A(n9440), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10691 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9452) );
  INV_X1 U10692 ( .A(n9625), .ZN(n9655) );
  AOI211_X1 U10693 ( .C1(n9443), .C2(n9442), .A(n9441), .B(n9644), .ZN(n9448)
         );
  AOI211_X1 U10694 ( .C1(n9446), .C2(n9445), .A(n9444), .B(n9649), .ZN(n9447)
         );
  AOI211_X1 U10695 ( .C1(n9655), .C2(n9449), .A(n9448), .B(n9447), .ZN(n9451)
         );
  NAND2_X1 U10696 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9450) );
  OAI211_X1 U10697 ( .C1(n9659), .C2(n9452), .A(n9451), .B(n9450), .ZN(
        P1_U3253) );
  INV_X1 U10698 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U10699 ( .A1(n9454), .A2(n9453), .ZN(n9457) );
  INV_X1 U10700 ( .A(n9455), .ZN(n9456) );
  NAND2_X1 U10701 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  OR2_X1 U10702 ( .A1(n9649), .A2(n9458), .ZN(n9466) );
  NAND2_X1 U10703 ( .A1(n9460), .A2(n9459), .ZN(n9463) );
  INV_X1 U10704 ( .A(n9461), .ZN(n9462) );
  NAND2_X1 U10705 ( .A1(n9463), .A2(n9462), .ZN(n9464) );
  OR2_X1 U10706 ( .A1(n9644), .A2(n9464), .ZN(n9465) );
  OAI211_X1 U10707 ( .C1(n9625), .C2(n9467), .A(n9466), .B(n9465), .ZN(n9468)
         );
  INV_X1 U10708 ( .A(n9468), .ZN(n9470) );
  NAND2_X1 U10709 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9469) );
  OAI211_X1 U10710 ( .C1(n9659), .C2(n9471), .A(n9470), .B(n9469), .ZN(
        P1_U3250) );
  INV_X1 U10711 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U10712 ( .A1(n9473), .A2(n9472), .ZN(n9475) );
  NAND2_X1 U10713 ( .A1(n9475), .A2(n9474), .ZN(n9476) );
  OR2_X1 U10714 ( .A1(n9649), .A2(n9476), .ZN(n9483) );
  NAND2_X1 U10715 ( .A1(n9478), .A2(n9477), .ZN(n9480) );
  NAND2_X1 U10716 ( .A1(n9480), .A2(n9479), .ZN(n9481) );
  OR2_X1 U10717 ( .A1(n9644), .A2(n9481), .ZN(n9482) );
  OAI211_X1 U10718 ( .C1(n9625), .C2(n9484), .A(n9483), .B(n9482), .ZN(n9485)
         );
  INV_X1 U10719 ( .A(n9485), .ZN(n9487) );
  NAND2_X1 U10720 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9486) );
  OAI211_X1 U10721 ( .C1(n9488), .C2(n9659), .A(n9487), .B(n9486), .ZN(
        P1_U3246) );
  INV_X1 U10722 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U10723 ( .A1(n9490), .A2(n9489), .ZN(n9493) );
  INV_X1 U10724 ( .A(n9491), .ZN(n9492) );
  NAND2_X1 U10725 ( .A1(n9493), .A2(n9492), .ZN(n9494) );
  OR2_X1 U10726 ( .A1(n9649), .A2(n9494), .ZN(n9502) );
  NAND2_X1 U10727 ( .A1(n9496), .A2(n9495), .ZN(n9499) );
  INV_X1 U10728 ( .A(n9497), .ZN(n9498) );
  NAND2_X1 U10729 ( .A1(n9499), .A2(n9498), .ZN(n9500) );
  OR2_X1 U10730 ( .A1(n9644), .A2(n9500), .ZN(n9501) );
  OAI211_X1 U10731 ( .C1(n9625), .C2(n9503), .A(n9502), .B(n9501), .ZN(n9504)
         );
  INV_X1 U10732 ( .A(n9504), .ZN(n9506) );
  OAI211_X1 U10733 ( .C1(n9659), .C2(n10217), .A(n9506), .B(n9505), .ZN(
        P1_U3251) );
  OAI211_X1 U10734 ( .C1(n9509), .C2(n9846), .A(n9508), .B(n9507), .ZN(n9510)
         );
  AOI21_X1 U10735 ( .B1(n9511), .B2(n9842), .A(n9510), .ZN(n9519) );
  AOI22_X1 U10736 ( .A1(n10233), .A2(n9519), .B1(n9093), .B2(n9878), .ZN(
        P1_U3539) );
  INV_X1 U10737 ( .A(n9512), .ZN(n9515) );
  OAI211_X1 U10738 ( .C1(n9515), .C2(n9846), .A(n9514), .B(n9513), .ZN(n9516)
         );
  AOI21_X1 U10739 ( .B1(n9517), .B2(n9842), .A(n9516), .ZN(n9521) );
  AOI22_X1 U10740 ( .A1(n10233), .A2(n9521), .B1(n9069), .B2(n9878), .ZN(
        P1_U3538) );
  INV_X1 U10741 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9518) );
  AOI22_X1 U10742 ( .A1(n9854), .A2(n9519), .B1(n9518), .B2(n9852), .ZN(
        P1_U3504) );
  INV_X1 U10743 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9520) );
  AOI22_X1 U10744 ( .A1(n9854), .A2(n9521), .B1(n9520), .B2(n9852), .ZN(
        P1_U3501) );
  XNOR2_X1 U10745 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10746 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U10747 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9522), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9540) );
  NAND2_X1 U10748 ( .A1(n9524), .A2(n9523), .ZN(n9527) );
  INV_X1 U10749 ( .A(n9525), .ZN(n9526) );
  NAND2_X1 U10750 ( .A1(n9527), .A2(n9526), .ZN(n9528) );
  OR2_X1 U10751 ( .A1(n9649), .A2(n9528), .ZN(n9536) );
  NAND2_X1 U10752 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9529) );
  NAND2_X1 U10753 ( .A1(n9530), .A2(n9529), .ZN(n9533) );
  INV_X1 U10754 ( .A(n9531), .ZN(n9532) );
  NAND2_X1 U10755 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  OR2_X1 U10756 ( .A1(n9644), .A2(n9534), .ZN(n9535) );
  OAI211_X1 U10757 ( .C1(n9625), .C2(n9537), .A(n9536), .B(n9535), .ZN(n9538)
         );
  INV_X1 U10758 ( .A(n9538), .ZN(n9539) );
  NAND2_X1 U10759 ( .A1(n9540), .A2(n9539), .ZN(P1_U3244) );
  INV_X1 U10760 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U10761 ( .A1(n9542), .A2(n9541), .ZN(n9543) );
  NAND2_X1 U10762 ( .A1(n9543), .A2(n4663), .ZN(n9544) );
  OR2_X1 U10763 ( .A1(n9649), .A2(n9544), .ZN(n9550) );
  OAI21_X1 U10764 ( .B1(n9547), .B2(n9546), .A(n9545), .ZN(n9548) );
  OR2_X1 U10765 ( .A1(n9644), .A2(n9548), .ZN(n9549) );
  OAI211_X1 U10766 ( .C1(n9625), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9552)
         );
  INV_X1 U10767 ( .A(n9552), .ZN(n9554) );
  NAND2_X1 U10768 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9553) );
  OAI211_X1 U10769 ( .C1(n10066), .C2(n9659), .A(n9554), .B(n9553), .ZN(
        P1_U3248) );
  INV_X1 U10770 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U10771 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  NAND2_X1 U10772 ( .A1(n4661), .A2(n9557), .ZN(n9558) );
  OR2_X1 U10773 ( .A1(n9649), .A2(n9558), .ZN(n9564) );
  NAND2_X1 U10774 ( .A1(n9560), .A2(n9559), .ZN(n9561) );
  NAND2_X1 U10775 ( .A1(n9561), .A2(n4442), .ZN(n9562) );
  OR2_X1 U10776 ( .A1(n9644), .A2(n9562), .ZN(n9563) );
  OAI211_X1 U10777 ( .C1(n9625), .C2(n9565), .A(n9564), .B(n9563), .ZN(n9566)
         );
  INV_X1 U10778 ( .A(n9566), .ZN(n9568) );
  NAND2_X1 U10779 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9567) );
  OAI211_X1 U10780 ( .C1(n9659), .C2(n9569), .A(n9568), .B(n9567), .ZN(
        P1_U3249) );
  INV_X1 U10781 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9588) );
  INV_X1 U10782 ( .A(n9570), .ZN(n9584) );
  NAND2_X1 U10783 ( .A1(n4440), .A2(n9571), .ZN(n9572) );
  NAND2_X1 U10784 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  OR2_X1 U10785 ( .A1(n9649), .A2(n9574), .ZN(n9583) );
  INV_X1 U10786 ( .A(n9575), .ZN(n9578) );
  INV_X1 U10787 ( .A(n9576), .ZN(n9577) );
  NAND2_X1 U10788 ( .A1(n9578), .A2(n9577), .ZN(n9579) );
  NAND2_X1 U10789 ( .A1(n9580), .A2(n9579), .ZN(n9581) );
  OR2_X1 U10790 ( .A1(n9644), .A2(n9581), .ZN(n9582) );
  OAI211_X1 U10791 ( .C1(n9625), .C2(n9584), .A(n9583), .B(n9582), .ZN(n9585)
         );
  INV_X1 U10792 ( .A(n9585), .ZN(n9587) );
  NAND2_X1 U10793 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9586) );
  OAI211_X1 U10794 ( .C1(n9659), .C2(n9588), .A(n9587), .B(n9586), .ZN(
        P1_U3254) );
  INV_X1 U10795 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9608) );
  INV_X1 U10796 ( .A(n9589), .ZN(n9604) );
  NAND2_X1 U10797 ( .A1(n9591), .A2(n9590), .ZN(n9594) );
  INV_X1 U10798 ( .A(n9592), .ZN(n9593) );
  NAND2_X1 U10799 ( .A1(n9594), .A2(n9593), .ZN(n9595) );
  OR2_X1 U10800 ( .A1(n9649), .A2(n9595), .ZN(n9603) );
  NAND2_X1 U10801 ( .A1(n9597), .A2(n9596), .ZN(n9600) );
  INV_X1 U10802 ( .A(n9598), .ZN(n9599) );
  NAND2_X1 U10803 ( .A1(n9600), .A2(n9599), .ZN(n9601) );
  OR2_X1 U10804 ( .A1(n9644), .A2(n9601), .ZN(n9602) );
  OAI211_X1 U10805 ( .C1(n9625), .C2(n9604), .A(n9603), .B(n9602), .ZN(n9605)
         );
  INV_X1 U10806 ( .A(n9605), .ZN(n9607) );
  NAND2_X1 U10807 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9606) );
  OAI211_X1 U10808 ( .C1(n9659), .C2(n9608), .A(n9607), .B(n9606), .ZN(
        P1_U3256) );
  INV_X1 U10809 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9629) );
  INV_X1 U10810 ( .A(n9609), .ZN(n9624) );
  NAND2_X1 U10811 ( .A1(n9611), .A2(n9610), .ZN(n9614) );
  INV_X1 U10812 ( .A(n9612), .ZN(n9613) );
  NAND2_X1 U10813 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  OR2_X1 U10814 ( .A1(n9649), .A2(n9615), .ZN(n9623) );
  NAND2_X1 U10815 ( .A1(n9617), .A2(n9616), .ZN(n9620) );
  INV_X1 U10816 ( .A(n9618), .ZN(n9619) );
  NAND2_X1 U10817 ( .A1(n9620), .A2(n9619), .ZN(n9621) );
  OR2_X1 U10818 ( .A1(n9644), .A2(n9621), .ZN(n9622) );
  OAI211_X1 U10819 ( .C1(n9625), .C2(n9624), .A(n9623), .B(n9622), .ZN(n9626)
         );
  INV_X1 U10820 ( .A(n9626), .ZN(n9628) );
  NAND2_X1 U10821 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9627) );
  OAI211_X1 U10822 ( .C1(n9659), .C2(n9629), .A(n9628), .B(n9627), .ZN(
        P1_U3257) );
  INV_X1 U10823 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9641) );
  AOI211_X1 U10824 ( .C1(n9632), .C2(n9631), .A(n9630), .B(n9644), .ZN(n9637)
         );
  AOI211_X1 U10825 ( .C1(n9635), .C2(n9634), .A(n9633), .B(n9649), .ZN(n9636)
         );
  AOI211_X1 U10826 ( .C1(n9655), .C2(n9638), .A(n9637), .B(n9636), .ZN(n9640)
         );
  NAND2_X1 U10827 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9639) );
  OAI211_X1 U10828 ( .C1(n9659), .C2(n9641), .A(n9640), .B(n9639), .ZN(
        P1_U3258) );
  INV_X1 U10829 ( .A(n9642), .ZN(n9643) );
  AOI211_X1 U10830 ( .C1(n9646), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9653)
         );
  INV_X1 U10831 ( .A(n9647), .ZN(n9648) );
  AOI211_X1 U10832 ( .C1(n9651), .C2(n9650), .A(n9649), .B(n9648), .ZN(n9652)
         );
  AOI211_X1 U10833 ( .C1(n9655), .C2(n9654), .A(n9653), .B(n9652), .ZN(n9658)
         );
  NAND2_X1 U10834 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9657) );
  OAI211_X1 U10835 ( .C1(n9659), .C2(n10015), .A(n9658), .B(n9657), .ZN(
        P1_U3261) );
  NAND2_X1 U10836 ( .A1(n9660), .A2(n9682), .ZN(n9661) );
  XNOR2_X1 U10837 ( .A(n9661), .B(n9667), .ZN(n9664) );
  INV_X1 U10838 ( .A(n9662), .ZN(n9663) );
  AOI21_X1 U10839 ( .B1(n9664), .B2(n9702), .A(n9663), .ZN(n9832) );
  AOI222_X1 U10840 ( .A1(n9665), .A2(n9739), .B1(n4962), .B2(n9749), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n9754), .ZN(n9672) );
  XNOR2_X1 U10841 ( .A(n9666), .B(n9667), .ZN(n9835) );
  OAI21_X1 U10842 ( .B1(n9687), .B2(n9833), .A(n9734), .ZN(n9668) );
  OR2_X1 U10843 ( .A1(n9669), .A2(n9668), .ZN(n9831) );
  INV_X1 U10844 ( .A(n9831), .ZN(n9670) );
  AOI22_X1 U10845 ( .A1(n9835), .A2(n9715), .B1(n9738), .B2(n9670), .ZN(n9671)
         );
  OAI211_X1 U10846 ( .C1(n9754), .C2(n9832), .A(n9672), .B(n9671), .ZN(
        P1_U3281) );
  NAND2_X1 U10847 ( .A1(n9673), .A2(n9705), .ZN(n9675) );
  NAND2_X1 U10848 ( .A1(n9675), .A2(n9674), .ZN(n9676) );
  XNOR2_X1 U10849 ( .A(n9676), .B(n9678), .ZN(n9829) );
  INV_X1 U10850 ( .A(n9677), .ZN(n9685) );
  INV_X1 U10851 ( .A(n9660), .ZN(n9683) );
  INV_X1 U10852 ( .A(n9678), .ZN(n9679) );
  OAI21_X1 U10853 ( .B1(n9680), .B2(n9679), .A(n9702), .ZN(n9681) );
  AOI21_X1 U10854 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n9684) );
  AOI211_X1 U10855 ( .C1(n9732), .C2(n9829), .A(n9685), .B(n9684), .ZN(n9826)
         );
  INV_X1 U10856 ( .A(n9686), .ZN(n9736) );
  INV_X1 U10857 ( .A(n9708), .ZN(n9689) );
  INV_X1 U10858 ( .A(n9687), .ZN(n9688) );
  OAI211_X1 U10859 ( .C1(n4769), .C2(n9689), .A(n9688), .B(n9734), .ZN(n9825)
         );
  AOI22_X1 U10860 ( .A1(n9754), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9690), .B2(
        n9749), .ZN(n9693) );
  NAND2_X1 U10861 ( .A1(n9691), .A2(n9739), .ZN(n9692) );
  OAI211_X1 U10862 ( .C1(n9825), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9695)
         );
  AOI21_X1 U10863 ( .B1(n9829), .B2(n9736), .A(n9695), .ZN(n9696) );
  OAI21_X1 U10864 ( .B1(n9754), .B2(n9826), .A(n9696), .ZN(P1_U3282) );
  OAI21_X1 U10865 ( .B1(n9699), .B2(n9698), .A(n9697), .ZN(n9703) );
  INV_X1 U10866 ( .A(n9700), .ZN(n9701) );
  AOI21_X1 U10867 ( .B1(n9703), .B2(n9702), .A(n9701), .ZN(n9820) );
  AOI222_X1 U10868 ( .A1(n9818), .A2(n9739), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n9754), .C1(n9749), .C2(n9704), .ZN(n9712) );
  XNOR2_X1 U10869 ( .A(n9673), .B(n9705), .ZN(n9823) );
  OAI21_X1 U10870 ( .B1(n9707), .B2(n4343), .A(n9818), .ZN(n9709) );
  NAND3_X1 U10871 ( .A1(n9709), .A2(n9734), .A3(n9708), .ZN(n9819) );
  INV_X1 U10872 ( .A(n9819), .ZN(n9710) );
  AOI22_X1 U10873 ( .A1(n9823), .A2(n9715), .B1(n9738), .B2(n9710), .ZN(n9711)
         );
  OAI211_X1 U10874 ( .C1(n9754), .C2(n9820), .A(n9712), .B(n9711), .ZN(
        P1_U3283) );
  INV_X1 U10875 ( .A(n9713), .ZN(n9714) );
  AOI22_X1 U10876 ( .A1(n9716), .A2(n9715), .B1(n9738), .B2(n9714), .ZN(n9725)
         );
  INV_X1 U10877 ( .A(n9717), .ZN(n9723) );
  AOI22_X1 U10878 ( .A1(n9754), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9718), .B2(
        n9749), .ZN(n9719) );
  OAI21_X1 U10879 ( .B1(n9721), .B2(n9720), .A(n9719), .ZN(n9722) );
  AOI21_X1 U10880 ( .B1(n9723), .B2(n9752), .A(n9722), .ZN(n9724) );
  NAND2_X1 U10881 ( .A1(n9725), .A2(n9724), .ZN(P1_U3287) );
  XNOR2_X1 U10882 ( .A(n9727), .B(n9726), .ZN(n9771) );
  XNOR2_X1 U10883 ( .A(n9728), .B(n9727), .ZN(n9729) );
  NOR2_X1 U10884 ( .A1(n9729), .A2(n9759), .ZN(n9730) );
  AOI211_X1 U10885 ( .C1(n9732), .C2(n9771), .A(n9731), .B(n9730), .ZN(n9768)
         );
  AOI22_X1 U10886 ( .A1(n9754), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9749), .ZN(n9742) );
  OAI211_X1 U10887 ( .C1(n9767), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9766)
         );
  INV_X1 U10888 ( .A(n9766), .ZN(n9737) );
  AOI222_X1 U10889 ( .A1(n9740), .A2(n9739), .B1(n9738), .B2(n9737), .C1(n9771), .C2(n9736), .ZN(n9741) );
  OAI211_X1 U10890 ( .C1(n9754), .C2(n9768), .A(n9742), .B(n9741), .ZN(
        P1_U3292) );
  INV_X1 U10891 ( .A(n9758), .ZN(n9744) );
  NAND3_X1 U10892 ( .A1(n9744), .A2(n9743), .A3(n9746), .ZN(n9751) );
  OAI21_X1 U10893 ( .B1(n9747), .B2(n9746), .A(n9745), .ZN(n9748) );
  AOI22_X1 U10894 ( .A1(n9749), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9762), .B2(
        n9748), .ZN(n9750) );
  AND3_X1 U10895 ( .A1(n9751), .A2(n9750), .A3(n9757), .ZN(n9753) );
  AOI22_X1 U10896 ( .A1(n9754), .A2(n6594), .B1(n9753), .B2(n9752), .ZN(
        P1_U3293) );
  AND2_X1 U10897 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9756), .ZN(P1_U3294) );
  AND2_X1 U10898 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9756), .ZN(P1_U3295) );
  AND2_X1 U10899 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9756), .ZN(P1_U3296) );
  AND2_X1 U10900 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9756), .ZN(P1_U3297) );
  AND2_X1 U10901 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9756), .ZN(P1_U3298) );
  AND2_X1 U10902 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9756), .ZN(P1_U3299) );
  AND2_X1 U10903 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9756), .ZN(P1_U3300) );
  INV_X1 U10904 ( .A(n9756), .ZN(n9755) );
  INV_X1 U10905 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10085) );
  NOR2_X1 U10906 ( .A1(n9755), .A2(n10085), .ZN(P1_U3301) );
  AND2_X1 U10907 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9756), .ZN(P1_U3302) );
  AND2_X1 U10908 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9756), .ZN(P1_U3303) );
  AND2_X1 U10909 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9756), .ZN(P1_U3304) );
  AND2_X1 U10910 ( .A1(n9756), .A2(P1_D_REG_20__SCAN_IN), .ZN(P1_U3305) );
  AND2_X1 U10911 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9756), .ZN(P1_U3306) );
  AND2_X1 U10912 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9756), .ZN(P1_U3307) );
  AND2_X1 U10913 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9756), .ZN(P1_U3308) );
  AND2_X1 U10914 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9756), .ZN(P1_U3309) );
  AND2_X1 U10915 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9756), .ZN(P1_U3310) );
  AND2_X1 U10916 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9756), .ZN(P1_U3311) );
  AND2_X1 U10917 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9756), .ZN(P1_U3312) );
  AND2_X1 U10918 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9756), .ZN(P1_U3313) );
  AND2_X1 U10919 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9756), .ZN(P1_U3314) );
  INV_X1 U10920 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U10921 ( .A1(n9755), .A2(n10219), .ZN(P1_U3315) );
  AND2_X1 U10922 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9756), .ZN(P1_U3316) );
  AND2_X1 U10923 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9756), .ZN(P1_U3317) );
  AND2_X1 U10924 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9756), .ZN(P1_U3318) );
  AND2_X1 U10925 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9756), .ZN(P1_U3319) );
  AND2_X1 U10926 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9756), .ZN(P1_U3320) );
  INV_X1 U10927 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10078) );
  NOR2_X1 U10928 ( .A1(n9755), .A2(n10078), .ZN(P1_U3321) );
  AND2_X1 U10929 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9756), .ZN(P1_U3322) );
  AND2_X1 U10930 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9756), .ZN(P1_U3323) );
  INV_X1 U10931 ( .A(n9757), .ZN(n9761) );
  AOI21_X1 U10932 ( .B1(n9759), .B2(n9791), .A(n9758), .ZN(n9760) );
  AOI211_X1 U10933 ( .C1(n9763), .C2(n9762), .A(n9761), .B(n9760), .ZN(n9856)
         );
  INV_X1 U10934 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9764) );
  AOI22_X1 U10935 ( .A1(n9854), .A2(n9856), .B1(n9764), .B2(n9852), .ZN(
        P1_U3453) );
  INV_X1 U10936 ( .A(n9765), .ZN(n9851) );
  OAI21_X1 U10937 ( .B1(n9767), .B2(n9846), .A(n9766), .ZN(n9770) );
  INV_X1 U10938 ( .A(n9768), .ZN(n9769) );
  AOI211_X1 U10939 ( .C1(n9851), .C2(n9771), .A(n9770), .B(n9769), .ZN(n9857)
         );
  INV_X1 U10940 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U10941 ( .A1(n9854), .A2(n9857), .B1(n9772), .B2(n9852), .ZN(
        P1_U3456) );
  OAI21_X1 U10942 ( .B1(n9774), .B2(n9846), .A(n9773), .ZN(n9776) );
  AOI211_X1 U10943 ( .C1(n9842), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9859)
         );
  INV_X1 U10944 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U10945 ( .A1(n9854), .A2(n9859), .B1(n9778), .B2(n9852), .ZN(
        P1_U3459) );
  OAI21_X1 U10946 ( .B1(n9780), .B2(n9846), .A(n9779), .ZN(n9782) );
  AOI211_X1 U10947 ( .C1(n9842), .C2(n9783), .A(n9782), .B(n9781), .ZN(n9861)
         );
  INV_X1 U10948 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U10949 ( .A1(n9854), .A2(n9861), .B1(n9784), .B2(n9852), .ZN(
        P1_U3462) );
  AOI21_X1 U10950 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n9788) );
  OAI211_X1 U10951 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9792)
         );
  INV_X1 U10952 ( .A(n9792), .ZN(n9863) );
  INV_X1 U10953 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10954 ( .A1(n9854), .A2(n9863), .B1(n9793), .B2(n9852), .ZN(
        P1_U3465) );
  OAI21_X1 U10955 ( .B1(n9795), .B2(n9846), .A(n9794), .ZN(n9797) );
  AOI211_X1 U10956 ( .C1(n9842), .C2(n9798), .A(n9797), .B(n9796), .ZN(n9865)
         );
  INV_X1 U10957 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U10958 ( .A1(n9854), .A2(n9865), .B1(n9799), .B2(n9852), .ZN(
        P1_U3468) );
  AND2_X1 U10959 ( .A1(n9800), .A2(n9842), .ZN(n9804) );
  OAI21_X1 U10960 ( .B1(n9802), .B2(n9846), .A(n9801), .ZN(n9803) );
  NOR3_X1 U10961 ( .A1(n9805), .A2(n9804), .A3(n9803), .ZN(n9867) );
  INV_X1 U10962 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9806) );
  AOI22_X1 U10963 ( .A1(n9854), .A2(n9867), .B1(n9806), .B2(n9852), .ZN(
        P1_U3474) );
  AND2_X1 U10964 ( .A1(n9807), .A2(n9842), .ZN(n9811) );
  OAI21_X1 U10965 ( .B1(n9809), .B2(n9846), .A(n9808), .ZN(n9810) );
  NOR3_X1 U10966 ( .A1(n9812), .A2(n9811), .A3(n9810), .ZN(n9869) );
  INV_X1 U10967 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10070) );
  AOI22_X1 U10968 ( .A1(n9854), .A2(n9869), .B1(n10070), .B2(n9852), .ZN(
        P1_U3477) );
  OAI21_X1 U10969 ( .B1(n4569), .B2(n9846), .A(n9813), .ZN(n9815) );
  AOI211_X1 U10970 ( .C1(n9842), .C2(n9816), .A(n9815), .B(n9814), .ZN(n9871)
         );
  INV_X1 U10971 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9817) );
  AOI22_X1 U10972 ( .A1(n9854), .A2(n9871), .B1(n9817), .B2(n9852), .ZN(
        P1_U3480) );
  INV_X1 U10973 ( .A(n9818), .ZN(n9821) );
  OAI211_X1 U10974 ( .C1(n9821), .C2(n9846), .A(n9820), .B(n9819), .ZN(n9822)
         );
  AOI21_X1 U10975 ( .B1(n9842), .B2(n9823), .A(n9822), .ZN(n9872) );
  INV_X1 U10976 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9824) );
  AOI22_X1 U10977 ( .A1(n9854), .A2(n9872), .B1(n9824), .B2(n9852), .ZN(
        P1_U3483) );
  OAI21_X1 U10978 ( .B1(n4769), .B2(n9846), .A(n9825), .ZN(n9828) );
  INV_X1 U10979 ( .A(n9826), .ZN(n9827) );
  AOI211_X1 U10980 ( .C1(n9851), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9874)
         );
  INV_X1 U10981 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9830) );
  AOI22_X1 U10982 ( .A1(n9854), .A2(n9874), .B1(n9830), .B2(n9852), .ZN(
        P1_U3486) );
  OAI211_X1 U10983 ( .C1(n9833), .C2(n9846), .A(n9832), .B(n9831), .ZN(n9834)
         );
  AOI21_X1 U10984 ( .B1(n9842), .B2(n9835), .A(n9834), .ZN(n9876) );
  INV_X1 U10985 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U10986 ( .A1(n9854), .A2(n9876), .B1(n9836), .B2(n9852), .ZN(
        P1_U3489) );
  OAI211_X1 U10987 ( .C1(n9839), .C2(n9846), .A(n9838), .B(n9837), .ZN(n9840)
         );
  AOI21_X1 U10988 ( .B1(n9842), .B2(n9841), .A(n9840), .ZN(n9877) );
  INV_X1 U10989 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U10990 ( .A1(n9854), .A2(n9877), .B1(n9843), .B2(n9852), .ZN(
        P1_U3492) );
  INV_X1 U10991 ( .A(n9844), .ZN(n9850) );
  OAI21_X1 U10992 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(n9849) );
  AOI211_X1 U10993 ( .C1(n9851), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9879)
         );
  INV_X1 U10994 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9853) );
  AOI22_X1 U10995 ( .A1(n9854), .A2(n9879), .B1(n9853), .B2(n9852), .ZN(
        P1_U3495) );
  AOI22_X1 U10996 ( .A1(n10233), .A2(n9856), .B1(n9855), .B2(n9878), .ZN(
        P1_U3522) );
  AOI22_X1 U10997 ( .A1(n10233), .A2(n9857), .B1(n6624), .B2(n9878), .ZN(
        P1_U3523) );
  INV_X1 U10998 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U10999 ( .A1(n10233), .A2(n9859), .B1(n9858), .B2(n9878), .ZN(
        P1_U3524) );
  INV_X1 U11000 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9860) );
  AOI22_X1 U11001 ( .A1(n10233), .A2(n9861), .B1(n9860), .B2(n9878), .ZN(
        P1_U3525) );
  AOI22_X1 U11002 ( .A1(n10233), .A2(n9863), .B1(n9862), .B2(n9878), .ZN(
        P1_U3526) );
  INV_X1 U11003 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9864) );
  AOI22_X1 U11004 ( .A1(n10233), .A2(n9865), .B1(n9864), .B2(n9878), .ZN(
        P1_U3527) );
  INV_X1 U11005 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9866) );
  AOI22_X1 U11006 ( .A1(n10233), .A2(n9867), .B1(n9866), .B2(n9878), .ZN(
        P1_U3529) );
  INV_X1 U11007 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U11008 ( .A1(n10233), .A2(n9869), .B1(n9868), .B2(n9878), .ZN(
        P1_U3530) );
  AOI22_X1 U11009 ( .A1(n10233), .A2(n9871), .B1(n9870), .B2(n9878), .ZN(
        P1_U3531) );
  AOI22_X1 U11010 ( .A1(n10233), .A2(n9872), .B1(n6998), .B2(n9878), .ZN(
        P1_U3532) );
  AOI22_X1 U11011 ( .A1(n10233), .A2(n9874), .B1(n9873), .B2(n9878), .ZN(
        P1_U3533) );
  AOI22_X1 U11012 ( .A1(n10233), .A2(n9876), .B1(n9875), .B2(n9878), .ZN(
        P1_U3534) );
  AOI22_X1 U11013 ( .A1(n10233), .A2(n9877), .B1(n9061), .B2(n9878), .ZN(
        P1_U3535) );
  AOI22_X1 U11014 ( .A1(n10233), .A2(n9879), .B1(n9064), .B2(n9878), .ZN(
        P1_U3536) );
  INV_X1 U11015 ( .A(n9880), .ZN(n9881) );
  AOI21_X1 U11016 ( .B1(n6692), .B2(n9882), .A(n9881), .ZN(n9888) );
  NAND2_X1 U11017 ( .A1(P2_U3151), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9887) );
  OAI211_X1 U11018 ( .C1(n9885), .C2(n9884), .A(n9883), .B(n9906), .ZN(n9886)
         );
  OAI211_X1 U11019 ( .C1(n9889), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9890)
         );
  AOI21_X1 U11020 ( .B1(n4592), .B2(n9891), .A(n9890), .ZN(n9898) );
  INV_X1 U11021 ( .A(n9892), .ZN(n9893) );
  AOI21_X1 U11022 ( .B1(n6955), .B2(n9894), .A(n9893), .ZN(n9895) );
  OR2_X1 U11023 ( .A1(n9896), .A2(n9895), .ZN(n9897) );
  OAI211_X1 U11024 ( .C1(n10013), .C2(n9899), .A(n9898), .B(n9897), .ZN(
        P2_U3183) );
  OAI21_X1 U11025 ( .B1(n9902), .B2(n9901), .A(n9900), .ZN(n9903) );
  AOI22_X1 U11026 ( .A1(n9905), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n9904), .B2(
        n9903), .ZN(n9911) );
  OAI211_X1 U11027 ( .C1(n9909), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9910)
         );
  OAI211_X1 U11028 ( .C1(n9913), .C2(n9912), .A(n9911), .B(n9910), .ZN(n9914)
         );
  INV_X1 U11029 ( .A(n9914), .ZN(n9921) );
  OAI21_X1 U11030 ( .B1(n9917), .B2(n9916), .A(n9915), .ZN(n9918) );
  NAND2_X1 U11031 ( .A1(n9919), .A2(n9918), .ZN(n9920) );
  OAI211_X1 U11032 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5791), .A(n9921), .B(
        n9920), .ZN(P2_U3184) );
  NAND2_X1 U11033 ( .A1(n9923), .A2(n9922), .ZN(n9925) );
  XNOR2_X1 U11034 ( .A(n9924), .B(n9938), .ZN(n9926) );
  XNOR2_X1 U11035 ( .A(n9925), .B(n9926), .ZN(n9966) );
  XNOR2_X1 U11036 ( .A(n9927), .B(n9926), .ZN(n9929) );
  NAND2_X1 U11037 ( .A1(n9929), .A2(n9928), .ZN(n9935) );
  AOI22_X1 U11038 ( .A1(n9933), .A2(n9932), .B1(n9931), .B2(n9930), .ZN(n9934)
         );
  NAND2_X1 U11039 ( .A1(n9935), .A2(n9934), .ZN(n9964) );
  MUX2_X1 U11040 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9964), .S(n8733), .Z(n9941)
         );
  OAI22_X1 U11041 ( .A1(n9939), .A2(n9938), .B1(n9937), .B2(n9936), .ZN(n9940)
         );
  NOR2_X1 U11042 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  OAI21_X1 U11043 ( .B1(n9943), .B2(n9966), .A(n9942), .ZN(P2_U3227) );
  INV_X1 U11044 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9947) );
  OAI22_X1 U11045 ( .A1(n9944), .A2(n9982), .B1(n4339), .B2(n9989), .ZN(n9945)
         );
  NOR2_X1 U11046 ( .A1(n9946), .A2(n9945), .ZN(n9998) );
  AOI22_X1 U11047 ( .A1(n9997), .A2(n9947), .B1(n9998), .B2(n9995), .ZN(
        P2_U3393) );
  AOI22_X1 U11048 ( .A1(n9950), .A2(n9949), .B1(n9987), .B2(n9948), .ZN(n9951)
         );
  AND2_X1 U11049 ( .A1(n9952), .A2(n9951), .ZN(n9999) );
  AOI22_X1 U11050 ( .A1(n9997), .A2(n5794), .B1(n9999), .B2(n9995), .ZN(
        P2_U3396) );
  INV_X1 U11051 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9958) );
  INV_X1 U11052 ( .A(n9953), .ZN(n9957) );
  OAI22_X1 U11053 ( .A1(n9955), .A2(n9965), .B1(n9954), .B2(n9989), .ZN(n9956)
         );
  NOR2_X1 U11054 ( .A1(n9957), .A2(n9956), .ZN(n10001) );
  AOI22_X1 U11055 ( .A1(n9997), .A2(n9958), .B1(n10001), .B2(n9995), .ZN(
        P2_U3399) );
  INV_X1 U11056 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9963) );
  OAI22_X1 U11057 ( .A1(n9960), .A2(n9982), .B1(n9959), .B2(n9989), .ZN(n9961)
         );
  NOR2_X1 U11058 ( .A1(n9962), .A2(n9961), .ZN(n10002) );
  AOI22_X1 U11059 ( .A1(n9997), .A2(n9963), .B1(n10002), .B2(n9995), .ZN(
        P2_U3405) );
  INV_X1 U11060 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9971) );
  INV_X1 U11061 ( .A(n9964), .ZN(n9970) );
  OR2_X1 U11062 ( .A1(n9966), .A2(n9965), .ZN(n9969) );
  NAND2_X1 U11063 ( .A1(n9987), .A2(n9967), .ZN(n9968) );
  AOI22_X1 U11064 ( .A1(n9997), .A2(n9971), .B1(n10003), .B2(n9995), .ZN(
        P2_U3408) );
  INV_X1 U11065 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9976) );
  OAI22_X1 U11066 ( .A1(n9973), .A2(n9982), .B1(n9972), .B2(n9989), .ZN(n9974)
         );
  NOR2_X1 U11067 ( .A1(n9975), .A2(n9974), .ZN(n10004) );
  AOI22_X1 U11068 ( .A1(n9997), .A2(n9976), .B1(n10004), .B2(n9995), .ZN(
        P2_U3411) );
  INV_X1 U11069 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U11070 ( .A1(n9977), .A2(n9982), .ZN(n9979) );
  AOI211_X1 U11071 ( .C1(n9987), .C2(n9980), .A(n9979), .B(n9978), .ZN(n10005)
         );
  AOI22_X1 U11072 ( .A1(n9997), .A2(n9981), .B1(n10005), .B2(n9995), .ZN(
        P2_U3417) );
  INV_X1 U11073 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9988) );
  NOR2_X1 U11074 ( .A1(n9983), .A2(n9982), .ZN(n9985) );
  AOI211_X1 U11075 ( .C1(n9987), .C2(n9986), .A(n9985), .B(n9984), .ZN(n10006)
         );
  AOI22_X1 U11076 ( .A1(n9997), .A2(n9988), .B1(n10006), .B2(n9995), .ZN(
        P2_U3420) );
  INV_X1 U11077 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U11078 ( .A1(n9990), .A2(n9989), .ZN(n9992) );
  AOI211_X1 U11079 ( .C1(n9994), .C2(n9993), .A(n9992), .B(n9991), .ZN(n10007)
         );
  AOI22_X1 U11080 ( .A1(n9997), .A2(n9996), .B1(n10007), .B2(n9995), .ZN(
        P2_U3423) );
  AOI22_X1 U11081 ( .A1(n10008), .A2(n9998), .B1(n6692), .B2(n6287), .ZN(
        P2_U3460) );
  AOI22_X1 U11082 ( .A1(n10008), .A2(n9999), .B1(n5792), .B2(n6287), .ZN(
        P2_U3461) );
  AOI22_X1 U11083 ( .A1(n10008), .A2(n10001), .B1(n10000), .B2(n6287), .ZN(
        P2_U3462) );
  AOI22_X1 U11084 ( .A1(n10008), .A2(n10002), .B1(n6793), .B2(n6287), .ZN(
        P2_U3464) );
  AOI22_X1 U11085 ( .A1(n10008), .A2(n10003), .B1(n5849), .B2(n6287), .ZN(
        P2_U3465) );
  AOI22_X1 U11086 ( .A1(n10008), .A2(n10004), .B1(n5864), .B2(n6287), .ZN(
        P2_U3466) );
  AOI22_X1 U11087 ( .A1(n10008), .A2(n10005), .B1(n5902), .B2(n6287), .ZN(
        P2_U3468) );
  AOI22_X1 U11088 ( .A1(n10008), .A2(n10006), .B1(n7361), .B2(n6287), .ZN(
        P2_U3469) );
  AOI22_X1 U11089 ( .A1(n10008), .A2(n10007), .B1(n5927), .B2(n6287), .ZN(
        P2_U3470) );
  OAI222_X1 U11090 ( .A1(n10013), .A2(n10012), .B1(n10013), .B2(n10011), .C1(
        n10010), .C2(n10009), .ZN(ADD_1068_U5) );
  XOR2_X1 U11091 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11092 ( .B1(n10016), .B2(n10015), .A(n10014), .ZN(n10018) );
  XNOR2_X1 U11093 ( .A(n10018), .B(n10017), .ZN(ADD_1068_U55) );
  OAI21_X1 U11094 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(ADD_1068_U56) );
  OAI21_X1 U11095 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(ADD_1068_U57) );
  OAI21_X1 U11096 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(ADD_1068_U58) );
  OAI21_X1 U11097 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(ADD_1068_U59) );
  OAI21_X1 U11098 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(ADD_1068_U60) );
  OAI21_X1 U11099 ( .B1(n10036), .B2(n10035), .A(n10034), .ZN(ADD_1068_U61) );
  OAI21_X1 U11100 ( .B1(n10039), .B2(n10038), .A(n10037), .ZN(ADD_1068_U62) );
  OAI21_X1 U11101 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(ADD_1068_U63) );
  AOI22_X1 U11102 ( .A1(n10208), .A2(keyinput120), .B1(keyinput122), .B2(n4573), .ZN(n10043) );
  OAI221_X1 U11103 ( .B1(n10208), .B2(keyinput120), .C1(n4573), .C2(
        keyinput122), .A(n10043), .ZN(n10051) );
  AOI22_X1 U11104 ( .A1(n6793), .A2(keyinput112), .B1(n10218), .B2(keyinput89), 
        .ZN(n10044) );
  OAI221_X1 U11105 ( .B1(n6793), .B2(keyinput112), .C1(n10218), .C2(keyinput89), .A(n10044), .ZN(n10050) );
  XNOR2_X1 U11106 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput119), .ZN(n10048)
         );
  XNOR2_X1 U11107 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput86), .ZN(n10047) );
  XNOR2_X1 U11108 ( .A(P2_REG0_REG_25__SCAN_IN), .B(keyinput65), .ZN(n10046)
         );
  XNOR2_X1 U11109 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput77), .ZN(n10045) );
  NAND4_X1 U11110 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10049) );
  NOR3_X1 U11111 ( .A1(n10051), .A2(n10050), .A3(n10049), .ZN(n10093) );
  AOI22_X1 U11112 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(keyinput93), .B1(n10195), 
        .B2(keyinput115), .ZN(n10052) );
  OAI221_X1 U11113 ( .B1(P1_REG1_REG_27__SCAN_IN), .B2(keyinput93), .C1(n10195), .C2(keyinput115), .A(n10052), .ZN(n10063) );
  AOI22_X1 U11114 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(keyinput97), .B1(
        P1_REG1_REG_20__SCAN_IN), .B2(keyinput100), .ZN(n10053) );
  OAI221_X1 U11115 ( .B1(P2_REG2_REG_24__SCAN_IN), .B2(keyinput97), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput100), .A(n10053), .ZN(n10062) );
  AOI22_X1 U11116 ( .A1(n10056), .A2(keyinput109), .B1(n10055), .B2(keyinput83), .ZN(n10054) );
  OAI221_X1 U11117 ( .B1(n10056), .B2(keyinput109), .C1(n10055), .C2(
        keyinput83), .A(n10054), .ZN(n10061) );
  AOI22_X1 U11118 ( .A1(n10059), .A2(keyinput70), .B1(keyinput71), .B2(n10058), 
        .ZN(n10057) );
  OAI221_X1 U11119 ( .B1(n10059), .B2(keyinput70), .C1(n10058), .C2(keyinput71), .A(n10057), .ZN(n10060) );
  NOR4_X1 U11120 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n10092) );
  AOI22_X1 U11121 ( .A1(n10200), .A2(keyinput92), .B1(n10167), .B2(keyinput118), .ZN(n10064) );
  OAI221_X1 U11122 ( .B1(n10200), .B2(keyinput92), .C1(n10167), .C2(
        keyinput118), .A(n10064), .ZN(n10075) );
  AOI22_X1 U11123 ( .A1(n10199), .A2(keyinput85), .B1(keyinput126), .B2(n10066), .ZN(n10065) );
  OAI221_X1 U11124 ( .B1(n10199), .B2(keyinput85), .C1(n10066), .C2(
        keyinput126), .A(n10065), .ZN(n10074) );
  INV_X1 U11125 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10068) );
  AOI22_X1 U11126 ( .A1(n10068), .A2(keyinput81), .B1(n6993), .B2(keyinput84), 
        .ZN(n10067) );
  OAI221_X1 U11127 ( .B1(n10068), .B2(keyinput81), .C1(n6993), .C2(keyinput84), 
        .A(n10067), .ZN(n10073) );
  AOI22_X1 U11128 ( .A1(n10071), .A2(keyinput106), .B1(n10070), .B2(keyinput95), .ZN(n10069) );
  OAI221_X1 U11129 ( .B1(n10071), .B2(keyinput106), .C1(n10070), .C2(
        keyinput95), .A(n10069), .ZN(n10072) );
  NOR4_X1 U11130 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n10091) );
  INV_X1 U11131 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U11132 ( .A1(n10187), .A2(keyinput75), .B1(n10077), .B2(keyinput67), 
        .ZN(n10076) );
  OAI221_X1 U11133 ( .B1(n10187), .B2(keyinput75), .C1(n10077), .C2(keyinput67), .A(n10076), .ZN(n10081) );
  XNOR2_X1 U11134 ( .A(n10078), .B(keyinput78), .ZN(n10080) );
  XOR2_X1 U11135 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput82), .Z(n10079) );
  OR3_X1 U11136 ( .A1(n10081), .A2(n10080), .A3(n10079), .ZN(n10089) );
  INV_X1 U11137 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10083) );
  AOI22_X1 U11138 ( .A1(n10083), .A2(keyinput105), .B1(n10219), .B2(keyinput88), .ZN(n10082) );
  OAI221_X1 U11139 ( .B1(n10083), .B2(keyinput105), .C1(n10219), .C2(
        keyinput88), .A(n10082), .ZN(n10088) );
  AOI22_X1 U11140 ( .A1(n10086), .A2(keyinput103), .B1(n10085), .B2(
        keyinput102), .ZN(n10084) );
  OAI221_X1 U11141 ( .B1(n10086), .B2(keyinput103), .C1(n10085), .C2(
        keyinput102), .A(n10084), .ZN(n10087) );
  NOR3_X1 U11142 ( .A1(n10089), .A2(n10088), .A3(n10087), .ZN(n10090) );
  AND4_X1 U11143 ( .A1(n10093), .A2(n10092), .A3(n10091), .A4(n10090), .ZN(
        n10230) );
  OAI22_X1 U11144 ( .A1(P2_D_REG_12__SCAN_IN), .A2(keyinput87), .B1(
        keyinput104), .B2(P2_REG0_REG_14__SCAN_IN), .ZN(n10094) );
  AOI221_X1 U11145 ( .B1(P2_D_REG_12__SCAN_IN), .B2(keyinput87), .C1(
        P2_REG0_REG_14__SCAN_IN), .C2(keyinput104), .A(n10094), .ZN(n10101) );
  OAI22_X1 U11146 ( .A1(P2_D_REG_28__SCAN_IN), .A2(keyinput99), .B1(keyinput66), .B2(P1_WR_REG_SCAN_IN), .ZN(n10095) );
  AOI221_X1 U11147 ( .B1(P2_D_REG_28__SCAN_IN), .B2(keyinput99), .C1(
        P1_WR_REG_SCAN_IN), .C2(keyinput66), .A(n10095), .ZN(n10100) );
  OAI22_X1 U11148 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(keyinput69), .B1(
        keyinput101), .B2(P1_REG1_REG_21__SCAN_IN), .ZN(n10096) );
  AOI221_X1 U11149 ( .B1(P1_REG2_REG_23__SCAN_IN), .B2(keyinput69), .C1(
        P1_REG1_REG_21__SCAN_IN), .C2(keyinput101), .A(n10096), .ZN(n10099) );
  OAI22_X1 U11150 ( .A1(P1_B_REG_SCAN_IN), .A2(keyinput124), .B1(
        P2_IR_REG_12__SCAN_IN), .B2(keyinput94), .ZN(n10097) );
  AOI221_X1 U11151 ( .B1(P1_B_REG_SCAN_IN), .B2(keyinput124), .C1(keyinput94), 
        .C2(P2_IR_REG_12__SCAN_IN), .A(n10097), .ZN(n10098) );
  NAND4_X1 U11152 ( .A1(n10101), .A2(n10100), .A3(n10099), .A4(n10098), .ZN(
        n10129) );
  OAI22_X1 U11153 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput113), .B1(
        keyinput96), .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n10102) );
  AOI221_X1 U11154 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput113), .C1(
        P1_DATAO_REG_16__SCAN_IN), .C2(keyinput96), .A(n10102), .ZN(n10109) );
  OAI22_X1 U11155 ( .A1(P1_D_REG_20__SCAN_IN), .A2(keyinput90), .B1(
        P2_REG0_REG_13__SCAN_IN), .B2(keyinput108), .ZN(n10103) );
  AOI221_X1 U11156 ( .B1(P1_D_REG_20__SCAN_IN), .B2(keyinput90), .C1(
        keyinput108), .C2(P2_REG0_REG_13__SCAN_IN), .A(n10103), .ZN(n10108) );
  OAI22_X1 U11157 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput73), .B1(
        keyinput127), .B2(P2_ADDR_REG_18__SCAN_IN), .ZN(n10104) );
  AOI221_X1 U11158 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput73), .C1(
        P2_ADDR_REG_18__SCAN_IN), .C2(keyinput127), .A(n10104), .ZN(n10107) );
  OAI22_X1 U11159 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput107), .B1(
        keyinput123), .B2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10105) );
  AOI221_X1 U11160 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput107), .C1(
        P1_ADDR_REG_8__SCAN_IN), .C2(keyinput123), .A(n10105), .ZN(n10106) );
  NAND4_X1 U11161 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n10128) );
  OAI22_X1 U11162 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput91), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput121), .ZN(n10110) );
  AOI221_X1 U11163 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput91), .C1(
        keyinput121), .C2(P2_DATAO_REG_15__SCAN_IN), .A(n10110), .ZN(n10117)
         );
  OAI22_X1 U11164 ( .A1(SI_0_), .A2(keyinput114), .B1(P1_ADDR_REG_6__SCAN_IN), 
        .B2(keyinput68), .ZN(n10111) );
  AOI221_X1 U11165 ( .B1(SI_0_), .B2(keyinput114), .C1(keyinput68), .C2(
        P1_ADDR_REG_6__SCAN_IN), .A(n10111), .ZN(n10116) );
  OAI22_X1 U11166 ( .A1(SI_8_), .A2(keyinput72), .B1(keyinput79), .B2(
        P2_D_REG_9__SCAN_IN), .ZN(n10112) );
  AOI221_X1 U11167 ( .B1(SI_8_), .B2(keyinput72), .C1(P2_D_REG_9__SCAN_IN), 
        .C2(keyinput79), .A(n10112), .ZN(n10115) );
  OAI22_X1 U11168 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput125), .B1(
        P2_REG1_REG_1__SCAN_IN), .B2(keyinput117), .ZN(n10113) );
  AOI221_X1 U11169 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput125), .C1(
        keyinput117), .C2(P2_REG1_REG_1__SCAN_IN), .A(n10113), .ZN(n10114) );
  NAND4_X1 U11170 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10127) );
  OAI22_X1 U11171 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(keyinput64), .B1(SI_30_), .B2(keyinput110), .ZN(n10118) );
  AOI221_X1 U11172 ( .B1(P1_DATAO_REG_10__SCAN_IN), .B2(keyinput64), .C1(
        keyinput110), .C2(SI_30_), .A(n10118), .ZN(n10125) );
  OAI22_X1 U11173 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(keyinput74), .B1(
        P2_D_REG_23__SCAN_IN), .B2(keyinput116), .ZN(n10119) );
  AOI221_X1 U11174 ( .B1(P2_IR_REG_22__SCAN_IN), .B2(keyinput74), .C1(
        keyinput116), .C2(P2_D_REG_23__SCAN_IN), .A(n10119), .ZN(n10124) );
  OAI22_X1 U11175 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput111), .B1(keyinput80), .B2(P1_ADDR_REG_12__SCAN_IN), .ZN(n10120) );
  AOI221_X1 U11176 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput111), .C1(
        P1_ADDR_REG_12__SCAN_IN), .C2(keyinput80), .A(n10120), .ZN(n10123) );
  OAI22_X1 U11177 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput98), .B1(keyinput76), .B2(P1_REG0_REG_6__SCAN_IN), .ZN(n10121) );
  AOI221_X1 U11178 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput98), .C1(
        P1_REG0_REG_6__SCAN_IN), .C2(keyinput76), .A(n10121), .ZN(n10122) );
  NAND4_X1 U11179 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10126) );
  NOR4_X1 U11180 ( .A1(n10129), .A2(n10128), .A3(n10127), .A4(n10126), .ZN(
        n10229) );
  AOI22_X1 U11181 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(keyinput0), .B1(
        P1_D_REG_24__SCAN_IN), .B2(keyinput38), .ZN(n10130) );
  OAI221_X1 U11182 ( .B1(P1_DATAO_REG_10__SCAN_IN), .B2(keyinput0), .C1(
        P1_D_REG_24__SCAN_IN), .C2(keyinput38), .A(n10130), .ZN(n10137) );
  AOI22_X1 U11183 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput55), .B1(
        P1_REG1_REG_21__SCAN_IN), .B2(keyinput37), .ZN(n10131) );
  OAI221_X1 U11184 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput55), .C1(
        P1_REG1_REG_21__SCAN_IN), .C2(keyinput37), .A(n10131), .ZN(n10136) );
  AOI22_X1 U11185 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(keyinput62), .B1(
        P1_REG3_REG_5__SCAN_IN), .B2(keyinput6), .ZN(n10132) );
  OAI221_X1 U11186 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(keyinput62), .C1(
        P1_REG3_REG_5__SCAN_IN), .C2(keyinput6), .A(n10132), .ZN(n10135) );
  AOI22_X1 U11187 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(keyinput44), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput27), .ZN(n10133) );
  OAI221_X1 U11188 ( .B1(P2_REG0_REG_13__SCAN_IN), .B2(keyinput44), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput27), .A(n10133), .ZN(n10134) );
  NOR4_X1 U11189 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10165) );
  AOI22_X1 U11190 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(keyinput4), .B1(SI_0_), 
        .B2(keyinput50), .ZN(n10138) );
  OAI221_X1 U11191 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(keyinput4), .C1(SI_0_), 
        .C2(keyinput50), .A(n10138), .ZN(n10145) );
  AOI22_X1 U11192 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput58), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(keyinput19), .ZN(n10139) );
  OAI221_X1 U11193 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput58), .C1(
        P1_DATAO_REG_24__SCAN_IN), .C2(keyinput19), .A(n10139), .ZN(n10144) );
  AOI22_X1 U11194 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(keyinput30), .B1(
        P1_D_REG_1__SCAN_IN), .B2(keyinput47), .ZN(n10140) );
  OAI221_X1 U11195 ( .B1(P2_IR_REG_12__SCAN_IN), .B2(keyinput30), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput47), .A(n10140), .ZN(n10143) );
  AOI22_X1 U11196 ( .A1(P1_REG1_REG_29__SCAN_IN), .A2(keyinput41), .B1(SI_28_), 
        .B2(keyinput45), .ZN(n10141) );
  OAI221_X1 U11197 ( .B1(P1_REG1_REG_29__SCAN_IN), .B2(keyinput41), .C1(SI_28_), .C2(keyinput45), .A(n10141), .ZN(n10142) );
  NOR4_X1 U11198 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10164) );
  AOI22_X1 U11199 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(keyinput40), .B1(
        P1_REG2_REG_2__SCAN_IN), .B2(keyinput7), .ZN(n10146) );
  OAI221_X1 U11200 ( .B1(P2_REG0_REG_14__SCAN_IN), .B2(keyinput40), .C1(
        P1_REG2_REG_2__SCAN_IN), .C2(keyinput7), .A(n10146), .ZN(n10153) );
  AOI22_X1 U11201 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput14), .B1(
        P1_D_REG_20__SCAN_IN), .B2(keyinput26), .ZN(n10147) );
  OAI221_X1 U11202 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput14), .C1(
        P1_D_REG_20__SCAN_IN), .C2(keyinput26), .A(n10147), .ZN(n10152) );
  AOI22_X1 U11203 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(keyinput39), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput22), .ZN(n10148) );
  OAI221_X1 U11204 ( .B1(P1_DATAO_REG_22__SCAN_IN), .B2(keyinput39), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput22), .A(n10148), .ZN(n10151) );
  AOI22_X1 U11205 ( .A1(P2_D_REG_23__SCAN_IN), .A2(keyinput52), .B1(
        P2_D_REG_9__SCAN_IN), .B2(keyinput15), .ZN(n10149) );
  OAI221_X1 U11206 ( .B1(P2_D_REG_23__SCAN_IN), .B2(keyinput52), .C1(
        P2_D_REG_9__SCAN_IN), .C2(keyinput15), .A(n10149), .ZN(n10150) );
  NOR4_X1 U11207 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10163) );
  AOI22_X1 U11208 ( .A1(P2_D_REG_12__SCAN_IN), .A2(keyinput23), .B1(
        P1_REG2_REG_23__SCAN_IN), .B2(keyinput5), .ZN(n10154) );
  OAI221_X1 U11209 ( .B1(P2_D_REG_12__SCAN_IN), .B2(keyinput23), .C1(
        P1_REG2_REG_23__SCAN_IN), .C2(keyinput5), .A(n10154), .ZN(n10161) );
  AOI22_X1 U11210 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput9), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput3), .ZN(n10155) );
  OAI221_X1 U11211 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput9), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput3), .A(n10155), .ZN(n10160) );
  AOI22_X1 U11212 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(keyinput53), .B1(
        P2_REG1_REG_17__SCAN_IN), .B2(keyinput42), .ZN(n10156) );
  OAI221_X1 U11213 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(keyinput53), .C1(
        P2_REG1_REG_17__SCAN_IN), .C2(keyinput42), .A(n10156), .ZN(n10159) );
  AOI22_X1 U11214 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput61), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(keyinput32), .ZN(n10157) );
  OAI221_X1 U11215 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput61), .C1(
        P1_DATAO_REG_16__SCAN_IN), .C2(keyinput32), .A(n10157), .ZN(n10158) );
  NOR4_X1 U11216 ( .A1(n10161), .A2(n10160), .A3(n10159), .A4(n10158), .ZN(
        n10162) );
  NAND4_X1 U11217 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10228) );
  AOI22_X1 U11218 ( .A1(n10167), .A2(keyinput54), .B1(keyinput48), .B2(n6793), 
        .ZN(n10166) );
  OAI221_X1 U11219 ( .B1(n10167), .B2(keyinput54), .C1(n6793), .C2(keyinput48), 
        .A(n10166), .ZN(n10178) );
  AOI22_X1 U11220 ( .A1(n10170), .A2(keyinput57), .B1(n10169), .B2(keyinput49), 
        .ZN(n10168) );
  OAI221_X1 U11221 ( .B1(n10170), .B2(keyinput57), .C1(n10169), .C2(keyinput49), .A(n10168), .ZN(n10177) );
  AOI22_X1 U11222 ( .A1(n5788), .A2(keyinput43), .B1(keyinput35), .B2(n10172), 
        .ZN(n10171) );
  OAI221_X1 U11223 ( .B1(n5788), .B2(keyinput43), .C1(n10172), .C2(keyinput35), 
        .A(n10171), .ZN(n10176) );
  INV_X1 U11224 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U11225 ( .A1(n8599), .A2(keyinput33), .B1(n10174), .B2(keyinput12), 
        .ZN(n10173) );
  OAI221_X1 U11226 ( .B1(n8599), .B2(keyinput33), .C1(n10174), .C2(keyinput12), 
        .A(n10173), .ZN(n10175) );
  NOR4_X1 U11227 ( .A1(n10178), .A2(n10177), .A3(n10176), .A4(n10175), .ZN(
        n10226) );
  AOI22_X1 U11228 ( .A1(P2_REG0_REG_4__SCAN_IN), .A2(keyinput17), .B1(
        P1_REG0_REG_8__SCAN_IN), .B2(keyinput31), .ZN(n10179) );
  OAI221_X1 U11229 ( .B1(P2_REG0_REG_4__SCAN_IN), .B2(keyinput17), .C1(
        P1_REG0_REG_8__SCAN_IN), .C2(keyinput31), .A(n10179), .ZN(n10180) );
  INV_X1 U11230 ( .A(n10180), .ZN(n10191) );
  AOI22_X1 U11231 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(keyinput63), .B1(
        P1_REG1_REG_20__SCAN_IN), .B2(keyinput36), .ZN(n10181) );
  OAI221_X1 U11232 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(keyinput63), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput36), .A(n10181), .ZN(n10182) );
  INV_X1 U11233 ( .A(n10182), .ZN(n10190) );
  XNOR2_X1 U11234 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput13), .ZN(n10185) );
  XNOR2_X1 U11235 ( .A(SI_8_), .B(keyinput8), .ZN(n10184) );
  XNOR2_X1 U11236 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput34), .ZN(n10183) );
  AND3_X1 U11237 ( .A1(n10185), .A2(n10184), .A3(n10183), .ZN(n10189) );
  INV_X1 U11238 ( .A(keyinput11), .ZN(n10186) );
  XNOR2_X1 U11239 ( .A(n10187), .B(n10186), .ZN(n10188) );
  AND4_X1 U11240 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n10225) );
  AOI22_X1 U11241 ( .A1(n10193), .A2(keyinput1), .B1(n6993), .B2(keyinput20), 
        .ZN(n10192) );
  OAI221_X1 U11242 ( .B1(n10193), .B2(keyinput1), .C1(n6993), .C2(keyinput20), 
        .A(n10192), .ZN(n10206) );
  AOI22_X1 U11243 ( .A1(n10196), .A2(keyinput16), .B1(n10195), .B2(keyinput51), 
        .ZN(n10194) );
  OAI221_X1 U11244 ( .B1(n10196), .B2(keyinput16), .C1(n10195), .C2(keyinput51), .A(n10194), .ZN(n10205) );
  INV_X1 U11245 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U11246 ( .A1(n10199), .A2(keyinput21), .B1(n10198), .B2(keyinput29), 
        .ZN(n10197) );
  OAI221_X1 U11247 ( .B1(n10199), .B2(keyinput21), .C1(n10198), .C2(keyinput29), .A(n10197), .ZN(n10204) );
  XOR2_X1 U11248 ( .A(n10200), .B(keyinput28), .Z(n10202) );
  XNOR2_X1 U11249 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput10), .ZN(n10201) );
  NAND2_X1 U11250 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  NOR4_X1 U11251 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10224) );
  INV_X1 U11252 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10209) );
  AOI22_X1 U11253 ( .A1(n10209), .A2(keyinput2), .B1(n10208), .B2(keyinput56), 
        .ZN(n10207) );
  OAI221_X1 U11254 ( .B1(n10209), .B2(keyinput2), .C1(n10208), .C2(keyinput56), 
        .A(n10207), .ZN(n10215) );
  AOI22_X1 U11255 ( .A1(n10212), .A2(keyinput46), .B1(n10211), .B2(keyinput60), 
        .ZN(n10210) );
  OAI221_X1 U11256 ( .B1(n10212), .B2(keyinput46), .C1(n10211), .C2(keyinput60), .A(n10210), .ZN(n10214) );
  XOR2_X1 U11257 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput18), .Z(n10213) );
  OR3_X1 U11258 ( .A1(n10215), .A2(n10214), .A3(n10213), .ZN(n10222) );
  AOI22_X1 U11259 ( .A1(n10218), .A2(keyinput25), .B1(keyinput59), .B2(n10217), 
        .ZN(n10216) );
  OAI221_X1 U11260 ( .B1(n10218), .B2(keyinput25), .C1(n10217), .C2(keyinput59), .A(n10216), .ZN(n10221) );
  XNOR2_X1 U11261 ( .A(n10219), .B(keyinput24), .ZN(n10220) );
  NOR3_X1 U11262 ( .A1(n10222), .A2(n10221), .A3(n10220), .ZN(n10223) );
  NAND4_X1 U11263 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10223), .ZN(
        n10227) );
  AOI211_X1 U11264 ( .C1(n10230), .C2(n10229), .A(n10228), .B(n10227), .ZN(
        n10235) );
  NAND2_X1 U11265 ( .A1(n10231), .A2(n10233), .ZN(n10232) );
  OAI21_X1 U11266 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10233), .A(n10232), .ZN(
        n10234) );
  XNOR2_X1 U11267 ( .A(n10235), .B(n10234), .ZN(P1_U3528) );
  OAI21_X1 U11268 ( .B1(n10238), .B2(n10237), .A(n10236), .ZN(ADD_1068_U51) );
  OAI21_X1 U11269 ( .B1(n10241), .B2(n10240), .A(n10239), .ZN(ADD_1068_U47) );
  OAI21_X1 U11270 ( .B1(n10244), .B2(n10243), .A(n10242), .ZN(ADD_1068_U50) );
  OAI21_X1 U11271 ( .B1(n10247), .B2(n10246), .A(n10245), .ZN(ADD_1068_U49) );
  OAI21_X1 U11272 ( .B1(n10250), .B2(n10249), .A(n10248), .ZN(ADD_1068_U48) );
  AOI21_X1 U11273 ( .B1(n10253), .B2(n10252), .A(n10251), .ZN(ADD_1068_U54) );
  AOI21_X1 U11274 ( .B1(n10256), .B2(n10255), .A(n10254), .ZN(ADD_1068_U53) );
  OAI21_X1 U11275 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4851 ( .A(n8244), .Z(n8245) );
  CLKBUF_X1 U4878 ( .A(n5151), .Z(n5520) );
  CLKBUF_X1 U4963 ( .A(n9706), .Z(n4343) );
  CLKBUF_X1 U9808 ( .A(n6429), .Z(n9740) );
endmodule

