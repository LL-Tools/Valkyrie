

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4269, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10293;

  NAND2_X1 U4774 ( .A1(n9449), .A2(n8053), .ZN(n9730) );
  AND2_X1 U4776 ( .A1(n8084), .A2(n8083), .ZN(n8147) );
  XNOR2_X1 U4777 ( .A(n7993), .B(n7988), .ZN(n8084) );
  NOR4_X1 U4778 ( .A1(n8410), .A2(n5936), .A3(n8435), .A4(n5861), .ZN(n5862)
         );
  NAND2_X1 U4779 ( .A1(n8036), .A2(n8035), .ZN(n9228) );
  AND2_X1 U4780 ( .A1(n9216), .A2(n9145), .ZN(n9530) );
  OR2_X1 U4781 ( .A1(n8438), .A2(n8017), .ZN(n5826) );
  NAND2_X1 U4782 ( .A1(n7839), .A2(n5851), .ZN(n7750) );
  NAND2_X2 U4783 ( .A1(n9982), .A2(n9353), .ZN(n9207) );
  INV_X1 U4784 ( .A(n6710), .ZN(n8880) );
  AND2_X1 U4785 ( .A1(n5304), .A2(n4287), .ZN(n7308) );
  INV_X4 U4786 ( .A(n6035), .ZN(n6091) );
  OAI211_X1 U4787 ( .C1(n5038), .C2(n6334), .A(n6332), .B(n6333), .ZN(n6754)
         );
  BUF_X1 U4788 ( .A(n5294), .Z(n4276) );
  INV_X1 U4790 ( .A(n8390), .ZN(n7373) );
  AND2_X2 U4791 ( .A1(n5988), .A2(n4670), .ZN(n6057) );
  NAND2_X1 U4792 ( .A1(n6650), .A2(n6005), .ZN(n5263) );
  INV_X1 U4793 ( .A(n5214), .ZN(n5494) );
  OR2_X1 U4794 ( .A1(n5067), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4419) );
  CLKBUF_X1 U4795 ( .A(n5276), .Z(n4269) );
  INV_X1 U4797 ( .A(n10293), .ZN(n4271) );
  INV_X1 U4798 ( .A(n5839), .ZN(n5837) );
  NAND2_X1 U4799 ( .A1(n7541), .A2(n8262), .ZN(n5738) );
  NOR2_X1 U4800 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5179) );
  INV_X1 U4801 ( .A(n5699), .ZN(n5670) );
  INV_X1 U4802 ( .A(n7936), .ZN(n5216) );
  NAND2_X1 U4803 ( .A1(n9818), .A2(n9095), .ZN(n9195) );
  NAND2_X1 U4804 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6038) );
  INV_X1 U4805 ( .A(n7124), .ZN(n7998) );
  INV_X1 U4806 ( .A(n5279), .ZN(n10043) );
  NAND2_X1 U4807 ( .A1(n8426), .A2(n5931), .ZN(n5932) );
  INV_X1 U4809 ( .A(n5900), .ZN(n7378) );
  INV_X1 U4810 ( .A(n8259), .ZN(n7474) );
  NAND2_X1 U4811 ( .A1(n5850), .A2(n7862), .ZN(n7850) );
  NAND2_X1 U4812 ( .A1(n5754), .A2(n5751), .ZN(n7690) );
  BUF_X1 U4813 ( .A(n5481), .Z(n5500) );
  INV_X1 U4814 ( .A(n7053), .ZN(n4860) );
  INV_X1 U4815 ( .A(n4807), .ZN(n9054) );
  AND4_X1 U4816 ( .A1(n5440), .A2(n5439), .A3(n5438), .A4(n5437), .ZN(n8172)
         );
  OAI211_X1 U4817 ( .C1(n6650), .C2(n6837), .A(n5278), .B(n5277), .ZN(n5279)
         );
  XNOR2_X1 U4818 ( .A(n4439), .B(n5313), .ZN(n6433) );
  OR2_X1 U4819 ( .A1(n4273), .A2(n7375), .ZN(n8620) );
  INV_X2 U4820 ( .A(n8645), .ZN(n4273) );
  AND2_X1 U4821 ( .A1(n6123), .A2(n6122), .ZN(n9902) );
  AND2_X1 U4822 ( .A1(n7690), .A2(n5910), .ZN(n4272) );
  AND2_X2 U4823 ( .A1(n9545), .A2(n9142), .ZN(n9566) );
  XNOR2_X1 U4824 ( .A(n8688), .B(n8519), .ZN(n8502) );
  INV_X1 U4825 ( .A(n7580), .ZN(n5943) );
  NAND2_X2 U4826 ( .A1(n8358), .A2(n8357), .ZN(n8374) );
  NAND2_X2 U4827 ( .A1(n6001), .A2(n6000), .ZN(n6613) );
  INV_X2 U4828 ( .A(n6335), .ZN(n9356) );
  OAI21_X2 U4829 ( .B1(n8865), .B2(n8866), .A(n8864), .ZN(n8908) );
  NAND2_X2 U4830 ( .A1(n5907), .A2(n5906), .ZN(n7657) );
  NAND2_X2 U4831 ( .A1(n7474), .A2(n5900), .ZN(n5848) );
  INV_X2 U4832 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10195) );
  INV_X1 U4833 ( .A(n7028), .ZN(n7268) );
  XNOR2_X2 U4834 ( .A(n5213), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7028) );
  XNOR2_X2 U4835 ( .A(n5061), .B(SI_3_), .ZN(n5256) );
  NAND2_X2 U4836 ( .A1(n4419), .A2(n5045), .ZN(n5061) );
  NAND2_X2 U4837 ( .A1(n6249), .A2(n6248), .ZN(n9571) );
  AOI22_X2 U4838 ( .A1(n9361), .A2(n9360), .B1(n9359), .B2(n9358), .ZN(n9374)
         );
  NOR2_X2 U4839 ( .A1(n5366), .A2(n5086), .ZN(n5386) );
  AOI211_X2 U4840 ( .C1(n9957), .C2(n9768), .A(n9767), .B(n9766), .ZN(n9769)
         );
  XNOR2_X2 U4841 ( .A(n9228), .B(n9462), .ZN(n9273) );
  AOI21_X2 U4842 ( .B1(n9486), .B2(n9315), .A(n9242), .ZN(n8043) );
  NAND2_X2 U4843 ( .A1(n6206), .A2(n6205), .ZN(n9624) );
  AOI21_X2 U4844 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10110), .ZN(n10109) );
  XOR2_X2 U4845 ( .A(n9883), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10269) );
  AOI21_X2 U4846 ( .B1(n9498), .B2(n9311), .A(n9147), .ZN(n9486) );
  NAND2_X1 U4847 ( .A1(n6294), .A2(n6293), .ZN(n9474) );
  OR2_X1 U4848 ( .A1(n8673), .A2(n8437), .ZN(n5817) );
  NAND2_X1 U4849 ( .A1(n9768), .A2(n9534), .ZN(n9531) );
  OAI21_X1 U4850 ( .B1(n5528), .B2(n5136), .A(n5139), .ZN(n5571) );
  NAND2_X1 U4851 ( .A1(n9299), .A2(n9070), .ZN(n6348) );
  INV_X1 U4853 ( .A(n9352), .ZN(n7568) );
  INV_X1 U4854 ( .A(n7073), .ZN(n9972) );
  INV_X1 U4855 ( .A(n8636), .ZN(n7156) );
  INV_X1 U4856 ( .A(n8761), .ZN(n7541) );
  INV_X2 U4857 ( .A(n5674), .ZN(n5282) );
  INV_X4 U4858 ( .A(n7991), .ZN(n8012) );
  CLKBUF_X3 U4859 ( .A(n6057), .Z(n9057) );
  OR2_X1 U4860 ( .A1(n7018), .A2(n5718), .ZN(n7991) );
  OR2_X1 U4861 ( .A1(n5203), .A2(n5270), .ZN(n5202) );
  INV_X1 U4862 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5449) );
  INV_X1 U4863 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n10129) );
  INV_X1 U4864 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5333) );
  INV_X1 U4865 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6698) );
  AOI21_X1 U4866 ( .B1(n5942), .B2(n8614), .A(n7937), .ZN(n7932) );
  NAND2_X1 U4867 ( .A1(n4719), .A2(n4932), .ZN(n9029) );
  AOI211_X1 U4868 ( .C1(n8762), .C2(n8673), .A(n8672), .B(n8671), .ZN(n8674)
         );
  NAND2_X1 U4869 ( .A1(n8875), .A2(n8952), .ZN(n4719) );
  AOI21_X1 U4870 ( .B1(n8660), .B2(n10066), .A(n8663), .ZN(n4441) );
  NAND2_X1 U4871 ( .A1(n4394), .A2(n7119), .ZN(n5868) );
  OAI21_X1 U4872 ( .B1(n4466), .B2(n8532), .A(n8614), .ZN(n4465) );
  OAI21_X1 U4873 ( .B1(n9546), .B2(n9547), .A(n9708), .ZN(n4479) );
  AND2_X1 U4874 ( .A1(n5841), .A2(n4310), .ZN(n4728) );
  AND2_X1 U4875 ( .A1(n4610), .A2(n4348), .ZN(n4609) );
  NAND2_X1 U4876 ( .A1(n4906), .A2(n9245), .ZN(n9529) );
  INV_X1 U4877 ( .A(n9443), .ZN(n9721) );
  NAND2_X1 U4878 ( .A1(n4928), .A2(n4324), .ZN(n9005) );
  CLKBUF_X1 U4879 ( .A(n5704), .Z(n8651) );
  NOR2_X1 U4880 ( .A1(n9489), .A2(n9474), .ZN(n4507) );
  NAND2_X1 U4881 ( .A1(n8834), .A2(n8833), .ZN(n9014) );
  XNOR2_X1 U4882 ( .A(n5689), .B(n5688), .ZN(n9055) );
  NAND2_X1 U4883 ( .A1(n9068), .A2(n9067), .ZN(n9725) );
  AND2_X1 U4884 ( .A1(n5195), .A2(n5194), .ZN(n8659) );
  AND2_X1 U4885 ( .A1(n5043), .A2(n5019), .ZN(n5018) );
  AND2_X1 U4886 ( .A1(n4907), .A2(n9121), .ZN(n4905) );
  AND2_X2 U4887 ( .A1(n9457), .A2(n9225), .ZN(n9316) );
  NAND2_X1 U4888 ( .A1(n9736), .A2(n8903), .ZN(n9226) );
  AND2_X1 U4889 ( .A1(n9530), .A2(n4498), .ZN(n4907) );
  OR2_X1 U4890 ( .A1(n4580), .A2(n4335), .ZN(n4707) );
  XNOR2_X1 U4891 ( .A(n5663), .B(n5666), .ZN(n8034) );
  NAND2_X2 U4892 ( .A1(n8031), .A2(n8030), .ZN(n9736) );
  INV_X1 U4893 ( .A(n9752), .ZN(n9501) );
  NAND2_X1 U4894 ( .A1(n5177), .A2(n5176), .ZN(n5663) );
  XNOR2_X1 U4895 ( .A(n5649), .B(n5648), .ZN(n9859) );
  NAND2_X2 U4896 ( .A1(n6266), .A2(n6265), .ZN(n9758) );
  NAND2_X1 U4897 ( .A1(n9665), .A2(n9797), .ZN(n9640) );
  CLKBUF_X1 U4898 ( .A(n8691), .Z(n4433) );
  CLKBUF_X1 U4899 ( .A(n7794), .Z(n4491) );
  NAND2_X1 U4900 ( .A1(n5624), .A2(n5625), .ZN(n5167) );
  NAND2_X1 U4901 ( .A1(n5585), .A2(n4513), .ZN(n7629) );
  AOI21_X1 U4902 ( .B1(n4914), .B2(n4916), .A(n4913), .ZN(n4912) );
  AOI21_X1 U4903 ( .B1(n7298), .B2(n6091), .A(n4367), .ZN(n9554) );
  XNOR2_X1 U4904 ( .A(n8842), .B(n8880), .ZN(n8991) );
  NAND2_X1 U4905 ( .A1(n5530), .A2(n5529), .ZN(n8698) );
  AND4_X2 U4906 ( .A1(n6300), .A2(n6299), .A3(n6298), .A4(n6297), .ZN(n9488)
         );
  OAI21_X1 U4907 ( .B1(n5571), .B2(n5570), .A(n5144), .ZN(n5587) );
  XNOR2_X1 U4908 ( .A(n5528), .B(n5527), .ZN(n7219) );
  NAND2_X1 U4909 ( .A1(n6232), .A2(n6231), .ZN(n9587) );
  NAND2_X1 U4910 ( .A1(n7438), .A2(n7439), .ZN(n7548) );
  NAND2_X1 U4911 ( .A1(n5518), .A2(n5517), .ZN(n8711) );
  NOR2_X1 U4912 ( .A1(n4857), .A2(n4856), .ZN(n4855) );
  NAND2_X2 U4913 ( .A1(n6218), .A2(n6217), .ZN(n9785) );
  NAND2_X1 U4914 ( .A1(n5453), .A2(n5452), .ZN(n8733) );
  AND2_X1 U4915 ( .A1(n5765), .A2(n5766), .ZN(n7864) );
  NAND2_X1 U4916 ( .A1(n4438), .A2(n6158), .ZN(n9814) );
  OR2_X1 U4917 ( .A1(n6886), .A2(n6887), .ZN(n6915) );
  NAND2_X1 U4918 ( .A1(n5417), .A2(n5416), .ZN(n8737) );
  NAND2_X1 U4919 ( .A1(n6343), .A2(n6342), .ZN(n7076) );
  NAND2_X1 U4920 ( .A1(n6149), .A2(n6148), .ZN(n9818) );
  NAND2_X1 U4921 ( .A1(n5490), .A2(n5489), .ZN(n8721) );
  XNOR2_X1 U4922 ( .A(n5447), .B(n5446), .ZN(n6479) );
  NAND2_X1 U4923 ( .A1(n5432), .A2(n5431), .ZN(n8743) );
  INV_X2 U4924 ( .A(n7106), .ZN(n4274) );
  XNOR2_X1 U4925 ( .A(n5368), .B(n5367), .ZN(n6452) );
  NAND2_X1 U4926 ( .A1(n5355), .A2(n5354), .ZN(n8627) );
  NAND2_X1 U4927 ( .A1(n7286), .A2(n9982), .ZN(n7285) );
  NOR2_X1 U4928 ( .A1(n9891), .A2(n10278), .ZN(n9892) );
  NAND2_X1 U4929 ( .A1(n6082), .A2(n6081), .ZN(n7414) );
  OR2_X1 U4930 ( .A1(n7561), .A2(n7423), .ZN(n9299) );
  CLKBUF_X1 U4931 ( .A(n5897), .Z(n7176) );
  INV_X1 U4932 ( .A(n7089), .ZN(n4520) );
  AND2_X1 U4933 ( .A1(n9202), .A2(n9291), .ZN(n9251) );
  CLKBUF_X1 U4934 ( .A(n7157), .Z(n4467) );
  NAND2_X1 U4935 ( .A1(n6055), .A2(n6054), .ZN(n7089) );
  NAND2_X1 U4936 ( .A1(n6069), .A2(n6068), .ZN(n7561) );
  INV_X1 U4937 ( .A(n6688), .ZN(n5891) );
  NAND2_X1 U4938 ( .A1(n6688), .A2(n7580), .ZN(n5890) );
  INV_X1 U4939 ( .A(n6993), .ZN(n6755) );
  INV_X1 U4940 ( .A(n7292), .ZN(n9982) );
  OR2_X2 U4941 ( .A1(n6484), .A2(P1_U3084), .ZN(n9336) );
  AND4_X1 U4942 ( .A1(n6116), .A2(n6115), .A3(n6114), .A4(n6113), .ZN(n7712)
         );
  INV_X1 U4943 ( .A(n5207), .ZN(n5699) );
  NAND2_X1 U4944 ( .A1(n6014), .A2(n4400), .ZN(n6993) );
  AND4_X1 U4945 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n7423)
         );
  NAND2_X1 U4946 ( .A1(n6051), .A2(n6052), .ZN(n7292) );
  OR2_X2 U4947 ( .A1(n7027), .A2(n8390), .ZN(n5839) );
  INV_X2 U4948 ( .A(n5321), .ZN(n5694) );
  NAND2_X1 U4949 ( .A1(n9884), .A2(n9885), .ZN(n9886) );
  BUF_X2 U4950 ( .A(n5283), .Z(n5207) );
  NAND4_X1 U4951 ( .A1(n6065), .A2(n6064), .A3(n6063), .A4(n6062), .ZN(n9352)
         );
  AND4_X1 U4952 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n7284)
         );
  OR2_X1 U4953 ( .A1(n5428), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5448) );
  NAND3_X1 U4954 ( .A1(n5262), .A2(n4471), .A3(n4470), .ZN(n8636) );
  OAI211_X1 U4955 ( .C1(n6439), .C2(n6035), .A(n4711), .B(n6024), .ZN(n7053)
         );
  NAND2_X2 U4956 ( .A1(n6396), .A2(n7876), .ZN(n6731) );
  NOR2_X2 U4957 ( .A1(n5986), .A2(n5987), .ZN(n6060) );
  NAND2_X1 U4958 ( .A1(n8791), .A2(n5206), .ZN(n7934) );
  NAND2_X1 U4959 ( .A1(n5544), .A2(n5543), .ZN(n8390) );
  NAND2_X1 U4960 ( .A1(n5998), .A2(n5997), .ZN(n6323) );
  OR2_X1 U4961 ( .A1(n5353), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U4962 ( .A1(n6308), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U4963 ( .A1(n4832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4831) );
  OR2_X1 U4964 ( .A1(n6395), .A2(n5993), .ZN(n4583) );
  NAND2_X1 U4965 ( .A1(n5082), .A2(n5081), .ZN(n5388) );
  NAND2_X1 U4966 ( .A1(n4460), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U4967 ( .A1(n5984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5983) );
  INV_X2 U4968 ( .A(n8795), .ZN(n4275) );
  NAND2_X1 U4969 ( .A1(n6388), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6395) );
  OAI21_X1 U4970 ( .B1(n5245), .B2(P1_DATAO_REG_10__SCAN_IN), .A(n4524), .ZN(
        n5082) );
  INV_X1 U4971 ( .A(n6084), .ZN(n4460) );
  NAND2_X2 U4972 ( .A1(n5245), .A2(P1_U3084), .ZN(n9866) );
  INV_X4 U4973 ( .A(n6005), .ZN(n4807) );
  INV_X1 U4974 ( .A(n6387), .ZN(n4595) );
  NAND2_X1 U4975 ( .A1(n4461), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6084) );
  NOR2_X1 U4976 ( .A1(n5980), .A2(n4695), .ZN(n4694) );
  INV_X1 U4977 ( .A(n6072), .ZN(n4461) );
  NAND3_X1 U4978 ( .A1(n5333), .A2(n5316), .A3(n4727), .ZN(n5483) );
  AND2_X1 U4979 ( .A1(n5975), .A2(n6168), .ZN(n6385) );
  INV_X1 U4980 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6587) );
  NOR2_X1 U4981 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5971) );
  NOR2_X1 U4982 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5972) );
  INV_X1 U4983 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5192) );
  INV_X1 U4984 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5409) );
  INV_X1 U4985 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4727) );
  NOR2_X1 U4986 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5977) );
  NOR2_X1 U4987 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5976) );
  NOR2_X1 U4988 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5181) );
  NOR2_X1 U4989 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5970) );
  CLKBUF_X1 U4990 ( .A(P1_IR_REG_8__SCAN_IN), .Z(n10238) );
  INV_X1 U4991 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6214) );
  NOR2_X1 U4992 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5183) );
  INV_X4 U4993 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4994 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5982) );
  INV_X2 U4995 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND2_X1 U4996 ( .A1(n8454), .A2(n5817), .ZN(n8434) );
  INV_X1 U4997 ( .A(n6800), .ZN(n9353) );
  NAND2_X1 U4998 ( .A1(n6800), .A2(n7292), .ZN(n9205) );
  AND2_X1 U4999 ( .A1(n8575), .A2(n8565), .ZN(n8561) );
  NOR2_X2 U5000 ( .A1(n5031), .A2(n8711), .ZN(n8575) );
  NAND2_X1 U5001 ( .A1(n7936), .A2(n5215), .ZN(n5674) );
  AND2_X2 U5002 ( .A1(n4898), .A2(n4899), .ZN(n9498) );
  INV_X1 U5004 ( .A(n5263), .ZN(n5294) );
  NOR2_X2 U5005 ( .A1(n10271), .A2(n9882), .ZN(n9883) );
  INV_X1 U5006 ( .A(n5207), .ZN(n4278) );
  AOI21_X1 U5007 ( .B1(n9132), .B2(n9221), .A(n4661), .ZN(n4660) );
  OR2_X1 U5008 ( .A1(n9814), .A2(n9098), .ZN(n9173) );
  NOR2_X1 U5009 ( .A1(n8417), .A2(n8017), .ZN(n4980) );
  OR2_X1 U5010 ( .A1(n9474), .A2(n9463), .ZN(n8032) );
  NOR2_X1 U5011 ( .A1(n9194), .A2(n4569), .ZN(n4568) );
  NAND2_X1 U5012 ( .A1(n4328), .A2(n4405), .ZN(n4567) );
  NAND2_X1 U5013 ( .A1(n9075), .A2(n4569), .ZN(n4691) );
  NAND2_X1 U5014 ( .A1(n5792), .A2(n5793), .ZN(n4751) );
  NOR2_X1 U5015 ( .A1(n9246), .A2(n4686), .ZN(n4685) );
  AND2_X1 U5016 ( .A1(n9138), .A2(n4330), .ZN(n4693) );
  OR2_X1 U5017 ( .A1(n5693), .A2(n5703), .ZN(n5838) );
  NOR2_X1 U5018 ( .A1(n5980), .A2(n4338), .ZN(n4640) );
  AND2_X1 U5019 ( .A1(n5105), .A2(n5446), .ZN(n5106) );
  AOI21_X1 U5020 ( .B1(n5104), .B2(n5406), .A(n5103), .ZN(n5105) );
  INV_X1 U5021 ( .A(n5444), .ZN(n5103) );
  INV_X1 U5022 ( .A(n5425), .ZN(n5099) );
  NAND2_X1 U5023 ( .A1(n4807), .A2(n6465), .ZN(n4524) );
  AND2_X1 U5024 ( .A1(n5080), .A2(n5075), .ZN(n4522) );
  INV_X1 U5025 ( .A(n5339), .ZN(n5080) );
  AND2_X1 U5027 ( .A1(n5614), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5628) );
  OR2_X1 U5028 ( .A1(n8701), .A2(n8536), .ZN(n8514) );
  AOI21_X1 U5029 ( .B1(n4839), .B2(n8595), .A(n4838), .ZN(n4837) );
  INV_X1 U5030 ( .A(n5788), .ZN(n4838) );
  OR2_X1 U5031 ( .A1(n5492), .A2(n5491), .ZN(n5508) );
  AND2_X1 U5032 ( .A1(n8608), .A2(n4285), .ZN(n4633) );
  OR2_X1 U5033 ( .A1(n8721), .A2(n8248), .ZN(n5778) );
  AOI21_X1 U5034 ( .B1(n4272), .B2(n7656), .A(n4332), .ZN(n5022) );
  NAND2_X1 U5035 ( .A1(n7535), .A2(n8636), .ZN(n7470) );
  NAND2_X1 U5036 ( .A1(n6935), .A2(n6936), .ZN(n7471) );
  OR2_X1 U5037 ( .A1(n7254), .A2(n7253), .ZN(n4713) );
  INV_X1 U5038 ( .A(n7675), .ZN(n4916) );
  AND2_X1 U5039 ( .A1(n8849), .A2(n4924), .ZN(n4923) );
  AND2_X1 U5040 ( .A1(n4281), .A2(n4314), .ZN(n4440) );
  OR3_X1 U5041 ( .A1(n9499), .A2(n9270), .A3(n9513), .ZN(n9271) );
  OAI21_X1 U5042 ( .B1(n9157), .B2(n4333), .A(n4579), .ZN(n4650) );
  NOR2_X1 U5043 ( .A1(n4652), .A2(n9163), .ZN(n4579) );
  NAND2_X1 U5044 ( .A1(n9443), .A2(n9337), .ZN(n9236) );
  OAI21_X1 U5045 ( .B1(n4884), .B2(n9273), .A(n4883), .ZN(n4882) );
  NAND2_X1 U5046 ( .A1(n9273), .A2(n9226), .ZN(n4883) );
  NOR2_X1 U5047 ( .A1(n5039), .A2(n4886), .ZN(n4884) );
  AND2_X1 U5048 ( .A1(n9742), .A2(n9500), .ZN(n9242) );
  OR2_X1 U5049 ( .A1(n9742), .A2(n9500), .ZN(n9315) );
  AOI21_X1 U5050 ( .B1(n4901), .B2(n4900), .A(n9148), .ZN(n4899) );
  OR2_X1 U5051 ( .A1(n6241), .A2(n4902), .ZN(n4898) );
  INV_X1 U5052 ( .A(n4905), .ZN(n4900) );
  OR2_X1 U5053 ( .A1(n9758), .A2(n9535), .ZN(n9218) );
  INV_X1 U5054 ( .A(n6370), .ZN(n4963) );
  NOR2_X1 U5055 ( .A1(n9566), .A2(n4966), .ZN(n4965) );
  INV_X1 U5056 ( .A(n4968), .ZN(n4966) );
  AND2_X1 U5057 ( .A1(n6117), .A2(n9087), .ZN(n9172) );
  OR2_X1 U5058 ( .A1(n6327), .A2(n7644), .ZN(n9087) );
  AND2_X1 U5059 ( .A1(n7314), .A2(n6348), .ZN(n6344) );
  AND2_X1 U5060 ( .A1(n4946), .A2(n4945), .ZN(n4944) );
  NOR2_X1 U5061 ( .A1(n9256), .A2(n6347), .ZN(n4945) );
  NAND2_X1 U5062 ( .A1(n6380), .A2(n6586), .ZN(n6710) );
  NOR2_X1 U5063 ( .A1(n6387), .A2(n5980), .ZN(n5999) );
  NAND2_X1 U5064 ( .A1(n4595), .A2(n4489), .ZN(n6000) );
  NOR2_X1 U5065 ( .A1(n5980), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4489) );
  AND2_X1 U5066 ( .A1(n5172), .A2(n5171), .ZN(n5638) );
  INV_X1 U5067 ( .A(n5527), .ZN(n5136) );
  XNOR2_X1 U5068 ( .A(n5122), .B(n10188), .ZN(n5498) );
  NAND2_X1 U5069 ( .A1(n5120), .A2(n5119), .ZN(n5499) );
  INV_X1 U5070 ( .A(n5352), .ZN(n5086) );
  AND2_X1 U5071 ( .A1(n8011), .A2(n8010), .ZN(n8059) );
  NAND2_X1 U5072 ( .A1(n4307), .A2(n4527), .ZN(n7996) );
  OR2_X1 U5073 ( .A1(n7994), .A2(n7995), .ZN(n4527) );
  AND2_X1 U5074 ( .A1(n4999), .A2(n8115), .ZN(n4998) );
  NAND2_X1 U5075 ( .A1(n5668), .A2(n5667), .ZN(n8417) );
  OR2_X1 U5076 ( .A1(n5641), .A2(n8065), .ZN(n5654) );
  CLKBUF_X1 U5077 ( .A(n5691), .Z(n4468) );
  AND2_X1 U5078 ( .A1(n8220), .A2(n8219), .ZN(n8457) );
  OR2_X1 U5079 ( .A1(n5602), .A2(n8155), .ZN(n5616) );
  AND2_X1 U5080 ( .A1(n8487), .A2(n4304), .ZN(n4851) );
  AOI21_X1 U5081 ( .B1(n8508), .B2(n4636), .A(n4345), .ZN(n5926) );
  OR2_X1 U5082 ( .A1(n8691), .A2(n8537), .ZN(n5802) );
  INV_X1 U5083 ( .A(n8246), .ZN(n8505) );
  NOR2_X1 U5084 ( .A1(n8533), .A2(n8534), .ZN(n8532) );
  NAND2_X1 U5085 ( .A1(n5028), .A2(n5027), .ZN(n7896) );
  AOI21_X1 U5086 ( .B1(n4280), .B2(n7864), .A(n4340), .ZN(n5027) );
  AND2_X1 U5087 ( .A1(n6473), .A2(n5940), .ZN(n8580) );
  NAND2_X2 U5088 ( .A1(n6650), .A2(n4410), .ZN(n5691) );
  NAND2_X1 U5089 ( .A1(n5542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4740) );
  AND2_X1 U5090 ( .A1(n4306), .A2(n4721), .ZN(n4720) );
  NAND2_X1 U5091 ( .A1(n4283), .A2(n4723), .ZN(n4721) );
  CLKBUF_X1 U5092 ( .A(n6060), .Z(n4448) );
  NAND2_X1 U5093 ( .A1(n4595), .A2(n4596), .ZN(n6397) );
  XNOR2_X1 U5094 ( .A(n9428), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U5095 ( .A1(n9925), .A2(n9427), .ZN(n9428) );
  XNOR2_X1 U5096 ( .A(n9434), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U5097 ( .A1(n9912), .A2(n9433), .ZN(n9434) );
  NOR2_X1 U5098 ( .A1(n9465), .A2(n9736), .ZN(n9468) );
  OR2_X1 U5099 ( .A1(n9742), .A2(n9339), .ZN(n6376) );
  OR2_X1 U5100 ( .A1(n9758), .A2(n9341), .ZN(n6374) );
  NAND2_X1 U5101 ( .A1(n6267), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6276) );
  BUF_X1 U5102 ( .A(n9066), .Z(n6286) );
  AND2_X2 U5103 ( .A1(n9592), .A2(n9201), .ZN(n6241) );
  AOI21_X1 U5104 ( .B1(n7794), .B2(n4955), .A(n4952), .ZN(n6359) );
  AND2_X1 U5105 ( .A1(n4353), .A2(n4282), .ZN(n4955) );
  INV_X1 U5106 ( .A(n4909), .ZN(n4908) );
  OAI21_X1 U5107 ( .B1(n4300), .B2(n4910), .A(n9173), .ZN(n4909) );
  NAND2_X1 U5108 ( .A1(n4911), .A2(n9195), .ZN(n4910) );
  NAND2_X1 U5109 ( .A1(n7333), .A2(n6353), .ZN(n7359) );
  NAND2_X1 U5110 ( .A1(n9056), .A2(n4410), .ZN(n6035) );
  NAND2_X2 U5111 ( .A1(n6323), .A2(n6613), .ZN(n9056) );
  INV_X1 U5112 ( .A(n9464), .ZN(n4399) );
  NAND2_X1 U5113 ( .A1(n9474), .A2(n9957), .ZN(n6329) );
  NAND2_X1 U5114 ( .A1(n5587), .A2(n5586), .ZN(n5585) );
  NAND2_X1 U5115 ( .A1(n6192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6204) );
  AND2_X1 U5116 ( .A1(n6156), .A2(n6147), .ZN(n9365) );
  NAND2_X1 U5117 ( .A1(n5597), .A2(n5596), .ZN(n8519) );
  OR2_X1 U5118 ( .A1(n8498), .A2(n5669), .ZN(n5597) );
  INV_X1 U5119 ( .A(n9340), .ZN(n9516) );
  AOI21_X1 U5120 ( .B1(n5763), .B2(n5850), .A(n4767), .ZN(n4766) );
  AOI21_X1 U5121 ( .B1(n4769), .B2(n7862), .A(n5839), .ZN(n4765) );
  INV_X1 U5122 ( .A(n7859), .ZN(n4769) );
  AOI21_X1 U5123 ( .B1(n4757), .B2(n4756), .A(n4755), .ZN(n5752) );
  NAND2_X1 U5124 ( .A1(n5750), .A2(n5751), .ZN(n4755) );
  INV_X1 U5125 ( .A(n4761), .ZN(n4759) );
  AOI21_X1 U5126 ( .B1(n4765), .B2(n7863), .A(n4762), .ZN(n4761) );
  NAND2_X1 U5127 ( .A1(n7864), .A2(n4763), .ZN(n4762) );
  NAND2_X1 U5128 ( .A1(n4766), .A2(n4764), .ZN(n4763) );
  NOR2_X1 U5129 ( .A1(n5768), .A2(n7885), .ZN(n4768) );
  NOR2_X1 U5130 ( .A1(n4690), .A2(n4689), .ZN(n4688) );
  INV_X1 U5131 ( .A(n9077), .ZN(n4689) );
  INV_X1 U5132 ( .A(n5791), .ZN(n4750) );
  OAI21_X1 U5133 ( .B1(n4663), .B2(n9115), .A(n4671), .ZN(n4673) );
  INV_X1 U5134 ( .A(n4672), .ZN(n4671) );
  NOR2_X1 U5135 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  AND2_X1 U5136 ( .A1(n8217), .A2(n8666), .ZN(n4560) );
  NAND2_X1 U5137 ( .A1(n4681), .A2(n4675), .ZN(n4674) );
  INV_X1 U5138 ( .A(n9189), .ZN(n4675) );
  INV_X1 U5139 ( .A(n4685), .ZN(n4680) );
  OR2_X1 U5140 ( .A1(n9122), .A2(n4684), .ZN(n4576) );
  OR2_X1 U5141 ( .A1(n9125), .A2(n4682), .ZN(n4575) );
  NOR2_X1 U5142 ( .A1(n9125), .A2(n4405), .ZN(n4644) );
  OAI21_X1 U5143 ( .B1(n9122), .B2(n4569), .A(n4676), .ZN(n4645) );
  INV_X1 U5144 ( .A(n4677), .ZN(n4676) );
  NOR4_X1 U5145 ( .A1(n8595), .A2(n5857), .A3(n8608), .A4(n5916), .ZN(n5858)
         );
  NAND2_X1 U5146 ( .A1(n4828), .A2(n4375), .ZN(n9240) );
  INV_X1 U5147 ( .A(n4564), .ZN(n4889) );
  NOR2_X1 U5148 ( .A1(n5665), .A2(SI_29_), .ZN(n4827) );
  NAND2_X1 U5149 ( .A1(n5665), .A2(SI_29_), .ZN(n4826) );
  NAND2_X1 U5150 ( .A1(n5096), .A2(n5095), .ZN(n5404) );
  NAND2_X1 U5151 ( .A1(n5077), .A2(n5076), .ZN(n5351) );
  OAI21_X1 U5152 ( .B1(n6005), .B2(n4485), .A(n4484), .ZN(n5293) );
  NAND2_X1 U5153 ( .A1(n6005), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4484) );
  AND2_X1 U5154 ( .A1(n4533), .A2(n7948), .ZN(n4532) );
  NAND2_X1 U5155 ( .A1(n5007), .A2(n4534), .ZN(n4533) );
  INV_X1 U5156 ( .A(n7909), .ZN(n4534) );
  INV_X1 U5157 ( .A(n5007), .ZN(n4535) );
  INV_X1 U5158 ( .A(n5508), .ZN(n5506) );
  NOR2_X1 U5159 ( .A1(n5519), .A2(n5507), .ZN(n4562) );
  NAND2_X1 U5160 ( .A1(n5838), .A2(n5833), .ZN(n5842) );
  NAND2_X1 U5161 ( .A1(n4395), .A2(n4319), .ZN(n4394) );
  NAND2_X1 U5162 ( .A1(n4729), .A2(n4728), .ZN(n4395) );
  OR2_X1 U5163 ( .A1(n8417), .A2(n7634), .ZN(n5831) );
  INV_X1 U5164 ( .A(n5562), .ZN(n5532) );
  NAND2_X1 U5165 ( .A1(n5418), .A2(n4295), .ZN(n5475) );
  OR2_X1 U5166 ( .A1(n8733), .A2(n8171), .ZN(n5769) );
  OR2_X1 U5167 ( .A1(n8737), .A2(n8071), .ZN(n5765) );
  OR2_X1 U5168 ( .A1(n7774), .A2(n7816), .ZN(n5756) );
  NAND2_X1 U5169 ( .A1(n5933), .A2(n7373), .ZN(n5939) );
  INV_X1 U5170 ( .A(n10030), .ZN(n5958) );
  NOR2_X1 U5171 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5011) );
  AND2_X1 U5172 ( .A1(n8857), .A2(n8856), .ZN(n8859) );
  OR2_X1 U5173 ( .A1(n9554), .A2(n8892), .ZN(n8857) );
  NOR2_X1 U5174 ( .A1(n4373), .A2(n6725), .ZN(n6797) );
  AND2_X1 U5175 ( .A1(n9235), .A2(n9228), .ZN(n4692) );
  AOI21_X1 U5176 ( .B1(n9378), .B2(n4486), .A(n9377), .ZN(n9394) );
  INV_X1 U5177 ( .A(n9541), .ZN(n9544) );
  NAND2_X1 U5178 ( .A1(n6241), .A2(n9121), .ZN(n4906) );
  OR2_X1 U5179 ( .A1(n6240), .A2(n9246), .ZN(n9576) );
  OR2_X1 U5180 ( .A1(n9624), .A2(n9632), .ZN(n9120) );
  OR2_X1 U5181 ( .A1(n9807), .A2(n9655), .ZN(n9181) );
  NAND2_X1 U5182 ( .A1(n4502), .A2(n4327), .ZN(n4501) );
  INV_X1 U5183 ( .A(n4871), .ZN(n4869) );
  OR2_X1 U5184 ( .A1(n9824), .A2(n7666), .ZN(n9112) );
  AND2_X1 U5185 ( .A1(n9081), .A2(n9078), .ZN(n9192) );
  NOR2_X1 U5186 ( .A1(n7336), .A2(n6327), .ZN(n4502) );
  AND2_X1 U5187 ( .A1(n9077), .A2(n9070), .ZN(n9194) );
  NOR2_X1 U5188 ( .A1(n9351), .A2(n7561), .ZN(n6347) );
  OR2_X1 U5189 ( .A1(n7414), .A2(n7570), .ZN(n9076) );
  AND2_X1 U5190 ( .A1(n9207), .A2(n4894), .ZN(n4887) );
  NOR2_X1 U5191 ( .A1(n7062), .A2(n4893), .ZN(n4476) );
  NAND2_X1 U5192 ( .A1(n9206), .A2(n9205), .ZN(n4893) );
  NAND2_X1 U5193 ( .A1(n6058), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U5194 ( .A1(n4889), .A2(n9205), .ZN(n4888) );
  NAND2_X1 U5195 ( .A1(n4520), .A2(n9352), .ZN(n4894) );
  NAND2_X1 U5196 ( .A1(n7568), .A2(n7089), .ZN(n9206) );
  NAND2_X1 U5197 ( .A1(n4564), .A2(n9295), .ZN(n7062) );
  NAND2_X1 U5198 ( .A1(n6339), .A2(n7053), .ZN(n9291) );
  NOR2_X1 U5199 ( .A1(n5988), .A2(n4669), .ZN(n4668) );
  NAND2_X1 U5200 ( .A1(n9956), .A2(n7092), .ZN(n4462) );
  OAI21_X1 U5201 ( .B1(n5663), .B2(n4827), .A(n4826), .ZN(n5680) );
  AND2_X1 U5202 ( .A1(n4809), .A2(n4814), .ZN(n4808) );
  AOI21_X1 U5203 ( .B1(n4816), .B2(n5154), .A(n4815), .ZN(n4814) );
  AND2_X1 U5204 ( .A1(n5166), .A2(n5165), .ZN(n5625) );
  NAND2_X1 U5205 ( .A1(n5585), .A2(n5150), .ZN(n5598) );
  AND2_X1 U5206 ( .A1(n5135), .A2(n5134), .ZN(n5555) );
  INV_X1 U5207 ( .A(n4821), .ZN(n4820) );
  AOI21_X1 U5208 ( .B1(n4821), .B2(n4819), .A(n4337), .ZN(n4818) );
  AND2_X1 U5209 ( .A1(n4822), .A2(n5124), .ZN(n4821) );
  NAND2_X1 U5210 ( .A1(n5130), .A2(n5129), .ZN(n5540) );
  XNOR2_X1 U5211 ( .A(n5125), .B(SI_18_), .ZN(n5513) );
  AOI21_X1 U5212 ( .B1(n5106), .B2(n4806), .A(n4342), .ZN(n4803) );
  NAND2_X1 U5213 ( .A1(n5113), .A2(n5112), .ZN(n5466) );
  XNOR2_X1 U5214 ( .A(n5107), .B(SI_14_), .ZN(n5446) );
  XNOR2_X1 U5215 ( .A(n5092), .B(SI_11_), .ZN(n5390) );
  NAND2_X1 U5216 ( .A1(n5388), .A2(n5084), .ZN(n5366) );
  NAND2_X1 U5217 ( .A1(n5292), .A2(n5291), .ZN(n5310) );
  NOR2_X1 U5218 ( .A1(n8168), .A2(n5008), .ZN(n5007) );
  INV_X1 U5219 ( .A(n7941), .ZN(n5008) );
  NAND2_X1 U5220 ( .A1(n5002), .A2(n5001), .ZN(n7993) );
  NAND2_X1 U5221 ( .A1(n5004), .A2(n4323), .ZN(n5001) );
  NAND2_X1 U5222 ( .A1(n8091), .A2(n5000), .ZN(n5002) );
  AOI21_X1 U5223 ( .B1(n4542), .B2(n4545), .A(n4541), .ZN(n4540) );
  INV_X1 U5224 ( .A(n7732), .ZN(n4541) );
  NOR2_X1 U5225 ( .A1(n4547), .A2(n7459), .ZN(n4543) );
  AND2_X1 U5226 ( .A1(n4548), .A2(n7592), .ZN(n4547) );
  NAND2_X1 U5227 ( .A1(n7451), .A2(n7455), .ZN(n4548) );
  OR2_X1 U5228 ( .A1(n8148), .A2(n8151), .ZN(n5033) );
  AND2_X1 U5229 ( .A1(n7119), .A2(n8390), .ZN(n7017) );
  NAND2_X1 U5230 ( .A1(n5418), .A2(n4561), .ZN(n5455) );
  NAND2_X1 U5231 ( .A1(n5573), .A2(n5572), .ZN(n8691) );
  NAND2_X1 U5232 ( .A1(n7035), .A2(n7033), .ZN(n4985) );
  AND2_X1 U5233 ( .A1(n7970), .A2(n7969), .ZN(n8196) );
  NOR2_X1 U5234 ( .A1(n4553), .A2(n5030), .ZN(n4552) );
  INV_X1 U5235 ( .A(n7182), .ZN(n4553) );
  NOR2_X1 U5236 ( .A1(n7039), .A2(n7016), .ZN(n7026) );
  INV_X1 U5237 ( .A(n7027), .ZN(n4504) );
  OAI21_X1 U5238 ( .B1(n8434), .B2(n4846), .A(n4844), .ZN(n8411) );
  INV_X1 U5239 ( .A(n4848), .ZN(n4846) );
  AND2_X1 U5240 ( .A1(n4847), .A2(n4845), .ZN(n4844) );
  NAND2_X1 U5241 ( .A1(n4848), .A2(n8435), .ZN(n4845) );
  NAND2_X1 U5242 ( .A1(n5813), .A2(n5814), .ZN(n8468) );
  INV_X1 U5243 ( .A(n8468), .ZN(n8465) );
  OR2_X1 U5244 ( .A1(n5926), .A2(n5020), .ZN(n8461) );
  NAND2_X1 U5245 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  AND2_X1 U5246 ( .A1(n5923), .A2(n5581), .ZN(n5582) );
  NOR2_X1 U5247 ( .A1(n8525), .A2(n4433), .ZN(n8509) );
  NAND2_X1 U5248 ( .A1(n5922), .A2(n5921), .ZN(n8508) );
  OR2_X1 U5249 ( .A1(n8698), .A2(n8543), .ZN(n5920) );
  NAND2_X1 U5250 ( .A1(n5532), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5574) );
  AOI21_X1 U5251 ( .B1(n8510), .B2(n5622), .A(n5579), .ZN(n8537) );
  AND2_X1 U5252 ( .A1(n5568), .A2(n5567), .ZN(n8536) );
  NAND2_X1 U5253 ( .A1(n4842), .A2(n4843), .ZN(n4841) );
  INV_X1 U5254 ( .A(n4425), .ZN(n4842) );
  INV_X1 U5255 ( .A(n4633), .ZN(n4632) );
  NAND2_X1 U5256 ( .A1(n4633), .A2(n4631), .ZN(n4630) );
  AND2_X1 U5257 ( .A1(n8595), .A2(n4303), .ZN(n5021) );
  NAND2_X1 U5258 ( .A1(n4634), .A2(n4633), .ZN(n8607) );
  OAI211_X1 U5259 ( .C1(n4621), .C2(n4622), .A(n4619), .B(n5913), .ZN(n7855)
         );
  OR2_X1 U5260 ( .A1(n7855), .A2(n7864), .ZN(n5029) );
  OR2_X1 U5261 ( .A1(n7819), .A2(n7919), .ZN(n7839) );
  OR2_X1 U5262 ( .A1(n5345), .A2(n5344), .ZN(n5356) );
  CLKBUF_X1 U5263 ( .A(n7649), .Z(n7691) );
  NAND2_X1 U5264 ( .A1(n7548), .A2(n4435), .ZN(n4854) );
  NOR2_X1 U5265 ( .A1(n5905), .A2(n5338), .ZN(n4435) );
  NAND2_X1 U5266 ( .A1(n10061), .A2(n8256), .ZN(n5747) );
  INV_X1 U5267 ( .A(n5903), .ZN(n4616) );
  NAND2_X1 U5268 ( .A1(n5281), .A2(n7471), .ZN(n4850) );
  NOR2_X1 U5269 ( .A1(n7528), .A2(n8636), .ZN(n7477) );
  OR2_X1 U5270 ( .A1(n7024), .A2(n5940), .ZN(n8605) );
  INV_X1 U5271 ( .A(n8580), .ZN(n8603) );
  OR2_X1 U5272 ( .A1(n10033), .A2(n5961), .ZN(n6692) );
  NAND2_X1 U5273 ( .A1(n8416), .A2(n8417), .ZN(n4981) );
  INV_X1 U5274 ( .A(n7558), .ZN(n10061) );
  OR2_X1 U5275 ( .A1(n7018), .A2(n5944), .ZN(n10052) );
  NOR2_X1 U5276 ( .A1(n10052), .A2(n8390), .ZN(n7037) );
  NAND2_X1 U5277 ( .A1(n7268), .A2(n7299), .ZN(n7018) );
  AND2_X1 U5279 ( .A1(n7042), .A2(n10037), .ZN(n10031) );
  INV_X1 U5280 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U5281 ( .A1(n5870), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U5282 ( .A1(n5212), .A2(n5011), .ZN(n5543) );
  NAND2_X1 U5283 ( .A1(n5212), .A2(n5211), .ZN(n5542) );
  INV_X1 U5284 ( .A(n7823), .ZN(n4593) );
  OAI22_X1 U5285 ( .A1(n8832), .A2(n6339), .B1(n4860), .B2(n6725), .ZN(n6726)
         );
  AND2_X1 U5286 ( .A1(n8900), .A2(n4341), .ZN(n4611) );
  NOR2_X1 U5287 ( .A1(n8848), .A2(n5041), .ZN(n8849) );
  NAND2_X1 U5288 ( .A1(n4710), .A2(n8876), .ZN(n8951) );
  NAND2_X1 U5289 ( .A1(n4582), .A2(n7092), .ZN(n6592) );
  AND2_X1 U5290 ( .A1(n9597), .A2(n8883), .ZN(n4581) );
  NAND2_X1 U5291 ( .A1(n6560), .A2(n4322), .ZN(n6606) );
  AND2_X1 U5292 ( .A1(n6767), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4772) );
  NOR2_X1 U5293 ( .A1(n7276), .A2(n7277), .ZN(n7386) );
  OR2_X1 U5294 ( .A1(n7386), .A2(n4784), .ZN(n4783) );
  AND2_X1 U5295 ( .A1(n7387), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U5296 ( .A1(n4783), .A2(n4782), .ZN(n4488) );
  INV_X1 U5297 ( .A(n7388), .ZN(n4782) );
  XNOR2_X1 U5298 ( .A(n9394), .B(n9393), .ZN(n9380) );
  NOR2_X1 U5299 ( .A1(n9394), .A2(n9393), .ZN(n9396) );
  NAND2_X1 U5300 ( .A1(n4882), .A2(n4885), .ZN(n4881) );
  OR2_X1 U5301 ( .A1(n9273), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U5302 ( .A1(n9243), .A2(n9315), .ZN(n9485) );
  INV_X1 U5303 ( .A(n9758), .ZN(n9517) );
  INV_X1 U5304 ( .A(n9216), .ZN(n4572) );
  INV_X1 U5305 ( .A(n9560), .ZN(n9534) );
  NAND2_X1 U5306 ( .A1(n4903), .A2(n4904), .ZN(n9532) );
  NAND2_X1 U5307 ( .A1(n6241), .A2(n4905), .ZN(n4903) );
  NOR2_X1 U5308 ( .A1(n9768), .A2(n4875), .ZN(n4381) );
  AOI21_X1 U5309 ( .B1(n4965), .B2(n6369), .A(n4301), .ZN(n4964) );
  OR2_X1 U5310 ( .A1(n9244), .A2(n4406), .ZN(n9541) );
  OR2_X1 U5311 ( .A1(n9587), .A2(n9598), .ZN(n4968) );
  OR2_X1 U5312 ( .A1(n9583), .A2(n6369), .ZN(n4967) );
  CLKBUF_X1 U5313 ( .A(n4965), .Z(n4388) );
  CLKBUF_X1 U5314 ( .A(n9581), .Z(n9583) );
  AOI21_X1 U5315 ( .B1(n4949), .B2(n6362), .A(n4288), .ZN(n4948) );
  AND2_X1 U5316 ( .A1(n9124), .A2(n9201), .ZN(n9607) );
  NAND2_X1 U5317 ( .A1(n9624), .A2(n9632), .ZN(n9594) );
  NAND2_X1 U5318 ( .A1(n6195), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6222) );
  NOR2_X1 U5319 ( .A1(n9618), .A2(n4950), .ZN(n4949) );
  INV_X1 U5320 ( .A(n6365), .ZN(n4950) );
  NAND2_X1 U5321 ( .A1(n6364), .A2(n6363), .ZN(n4951) );
  AND2_X1 U5322 ( .A1(n9120), .A2(n9594), .ZN(n9618) );
  AND2_X1 U5323 ( .A1(n4443), .A2(n4442), .ZN(n9665) );
  NAND2_X1 U5324 ( .A1(n4958), .A2(n4282), .ZN(n4956) );
  AND2_X1 U5325 ( .A1(n9181), .A2(n9178), .ZN(n9684) );
  NAND2_X1 U5326 ( .A1(n7603), .A2(n4300), .ZN(n7786) );
  NOR2_X1 U5327 ( .A1(n7361), .A2(n7681), .ZN(n4877) );
  NAND2_X1 U5328 ( .A1(n7244), .A2(n7248), .ZN(n7336) );
  AND2_X1 U5329 ( .A1(n7334), .A2(n6351), .ZN(n6352) );
  INV_X1 U5330 ( .A(n6347), .ZN(n4943) );
  NAND2_X1 U5331 ( .A1(n4944), .A2(n4941), .ZN(n7242) );
  AND2_X1 U5332 ( .A1(n9076), .A2(n9077), .ZN(n9256) );
  INV_X1 U5333 ( .A(n7062), .ZN(n4897) );
  NAND2_X1 U5334 ( .A1(n7050), .A2(n4860), .ZN(n7069) );
  NAND2_X1 U5335 ( .A1(n9859), .A2(n6091), .ZN(n8031) );
  INV_X1 U5336 ( .A(n9479), .ZN(n6330) );
  NOR2_X1 U5337 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  AND2_X1 U5338 ( .A1(n9742), .A2(n9957), .ZN(n9743) );
  AND2_X1 U5339 ( .A1(n9689), .A2(n9811), .ZN(n9961) );
  AND2_X1 U5340 ( .A1(n7301), .A2(n9165), .ZN(n6984) );
  AND2_X1 U5341 ( .A1(n6731), .A2(n6400), .ZN(n6577) );
  AND2_X1 U5342 ( .A1(n5978), .A2(n5979), .ZN(n4641) );
  NAND2_X1 U5343 ( .A1(n4415), .A2(n4414), .ZN(n5985) );
  NAND2_X1 U5344 ( .A1(n4417), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4414) );
  AOI21_X1 U5345 ( .B1(n5638), .B2(n4801), .A(n4800), .ZN(n4799) );
  INV_X1 U5346 ( .A(n5172), .ZN(n4800) );
  INV_X1 U5347 ( .A(n5166), .ZN(n4801) );
  INV_X1 U5348 ( .A(n5638), .ZN(n4802) );
  CLKBUF_X1 U5349 ( .A(n6323), .Z(n6729) );
  XNOR2_X1 U5350 ( .A(n5611), .B(n5610), .ZN(n7798) );
  OAI21_X1 U5351 ( .B1(n5598), .B2(n5154), .A(n5153), .ZN(n5611) );
  XNOR2_X1 U5352 ( .A(n5598), .B(n5599), .ZN(n7757) );
  AND2_X1 U5353 ( .A1(n5150), .A2(n5149), .ZN(n5586) );
  AND2_X1 U5354 ( .A1(n6312), .A2(n6582), .ZN(n9284) );
  XNOR2_X1 U5355 ( .A(n6023), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U5356 ( .A1(n9888), .A2(n9889), .ZN(n9890) );
  NAND2_X1 U5357 ( .A1(n7305), .A2(n7304), .ZN(n7452) );
  OAI21_X1 U5358 ( .B1(n4991), .B2(n4990), .A(n4994), .ZN(n8062) );
  INV_X1 U5359 ( .A(n4995), .ZN(n4994) );
  NAND2_X1 U5360 ( .A1(n7996), .A2(n4992), .ZN(n4991) );
  AND2_X1 U5361 ( .A1(n5654), .A2(n5642), .ZN(n8431) );
  INV_X1 U5362 ( .A(n7992), .ZN(n7988) );
  NAND2_X2 U5363 ( .A1(n5589), .A2(n5588), .ZN(n8688) );
  NAND2_X1 U5364 ( .A1(n7910), .A2(n7909), .ZN(n7942) );
  AOI21_X1 U5365 ( .B1(n7167), .B2(n7166), .A(n7165), .ZN(n7183) );
  OR2_X1 U5366 ( .A1(n5263), .A2(n6446), .ZN(n5248) );
  AND3_X1 U5367 ( .A1(n5512), .A2(n5511), .A3(n5510), .ZN(n8606) );
  AND2_X1 U5368 ( .A1(n5554), .A2(n5553), .ZN(n8203) );
  AND4_X1 U5369 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n7653)
         );
  AOI21_X1 U5370 ( .B1(n8475), .B2(n5647), .A(n5621), .ZN(n8218) );
  NAND2_X1 U5371 ( .A1(n5609), .A2(n5608), .ZN(n8246) );
  AND3_X1 U5372 ( .A1(n5497), .A2(n5496), .A3(n5495), .ZN(n8248) );
  AND2_X1 U5373 ( .A1(n6660), .A2(n6659), .ZN(n8388) );
  INV_X1 U5374 ( .A(n8383), .ZN(n8386) );
  AOI21_X1 U5375 ( .B1(n8520), .B2(n8614), .A(n4444), .ZN(n8694) );
  NAND2_X1 U5376 ( .A1(n4446), .A2(n4445), .ZN(n4444) );
  NAND2_X1 U5377 ( .A1(n8543), .A2(n8580), .ZN(n4445) );
  AND2_X1 U5378 ( .A1(n10031), .A2(n7037), .ZN(n8641) );
  INV_X1 U5379 ( .A(n8630), .ZN(n8643) );
  NAND2_X1 U5380 ( .A1(n8799), .A2(n6091), .ZN(n6294) );
  AND4_X1 U5381 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n9095)
         );
  AND2_X1 U5382 ( .A1(n6273), .A2(n6272), .ZN(n9535) );
  NAND2_X1 U5383 ( .A1(n7629), .A2(n6091), .ZN(n6256) );
  NAND2_X1 U5384 ( .A1(n8952), .A2(n4935), .ZN(n4934) );
  NAND2_X1 U5385 ( .A1(n4718), .A2(n4717), .ZN(n4716) );
  INV_X1 U5386 ( .A(n8937), .ZN(n4718) );
  NOR2_X1 U5387 ( .A1(n8936), .A2(n9024), .ZN(n4717) );
  NOR2_X1 U5388 ( .A1(n4719), .A2(n4607), .ZN(n4606) );
  INV_X1 U5389 ( .A(n4611), .ZN(n4607) );
  NAND2_X1 U5390 ( .A1(n6194), .A2(n6193), .ZN(n9642) );
  AND2_X1 U5391 ( .A1(n6229), .A2(n6228), .ZN(n9615) );
  AND2_X1 U5392 ( .A1(n6264), .A2(n6263), .ZN(n9548) );
  INV_X1 U5393 ( .A(n9554), .ZN(n9768) );
  INV_X1 U5394 ( .A(n9043), .ZN(n9024) );
  OR2_X1 U5395 ( .A1(n4653), .A2(n4649), .ZN(n4495) );
  INV_X1 U5396 ( .A(n9335), .ZN(n4404) );
  NAND4_X2 U5397 ( .A1(n8041), .A2(n8040), .A3(n8039), .A4(n8038), .ZN(n9462)
         );
  NAND2_X1 U5398 ( .A1(n6285), .A2(n6284), .ZN(n9340) );
  OR2_X1 U5399 ( .A1(n9505), .A2(n6278), .ZN(n6285) );
  INV_X1 U5400 ( .A(n9562), .ZN(n9598) );
  INV_X1 U5401 ( .A(n9657), .ZN(n9345) );
  INV_X1 U5402 ( .A(n9095), .ZN(n9706) );
  AND2_X1 U5403 ( .A1(n9375), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9388) );
  INV_X1 U5404 ( .A(n4781), .ZN(n4780) );
  OAI21_X1 U5405 ( .B1(n9436), .B2(n9923), .A(n9918), .ZN(n4781) );
  OAI22_X1 U5406 ( .A1(n9439), .A2(n9438), .B1(n9923), .B2(n9437), .ZN(n4778)
         );
  NOR2_X1 U5407 ( .A1(n9442), .A2(n9898), .ZN(n4776) );
  CLKBUF_X1 U5408 ( .A(n8033), .Z(n6378) );
  CLKBUF_X1 U5409 ( .A(n9661), .Z(n9662) );
  INV_X1 U5410 ( .A(n4401), .ZN(n4400) );
  OAI21_X1 U5411 ( .B1(n6035), .B2(n6446), .A(n6013), .ZN(n4401) );
  NOR2_X1 U5412 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  INV_X2 U5413 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9898) );
  NOR2_X1 U5414 ( .A1(n4849), .A2(n5730), .ZN(n5733) );
  NAND2_X1 U5415 ( .A1(n4753), .A2(n4752), .ZN(n4757) );
  AND2_X1 U5416 ( .A1(n4312), .A2(n7549), .ZN(n4752) );
  AND2_X1 U5417 ( .A1(n5748), .A2(n7656), .ZN(n4756) );
  INV_X1 U5418 ( .A(n5850), .ZN(n4764) );
  NAND2_X1 U5419 ( .A1(n4768), .A2(n4315), .ZN(n4760) );
  NAND2_X1 U5420 ( .A1(n4759), .A2(n4768), .ZN(n4758) );
  INV_X1 U5421 ( .A(n4568), .ZN(n4566) );
  OAI21_X1 U5422 ( .B1(n9110), .B2(n9094), .A(n9093), .ZN(n4666) );
  NOR2_X1 U5423 ( .A1(n9650), .A2(n4665), .ZN(n4664) );
  OAI21_X1 U5424 ( .B1(n9650), .B2(n9114), .A(n9116), .ZN(n4672) );
  NOR2_X1 U5425 ( .A1(n4747), .A2(n4751), .ZN(n4744) );
  NOR2_X1 U5426 ( .A1(n4749), .A2(n4748), .ZN(n4747) );
  NOR2_X1 U5427 ( .A1(n5791), .A2(n5797), .ZN(n4748) );
  INV_X1 U5428 ( .A(n5790), .ZN(n4749) );
  INV_X1 U5429 ( .A(n5802), .ZN(n4743) );
  NOR2_X1 U5430 ( .A1(n4751), .A2(n4746), .ZN(n4745) );
  NAND2_X1 U5431 ( .A1(n4750), .A2(n5788), .ZN(n4746) );
  OAI21_X1 U5432 ( .B1(n5810), .B2(n5809), .A(n5808), .ZN(n4432) );
  OAI22_X1 U5433 ( .A1(n4685), .A2(n4569), .B1(n9189), .B2(n4405), .ZN(n4677)
         );
  AOI21_X1 U5434 ( .B1(n4683), .B2(n4680), .A(n4679), .ZN(n4678) );
  AND2_X1 U5435 ( .A1(n4674), .A2(n9217), .ZN(n4387) );
  AND2_X1 U5436 ( .A1(n9281), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U5437 ( .A1(n9128), .A2(n4572), .ZN(n4571) );
  OAI21_X1 U5438 ( .B1(n9311), .B2(n9339), .A(n9494), .ZN(n9150) );
  INV_X1 U5439 ( .A(n9202), .ZN(n4563) );
  AOI21_X1 U5440 ( .B1(n4643), .B2(n9142), .A(n9127), .ZN(n4642) );
  NAND2_X1 U5441 ( .A1(n9134), .A2(n4662), .ZN(n4661) );
  AND2_X1 U5442 ( .A1(n9457), .A2(n9160), .ZN(n4662) );
  INV_X1 U5443 ( .A(n4894), .ZN(n9203) );
  INV_X1 U5444 ( .A(n5150), .ZN(n4813) );
  NOR2_X1 U5445 ( .A1(n4732), .A2(n4731), .ZN(n4730) );
  INV_X1 U5446 ( .A(n5832), .ZN(n4732) );
  INV_X1 U5447 ( .A(n5773), .ZN(n4856) );
  INV_X1 U5448 ( .A(n5285), .ZN(n4558) );
  NAND2_X1 U5449 ( .A1(n4920), .A2(n8859), .ZN(n4919) );
  AOI21_X1 U5450 ( .B1(n4923), .B2(n4922), .A(n8940), .ZN(n4921) );
  INV_X1 U5451 ( .A(n4306), .ZN(n4922) );
  NAND2_X1 U5452 ( .A1(n4923), .A2(n8859), .ZN(n4918) );
  OAI21_X1 U5453 ( .B1(n8959), .B2(n4335), .A(n4437), .ZN(n4436) );
  NOR2_X1 U5454 ( .A1(n8824), .A2(n8974), .ZN(n4437) );
  NAND2_X1 U5455 ( .A1(n4938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4937) );
  INV_X1 U5456 ( .A(n9235), .ZN(n4652) );
  OR2_X1 U5457 ( .A1(n9228), .A2(n9227), .ZN(n9167) );
  AND2_X1 U5458 ( .A1(n9217), .A2(n9545), .ZN(n9126) );
  NOR2_X1 U5459 ( .A1(n4499), .A2(n4406), .ZN(n4498) );
  NOR2_X1 U5460 ( .A1(n9244), .A2(n9142), .ZN(n4499) );
  AOI21_X1 U5461 ( .B1(n4799), .B2(n4802), .A(n4797), .ZN(n4796) );
  INV_X1 U5462 ( .A(n5648), .ZN(n4797) );
  NOR2_X1 U5463 ( .A1(n5610), .A2(n4817), .ZN(n4816) );
  INV_X1 U5464 ( .A(n5153), .ZN(n4817) );
  INV_X1 U5465 ( .A(n5160), .ZN(n4815) );
  INV_X1 U5466 ( .A(n4812), .ZN(n4811) );
  OAI21_X1 U5467 ( .B1(n5586), .B2(n4813), .A(n4816), .ZN(n4812) );
  NAND2_X1 U5468 ( .A1(n4811), .A2(n4813), .ZN(n4809) );
  NAND2_X1 U5469 ( .A1(n5121), .A2(n5123), .ZN(n4822) );
  INV_X1 U5470 ( .A(n5123), .ZN(n4819) );
  NAND2_X1 U5471 ( .A1(n5099), .A2(n5406), .ZN(n4806) );
  NAND2_X1 U5472 ( .A1(n5110), .A2(n5109), .ZN(n5113) );
  NAND2_X1 U5473 ( .A1(n5245), .A2(n6463), .ZN(n4519) );
  INV_X1 U5474 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n4493) );
  OAI21_X1 U5475 ( .B1(n5245), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n4523), .ZN(
        n5077) );
  NAND2_X1 U5476 ( .A1(n4807), .A2(n6449), .ZN(n4523) );
  AND2_X1 U5477 ( .A1(n5311), .A2(n5291), .ZN(n4512) );
  OAI21_X1 U5478 ( .B1(n5067), .B2(n4515), .A(n4514), .ZN(n5066) );
  NAND2_X1 U5479 ( .A1(n5067), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4514) );
  INV_X1 U5480 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4793) );
  NAND2_X1 U5481 ( .A1(n4997), .A2(n8005), .ZN(n4996) );
  AND2_X1 U5482 ( .A1(n5003), .A2(n7975), .ZN(n5000) );
  AND2_X1 U5483 ( .A1(n5004), .A2(n5005), .ZN(n5003) );
  AOI21_X1 U5484 ( .B1(n4532), .B2(n4535), .A(n4531), .ZN(n4530) );
  INV_X1 U5485 ( .A(n7953), .ZN(n4531) );
  INV_X1 U5486 ( .A(n8163), .ZN(n5005) );
  NOR2_X1 U5487 ( .A1(n6968), .A2(n5433), .ZN(n4561) );
  AND2_X1 U5488 ( .A1(n5397), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5418) );
  INV_X1 U5489 ( .A(n5398), .ZN(n5397) );
  INV_X1 U5490 ( .A(n8211), .ZN(n4999) );
  NAND2_X1 U5491 ( .A1(n5506), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U5492 ( .A1(n5506), .A2(n4562), .ZN(n5548) );
  AND2_X1 U5493 ( .A1(n5826), .A2(n5824), .ZN(n4848) );
  NAND2_X1 U5494 ( .A1(n5936), .A2(n5826), .ZN(n4847) );
  NAND2_X1 U5495 ( .A1(n5927), .A2(n8487), .ZN(n5019) );
  NAND2_X1 U5496 ( .A1(n5817), .A2(n5818), .ZN(n5928) );
  OR2_X1 U5497 ( .A1(n8678), .A2(n8218), .ZN(n5813) );
  INV_X1 U5498 ( .A(n8519), .ZN(n5924) );
  NAND2_X1 U5499 ( .A1(n4976), .A2(n8486), .ZN(n4975) );
  INV_X1 U5500 ( .A(n5036), .ZN(n4635) );
  NOR2_X1 U5501 ( .A1(n8190), .A2(n5533), .ZN(n4559) );
  NOR2_X1 U5502 ( .A1(n8688), .A2(n4433), .ZN(n4976) );
  AND2_X1 U5503 ( .A1(n5569), .A2(n4835), .ZN(n4834) );
  NAND2_X1 U5504 ( .A1(n4837), .A2(n4840), .ZN(n4835) );
  INV_X1 U5505 ( .A(n4837), .ZN(n4836) );
  NOR2_X1 U5506 ( .A1(n8502), .A2(n4638), .ZN(n4636) );
  AND2_X1 U5507 ( .A1(n5802), .A2(n5793), .ZN(n5923) );
  NAND2_X1 U5508 ( .A1(n5473), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5492) );
  INV_X1 U5509 ( .A(n5475), .ZN(n5473) );
  OR2_X1 U5510 ( .A1(n8728), .A2(n8604), .ZN(n5773) );
  AND2_X1 U5511 ( .A1(n5765), .A2(n7859), .ZN(n5441) );
  OR2_X1 U5512 ( .A1(n5914), .A2(n4618), .ZN(n4621) );
  INV_X1 U5513 ( .A(n4625), .ZN(n4618) );
  INV_X1 U5514 ( .A(n4621), .ZN(n4617) );
  NAND2_X1 U5515 ( .A1(n7774), .A2(n4626), .ZN(n4625) );
  NOR2_X1 U5516 ( .A1(n4978), .A2(n7774), .ZN(n4977) );
  NOR2_X1 U5517 ( .A1(n8627), .A2(n7658), .ZN(n4979) );
  INV_X1 U5518 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U5519 ( .A1(n4558), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U5520 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5285) );
  AND2_X2 U5521 ( .A1(n5738), .A2(n5737), .ZN(n5894) );
  NAND2_X1 U5522 ( .A1(n5237), .A2(n7434), .ZN(n6777) );
  NOR2_X1 U5523 ( .A1(n5197), .A2(n5025), .ZN(n5023) );
  NAND2_X1 U5524 ( .A1(n5198), .A2(n5196), .ZN(n5025) );
  NOR2_X1 U5525 ( .A1(n5197), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5024) );
  CLKBUF_X1 U5526 ( .A(n5877), .Z(n5878) );
  INV_X1 U5527 ( .A(n9017), .ZN(n4725) );
  NAND2_X1 U5528 ( .A1(n4724), .A2(n9017), .ZN(n4723) );
  NOR2_X1 U5529 ( .A1(n4918), .A2(n4724), .ZN(n4600) );
  NAND2_X1 U5530 ( .A1(n8834), .A2(n4602), .ZN(n4598) );
  INV_X1 U5531 ( .A(n4918), .ZN(n4602) );
  INV_X1 U5532 ( .A(n8812), .ZN(n4590) );
  INV_X1 U5533 ( .A(n6386), .ZN(n4596) );
  NAND2_X1 U5534 ( .A1(n9365), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4487) );
  NAND2_X1 U5535 ( .A1(n9054), .A2(n5686), .ZN(n4829) );
  OR2_X1 U5536 ( .A1(n9055), .A2(n9054), .ZN(n4828) );
  OR2_X1 U5537 ( .A1(n9228), .A2(n9736), .ZN(n4867) );
  AND2_X1 U5538 ( .A1(n9459), .A2(n9457), .ZN(n5039) );
  INV_X1 U5539 ( .A(n9226), .ZN(n4886) );
  NAND2_X1 U5540 ( .A1(n9474), .A2(n9488), .ZN(n9225) );
  INV_X1 U5541 ( .A(n9477), .ZN(n6296) );
  INV_X1 U5542 ( .A(n9147), .ZN(n9223) );
  NAND2_X1 U5543 ( .A1(n4876), .A2(n9772), .ZN(n4875) );
  NOR2_X1 U5544 ( .A1(n9587), .A2(n9785), .ZN(n4876) );
  AND2_X1 U5545 ( .A1(n9120), .A2(n9611), .ZN(n9187) );
  INV_X1 U5546 ( .A(n6357), .ZN(n4954) );
  NAND2_X1 U5547 ( .A1(n6150), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U5548 ( .A1(n7792), .A2(n4872), .ZN(n4871) );
  NOR2_X1 U5549 ( .A1(n9824), .A2(n7361), .ZN(n4872) );
  NOR2_X2 U5550 ( .A1(n6038), .A2(n6698), .ZN(n6058) );
  AND2_X1 U5551 ( .A1(n7318), .A2(n9999), .ZN(n7244) );
  NAND2_X1 U5552 ( .A1(n4825), .A2(n4823), .ZN(n5683) );
  AOI21_X1 U5553 ( .B1(n4827), .B2(n4826), .A(n4824), .ZN(n4823) );
  AOI21_X1 U5554 ( .B1(n5994), .B2(P1_IR_REG_31__SCAN_IN), .A(n4417), .ZN(
        n4416) );
  NAND2_X1 U5555 ( .A1(n6000), .A2(n4290), .ZN(n5998) );
  INV_X1 U5556 ( .A(n5599), .ZN(n5154) );
  XNOR2_X1 U5557 ( .A(n5137), .B(SI_21_), .ZN(n5527) );
  NAND2_X1 U5558 ( .A1(n4794), .A2(n5135), .ZN(n5528) );
  NAND2_X1 U5559 ( .A1(n6203), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U5560 ( .A1(n5102), .A2(n5101), .ZN(n5444) );
  OR2_X1 U5561 ( .A1(n6130), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U5562 ( .A1(n5404), .A2(n5098), .ZN(n5425) );
  AOI211_X1 U5563 ( .C1(n5386), .C2(n5384), .A(n5089), .B(n5390), .ZN(n5090)
         );
  XNOR2_X1 U5564 ( .A(n5074), .B(SI_7_), .ZN(n5329) );
  NAND2_X1 U5565 ( .A1(n4786), .A2(n6587), .ZN(n6030) );
  NAND2_X1 U5566 ( .A1(n6030), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6021) );
  NOR2_X1 U5567 ( .A1(n4996), .A2(n4993), .ZN(n4992) );
  INV_X1 U5568 ( .A(n5033), .ZN(n4993) );
  OAI21_X1 U5569 ( .B1(n4998), .B2(n4996), .A(n8059), .ZN(n4995) );
  NAND2_X1 U5570 ( .A1(n4529), .A2(n4532), .ZN(n8077) );
  OR2_X1 U5571 ( .A1(n7910), .A2(n4535), .ZN(n4529) );
  NAND2_X1 U5572 ( .A1(n4556), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5398) );
  INV_X1 U5573 ( .A(n5376), .ZN(n4556) );
  NAND2_X1 U5574 ( .A1(n4557), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5376) );
  INV_X1 U5575 ( .A(n5356), .ZN(n4557) );
  NAND2_X1 U5576 ( .A1(n5506), .A2(n4294), .ZN(n5560) );
  NAND2_X1 U5577 ( .A1(n5006), .A2(n5005), .ZN(n8160) );
  INV_X1 U5578 ( .A(n8162), .ZN(n5006) );
  NAND2_X1 U5579 ( .A1(n5418), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5436) );
  XNOR2_X1 U5580 ( .A(n7541), .B(n7124), .ZN(n7149) );
  NAND2_X1 U5581 ( .A1(n8138), .A2(n8139), .ZN(n8198) );
  NAND2_X1 U5582 ( .A1(n4999), .A2(n8000), .ZN(n4997) );
  AND2_X1 U5583 ( .A1(n7367), .A2(n7015), .ZN(n7021) );
  OR2_X1 U5584 ( .A1(n4278), .A2(n4418), .ZN(n5400) );
  NAND2_X1 U5585 ( .A1(n6915), .A2(n6914), .ZN(n6958) );
  OR2_X1 U5586 ( .A1(n6958), .A2(n6957), .ZN(n6955) );
  OR2_X1 U5587 ( .A1(n6966), .A2(n6967), .ZN(n6964) );
  OAI21_X1 U5588 ( .B1(n7615), .B2(n7614), .A(n7616), .ZN(n7618) );
  AOI21_X1 U5589 ( .B1(n9055), .B2(n4277), .A(n5692), .ZN(n5704) );
  INV_X1 U5590 ( .A(n8659), .ZN(n8402) );
  NOR2_X1 U5591 ( .A1(n5662), .A2(n5820), .ZN(n5014) );
  NAND2_X1 U5592 ( .A1(n5936), .A2(n5016), .ZN(n5015) );
  INV_X1 U5593 ( .A(n5931), .ZN(n5016) );
  AND2_X1 U5594 ( .A1(n5636), .A2(n5635), .ZN(n8437) );
  OR2_X1 U5595 ( .A1(n8451), .A2(n5669), .ZN(n5636) );
  AND2_X1 U5596 ( .A1(n5660), .A2(n5659), .ZN(n8438) );
  OR2_X1 U5597 ( .A1(n8025), .A2(n5669), .ZN(n5660) );
  NAND2_X1 U5598 ( .A1(n5628), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U5599 ( .A1(n4429), .A2(n4428), .ZN(n8473) );
  NOR2_X1 U5600 ( .A1(n4975), .A2(n8678), .ZN(n4428) );
  AND2_X1 U5601 ( .A1(n8502), .A2(n5802), .ZN(n4853) );
  NAND2_X1 U5602 ( .A1(n8493), .A2(n5036), .ZN(n8481) );
  NAND2_X1 U5603 ( .A1(n5532), .A2(n4559), .ZN(n5591) );
  NOR2_X1 U5604 ( .A1(n8525), .A2(n4974), .ZN(n8495) );
  INV_X1 U5605 ( .A(n4976), .ZN(n4974) );
  NAND2_X1 U5606 ( .A1(n8519), .A2(n8582), .ZN(n4446) );
  NAND2_X1 U5607 ( .A1(n5531), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5562) );
  INV_X1 U5608 ( .A(n5560), .ZN(n5531) );
  NAND2_X1 U5609 ( .A1(n4425), .A2(n4839), .ZN(n4833) );
  AOI21_X1 U5610 ( .B1(n4279), .B2(n4632), .A(n4339), .ZN(n4628) );
  NAND2_X1 U5611 ( .A1(n4385), .A2(n4384), .ZN(n5031) );
  INV_X1 U5612 ( .A(n8717), .ZN(n4384) );
  NAND2_X1 U5613 ( .A1(n4386), .A2(n5773), .ZN(n8602) );
  CLKBUF_X1 U5614 ( .A(n7897), .Z(n4386) );
  INV_X1 U5615 ( .A(n4970), .ZN(n7887) );
  NAND2_X1 U5616 ( .A1(n5382), .A2(n4858), .ZN(n7860) );
  NOR2_X1 U5617 ( .A1(n5763), .A2(n4859), .ZN(n4858) );
  INV_X1 U5618 ( .A(n5758), .ZN(n4859) );
  NAND2_X1 U5619 ( .A1(n4624), .A2(n5022), .ZN(n7761) );
  NAND2_X1 U5620 ( .A1(n7654), .A2(n4979), .ZN(n7775) );
  OR2_X1 U5621 ( .A1(n5323), .A2(n5322), .ZN(n5345) );
  INV_X1 U5622 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U5623 ( .A1(n7654), .A2(n10071), .ZN(n7686) );
  NAND2_X1 U5624 ( .A1(n7308), .A2(n7448), .ZN(n7547) );
  AND2_X1 U5625 ( .A1(n7547), .A2(n5741), .ZN(n7439) );
  NAND2_X1 U5626 ( .A1(n5299), .A2(n5848), .ZN(n7438) );
  NAND2_X1 U5627 ( .A1(n4971), .A2(n4284), .ZN(n7442) );
  INV_X1 U5628 ( .A(n5894), .ZN(n7540) );
  CLKBUF_X1 U5629 ( .A(n6688), .Z(n7534) );
  AND2_X1 U5630 ( .A1(n4483), .A2(n7434), .ZN(n6776) );
  NAND2_X1 U5631 ( .A1(n6774), .A2(n6776), .ZN(n6775) );
  NAND2_X1 U5632 ( .A1(n5640), .A2(n5639), .ZN(n8666) );
  NAND2_X1 U5633 ( .A1(n5627), .A2(n5626), .ZN(n8673) );
  NAND2_X1 U5634 ( .A1(n5601), .A2(n5600), .ZN(n8681) );
  NAND2_X1 U5635 ( .A1(n5558), .A2(n5557), .ZN(n8701) );
  NAND2_X1 U5636 ( .A1(n5547), .A2(n5546), .ZN(n8707) );
  OR2_X1 U5637 ( .A1(n5691), .A2(n6430), .ZN(n4471) );
  OR2_X1 U5638 ( .A1(n5263), .A2(n6439), .ZN(n4470) );
  INV_X1 U5639 ( .A(n10052), .ZN(n8763) );
  CLKBUF_X1 U5640 ( .A(n10129), .Z(n10157) );
  OAI21_X1 U5641 ( .B1(n5716), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5869) );
  INV_X1 U5642 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U5643 ( .A1(n5716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U5644 ( .A1(n5212), .A2(n5009), .ZN(n5716) );
  AND2_X1 U5645 ( .A1(n5011), .A2(n5010), .ZN(n5009) );
  INV_X1 U5646 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5010) );
  AND2_X1 U5647 ( .A1(n5415), .A2(n5448), .ZN(n6919) );
  OR2_X1 U5648 ( .A1(n5411), .A2(n5410), .ZN(n5426) );
  INV_X2 U5649 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5316) );
  OR2_X1 U5650 ( .A1(n5485), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5315) );
  NOR2_X1 U5651 ( .A1(n8899), .A2(n8898), .ZN(n8900) );
  OR2_X1 U5652 ( .A1(n8900), .A2(n4716), .ZN(n4610) );
  AND2_X1 U5653 ( .A1(n6188), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6195) );
  CLKBUF_X1 U5654 ( .A(n6797), .Z(n8924) );
  INV_X1 U5655 ( .A(n7259), .ZN(n4508) );
  INV_X1 U5656 ( .A(n8984), .ZN(n4587) );
  NAND3_X1 U5657 ( .A1(n6749), .A2(n6791), .A3(n6748), .ZN(n4715) );
  NAND2_X1 U5658 ( .A1(n8841), .A2(n8840), .ZN(n8842) );
  AOI21_X1 U5659 ( .B1(n9785), .B2(n8883), .A(n8843), .ZN(n8992) );
  INV_X1 U5660 ( .A(n7720), .ZN(n4913) );
  INV_X1 U5661 ( .A(n4915), .ZN(n4914) );
  NOR2_X1 U5662 ( .A1(n4915), .A2(n4702), .ZN(n4701) );
  INV_X1 U5663 ( .A(n7493), .ZN(n4702) );
  NOR2_X1 U5664 ( .A1(n4915), .A2(n4700), .ZN(n4699) );
  INV_X1 U5665 ( .A(n7509), .ZN(n4700) );
  INV_X1 U5666 ( .A(n8859), .ZN(n8860) );
  OAI22_X1 U5667 ( .A1(n9902), .A2(n6725), .B1(n7681), .B2(n8832), .ZN(n7514)
         );
  NAND2_X1 U5668 ( .A1(n7510), .A2(n7509), .ZN(n4703) );
  NAND2_X1 U5669 ( .A1(n7494), .A2(n7493), .ZN(n4704) );
  NAND2_X1 U5670 ( .A1(n8951), .A2(n8952), .ZN(n8950) );
  NOR2_X2 U5671 ( .A1(n4297), .A2(n10234), .ZN(n6188) );
  MUX2_X1 U5672 ( .A(n9275), .B(n9274), .S(n4302), .Z(n9279) );
  NAND2_X1 U5673 ( .A1(n9278), .A2(n6983), .ZN(n4647) );
  INV_X1 U5674 ( .A(n4650), .ZN(n4651) );
  NAND2_X1 U5675 ( .A1(n4650), .A2(n4308), .ZN(n4649) );
  NOR2_X1 U5676 ( .A1(n9158), .A2(n4405), .ZN(n4655) );
  AND4_X1 U5677 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n7666)
         );
  NAND2_X1 U5678 ( .A1(n6061), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U5679 ( .A1(n6486), .A2(n4331), .ZN(n6510) );
  NAND2_X1 U5680 ( .A1(n6510), .A2(n4424), .ZN(n6623) );
  NAND2_X1 U5681 ( .A1(n6518), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4424) );
  NAND2_X1 U5682 ( .A1(n6561), .A2(n6562), .ZN(n6560) );
  NOR2_X1 U5683 ( .A1(n6605), .A2(n4305), .ZN(n6702) );
  NAND2_X1 U5684 ( .A1(n6702), .A2(n6703), .ZN(n6701) );
  NAND2_X1 U5685 ( .A1(n6601), .A2(n4325), .ZN(n6699) );
  AOI21_X1 U5686 ( .B1(n6699), .B2(n6700), .A(n4773), .ZN(n6680) );
  AND2_X1 U5687 ( .A1(n6522), .A2(n7290), .ZN(n4773) );
  NOR2_X1 U5688 ( .A1(n6534), .A2(n6535), .ZN(n6533) );
  AOI21_X1 U5689 ( .B1(n7321), .B2(n6532), .A(n6533), .ZN(n6548) );
  AND2_X1 U5690 ( .A1(n6816), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4771) );
  NAND2_X1 U5691 ( .A1(n7274), .A2(n4785), .ZN(n7276) );
  OR2_X1 U5692 ( .A1(n7275), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4785) );
  NOR2_X1 U5693 ( .A1(n9380), .A2(n9379), .ZN(n9395) );
  NAND2_X1 U5694 ( .A1(n4866), .A2(n4865), .ZN(n4864) );
  INV_X1 U5695 ( .A(n9725), .ZN(n4865) );
  INV_X1 U5696 ( .A(n4867), .ZN(n4866) );
  NAND2_X1 U5697 ( .A1(n4828), .A2(n4372), .ZN(n9443) );
  INV_X1 U5698 ( .A(n8037), .ZN(n8054) );
  NAND2_X1 U5699 ( .A1(n6288), .A2(n6287), .ZN(n9742) );
  NAND2_X1 U5700 ( .A1(n7875), .A2(n6091), .ZN(n6288) );
  XNOR2_X1 U5701 ( .A(n9498), .B(n9499), .ZN(n4392) );
  AND2_X1 U5702 ( .A1(n9761), .A2(n9342), .ZN(n6371) );
  NAND2_X1 U5703 ( .A1(n4421), .A2(n9548), .ZN(n6372) );
  NOR2_X2 U5704 ( .A1(n4296), .A2(n8944), .ZN(n6251) );
  INV_X1 U5705 ( .A(n9529), .ZN(n9559) );
  NOR2_X1 U5706 ( .A1(n5044), .A2(n4874), .ZN(n9585) );
  INV_X1 U5707 ( .A(n4876), .ZN(n4874) );
  NOR2_X1 U5708 ( .A1(n5044), .A2(n9785), .ZN(n9600) );
  INV_X1 U5709 ( .A(n4382), .ZN(n5044) );
  NAND2_X1 U5710 ( .A1(n9649), .A2(n9168), .ZN(n9629) );
  NAND2_X1 U5711 ( .A1(n6479), .A2(n6091), .ZN(n4438) );
  AND2_X1 U5712 ( .A1(n9174), .A2(n9195), .ZN(n9265) );
  NOR2_X1 U5713 ( .A1(n7360), .A2(n7361), .ZN(n7605) );
  NOR2_X1 U5714 ( .A1(n7360), .A2(n4870), .ZN(n7788) );
  INV_X1 U5715 ( .A(n4872), .ZN(n4870) );
  INV_X1 U5716 ( .A(n4475), .ZN(n6135) );
  INV_X1 U5717 ( .A(n9192), .ZN(n6118) );
  NAND2_X1 U5718 ( .A1(n6452), .A2(n6091), .ZN(n6096) );
  INV_X1 U5719 ( .A(n4502), .ZN(n7360) );
  NAND2_X1 U5720 ( .A1(n6108), .A2(n6107), .ZN(n7640) );
  NAND2_X1 U5721 ( .A1(n4887), .A2(n4888), .ZN(n4891) );
  NAND2_X1 U5722 ( .A1(n4521), .A2(n4520), .ZN(n7316) );
  INV_X1 U5723 ( .A(n7285), .ZN(n4521) );
  NOR2_X2 U5724 ( .A1(n7316), .A2(n7561), .ZN(n7318) );
  AND2_X1 U5725 ( .A1(n9073), .A2(n7078), .ZN(n7314) );
  INV_X1 U5726 ( .A(n6348), .ZN(n9255) );
  NOR2_X2 U5727 ( .A1(n7069), .A2(n7073), .ZN(n7286) );
  INV_X1 U5728 ( .A(n4578), .ZN(n7063) );
  NAND2_X1 U5729 ( .A1(n4670), .A2(n4668), .ZN(n4667) );
  AND4_X2 U5730 ( .A1(n5991), .A2(n5989), .A3(n5990), .A4(n4480), .ZN(n7004)
         );
  NAND2_X1 U5731 ( .A1(n6060), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4480) );
  AND3_X1 U5732 ( .A1(n9503), .A2(n10008), .A3(n9502), .ZN(n9751) );
  INV_X1 U5733 ( .A(n9571), .ZN(n9772) );
  NAND2_X1 U5734 ( .A1(n6176), .A2(n6175), .ZN(n9807) );
  INV_X1 U5735 ( .A(n7050), .ZN(n7049) );
  AND2_X1 U5736 ( .A1(n6733), .A2(n6577), .ZN(n6980) );
  AND2_X1 U5737 ( .A1(n6981), .A2(n6414), .ZN(n6638) );
  INV_X1 U5738 ( .A(n4462), .ZN(n7007) );
  XNOR2_X1 U5739 ( .A(n5680), .B(n5178), .ZN(n9065) );
  NAND2_X1 U5740 ( .A1(n4709), .A2(n4708), .ZN(n6001) );
  NAND2_X1 U5741 ( .A1(n5981), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4708) );
  XNOR2_X1 U5742 ( .A(n5637), .B(n5638), .ZN(n8799) );
  NAND2_X1 U5743 ( .A1(n5167), .A2(n5166), .ZN(n5637) );
  INV_X1 U5744 ( .A(n4586), .ZN(n4585) );
  OAI21_X1 U5745 ( .B1(n6394), .B2(n5993), .A(n6390), .ZN(n4586) );
  XNOR2_X1 U5746 ( .A(n5624), .B(n5625), .ZN(n7875) );
  OAI21_X1 U5747 ( .B1(n5499), .B2(n5121), .A(n5123), .ZN(n5514) );
  XNOR2_X1 U5748 ( .A(n5499), .B(n5498), .ZN(n6570) );
  AND2_X1 U5749 ( .A1(n6168), .A2(n6167), .ZN(n6170) );
  INV_X1 U5750 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6167) );
  INV_X1 U5751 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6181) );
  XNOR2_X1 U5752 ( .A(n5392), .B(n5391), .ZN(n6454) );
  NAND2_X1 U5753 ( .A1(n5312), .A2(n5311), .ZN(n4439) );
  OR2_X1 U5754 ( .A1(n6045), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U5755 ( .A1(n5226), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4412) );
  NOR2_X1 U5756 ( .A1(n9880), .A2(n9879), .ZN(n9881) );
  NOR2_X1 U5757 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10270), .ZN(n9882) );
  AND4_X1 U5758 ( .A1(n5350), .A2(n5349), .A3(n5348), .A4(n5347), .ZN(n7694)
         );
  AOI21_X1 U5759 ( .B1(n8213), .B2(n8060), .A(n8230), .ZN(n8064) );
  OR2_X1 U5760 ( .A1(n8230), .A2(n8012), .ZN(n8209) );
  NAND2_X1 U5761 ( .A1(n4538), .A2(n4537), .ZN(n7808) );
  AOI21_X1 U5762 ( .B1(n4540), .B2(n4543), .A(n4344), .ZN(n4537) );
  NAND2_X1 U5763 ( .A1(n7735), .A2(n7734), .ZN(n7740) );
  NAND2_X1 U5764 ( .A1(n4536), .A2(n4540), .ZN(n7735) );
  OR2_X1 U5765 ( .A1(n7452), .A2(n4543), .ZN(n4536) );
  NAND2_X1 U5766 ( .A1(n8090), .A2(n7971), .ZN(n8091) );
  OR2_X1 U5767 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  NAND2_X1 U5768 ( .A1(n4546), .A2(n7455), .ZN(n7591) );
  OR2_X1 U5769 ( .A1(n7452), .A2(n7451), .ZN(n4546) );
  NAND2_X1 U5770 ( .A1(n7097), .A2(n7434), .ZN(n4987) );
  NAND2_X1 U5771 ( .A1(n7124), .A2(n7102), .ZN(n4986) );
  AND2_X1 U5772 ( .A1(n7122), .A2(n7033), .ZN(n7036) );
  AND4_X1 U5773 ( .A1(n5423), .A2(n5422), .A3(n5421), .A4(n5420), .ZN(n8071)
         );
  AND2_X1 U5774 ( .A1(n7996), .A2(n5033), .ZN(n4989) );
  NAND2_X1 U5775 ( .A1(n8116), .A2(n8115), .ZN(n8212) );
  NAND2_X1 U5776 ( .A1(n7181), .A2(n7173), .ZN(n7193) );
  AND2_X1 U5777 ( .A1(n5616), .A2(n5603), .ZN(n8484) );
  NAND2_X1 U5778 ( .A1(n7183), .A2(n7182), .ZN(n7181) );
  NAND2_X1 U5779 ( .A1(n7452), .A2(n4544), .ZN(n4539) );
  NAND2_X1 U5780 ( .A1(n8091), .A2(n7975), .ZN(n8162) );
  AND4_X1 U5781 ( .A1(n5460), .A2(n5459), .A3(n5458), .A4(n5457), .ZN(n8171)
         );
  NAND2_X1 U5782 ( .A1(n7942), .A2(n7941), .ZN(n8169) );
  XNOR2_X1 U5783 ( .A(n7148), .B(n7149), .ZN(n7153) );
  NAND2_X1 U5784 ( .A1(n4525), .A2(n8196), .ZN(n8090) );
  NAND2_X1 U5785 ( .A1(n8198), .A2(n7965), .ZN(n4525) );
  OR2_X1 U5786 ( .A1(n8221), .A2(n8605), .ZN(n8204) );
  OR2_X1 U5787 ( .A1(n8221), .A2(n8603), .ZN(n8205) );
  NAND2_X1 U5788 ( .A1(n4551), .A2(n4550), .ZN(n7199) );
  OAI21_X1 U5789 ( .B1(n7194), .B2(n4554), .A(n4555), .ZN(n4550) );
  INV_X1 U5790 ( .A(n7173), .ZN(n4554) );
  INV_X1 U5791 ( .A(n8230), .ZN(n8184) );
  AOI21_X1 U5792 ( .B1(n8116), .B2(n4998), .A(n4526), .ZN(n8213) );
  INV_X1 U5793 ( .A(n4997), .ZN(n4526) );
  INV_X1 U5794 ( .A(n7299), .ZN(n5933) );
  AND2_X1 U5795 ( .A1(n4431), .A2(n4430), .ZN(n4503) );
  NAND2_X1 U5796 ( .A1(n4505), .A2(n4504), .ZN(n4431) );
  AND2_X1 U5797 ( .A1(n5678), .A2(n5677), .ZN(n7634) );
  AOI21_X1 U5798 ( .B1(n8431), .B2(n5647), .A(n5646), .ZN(n8217) );
  NAND2_X1 U5799 ( .A1(n5539), .A2(n5538), .ZN(n8543) );
  OR2_X1 U5800 ( .A1(n8528), .A2(n5669), .ZN(n5539) );
  NAND4_X2 U5801 ( .A1(n5290), .A2(n5289), .A3(n5288), .A4(n5287), .ZN(n8259)
         );
  INV_X1 U5802 ( .A(n7535), .ZN(n8261) );
  CLKBUF_X1 U5803 ( .A(n7034), .Z(n4483) );
  NAND2_X1 U5804 ( .A1(n8276), .A2(n8275), .ZN(n8288) );
  NAND2_X1 U5805 ( .A1(n6669), .A2(n6668), .ZN(n6841) );
  NAND2_X1 U5806 ( .A1(n6860), .A2(n6859), .ZN(n8320) );
  NAND2_X1 U5807 ( .A1(n6881), .A2(n6880), .ZN(n8347) );
  AND2_X1 U5808 ( .A1(n5467), .A2(n5451), .ZN(n7136) );
  AND2_X1 U5809 ( .A1(n6475), .A2(n6474), .ZN(n8395) );
  INV_X1 U5810 ( .A(n8391), .ZN(n4451) );
  INV_X1 U5811 ( .A(n8666), .ZN(n8433) );
  AND2_X1 U5812 ( .A1(n5630), .A2(n5617), .ZN(n8475) );
  AOI21_X1 U5813 ( .B1(n8465), .B2(n8464), .A(n8463), .ZN(n8680) );
  NAND2_X1 U5814 ( .A1(n5584), .A2(n5802), .ZN(n8503) );
  INV_X1 U5815 ( .A(n4464), .ZN(n4463) );
  OAI22_X1 U5816 ( .A1(n8537), .A2(n8605), .B1(n8603), .B2(n8536), .ZN(n4464)
         );
  INV_X1 U5817 ( .A(n8701), .ZN(n8553) );
  INV_X1 U5818 ( .A(n8707), .ZN(n8565) );
  NAND2_X1 U5819 ( .A1(n4841), .A2(n4839), .ZN(n8579) );
  NAND2_X1 U5820 ( .A1(n8607), .A2(n4303), .ZN(n8596) );
  OR2_X1 U5821 ( .A1(n7896), .A2(n4632), .ZN(n4627) );
  AND2_X1 U5822 ( .A1(n4634), .A2(n4285), .ZN(n8609) );
  NAND2_X1 U5823 ( .A1(n5029), .A2(n4280), .ZN(n7884) );
  AND2_X1 U5824 ( .A1(n5029), .A2(n4347), .ZN(n7886) );
  INV_X1 U5825 ( .A(n8743), .ZN(n7847) );
  NAND2_X1 U5826 ( .A1(n5382), .A2(n5758), .ZN(n7747) );
  NAND2_X1 U5827 ( .A1(n7655), .A2(n4272), .ZN(n7685) );
  NAND2_X1 U5828 ( .A1(n4854), .A2(n5747), .ZN(n7651) );
  CLKBUF_X1 U5829 ( .A(n7545), .Z(n7546) );
  NAND2_X1 U5830 ( .A1(n4850), .A2(n5729), .ZN(n7108) );
  INV_X1 U5831 ( .A(n8597), .ZN(n8555) );
  OAI211_X1 U5832 ( .C1(n5943), .C2(n7102), .A(n7530), .B(n8763), .ZN(n7576)
         );
  INV_X1 U5833 ( .A(n8641), .ZN(n8527) );
  OR2_X1 U5834 ( .A1(n7367), .A2(n6696), .ZN(n10081) );
  INV_X1 U5835 ( .A(n8664), .ZN(n4490) );
  AND2_X1 U5836 ( .A1(n7927), .A2(n4343), .ZN(n4510) );
  AND2_X2 U5837 ( .A1(n5964), .A2(n5963), .ZN(n10076) );
  INV_X1 U5838 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U5839 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  XNOR2_X1 U5840 ( .A(n5869), .B(n5717), .ZN(n7299) );
  NAND2_X1 U5841 ( .A1(n4739), .A2(n4737), .ZN(n5544) );
  NAND2_X1 U5842 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4738), .ZN(n4737) );
  NAND2_X1 U5843 ( .A1(n4740), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n4739) );
  INV_X1 U5844 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6478) );
  INV_X1 U5845 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10183) );
  INV_X1 U5846 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6459) );
  AND2_X1 U5847 ( .A1(n5393), .A2(n5372), .ZN(n8344) );
  XNOR2_X1 U5848 ( .A(n5258), .B(n5257), .ZN(n6661) );
  AND4_X1 U5849 ( .A1(n6090), .A2(n6089), .A3(n6088), .A4(n6087), .ZN(n7570)
         );
  AND4_X1 U5850 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(n9500)
         );
  AND2_X1 U5851 ( .A1(n9029), .A2(n8900), .ZN(n8931) );
  CLKBUF_X1 U5852 ( .A(n9814), .Z(n4411) );
  NAND2_X1 U5853 ( .A1(n6748), .A2(n6749), .ZN(n4930) );
  AND2_X1 U5854 ( .A1(n6239), .A2(n6238), .ZN(n9562) );
  NAND2_X1 U5855 ( .A1(n4925), .A2(n8849), .ZN(n8943) );
  NAND2_X1 U5856 ( .A1(n7676), .A2(n7675), .ZN(n7719) );
  AND2_X1 U5857 ( .A1(n6212), .A2(n6211), .ZN(n9632) );
  NAND2_X1 U5858 ( .A1(n7757), .A2(n6091), .ZN(n6266) );
  OR2_X1 U5859 ( .A1(n4714), .A2(n4712), .ZN(n7256) );
  INV_X1 U5860 ( .A(n4929), .ZN(n4712) );
  NAND2_X1 U5861 ( .A1(n4715), .A2(n6796), .ZN(n4714) );
  AND3_X1 U5862 ( .A1(n6166), .A2(n6165), .A3(n6164), .ZN(n9098) );
  AND4_X1 U5863 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n7644)
         );
  NAND2_X1 U5864 ( .A1(n7519), .A2(n7518), .ZN(n7676) );
  AND2_X1 U5865 ( .A1(n6201), .A2(n6200), .ZN(n9657) );
  NOR2_X1 U5866 ( .A1(n8834), .A2(n8833), .ZN(n9016) );
  AND2_X1 U5867 ( .A1(n7646), .A2(n9957), .ZN(n9022) );
  OR2_X1 U5868 ( .A1(n6730), .A2(n6729), .ZN(n9032) );
  OR2_X1 U5869 ( .A1(n6730), .A2(n6579), .ZN(n9048) );
  AND2_X1 U5870 ( .A1(n6598), .A2(n6597), .ZN(n9043) );
  INV_X1 U5871 ( .A(n9032), .ZN(n9050) );
  INV_X1 U5872 ( .A(n9022), .ZN(n9053) );
  INV_X1 U5873 ( .A(n9535), .ZN(n9341) );
  INV_X1 U5874 ( .A(n9548), .ZN(n9342) );
  OAI21_X1 U5875 ( .B1(n9550), .B2(n6278), .A(n6247), .ZN(n9560) );
  INV_X1 U5876 ( .A(n9615), .ZN(n9344) );
  INV_X1 U5877 ( .A(n9632), .ZN(n9597) );
  INV_X1 U5878 ( .A(n7666), .ZN(n9346) );
  INV_X1 U5879 ( .A(n6339), .ZN(n9355) );
  INV_X1 U5880 ( .A(n7004), .ZN(n6334) );
  AOI21_X1 U5881 ( .B1(n10116), .B2(n6523), .A(n6675), .ZN(n6530) );
  AOI22_X1 U5882 ( .A1(n6812), .A2(n6811), .B1(n6810), .B2(n6809), .ZN(n6813)
         );
  INV_X1 U5883 ( .A(n4783), .ZN(n7389) );
  INV_X1 U5884 ( .A(n4488), .ZN(n9364) );
  OAI21_X1 U5885 ( .B1(n9380), .B2(n4788), .A(n4787), .ZN(n9413) );
  NAND2_X1 U5886 ( .A1(n4789), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4788) );
  INV_X1 U5887 ( .A(n9398), .ZN(n4789) );
  NOR2_X1 U5888 ( .A1(n9388), .A2(n4423), .ZN(n9392) );
  AND2_X1 U5889 ( .A1(n9390), .A2(n9389), .ZN(n4423) );
  OR2_X1 U5890 ( .A1(n9922), .A2(n9921), .ZN(n9925) );
  INV_X1 U5891 ( .A(n9441), .ZN(n4775) );
  OAI21_X1 U5892 ( .B1(n9465), .B2(n4862), .A(n4861), .ZN(n9723) );
  NAND2_X1 U5893 ( .A1(n9443), .A2(n4863), .ZN(n4862) );
  OAI21_X1 U5894 ( .B1(n9465), .B2(n4864), .A(n9721), .ZN(n4861) );
  INV_X1 U5895 ( .A(n4864), .ZN(n4863) );
  AOI21_X1 U5896 ( .B1(n8051), .B2(n9705), .A(n8050), .ZN(n8052) );
  NAND2_X1 U5897 ( .A1(n4881), .A2(n9708), .ZN(n4880) );
  NOR2_X1 U5898 ( .A1(n4473), .A2(n8903), .ZN(n4472) );
  NAND2_X1 U5899 ( .A1(n6316), .A2(n4459), .ZN(n9477) );
  OR2_X1 U5900 ( .A1(n6295), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n4459) );
  INV_X1 U5901 ( .A(n9742), .ZN(n9494) );
  NAND2_X1 U5902 ( .A1(n6275), .A2(n6274), .ZN(n9752) );
  NAND2_X1 U5903 ( .A1(n4391), .A2(n4389), .ZN(n9750) );
  INV_X1 U5904 ( .A(n4390), .ZN(n4389) );
  NAND2_X1 U5905 ( .A1(n4392), .A2(n9708), .ZN(n4391) );
  OAI22_X1 U5906 ( .A1(n9500), .A2(n9656), .B1(n9654), .B2(n9535), .ZN(n4390)
         );
  AND2_X1 U5907 ( .A1(n6268), .A2(n6276), .ZN(n9520) );
  NOR2_X1 U5908 ( .A1(n9532), .A2(n4572), .ZN(n9514) );
  INV_X1 U5909 ( .A(n6373), .ZN(n9525) );
  NAND2_X1 U5910 ( .A1(n4479), .A2(n4477), .ZN(n9766) );
  INV_X1 U5911 ( .A(n4478), .ZN(n4477) );
  OAI22_X1 U5912 ( .A1(n9548), .A2(n9656), .B1(n9654), .B2(n9578), .ZN(n4478)
         );
  NAND2_X1 U5913 ( .A1(n4964), .A2(n4961), .ZN(n9542) );
  NAND2_X1 U5914 ( .A1(n4388), .A2(n9583), .ZN(n4961) );
  NAND2_X1 U5915 ( .A1(n4388), .A2(n4967), .ZN(n9569) );
  NAND2_X1 U5916 ( .A1(n4967), .A2(n4968), .ZN(n9567) );
  INV_X1 U5917 ( .A(n6241), .ZN(n9577) );
  CLKBUF_X1 U5918 ( .A(n9605), .Z(n9606) );
  NAND2_X1 U5919 ( .A1(n4951), .A2(n4949), .ZN(n9621) );
  NAND2_X1 U5920 ( .A1(n4951), .A2(n6365), .ZN(n9619) );
  NAND2_X1 U5921 ( .A1(n4953), .A2(n4956), .ZN(n9681) );
  NAND2_X1 U5922 ( .A1(n4491), .A2(n4368), .ZN(n4953) );
  NAND2_X1 U5923 ( .A1(n4957), .A2(n6356), .ZN(n9715) );
  OR2_X1 U5924 ( .A1(n4491), .A2(n6355), .ZN(n4957) );
  NAND2_X1 U5925 ( .A1(n7786), .A2(n9195), .ZN(n9702) );
  NAND2_X1 U5926 ( .A1(n4941), .A2(n4942), .ZN(n7222) );
  AND2_X1 U5927 ( .A1(n4946), .A2(n4943), .ZN(n4942) );
  INV_X1 U5928 ( .A(n9716), .ZN(n9677) );
  NAND2_X1 U5929 ( .A1(n9066), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4711) );
  OR2_X1 U5930 ( .A1(n6981), .A2(n9849), .ZN(n9667) );
  NAND2_X1 U5931 ( .A1(n9066), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6008) );
  INV_X1 U5932 ( .A(n9667), .ZN(n9710) );
  INV_X1 U5933 ( .A(n9714), .ZN(n9672) );
  INV_X1 U5934 ( .A(n10029), .ZN(n10026) );
  OR2_X1 U5935 ( .A1(n9739), .A2(n9961), .ZN(n4379) );
  NOR2_X1 U5936 ( .A1(n9480), .A2(n6331), .ZN(n6383) );
  NAND2_X1 U5937 ( .A1(n6330), .A2(n6329), .ZN(n6331) );
  NAND2_X1 U5938 ( .A1(n9749), .A2(n9748), .ZN(n9832) );
  INV_X1 U5939 ( .A(n9747), .ZN(n9748) );
  INV_X1 U5940 ( .A(n9741), .ZN(n9749) );
  OR2_X1 U5941 ( .A1(n9806), .A2(n9805), .ZN(n9843) );
  INV_X1 U5942 ( .A(n10017), .ZN(n10015) );
  NAND2_X1 U5944 ( .A1(n4960), .A2(n5981), .ZN(n4695) );
  NOR2_X1 U5945 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4960) );
  OAI21_X1 U5946 ( .B1(n5167), .B2(n4802), .A(n4799), .ZN(n5649) );
  NAND2_X1 U5947 ( .A1(n4497), .A2(n4496), .ZN(n4513) );
  INV_X1 U5948 ( .A(n5586), .ZN(n4496) );
  NAND2_X1 U5949 ( .A1(n6204), .A2(n6203), .ZN(n6213) );
  INV_X1 U5950 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6556) );
  INV_X1 U5951 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6481) );
  INV_X1 U5952 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6457) );
  INV_X1 U5953 ( .A(n6684), .ZN(n6523) );
  OAI21_X1 U5954 ( .B1(n5245), .B2(n6432), .A(n5046), .ZN(n5246) );
  NAND2_X1 U5955 ( .A1(n4410), .A2(SI_0_), .ZN(n5992) );
  INV_X1 U5956 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10219) );
  AND2_X1 U5957 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9881), .ZN(n10270) );
  XNOR2_X1 U5958 ( .A(n9886), .B(n9887), .ZN(n10273) );
  XNOR2_X1 U5959 ( .A(n9890), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n10280) );
  NOR2_X1 U5960 ( .A1(n9893), .A2(n10281), .ZN(n10112) );
  NOR2_X1 U5961 ( .A1(n10107), .A2(n4377), .ZN(n10106) );
  NAND2_X1 U5962 ( .A1(n10106), .A2(n10105), .ZN(n10104) );
  OAI21_X1 U5963 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10104), .ZN(n10102) );
  NAND2_X1 U5964 ( .A1(n10102), .A2(n10103), .ZN(n10101) );
  NAND2_X1 U5965 ( .A1(n10101), .A2(n4453), .ZN(n10099) );
  NAND2_X1 U5966 ( .A1(n4455), .A2(n4454), .ZN(n4453) );
  INV_X1 U5967 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n4455) );
  INV_X1 U5968 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n4454) );
  OAI21_X1 U5969 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10098), .ZN(n10096) );
  NAND2_X1 U5970 ( .A1(n10096), .A2(n10097), .ZN(n10095) );
  NAND2_X1 U5971 ( .A1(n10095), .A2(n4456), .ZN(n10093) );
  NAND2_X1 U5972 ( .A1(n4458), .A2(n4457), .ZN(n4456) );
  INV_X1 U5973 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n4458) );
  INV_X1 U5974 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n4457) );
  NAND2_X1 U5975 ( .A1(n4452), .A2(n4449), .ZN(P2_U3264) );
  AOI21_X1 U5976 ( .B1(n4451), .B2(n8390), .A(n4450), .ZN(n4449) );
  OR2_X1 U5977 ( .A1(n8392), .A2(n8390), .ZN(n4452) );
  OAI21_X1 U5978 ( .B1(n8394), .B2(n8395), .A(n8393), .ZN(n4450) );
  NOR2_X1 U5979 ( .A1(n8694), .A2(n4273), .ZN(n8521) );
  NAND2_X1 U5980 ( .A1(n4719), .A2(n4608), .ZN(n4612) );
  NOR2_X1 U5981 ( .A1(n4716), .A2(n4933), .ZN(n4608) );
  OR2_X1 U5982 ( .A1(n9334), .A2(n9333), .ZN(n4402) );
  AND4_X1 U5983 ( .A1(n9422), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(n9423)
         );
  NOR2_X1 U5984 ( .A1(n4776), .A2(n4775), .ZN(n4774) );
  OAI21_X1 U5985 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9897), .A(n10274), .ZN(
        n9900) );
  NOR2_X1 U5986 ( .A1(n6379), .A2(n9440), .ZN(n9160) );
  AND2_X1 U5987 ( .A1(n5021), .A2(n4630), .ZN(n4279) );
  AND2_X1 U5988 ( .A1(n7885), .A2(n4347), .ZN(n4280) );
  AND2_X1 U5989 ( .A1(n9240), .A2(n9239), .ZN(n4281) );
  BUF_X2 U5990 ( .A(n6715), .Z(n8892) );
  INV_X1 U5991 ( .A(n9902), .ZN(n7361) );
  OR2_X1 U5992 ( .A1(n9814), .A2(n9685), .ZN(n4282) );
  AND2_X1 U5993 ( .A1(n8833), .A2(n4725), .ZN(n4283) );
  INV_X1 U5994 ( .A(n9201), .ZN(n4686) );
  INV_X1 U5995 ( .A(n4543), .ZN(n4542) );
  NAND2_X1 U5996 ( .A1(n8259), .A2(n7378), .ZN(n5847) );
  AND2_X1 U5997 ( .A1(n4972), .A2(n7378), .ZN(n4284) );
  OR2_X1 U5998 ( .A1(n8728), .A2(n5915), .ZN(n4285) );
  AND2_X1 U5999 ( .A1(n4977), .A2(n8748), .ZN(n4286) );
  AND2_X1 U6000 ( .A1(n5307), .A2(n4357), .ZN(n4287) );
  AND2_X1 U6001 ( .A1(n5749), .A2(n7689), .ZN(n7656) );
  AND2_X1 U6002 ( .A1(n9624), .A2(n9597), .ZN(n4288) );
  AND2_X1 U6003 ( .A1(n4432), .A2(n4355), .ZN(n4289) );
  AND2_X1 U6004 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4290) );
  INV_X1 U6005 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10137) );
  INV_X1 U6006 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6007 ( .A1(n5374), .A2(n5373), .ZN(n7774) );
  AND2_X1 U6008 ( .A1(n5796), .A2(n5788), .ZN(n4291) );
  AND2_X1 U6009 ( .A1(n4882), .A2(n4326), .ZN(n4292) );
  OR2_X1 U6010 ( .A1(n8487), .A2(n4635), .ZN(n4293) );
  INV_X1 U6011 ( .A(n8595), .ZN(n4843) );
  AND2_X1 U6012 ( .A1(n4562), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n4294) );
  AND2_X1 U6013 ( .A1(n4561), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n4295) );
  INV_X1 U6014 ( .A(n4501), .ZN(n4868) );
  OR2_X2 U6015 ( .A1(n6233), .A2(n8999), .ZN(n4296) );
  OR2_X1 U6016 ( .A1(n6160), .A2(n6159), .ZN(n4297) );
  INV_X1 U6017 ( .A(n8892), .ZN(n8883) );
  OR2_X1 U6018 ( .A1(n6276), .A2(n8954), .ZN(n4298) );
  INV_X1 U6019 ( .A(n8833), .ZN(n4724) );
  INV_X2 U6020 ( .A(n6797), .ZN(n6727) );
  AND2_X1 U6021 ( .A1(n5356), .A2(n5346), .ZN(n4299) );
  NAND2_X1 U6022 ( .A1(n9752), .A2(n9516), .ZN(n9311) );
  INV_X1 U6023 ( .A(n7434), .ZN(n7102) );
  INV_X1 U6024 ( .A(n9814), .ZN(n4873) );
  INV_X1 U6025 ( .A(n6056), .ZN(n6086) );
  NAND2_X1 U6026 ( .A1(n4291), .A2(n5783), .ZN(n4840) );
  AND2_X1 U6027 ( .A1(n9265), .A2(n9175), .ZN(n4300) );
  OR2_X1 U6028 ( .A1(n8707), .A2(n8203), .ZN(n5797) );
  OR2_X1 U6029 ( .A1(n9761), .A2(n9548), .ZN(n9216) );
  INV_X1 U6030 ( .A(n4380), .ZN(n4422) );
  NAND2_X1 U6031 ( .A1(n4382), .A2(n4381), .ZN(n4380) );
  NOR2_X1 U6032 ( .A1(n9772), .A2(n9578), .ZN(n4301) );
  AND3_X1 U6033 ( .A1(n9236), .A2(n9272), .A3(n4440), .ZN(n4302) );
  OR2_X1 U6034 ( .A1(n8621), .A2(n8248), .ZN(n4303) );
  NAND2_X1 U6035 ( .A1(n8688), .A2(n5924), .ZN(n4304) );
  AND2_X1 U6036 ( .A1(n6521), .A2(n6515), .ZN(n4305) );
  AND2_X1 U6037 ( .A1(n8845), .A2(n8844), .ZN(n4306) );
  AND2_X1 U6038 ( .A1(n7993), .A2(n7992), .ZN(n4307) );
  INV_X1 U6039 ( .A(n5927), .ZN(n5020) );
  INV_X1 U6040 ( .A(n4926), .ZN(n8917) );
  AND4_X1 U6041 ( .A1(n9236), .A2(n9284), .A3(n9164), .A4(n6379), .ZN(n4308)
         );
  INV_X1 U6042 ( .A(n5916), .ZN(n4631) );
  OR2_X1 U6043 ( .A1(n6650), .A2(n6663), .ZN(n4309) );
  OR2_X1 U6044 ( .A1(n5864), .A2(n5837), .ZN(n4310) );
  XNOR2_X1 U6045 ( .A(n8666), .B(n8217), .ZN(n8435) );
  INV_X1 U6046 ( .A(n9531), .ZN(n4406) );
  NAND2_X1 U6047 ( .A1(n5298), .A2(n5297), .ZN(n5900) );
  INV_X1 U6048 ( .A(n9228), .ZN(n9729) );
  OAI21_X1 U6049 ( .B1(n8834), .B2(n4283), .A(n4723), .ZN(n4926) );
  INV_X1 U6050 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6309) );
  INV_X1 U6051 ( .A(n4429), .ZN(n8525) );
  NOR2_X1 U6052 ( .A1(n8549), .A2(n8698), .ZN(n4429) );
  OR2_X1 U6053 ( .A1(n5044), .A2(n4875), .ZN(n4311) );
  AND4_X1 U6054 ( .A1(n6129), .A2(n6128), .A3(n6127), .A4(n6126), .ZN(n7681)
         );
  INV_X1 U6055 ( .A(n7681), .ZN(n9347) );
  OR2_X1 U6056 ( .A1(n7547), .A2(n5839), .ZN(n4312) );
  NOR2_X1 U6057 ( .A1(n9395), .A2(n9396), .ZN(n4313) );
  AND4_X1 U6058 ( .A1(n9273), .A2(n9317), .A3(n9316), .A4(n9459), .ZN(n4314)
         );
  NAND2_X1 U6059 ( .A1(n6133), .A2(n6132), .ZN(n9824) );
  OR2_X1 U6060 ( .A1(n4765), .A2(n4766), .ZN(n4315) );
  NAND2_X1 U6061 ( .A1(n4833), .A2(n4837), .ZN(n8513) );
  INV_X1 U6062 ( .A(n9736), .ZN(n4473) );
  AND2_X1 U6063 ( .A1(n4636), .A2(n5923), .ZN(n4316) );
  AND2_X1 U6064 ( .A1(n4841), .A2(n5783), .ZN(n4317) );
  OR2_X1 U6065 ( .A1(n6650), .A2(n6661), .ZN(n4318) );
  INV_X1 U6066 ( .A(n4545), .ZN(n4544) );
  NAND2_X1 U6067 ( .A1(n4549), .A2(n7455), .ZN(n4545) );
  NAND2_X1 U6068 ( .A1(n5840), .A2(n5839), .ZN(n4319) );
  AND2_X1 U6069 ( .A1(n4639), .A2(n4637), .ZN(n4320) );
  AND2_X1 U6070 ( .A1(n9587), .A2(n9562), .ZN(n9246) );
  INV_X1 U6071 ( .A(n8876), .ZN(n4935) );
  AND2_X1 U6072 ( .A1(n9216), .A2(n9218), .ZN(n4321) );
  OR2_X1 U6073 ( .A1(n6564), .A2(n6514), .ZN(n4322) );
  INV_X1 U6074 ( .A(n4840), .ZN(n4839) );
  OR2_X1 U6075 ( .A1(n7986), .A2(n7981), .ZN(n4323) );
  INV_X1 U6076 ( .A(n8688), .ZN(n8497) );
  AND2_X1 U6077 ( .A1(n4927), .A2(n8860), .ZN(n4324) );
  OR2_X1 U6078 ( .A1(n6612), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4325) );
  NAND2_X1 U6079 ( .A1(n9273), .A2(n5039), .ZN(n4326) );
  NAND2_X1 U6080 ( .A1(n5100), .A2(SI_13_), .ZN(n5406) );
  AND2_X1 U6081 ( .A1(n4869), .A2(n4873), .ZN(n4327) );
  AND3_X1 U6082 ( .A1(n9074), .A2(n4894), .A3(n9299), .ZN(n4328) );
  AND2_X1 U6083 ( .A1(n9642), .A2(n9657), .ZN(n9170) );
  NAND2_X1 U6084 ( .A1(n4852), .A2(n4304), .ZN(n4329) );
  AND4_X1 U6085 ( .A1(n9140), .A2(n9141), .A3(n9459), .A4(n9139), .ZN(n4330)
         );
  AND2_X1 U6086 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4331) );
  NOR2_X1 U6087 ( .A1(n8627), .A2(n8254), .ZN(n4332) );
  INV_X1 U6088 ( .A(n4973), .ZN(n8482) );
  NOR2_X1 U6089 ( .A1(n8525), .A2(n4975), .ZN(n4973) );
  OR2_X1 U6090 ( .A1(n9228), .A2(n9462), .ZN(n4333) );
  AND2_X1 U6091 ( .A1(n4279), .A2(n4627), .ZN(n4334) );
  INV_X1 U6092 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6071) );
  INV_X1 U6093 ( .A(n8017), .ZN(n8406) );
  NAND2_X1 U6094 ( .A1(n5651), .A2(n5650), .ZN(n8017) );
  NAND2_X1 U6095 ( .A1(n8972), .A2(n9040), .ZN(n4335) );
  INV_X1 U6096 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10148) );
  INV_X1 U6097 ( .A(n4638), .ZN(n4637) );
  NOR2_X1 U6098 ( .A1(n8247), .A2(n4433), .ZN(n4638) );
  AND2_X1 U6099 ( .A1(n4919), .A2(n9017), .ZN(n4336) );
  NAND2_X1 U6100 ( .A1(n5320), .A2(n5319), .ZN(n7448) );
  AND2_X1 U6101 ( .A1(n5125), .A2(SI_18_), .ZN(n4337) );
  NAND2_X1 U6102 ( .A1(n5981), .A2(n10137), .ZN(n4338) );
  NOR2_X1 U6103 ( .A1(n8717), .A2(n8581), .ZN(n4339) );
  NOR2_X1 U6104 ( .A1(n8733), .A2(n8250), .ZN(n4340) );
  AND2_X1 U6105 ( .A1(n8936), .A2(n9043), .ZN(n4341) );
  INV_X1 U6106 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4738) );
  NAND2_X1 U6107 ( .A1(n5661), .A2(n5826), .ZN(n5936) );
  INV_X1 U6108 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U6109 ( .A1(n9173), .A2(n9177), .ZN(n9247) );
  INV_X1 U6110 ( .A(n9247), .ZN(n4911) );
  AND2_X1 U6111 ( .A1(n5108), .A2(SI_14_), .ZN(n4342) );
  OR2_X1 U6112 ( .A1(n8406), .A2(n10070), .ZN(n4343) );
  INV_X1 U6113 ( .A(n5030), .ZN(n4555) );
  NAND2_X1 U6114 ( .A1(n7742), .A2(n7734), .ZN(n4344) );
  AND2_X1 U6115 ( .A1(n9758), .A2(n9535), .ZN(n9148) );
  AND2_X1 U6116 ( .A1(n8855), .A2(n8854), .ZN(n8940) );
  INV_X1 U6117 ( .A(n8940), .ZN(n4927) );
  OR2_X1 U6118 ( .A1(n4293), .A2(n4316), .ZN(n4345) );
  NAND2_X1 U6119 ( .A1(n5831), .A2(n5830), .ZN(n8410) );
  AND2_X1 U6120 ( .A1(n6520), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4346) );
  NAND2_X1 U6121 ( .A1(n8737), .A2(n8251), .ZN(n4347) );
  AND2_X1 U6122 ( .A1(n8938), .A2(n8939), .ZN(n4348) );
  AND2_X1 U6123 ( .A1(n6518), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4349) );
  NAND2_X2 U6124 ( .A1(n6256), .A2(n6255), .ZN(n9761) );
  INV_X1 U6125 ( .A(n9761), .ZN(n4421) );
  AND2_X1 U6126 ( .A1(n4965), .A2(n6370), .ZN(n4350) );
  NOR2_X1 U6127 ( .A1(n9472), .A2(n4397), .ZN(n4351) );
  INV_X1 U6128 ( .A(n4500), .ZN(n8826) );
  NOR2_X1 U6129 ( .A1(n4568), .A2(n9079), .ZN(n4352) );
  AND2_X1 U6130 ( .A1(n6357), .A2(n6356), .ZN(n4353) );
  AND2_X1 U6131 ( .A1(n9554), .A2(n9560), .ZN(n9244) );
  AND2_X1 U6132 ( .A1(n5829), .A2(n5828), .ZN(n4354) );
  AND2_X1 U6133 ( .A1(n8465), .A2(n5812), .ZN(n4355) );
  AND2_X1 U6134 ( .A1(n7656), .A2(n5747), .ZN(n4356) );
  AND2_X1 U6135 ( .A1(n5305), .A2(n5306), .ZN(n4357) );
  NAND2_X1 U6136 ( .A1(n5396), .A2(n5395), .ZN(n7819) );
  NAND2_X1 U6137 ( .A1(n9768), .A2(n9560), .ZN(n4358) );
  AND2_X1 U6138 ( .A1(n4888), .A2(n9207), .ZN(n4359) );
  INV_X1 U6139 ( .A(n4682), .ZN(n4681) );
  NAND2_X1 U6140 ( .A1(n4687), .A2(n4569), .ZN(n4682) );
  AND2_X1 U6141 ( .A1(n4937), .A2(n6303), .ZN(n4360) );
  AND2_X1 U6142 ( .A1(n5015), .A2(n8407), .ZN(n4361) );
  INV_X1 U6143 ( .A(n4933), .ZN(n4932) );
  NAND2_X1 U6144 ( .A1(n8886), .A2(n4934), .ZN(n4933) );
  NAND2_X1 U6145 ( .A1(n9126), .A2(n9245), .ZN(n4362) );
  INV_X1 U6146 ( .A(n4684), .ZN(n4683) );
  NAND2_X1 U6147 ( .A1(n4687), .A2(n4405), .ZN(n4684) );
  INV_X1 U6148 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6134) );
  AND2_X1 U6149 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .ZN(n4363) );
  INV_X1 U6150 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4417) );
  CLKBUF_X3 U6151 ( .A(n4807), .Z(n4410) );
  NAND2_X1 U6152 ( .A1(n7657), .A2(n4272), .ZN(n4624) );
  NAND2_X1 U6153 ( .A1(n4620), .A2(n4625), .ZN(n7749) );
  NAND2_X1 U6154 ( .A1(n7324), .A2(n9194), .ZN(n7236) );
  INV_X1 U6155 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4413) );
  AND2_X1 U6156 ( .A1(n7942), .A2(n5007), .ZN(n4364) );
  NAND2_X1 U6157 ( .A1(n5909), .A2(n5908), .ZN(n7655) );
  NAND2_X1 U6158 ( .A1(n6184), .A2(n6181), .ZN(n4365) );
  NAND2_X1 U6159 ( .A1(n4704), .A2(n4703), .ZN(n7519) );
  AND2_X1 U6160 ( .A1(n7654), .A2(n4977), .ZN(n4366) );
  AND2_X1 U6161 ( .A1(n6286), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n4367) );
  INV_X1 U6162 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5270) );
  INV_X1 U6163 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U6164 ( .A1(n4539), .A2(n4542), .ZN(n7733) );
  AND2_X1 U6165 ( .A1(n5756), .A2(n5758), .ZN(n7765) );
  INV_X1 U6166 ( .A(n7765), .ZN(n4623) );
  INV_X1 U6167 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4939) );
  AND2_X1 U6168 ( .A1(n5026), .A2(n5024), .ZN(n5880) );
  INV_X1 U6169 ( .A(n8616), .ZN(n4385) );
  NAND2_X1 U6170 ( .A1(n5783), .A2(n5782), .ZN(n8595) );
  AND2_X1 U6171 ( .A1(n4282), .A2(n6356), .ZN(n4368) );
  INV_X1 U6172 ( .A(n4443), .ZN(n9691) );
  NOR2_X1 U6173 ( .A1(n4501), .A2(n9807), .ZN(n4443) );
  INV_X1 U6174 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5196) );
  OR2_X1 U6175 ( .A1(n7360), .A2(n4871), .ZN(n4369) );
  INV_X1 U6176 ( .A(n9207), .ZN(n4895) );
  AND2_X1 U6177 ( .A1(n7603), .A2(n9175), .ZN(n4370) );
  AND2_X1 U6178 ( .A1(n7655), .A2(n5910), .ZN(n4371) );
  INV_X1 U6179 ( .A(n4569), .ZN(n4405) );
  AND4_X1 U6180 ( .A1(n5381), .A2(n5380), .A3(n5379), .A4(n5378), .ZN(n7816)
         );
  INV_X1 U6181 ( .A(n7816), .ZN(n4626) );
  NAND2_X1 U6182 ( .A1(n6187), .A2(n6186), .ZN(n9673) );
  INV_X1 U6183 ( .A(n9673), .ZN(n4442) );
  NAND2_X1 U6184 ( .A1(n4971), .A2(n4972), .ZN(n7110) );
  AND2_X1 U6185 ( .A1(n9056), .A2(n4829), .ZN(n4372) );
  NAND2_X1 U6186 ( .A1(n4985), .A2(n7122), .ZN(n7154) );
  AND4_X1 U6187 ( .A1(n9276), .A2(n6584), .A3(n9440), .A4(n6583), .ZN(n4373)
         );
  OR2_X1 U6188 ( .A1(n7640), .A2(n9349), .ZN(n4374) );
  INV_X1 U6189 ( .A(n8733), .ZN(n4969) );
  INV_X1 U6190 ( .A(n9078), .ZN(n4690) );
  AND2_X1 U6191 ( .A1(n9444), .A2(n4372), .ZN(n4375) );
  OR2_X1 U6192 ( .A1(n7530), .A2(n8761), .ZN(n7528) );
  AND3_X1 U6193 ( .A1(n5479), .A2(n5478), .A3(n5477), .ZN(n8604) );
  INV_X1 U6194 ( .A(n8604), .ZN(n5915) );
  AND2_X1 U6195 ( .A1(n4559), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4376) );
  INV_X1 U6196 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n4418) );
  NAND2_X1 U6197 ( .A1(n6308), .A2(n6216), .ZN(n9440) );
  AND2_X1 U6198 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4377) );
  INV_X1 U6199 ( .A(SI_30_), .ZN(n4824) );
  INV_X1 U6200 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n4669) );
  INV_X1 U6201 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4485) );
  INV_X1 U6202 ( .A(n9160), .ZN(n4569) );
  NAND2_X1 U6203 ( .A1(n8470), .A2(n5813), .ZN(n8456) );
  NAND2_X1 U6204 ( .A1(n5249), .A2(n5894), .ZN(n7533) );
  AOI21_X1 U6205 ( .B1(n8411), .B2(n5829), .A(n5679), .ZN(n5707) );
  OR2_X1 U6206 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  XNOR2_X2 U6207 ( .A(n5202), .B(n5201), .ZN(n7936) );
  NAND2_X1 U6208 ( .A1(n4852), .A2(n4851), .ZN(n8466) );
  NAND2_X1 U6209 ( .A1(n8456), .A2(n8455), .ZN(n8454) );
  NAND2_X1 U6210 ( .A1(n7693), .A2(n5751), .ZN(n7766) );
  NAND2_X1 U6211 ( .A1(n5464), .A2(n5463), .ZN(n7880) );
  NAND2_X1 U6212 ( .A1(n4378), .A2(n5779), .ZN(n8588) );
  NAND2_X2 U6213 ( .A1(n5890), .A2(n6777), .ZN(n6779) );
  NAND2_X1 U6214 ( .A1(n7897), .A2(n4855), .ZN(n4378) );
  AOI21_X1 U6215 ( .B1(n9497), .B2(n9499), .A(n5040), .ZN(n9484) );
  NAND2_X1 U6216 ( .A1(n5072), .A2(n5071), .ZN(n5330) );
  AOI21_X2 U6217 ( .B1(n6373), .B2(n6372), .A(n6371), .ZN(n9512) );
  NAND2_X1 U6218 ( .A1(n5094), .A2(n5093), .ZN(n5424) );
  NOR2_X1 U6219 ( .A1(n9455), .A2(n9459), .ZN(n9454) );
  NAND3_X1 U6220 ( .A1(n9737), .A2(n9738), .A3(n4379), .ZN(n9831) );
  NAND2_X1 U6221 ( .A1(n5276), .A2(n5065), .ZN(n5292) );
  NOR2_X1 U6222 ( .A1(n9454), .A2(n4472), .ZN(n8042) );
  NOR2_X2 U6223 ( .A1(n9640), .A2(n9624), .ZN(n4382) );
  OAI21_X1 U6224 ( .B1(n8033), .B2(n9316), .A(n8032), .ZN(n9455) );
  NAND2_X1 U6225 ( .A1(n4795), .A2(n4522), .ZN(n5383) );
  NAND2_X1 U6226 ( .A1(n4383), .A2(n4404), .ZN(n4403) );
  NAND3_X1 U6227 ( .A1(n4646), .A2(n4495), .A3(n4494), .ZN(n4383) );
  NAND2_X1 U6228 ( .A1(n4393), .A2(n4824), .ZN(n5685) );
  NAND2_X1 U6229 ( .A1(n5330), .A2(n5073), .ZN(n4795) );
  OAI21_X1 U6230 ( .B1(n5383), .B2(n5091), .A(n5090), .ZN(n5094) );
  INV_X1 U6231 ( .A(n4979), .ZN(n4978) );
  NOR2_X2 U6232 ( .A1(n8473), .A2(n8673), .ZN(n8448) );
  NAND2_X1 U6233 ( .A1(n4804), .A2(n4803), .ZN(n5465) );
  NAND2_X1 U6234 ( .A1(n7533), .A2(n5737), .ZN(n6935) );
  NAND2_X1 U6235 ( .A1(n5623), .A2(n8465), .ZN(n8470) );
  OAI21_X1 U6236 ( .B1(n8588), .B2(n4836), .A(n4834), .ZN(n5583) );
  NAND2_X1 U6237 ( .A1(n7898), .A2(n4631), .ZN(n7897) );
  NAND4_X1 U6238 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5232), .ZN(n7034)
         );
  NAND2_X1 U6239 ( .A1(n5584), .A2(n4853), .ZN(n4852) );
  INV_X1 U6240 ( .A(n5674), .ZN(n5250) );
  AND4_X2 U6241 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n7157)
         );
  OAI22_X2 U6242 ( .A1(n7357), .A2(n4877), .B1(n9902), .B2(n9347), .ZN(n7601)
         );
  NAND3_X1 U6243 ( .A1(n8868), .A2(n9005), .A3(n8867), .ZN(n8909) );
  NAND2_X1 U6244 ( .A1(n9006), .A2(n9008), .ZN(n8868) );
  NAND2_X2 U6245 ( .A1(n8043), .A2(n9316), .ZN(n9458) );
  AND2_X2 U6246 ( .A1(n4892), .A2(n4890), .ZN(n9072) );
  NAND2_X1 U6247 ( .A1(n9972), .A2(n9354), .ZN(n4564) );
  NAND2_X1 U6248 ( .A1(n6230), .A2(n9607), .ZN(n9592) );
  INV_X1 U6249 ( .A(n4919), .ZN(n4601) );
  INV_X1 U6250 ( .A(n4710), .ZN(n8875) );
  INV_X1 U6251 ( .A(n4921), .ZN(n4920) );
  NAND2_X1 U6252 ( .A1(n9682), .A2(n9181), .ZN(n9651) );
  INV_X1 U6253 ( .A(n8941), .ZN(n4924) );
  NAND2_X1 U6254 ( .A1(n4396), .A2(n9663), .ZN(n9649) );
  NAND2_X1 U6255 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  INV_X1 U6256 ( .A(n9306), .ZN(n4687) );
  NAND4_X1 U6257 ( .A1(n4575), .A2(n4576), .A3(n4678), .A4(n4387), .ZN(n4574)
         );
  NOR2_X1 U6258 ( .A1(n9306), .A2(n9545), .ZN(n4679) );
  NAND2_X1 U6259 ( .A1(n9157), .A2(n4692), .ZN(n9159) );
  NAND2_X1 U6260 ( .A1(n4573), .A2(n4570), .ZN(n9152) );
  INV_X1 U6261 ( .A(n5587), .ZN(n4497) );
  INV_X1 U6262 ( .A(n4902), .ZN(n4901) );
  NAND2_X1 U6263 ( .A1(n4810), .A2(n4808), .ZN(n5624) );
  INV_X1 U6264 ( .A(n9236), .ZN(n9321) );
  INV_X1 U6265 ( .A(n5680), .ZN(n4393) );
  NAND2_X1 U6266 ( .A1(n5064), .A2(n5063), .ZN(n5276) );
  NOR2_X1 U6267 ( .A1(n5704), .A2(n8398), .ZN(n5835) );
  NAND2_X1 U6268 ( .A1(n5864), .A2(n5833), .ZN(n4731) );
  INV_X1 U6269 ( .A(n5054), .ZN(n5226) );
  NAND2_X1 U6270 ( .A1(n5480), .A2(n5032), .ZN(n5120) );
  NAND2_X1 U6271 ( .A1(n4694), .A2(n4696), .ZN(n5984) );
  INV_X1 U6272 ( .A(n9651), .ZN(n4396) );
  NAND2_X1 U6273 ( .A1(n4398), .A2(n4351), .ZN(P1_U3263) );
  NOR2_X1 U6274 ( .A1(n9739), .A2(n9716), .ZN(n4397) );
  NAND2_X1 U6275 ( .A1(n9473), .A2(n9670), .ZN(n4398) );
  AOI21_X2 U6276 ( .B1(n4481), .B2(n9708), .A(n4399), .ZN(n9738) );
  NAND2_X1 U6277 ( .A1(n4578), .A2(n4476), .ZN(n4892) );
  NAND2_X1 U6278 ( .A1(n4403), .A2(n4402), .ZN(P1_U3240) );
  NAND3_X1 U6279 ( .A1(n4567), .A2(n4691), .A3(n4566), .ZN(n9086) );
  OR2_X1 U6280 ( .A1(n4642), .A2(n4406), .ZN(n9129) );
  INV_X1 U6281 ( .A(n6387), .ZN(n4696) );
  NAND2_X1 U6282 ( .A1(n9159), .A2(n9232), .ZN(n4656) );
  NAND2_X1 U6283 ( .A1(n4657), .A2(n4654), .ZN(n4653) );
  NAND2_X1 U6284 ( .A1(n4925), .A2(n4923), .ZN(n4928) );
  NAND2_X1 U6285 ( .A1(n7825), .A2(n4591), .ZN(n8813) );
  NAND2_X1 U6286 ( .A1(n4359), .A2(n4577), .ZN(n7080) );
  NAND2_X1 U6287 ( .A1(n7080), .A2(n9257), .ZN(n9074) );
  OAI21_X2 U6288 ( .B1(n4660), .B2(n4659), .A(n9154), .ZN(n9157) );
  NAND2_X1 U6289 ( .A1(n9435), .A2(n4780), .ZN(n4482) );
  NOR2_X1 U6290 ( .A1(n6517), .A2(n4349), .ZN(n6621) );
  NOR2_X1 U6291 ( .A1(n6557), .A2(n4346), .ZN(n6602) );
  NOR2_X1 U6292 ( .A1(n6815), .A2(n4771), .ZN(n6817) );
  NAND2_X1 U6293 ( .A1(n9439), .A2(n9913), .ZN(n9435) );
  NAND2_X1 U6294 ( .A1(n4488), .A2(n4487), .ZN(n4486) );
  NAND2_X1 U6295 ( .A1(n4482), .A2(n9164), .ZN(n4779) );
  AND2_X1 U6296 ( .A1(n5895), .A2(n5903), .ZN(n4615) );
  NOR2_X1 U6297 ( .A1(n6769), .A2(n6768), .ZN(n6815) );
  INV_X1 U6298 ( .A(n9636), .ZN(n6364) );
  NAND2_X1 U6299 ( .A1(n4407), .A2(n4948), .ZN(n9605) );
  NAND2_X1 U6300 ( .A1(n9636), .A2(n4949), .ZN(n4407) );
  NAND2_X1 U6301 ( .A1(n6361), .A2(n6360), .ZN(n9636) );
  NOR2_X2 U6302 ( .A1(n9956), .A2(n7092), .ZN(n7008) );
  NAND2_X2 U6303 ( .A1(n4408), .A2(n6008), .ZN(n9956) );
  INV_X1 U6304 ( .A(n4409), .ZN(n4408) );
  OAI21_X1 U6305 ( .B1(n6444), .B2(n6035), .A(n6007), .ZN(n4409) );
  NAND2_X1 U6306 ( .A1(n7313), .A2(n6348), .ZN(n4946) );
  AND2_X4 U6307 ( .A1(n9056), .A2(n6005), .ZN(n9066) );
  NAND2_X1 U6308 ( .A1(n4519), .A2(n4492), .ZN(n5088) );
  AND2_X2 U6309 ( .A1(n4422), .A2(n4421), .ZN(n9526) );
  XNOR2_X1 U6310 ( .A(n5227), .B(n5224), .ZN(n4420) );
  OAI21_X1 U6311 ( .B1(n4964), .B2(n4963), .A(n4358), .ZN(n4962) );
  AOI21_X2 U6312 ( .B1(n7359), .B2(n7354), .A(n7356), .ZN(n7610) );
  NAND3_X1 U6313 ( .A1(n4944), .A2(n4374), .A3(n4947), .ZN(n4940) );
  NOR2_X1 U6314 ( .A1(n4601), .A2(n4600), .ZN(n4599) );
  NAND2_X1 U6315 ( .A1(n4653), .A2(n9280), .ZN(n4494) );
  NAND2_X1 U6316 ( .A1(n4658), .A2(n4405), .ZN(n4657) );
  NAND2_X1 U6317 ( .A1(n6341), .A2(n6340), .ZN(n7061) );
  OAI21_X1 U6318 ( .B1(n4807), .B2(n4413), .A(n4412), .ZN(n5227) );
  INV_X1 U6319 ( .A(n7601), .ZN(n6142) );
  NAND2_X1 U6320 ( .A1(n4462), .A2(n6633), .ZN(n6333) );
  NAND2_X1 U6321 ( .A1(n7054), .A2(n9251), .ZN(n7055) );
  NAND2_X1 U6322 ( .A1(n9288), .A2(n9287), .ZN(n6756) );
  INV_X1 U6323 ( .A(n4416), .ZN(n4415) );
  NAND2_X1 U6324 ( .A1(n5867), .A2(n5868), .ZN(n4430) );
  INV_X1 U6325 ( .A(n5868), .ZN(n4505) );
  INV_X1 U6326 ( .A(n5321), .ZN(n5671) );
  NAND2_X1 U6327 ( .A1(n4798), .A2(n4796), .ZN(n5177) );
  INV_X1 U6328 ( .A(n4436), .ZN(n4706) );
  NOR2_X1 U6329 ( .A1(n5835), .A2(n5834), .ZN(n5864) );
  NAND2_X1 U6330 ( .A1(n5405), .A2(n5404), .ZN(n5443) );
  NAND2_X1 U6331 ( .A1(n6355), .A2(n6356), .ZN(n4959) );
  XNOR2_X1 U6332 ( .A(n4420), .B(n5225), .ZN(n6444) );
  NAND2_X1 U6333 ( .A1(n4426), .A2(n8415), .ZN(n8664) );
  NAND2_X1 U6334 ( .A1(n4427), .A2(n8614), .ZN(n4426) );
  XNOR2_X1 U6335 ( .A(n8411), .B(n5829), .ZN(n4427) );
  NAND3_X1 U6336 ( .A1(n5482), .A2(n5273), .A3(n5184), .ZN(n5481) );
  NAND2_X1 U6337 ( .A1(n7766), .A2(n5756), .ZN(n5382) );
  NAND2_X1 U6338 ( .A1(n7880), .A2(n5769), .ZN(n7898) );
  NAND2_X1 U6339 ( .A1(n4434), .A2(n5722), .ZN(n7693) );
  NAND2_X1 U6340 ( .A1(n7649), .A2(n7689), .ZN(n4434) );
  OAI211_X2 U6341 ( .C1(n6432), .C2(n5691), .A(n5248), .B(n4318), .ZN(n8761)
         );
  INV_X1 U6342 ( .A(n7260), .ZN(n4509) );
  NAND2_X1 U6343 ( .A1(n6594), .A2(n6711), .ZN(n6712) );
  NAND2_X2 U6344 ( .A1(n8813), .A2(n8812), .ZN(n8959) );
  INV_X1 U6345 ( .A(n6070), .ZN(n9058) );
  NAND2_X2 U6346 ( .A1(n5985), .A2(n5984), .ZN(n5987) );
  NAND2_X1 U6347 ( .A1(n4517), .A2(n4518), .ZN(n6373) );
  INV_X1 U6348 ( .A(n6731), .ZN(n6585) );
  OR2_X2 U6349 ( .A1(n8508), .A2(n5923), .ZN(n4639) );
  NAND2_X1 U6350 ( .A1(n4490), .A2(n4441), .ZN(n8771) );
  NOR2_X2 U6351 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6168) );
  NAND2_X1 U6352 ( .A1(n4584), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6391) );
  NOR2_X1 U6353 ( .A1(n6386), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U6354 ( .A1(n4598), .A2(n4599), .ZN(n4597) );
  NAND2_X1 U6355 ( .A1(n5292), .A2(n4512), .ZN(n4511) );
  NAND2_X1 U6356 ( .A1(n4509), .A2(n4508), .ZN(n7407) );
  XNOR2_X1 U6357 ( .A(n6795), .B(n6793), .ZN(n6791) );
  NAND2_X2 U6358 ( .A1(n4447), .A2(n8975), .ZN(n8834) );
  NAND3_X1 U6359 ( .A1(n4705), .A2(n4707), .A3(n4706), .ZN(n4447) );
  NAND2_X1 U6360 ( .A1(n4474), .A2(n7255), .ZN(n7260) );
  NAND2_X1 U6361 ( .A1(n4722), .A2(n4720), .ZN(n4925) );
  NAND3_X1 U6362 ( .A1(n9073), .A2(n7287), .A3(n7078), .ZN(n6346) );
  NOR2_X1 U6363 ( .A1(n10283), .A2(n10282), .ZN(n10281) );
  NAND2_X1 U6364 ( .A1(n6112), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U6365 ( .A1(n4609), .A2(n4605), .ZN(n4604) );
  AND2_X2 U6366 ( .A1(n4475), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6150) );
  NAND3_X1 U6367 ( .A1(n4698), .A2(n4697), .A3(n4912), .ZN(n7824) );
  NAND3_X1 U6368 ( .A1(n5945), .A2(n4510), .A3(n7932), .ZN(n8665) );
  NAND2_X1 U6369 ( .A1(n9581), .A2(n4350), .ZN(n4517) );
  NAND2_X1 U6370 ( .A1(n4894), .A2(n9206), .ZN(n9073) );
  NAND2_X1 U6371 ( .A1(n7609), .A2(n6354), .ZN(n7794) );
  INV_X1 U6372 ( .A(n5386), .ZN(n5091) );
  NAND2_X1 U6373 ( .A1(n5244), .A2(n5057), .ZN(n5060) );
  NAND2_X1 U6374 ( .A1(n5055), .A2(n5056), .ZN(n5244) );
  INV_X1 U6375 ( .A(n4962), .ZN(n4518) );
  NAND2_X1 U6376 ( .A1(n4465), .A2(n4463), .ZN(n8696) );
  AND2_X1 U6377 ( .A1(n8533), .A2(n8534), .ZN(n4466) );
  INV_X1 U6378 ( .A(n8260), .ZN(n5897) );
  NOR2_X1 U6379 ( .A1(n4292), .A2(n9557), .ZN(n4879) );
  INV_X2 U6380 ( .A(n7308), .ZN(n8258) );
  NAND3_X2 U6381 ( .A1(n5228), .A2(n4309), .A3(n4469), .ZN(n7580) );
  OR2_X2 U6382 ( .A1(n5691), .A2(n4413), .ZN(n4469) );
  INV_X1 U6383 ( .A(n5847), .ZN(n4849) );
  NAND2_X1 U6384 ( .A1(n6779), .A2(n5889), .ZN(n7531) );
  NAND2_X1 U6385 ( .A1(n4830), .A2(n4832), .ZN(n8800) );
  NAND2_X4 U6386 ( .A1(n5884), .A2(n8800), .ZN(n6650) );
  NAND2_X1 U6387 ( .A1(n9247), .A2(n4959), .ZN(n4958) );
  NOR2_X1 U6388 ( .A1(n4956), .A2(n4954), .ZN(n4952) );
  INV_X1 U6389 ( .A(n5424), .ZN(n4805) );
  NAND2_X1 U6390 ( .A1(n4805), .A2(n5099), .ZN(n5405) );
  NAND3_X1 U6391 ( .A1(n6171), .A2(n6170), .A3(n6169), .ZN(n6173) );
  AND4_X2 U6392 ( .A1(n5970), .A2(n5967), .A3(n5969), .A4(n5968), .ZN(n6171)
         );
  NAND4_X1 U6393 ( .A1(n4715), .A2(n4929), .A3(n6796), .A4(n4713), .ZN(n4474)
         );
  NAND2_X1 U6394 ( .A1(n6317), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8037) );
  NOR2_X2 U6395 ( .A1(n6124), .A2(n6820), .ZN(n4475) );
  NAND2_X1 U6396 ( .A1(n4588), .A2(n4587), .ZN(n4710) );
  AOI21_X2 U6397 ( .B1(n9231), .B2(n9230), .A(n9229), .ZN(n9318) );
  INV_X1 U6398 ( .A(n9279), .ZN(n4648) );
  NOR2_X2 U6399 ( .A1(n6110), .A2(n6109), .ZN(n6112) );
  AND2_X2 U6400 ( .A1(n7055), .A2(n9291), .ZN(n4578) );
  NAND2_X2 U6401 ( .A1(n9072), .A2(n9255), .ZN(n7324) );
  AND4_X2 U6402 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5220), .ZN(n6688)
         );
  NAND2_X1 U6403 ( .A1(n9460), .A2(n9461), .ZN(n4481) );
  NAND3_X2 U6404 ( .A1(n6385), .A2(n6169), .A3(n4641), .ZN(n5980) );
  INV_X1 U6405 ( .A(n4486), .ZN(n9376) );
  NAND2_X1 U6406 ( .A1(n9396), .A2(n4789), .ZN(n4787) );
  NOR2_X1 U6407 ( .A1(n6766), .A2(n4772), .ZN(n6769) );
  AOI21_X1 U6408 ( .B1(n6519), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6619), .ZN(
        n6559) );
  XNOR2_X2 U6409 ( .A(n6006), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6518) );
  INV_X1 U6410 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4791) );
  NAND2_X1 U6411 ( .A1(n4795), .A2(n5075), .ZN(n5340) );
  NAND2_X1 U6412 ( .A1(n4970), .A2(n4969), .ZN(n7901) );
  NAND2_X1 U6413 ( .A1(n8615), .A2(n8621), .ZN(n8616) );
  NAND2_X1 U6414 ( .A1(n4891), .A2(n9206), .ZN(n4890) );
  NAND2_X1 U6415 ( .A1(n4666), .A2(n4664), .ZN(n4663) );
  OAI21_X2 U6416 ( .B1(n7518), .B2(n4916), .A(n7718), .ZN(n4915) );
  INV_X1 U6417 ( .A(n5481), .ZN(n5026) );
  NAND2_X1 U6418 ( .A1(n4639), .A2(n4636), .ZN(n8493) );
  NAND2_X1 U6419 ( .A1(n4629), .A2(n4628), .ZN(n8574) );
  NAND2_X1 U6420 ( .A1(n5932), .A2(n5936), .ZN(n8408) );
  NAND2_X1 U6421 ( .A1(n6602), .A2(n6603), .ZN(n6601) );
  NOR2_X1 U6422 ( .A1(n6549), .A2(n6550), .ZN(n6766) );
  OAI21_X2 U6423 ( .B1(n5499), .B2(n4820), .A(n4818), .ZN(n5541) );
  NOR2_X1 U6424 ( .A1(n6621), .A2(n6620), .ZN(n6619) );
  AND2_X2 U6425 ( .A1(n7008), .A2(n6755), .ZN(n7050) );
  OAI21_X1 U6426 ( .B1(n5999), .B2(n5993), .A(P1_IR_REG_27__SCAN_IN), .ZN(
        n4709) );
  INV_X1 U6427 ( .A(n5088), .ZN(n5085) );
  NAND2_X1 U6428 ( .A1(n6005), .A2(n4493), .ZN(n4492) );
  NAND2_X1 U6429 ( .A1(n9156), .A2(n9235), .ZN(n4658) );
  NAND2_X1 U6430 ( .A1(n9153), .A2(n4693), .ZN(n4659) );
  NAND2_X1 U6431 ( .A1(n4904), .A2(n4321), .ZN(n4902) );
  AOI21_X1 U6432 ( .B1(n9458), .B2(n9457), .A(n9459), .ZN(n4516) );
  INV_X1 U6433 ( .A(n4516), .ZN(n9460) );
  NAND2_X1 U6434 ( .A1(n9014), .A2(n4336), .ZN(n4917) );
  NAND2_X1 U6435 ( .A1(n8909), .A2(n8911), .ZN(n4589) );
  NAND2_X1 U6436 ( .A1(n4500), .A2(n8804), .ZN(n4580) );
  NAND3_X1 U6437 ( .A1(n7825), .A2(n4590), .A3(n4591), .ZN(n4500) );
  NAND2_X1 U6438 ( .A1(n4506), .A2(n4503), .ZN(n4770) );
  OAI22_X1 U6439 ( .A1(n5721), .A2(n5720), .B1(n5719), .B2(n8012), .ZN(n4506)
         );
  NAND2_X1 U6440 ( .A1(n9518), .A2(n9501), .ZN(n9503) );
  INV_X1 U6441 ( .A(n4507), .ZN(n9465) );
  INV_X1 U6442 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4786) );
  NAND2_X1 U6443 ( .A1(n4778), .A2(n9440), .ZN(n4777) );
  INV_X1 U6444 ( .A(n8983), .ZN(n4588) );
  NAND2_X1 U6445 ( .A1(n4589), .A2(n8908), .ZN(n8983) );
  NAND2_X1 U6446 ( .A1(n6393), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6389) );
  OAI22_X1 U6447 ( .A1(n8832), .A2(n6633), .B1(n6725), .B2(n6716), .ZN(n6714)
         );
  OAI22_X1 U6448 ( .A1(n8832), .A2(n6335), .B1(n6725), .B2(n6755), .ZN(n6720)
         );
  XNOR2_X1 U6449 ( .A(n6723), .B(n6721), .ZN(n6749) );
  NAND2_X1 U6450 ( .A1(n6719), .A2(n6718), .ZN(n6748) );
  NAND3_X1 U6451 ( .A1(n5272), .A2(n5449), .A3(n10129), .ZN(n5182) );
  NAND2_X1 U6452 ( .A1(n4907), .A2(n4362), .ZN(n4904) );
  NAND2_X1 U6453 ( .A1(n4511), .A2(n5069), .ZN(n5072) );
  NAND3_X2 U6454 ( .A1(n9898), .A2(n8394), .A3(n4793), .ZN(n4792) );
  NAND2_X1 U6455 ( .A1(n5085), .A2(SI_9_), .ZN(n5352) );
  NAND2_X2 U6456 ( .A1(n6142), .A2(n6141), .ZN(n7603) );
  INV_X1 U6457 ( .A(n9251), .ZN(n6338) );
  NAND2_X1 U6458 ( .A1(n4696), .A2(n4640), .ZN(n5994) );
  NAND2_X1 U6459 ( .A1(n5556), .A2(n5555), .ZN(n4794) );
  XNOR2_X1 U6460 ( .A(n8042), .B(n9273), .ZN(n9734) );
  NAND2_X1 U6461 ( .A1(n4528), .A2(n4530), .ZN(n7960) );
  NAND2_X1 U6462 ( .A1(n7910), .A2(n4532), .ZN(n4528) );
  NAND2_X1 U6463 ( .A1(n7452), .A2(n4540), .ZN(n4538) );
  INV_X1 U6464 ( .A(n7459), .ZN(n4549) );
  NAND2_X1 U6465 ( .A1(n4552), .A2(n7183), .ZN(n4551) );
  NAND2_X1 U6466 ( .A1(n4558), .A2(n4363), .ZN(n5323) );
  NAND2_X1 U6467 ( .A1(n5532), .A2(n4376), .ZN(n5602) );
  OAI21_X1 U6468 ( .B1(n5936), .B2(n4560), .A(n5839), .ZN(n5822) );
  NOR2_X1 U6469 ( .A1(n4889), .A2(n4563), .ZN(n9293) );
  NAND3_X1 U6470 ( .A1(n9208), .A2(n9207), .A3(n4564), .ZN(n9209) );
  NAND2_X1 U6471 ( .A1(n4896), .A2(n4564), .ZN(n7282) );
  NAND3_X1 U6472 ( .A1(n4691), .A2(n4567), .A3(n4352), .ZN(n4565) );
  NAND2_X1 U6473 ( .A1(n4565), .A2(n4688), .ZN(n9084) );
  NAND3_X1 U6474 ( .A1(n4574), .A2(n9511), .A3(n9145), .ZN(n4573) );
  NAND3_X1 U6475 ( .A1(n4897), .A2(n4578), .A3(n9205), .ZN(n4577) );
  NAND3_X1 U6476 ( .A1(n4580), .A2(n8959), .A3(n8960), .ZN(n9039) );
  NAND2_X4 U6477 ( .A1(n6731), .A2(n6586), .ZN(n6725) );
  NAND2_X1 U6478 ( .A1(n7561), .A2(n4582), .ZN(n7395) );
  NAND2_X1 U6479 ( .A1(n7292), .A2(n4582), .ZN(n7257) );
  NAND2_X1 U6480 ( .A1(n7414), .A2(n4582), .ZN(n7416) );
  NAND2_X1 U6481 ( .A1(n7640), .A2(n4582), .ZN(n7489) );
  NAND2_X1 U6482 ( .A1(n9824), .A2(n4582), .ZN(n7664) );
  NAND2_X1 U6483 ( .A1(n6327), .A2(n4582), .ZN(n7496) );
  NAND2_X1 U6484 ( .A1(n9807), .A2(n4582), .ZN(n8819) );
  NAND2_X1 U6485 ( .A1(n9818), .A2(n4582), .ZN(n7724) );
  NAND2_X1 U6486 ( .A1(n9673), .A2(n4582), .ZN(n8806) );
  NAND2_X1 U6487 ( .A1(n4411), .A2(n4582), .ZN(n7827) );
  NAND2_X1 U6488 ( .A1(n9642), .A2(n4582), .ZN(n8815) );
  AOI21_X1 U6489 ( .B1(n9624), .B2(n4582), .A(n4581), .ZN(n8831) );
  NAND2_X1 U6490 ( .A1(n9785), .A2(n4582), .ZN(n8841) );
  NAND2_X1 U6491 ( .A1(n9587), .A2(n4582), .ZN(n8836) );
  NAND2_X1 U6492 ( .A1(n9571), .A2(n4582), .ZN(n8851) );
  NAND2_X1 U6493 ( .A1(n9761), .A2(n4582), .ZN(n8862) );
  NAND2_X1 U6494 ( .A1(n9742), .A2(n4582), .ZN(n8879) );
  NAND2_X1 U6495 ( .A1(n9758), .A2(n4582), .ZN(n8870) );
  AOI22_X1 U6496 ( .A1(n9463), .A2(n8883), .B1(n4582), .B2(n9474), .ZN(n8891)
         );
  AOI22_X1 U6497 ( .A1(n8883), .A2(n8051), .B1(n9736), .B2(n4582), .ZN(n8929)
         );
  INV_X4 U6498 ( .A(n6725), .ZN(n4582) );
  NAND2_X1 U6499 ( .A1(n6395), .A2(n6394), .ZN(n4584) );
  NAND2_X1 U6500 ( .A1(n4583), .A2(n4585), .ZN(n6393) );
  NAND2_X1 U6501 ( .A1(n4592), .A2(n7822), .ZN(n4591) );
  NAND4_X1 U6502 ( .A1(n4698), .A2(n4697), .A3(n4912), .A4(n4593), .ZN(n4592)
         );
  NAND2_X1 U6503 ( .A1(n4595), .A2(n4594), .ZN(n6388) );
  NAND2_X1 U6504 ( .A1(n4917), .A2(n4597), .ZN(n9006) );
  NAND2_X1 U6505 ( .A1(n4612), .A2(n4603), .ZN(P1_U3218) );
  NOR2_X1 U6506 ( .A1(n4606), .A2(n4604), .ZN(n4603) );
  NAND2_X1 U6507 ( .A1(n4611), .A2(n4933), .ZN(n4605) );
  INV_X2 U6508 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5272) );
  NAND3_X1 U6509 ( .A1(n4615), .A2(n6932), .A3(n4274), .ZN(n4613) );
  OAI211_X1 U6510 ( .C1(n5902), .C2(n4616), .A(n4613), .B(n5904), .ZN(n7545)
         );
  NAND2_X1 U6511 ( .A1(n5902), .A2(n4614), .ZN(n7437) );
  NAND3_X1 U6512 ( .A1(n6932), .A2(n4274), .A3(n5895), .ZN(n4614) );
  NAND3_X1 U6513 ( .A1(n7657), .A2(n4617), .A3(n4272), .ZN(n4619) );
  AND2_X1 U6514 ( .A1(n5022), .A2(n4623), .ZN(n4622) );
  NAND2_X1 U6515 ( .A1(n4624), .A2(n4622), .ZN(n4620) );
  INV_X1 U6516 ( .A(n7657), .ZN(n5909) );
  NAND2_X1 U6517 ( .A1(n7896), .A2(n4279), .ZN(n4629) );
  NAND2_X1 U6518 ( .A1(n7896), .A2(n5916), .ZN(n4634) );
  NAND2_X2 U6519 ( .A1(n5943), .A2(n5891), .ZN(n5889) );
  AND2_X2 U6520 ( .A1(n5976), .A2(n5977), .ZN(n6169) );
  OAI21_X1 U6521 ( .B1(n4645), .B2(n4644), .A(n9245), .ZN(n4643) );
  AOI211_X2 U6522 ( .C1(n4651), .C2(n9280), .A(n4648), .B(n4647), .ZN(n4646)
         );
  NAND3_X1 U6523 ( .A1(n9107), .A2(n9106), .A3(n9684), .ZN(n4665) );
  AND4_X2 U6524 ( .A1(n6010), .A2(n6011), .A3(n6012), .A4(n4667), .ZN(n6335)
         );
  INV_X2 U6525 ( .A(n5987), .ZN(n4670) );
  OAI21_X2 U6526 ( .B1(n6756), .B2(n9249), .A(n9290), .ZN(n7054) );
  NAND2_X2 U6527 ( .A1(n9286), .A2(n9290), .ZN(n9249) );
  INV_X1 U6528 ( .A(n5986), .ZN(n9854) );
  NAND2_X1 U6529 ( .A1(n4673), .A2(n9637), .ZN(n9119) );
  NAND2_X1 U6530 ( .A1(n6791), .A2(n4931), .ZN(n4929) );
  NAND2_X1 U6531 ( .A1(n7510), .A2(n4699), .ZN(n4697) );
  NAND2_X1 U6532 ( .A1(n7494), .A2(n4701), .ZN(n4698) );
  NAND2_X1 U6533 ( .A1(n8964), .A2(n8828), .ZN(n4705) );
  NAND2_X1 U6534 ( .A1(n7260), .A2(n7259), .ZN(n7403) );
  NAND2_X1 U6535 ( .A1(n8834), .A2(n4723), .ZN(n4722) );
  NAND4_X2 U6536 ( .A1(n6002), .A2(n6004), .A3(n6003), .A4(n4726), .ZN(n6009)
         );
  NAND3_X1 U6537 ( .A1(n9854), .A2(P1_REG3_REG_1__SCAN_IN), .A3(n4670), .ZN(
        n4726) );
  INV_X2 U6538 ( .A(n6009), .ZN(n6633) );
  NAND2_X1 U6539 ( .A1(n4733), .A2(n4730), .ZN(n4729) );
  NAND2_X1 U6540 ( .A1(n4734), .A2(n4354), .ZN(n4733) );
  NAND2_X1 U6541 ( .A1(n4736), .A2(n4735), .ZN(n4734) );
  INV_X1 U6542 ( .A(n5825), .ZN(n4735) );
  NAND2_X1 U6543 ( .A1(n5827), .A2(n5826), .ZN(n4736) );
  NAND2_X1 U6544 ( .A1(n4741), .A2(n4742), .ZN(n5794) );
  NAND2_X1 U6545 ( .A1(n5789), .A2(n4745), .ZN(n4741) );
  NAND2_X1 U6546 ( .A1(n5744), .A2(n4754), .ZN(n4753) );
  OR2_X1 U6547 ( .A1(n5745), .A2(n5839), .ZN(n4754) );
  OAI21_X1 U6548 ( .B1(n5764), .B2(n4760), .A(n4758), .ZN(n5777) );
  NAND2_X1 U6549 ( .A1(n7862), .A2(n5839), .ZN(n4767) );
  NAND2_X1 U6550 ( .A1(n4770), .A2(n5871), .ZN(n5888) );
  NAND4_X1 U6551 ( .A1(n5184), .A2(n5482), .A3(n5273), .A4(n5196), .ZN(n5502)
         );
  NAND3_X1 U6552 ( .A1(n4779), .A2(n4777), .A3(n4774), .ZN(P1_U3260) );
  XNOR2_X2 U6553 ( .A(n6021), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6519) );
  NAND2_X4 U6554 ( .A1(n4792), .A2(n4790), .ZN(n5067) );
  NAND3_X1 U6555 ( .A1(n4791), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4790) );
  INV_X2 U6556 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U6557 ( .A1(n5167), .A2(n4799), .ZN(n4798) );
  NAND2_X1 U6558 ( .A1(n5424), .A2(n5106), .ZN(n4804) );
  MUX2_X1 U6559 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6005), .Z(n5074) );
  MUX2_X1 U6560 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n6005), .Z(n5092) );
  MUX2_X1 U6561 ( .A(n6481), .B(n10183), .S(n6005), .Z(n5107) );
  MUX2_X1 U6562 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n6005), .Z(n5122) );
  NAND2_X1 U6563 ( .A1(n5587), .A2(n4811), .ZN(n4810) );
  NAND2_X1 U6564 ( .A1(n5663), .A2(n4826), .ZN(n4825) );
  OR2_X1 U6565 ( .A1(n5193), .A2(n5191), .ZN(n4830) );
  XNOR2_X2 U6566 ( .A(n4831), .B(n5192), .ZN(n5884) );
  NAND2_X1 U6567 ( .A1(n5193), .A2(n5191), .ZN(n4832) );
  NAND2_X1 U6568 ( .A1(n8434), .A2(n5820), .ZN(n8440) );
  NAND2_X1 U6569 ( .A1(n8440), .A2(n5824), .ZN(n5937) );
  NAND2_X1 U6570 ( .A1(n4850), .A2(n5733), .ZN(n5299) );
  NAND2_X1 U6571 ( .A1(n4854), .A2(n4356), .ZN(n7649) );
  INV_X1 U6572 ( .A(n5778), .ZN(n4857) );
  NAND2_X1 U6573 ( .A1(n7860), .A2(n5441), .ZN(n5464) );
  OR2_X2 U6574 ( .A1(n9465), .A2(n4867), .ZN(n9449) );
  INV_X1 U6575 ( .A(n4868), .ZN(n9709) );
  NAND2_X1 U6576 ( .A1(n9649), .A2(n9199), .ZN(n9612) );
  NAND2_X1 U6577 ( .A1(n9458), .A2(n4879), .ZN(n4878) );
  OAI211_X1 U6578 ( .C1(n9458), .C2(n4880), .A(n4878), .B(n8052), .ZN(n9728)
         );
  NAND2_X1 U6579 ( .A1(n9458), .A2(n5039), .ZN(n9461) );
  NAND2_X1 U6580 ( .A1(n4578), .A2(n4897), .ZN(n4896) );
  OAI21_X2 U6581 ( .B1(n7603), .B2(n4910), .A(n4908), .ZN(n9683) );
  NAND2_X1 U6582 ( .A1(n6385), .A2(n6169), .ZN(n6386) );
  NAND2_X1 U6583 ( .A1(n4930), .A2(n6724), .ZN(n6792) );
  INV_X1 U6584 ( .A(n6724), .ZN(n4931) );
  NAND2_X1 U6585 ( .A1(n6192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4936) );
  OAI21_X1 U6586 ( .B1(n6192), .B2(n4938), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6304) );
  NAND2_X1 U6587 ( .A1(n4936), .A2(n4360), .ZN(n6311) );
  NAND2_X1 U6588 ( .A1(n4940), .A2(n6352), .ZN(n7333) );
  NAND2_X1 U6589 ( .A1(n7076), .A2(n6344), .ZN(n4947) );
  CLKBUF_X1 U6590 ( .A(n4947), .Z(n4941) );
  NOR2_X2 U6591 ( .A1(n7901), .A2(n8728), .ZN(n8615) );
  NOR2_X2 U6592 ( .A1(n7843), .A2(n8737), .ZN(n4970) );
  CLKBUF_X1 U6593 ( .A(n7529), .Z(n4971) );
  AND3_X2 U6594 ( .A1(n7529), .A2(n4284), .A3(n10051), .ZN(n7554) );
  AND2_X1 U6595 ( .A1(n10043), .A2(n7156), .ZN(n4972) );
  AND2_X2 U6596 ( .A1(n7654), .A2(n4286), .ZN(n7842) );
  NAND2_X1 U6597 ( .A1(n8429), .A2(n4980), .ZN(n8418) );
  NAND2_X1 U6598 ( .A1(n8429), .A2(n8406), .ZN(n8416) );
  INV_X1 U6599 ( .A(n8418), .ZN(n8401) );
  NAND2_X1 U6600 ( .A1(n4981), .A2(n8418), .ZN(n8662) );
  NAND2_X1 U6601 ( .A1(n4982), .A2(n7152), .ZN(n7167) );
  NAND3_X1 U6602 ( .A1(n4983), .A2(n7122), .A3(n4985), .ZN(n4982) );
  INV_X1 U6603 ( .A(n7153), .ZN(n4983) );
  NAND2_X1 U6604 ( .A1(n4984), .A2(n7122), .ZN(n7123) );
  INV_X1 U6605 ( .A(n4985), .ZN(n4984) );
  NAND2_X1 U6606 ( .A1(n4986), .A2(n4987), .ZN(n7035) );
  NAND2_X1 U6607 ( .A1(n5939), .A2(n7018), .ZN(n7027) );
  NAND3_X1 U6608 ( .A1(n5939), .A2(n7268), .A3(n7018), .ZN(n4988) );
  NAND2_X4 U6609 ( .A1(n4988), .A2(n7369), .ZN(n7124) );
  NAND2_X1 U6610 ( .A1(n7808), .A2(n7807), .ZN(n7810) );
  INV_X1 U6611 ( .A(n7997), .ZN(n4990) );
  NAND2_X1 U6612 ( .A1(n4989), .A2(n7997), .ZN(n8116) );
  INV_X1 U6613 ( .A(n7987), .ZN(n5004) );
  NAND2_X1 U6614 ( .A1(n6932), .A2(n5895), .ZN(n5012) );
  NAND2_X1 U6615 ( .A1(n5012), .A2(n7105), .ZN(n7107) );
  NAND2_X1 U6616 ( .A1(n8427), .A2(n8435), .ZN(n8426) );
  NAND2_X1 U6617 ( .A1(n5013), .A2(n4361), .ZN(n8409) );
  NAND2_X1 U6618 ( .A1(n8427), .A2(n5014), .ZN(n5013) );
  NAND2_X1 U6619 ( .A1(n5017), .A2(n5018), .ZN(n5930) );
  NAND2_X1 U6620 ( .A1(n8481), .A2(n5927), .ZN(n5017) );
  NAND2_X1 U6621 ( .A1(n5026), .A2(n5023), .ZN(n5877) );
  NAND2_X1 U6622 ( .A1(n7855), .A2(n4280), .ZN(n5028) );
  INV_X1 U6623 ( .A(n5029), .ZN(n7856) );
  NAND2_X1 U6624 ( .A1(n6383), .A2(n6382), .ZN(n9740) );
  OR2_X1 U6625 ( .A1(n9483), .A2(n9961), .ZN(n6382) );
  NAND2_X1 U6626 ( .A1(n8654), .A2(n8653), .ZN(n8769) );
  NAND2_X1 U6627 ( .A1(n8650), .A2(n8763), .ZN(n8654) );
  NAND2_X1 U6628 ( .A1(n8561), .A2(n8553), .ZN(n8549) );
  NAND2_X1 U6629 ( .A1(n8401), .A2(n8659), .ZN(n8655) );
  NAND2_X1 U6630 ( .A1(n8665), .A2(n10076), .ZN(n5966) );
  CLKBUF_X1 U6631 ( .A(n6009), .Z(n9357) );
  CLKBUF_X1 U6632 ( .A(n9636), .Z(n9638) );
  NAND2_X1 U6633 ( .A1(n7924), .A2(n10066), .ZN(n5945) );
  NAND2_X1 U6634 ( .A1(n6304), .A2(n6214), .ZN(n6308) );
  INV_X1 U6635 ( .A(n5502), .ZN(n5212) );
  INV_X1 U6636 ( .A(n9284), .ZN(n9165) );
  NAND2_X1 U6637 ( .A1(n8084), .A2(n7990), .ZN(n7997) );
  CLKBUF_X1 U6638 ( .A(n5884), .Z(n6658) );
  NAND2_X1 U6639 ( .A1(n5622), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5219) );
  AND2_X1 U6640 ( .A1(n7198), .A2(n7197), .ZN(n5030) );
  INV_X1 U6641 ( .A(n8903), .ZN(n8051) );
  AND2_X1 U6642 ( .A1(n5119), .A2(n5118), .ZN(n5032) );
  OR2_X1 U6643 ( .A1(n8565), .A2(n8203), .ZN(n5034) );
  OR2_X1 U6644 ( .A1(n8553), .A2(n8536), .ZN(n5035) );
  OR2_X1 U6645 ( .A1(n8497), .A2(n5924), .ZN(n5036) );
  OR2_X1 U6646 ( .A1(n9494), .A2(n9500), .ZN(n5037) );
  AND2_X1 U6647 ( .A1(n6009), .A2(n9956), .ZN(n5038) );
  INV_X1 U6648 ( .A(n7630), .ZN(n5871) );
  AND2_X1 U6649 ( .A1(n6314), .A2(n6313), .ZN(n9557) );
  NAND2_X1 U6650 ( .A1(n7842), .A2(n7847), .ZN(n7843) );
  INV_X1 U6651 ( .A(n9170), .ZN(n6202) );
  AND2_X1 U6652 ( .A1(n9501), .A2(n9516), .ZN(n5040) );
  NAND2_X1 U6653 ( .A1(n6595), .A2(n6579), .ZN(n9654) );
  AND2_X1 U6654 ( .A1(n8847), .A2(n8996), .ZN(n5041) );
  INV_X1 U6655 ( .A(n9245), .ZN(n6240) );
  AND2_X1 U6656 ( .A1(n8567), .A2(n8514), .ZN(n5042) );
  AND2_X1 U6657 ( .A1(n5928), .A2(n8468), .ZN(n5043) );
  INV_X1 U6658 ( .A(n8487), .ZN(n5925) );
  INV_X1 U6659 ( .A(n9248), .ZN(n6141) );
  INV_X1 U6660 ( .A(n5729), .ZN(n5730) );
  OAI21_X1 U6661 ( .B1(n5837), .B2(n5731), .A(n6933), .ZN(n5732) );
  NOR2_X1 U6662 ( .A1(n5762), .A2(n5761), .ZN(n5764) );
  NOR2_X1 U6663 ( .A1(n5787), .A2(n5786), .ZN(n5799) );
  AND2_X1 U6664 ( .A1(n8487), .A2(n5807), .ZN(n5808) );
  AND2_X1 U6665 ( .A1(n5843), .A2(n5042), .ZN(n5569) );
  INV_X1 U6666 ( .A(n7656), .ZN(n5908) );
  INV_X1 U6667 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5198) );
  AND2_X1 U6668 ( .A1(n7705), .A2(n7504), .ZN(n7505) );
  INV_X1 U6669 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U6670 ( .B1(n7994), .B2(n8246), .A(n8083), .ZN(n7989) );
  INV_X1 U6671 ( .A(n5616), .ZN(n5614) );
  INV_X1 U6672 ( .A(n6692), .ZN(n7013) );
  NOR3_X1 U6673 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .A3(
        P2_IR_REG_28__SCAN_IN), .ZN(n5199) );
  INV_X1 U6674 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6083) );
  NOR2_X1 U6675 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5995) );
  INV_X1 U6676 ( .A(n9316), .ZN(n6301) );
  INV_X1 U6677 ( .A(n5513), .ZN(n5124) );
  INV_X1 U6678 ( .A(n5329), .ZN(n5073) );
  OR2_X1 U6679 ( .A1(n7190), .A2(n7191), .ZN(n7304) );
  INV_X1 U6680 ( .A(n9057), .ZN(n6282) );
  OR2_X1 U6681 ( .A1(n9468), .A2(n9729), .ZN(n8053) );
  AND2_X1 U6682 ( .A1(n6143), .A2(n9112), .ZN(n9175) );
  INV_X1 U6683 ( .A(n9440), .ZN(n9164) );
  NAND2_X1 U6684 ( .A1(n5685), .A2(n5684), .ZN(n5689) );
  NAND2_X1 U6685 ( .A1(n5127), .A2(n5126), .ZN(n5130) );
  AND2_X1 U6686 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  NAND2_X1 U6687 ( .A1(n5067), .A2(n6440), .ZN(n5045) );
  INV_X1 U6688 ( .A(n7021), .ZN(n7039) );
  INV_X1 U6689 ( .A(n7934), .ZN(n5215) );
  INV_X1 U6690 ( .A(n5647), .ZN(n5669) );
  OR2_X1 U6691 ( .A1(n6952), .A2(n6953), .ZN(n6950) );
  AND2_X1 U6692 ( .A1(n7141), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7208) );
  NOR2_X1 U6693 ( .A1(n8711), .A2(n8568), .ZN(n5918) );
  INV_X1 U6694 ( .A(n8721), .ZN(n8621) );
  AOI21_X1 U6695 ( .B1(n7104), .B2(n4274), .A(n5901), .ZN(n5902) );
  OAI21_X1 U6696 ( .B1(n8651), .B2(n10070), .A(n8657), .ZN(n8652) );
  INV_X1 U6697 ( .A(n10070), .ZN(n8762) );
  OR2_X1 U6698 ( .A1(n5949), .A2(n5946), .ZN(n5947) );
  INV_X1 U6699 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6820) );
  OR2_X1 U6700 ( .A1(n6506), .A2(n6492), .ZN(n9918) );
  AOI21_X1 U6701 ( .B1(n8051), .B2(n9703), .A(n6324), .ZN(n6325) );
  INV_X1 U6702 ( .A(n9576), .ZN(n9582) );
  AND2_X1 U6703 ( .A1(n6202), .A2(n9611), .ZN(n9637) );
  AND2_X1 U6704 ( .A1(n6379), .A2(n9284), .ZN(n6595) );
  NAND2_X1 U6705 ( .A1(n6009), .A2(n6716), .ZN(n9287) );
  OAI21_X1 U6706 ( .B1(n9746), .B2(n9961), .A(n9745), .ZN(n9747) );
  INV_X1 U6707 ( .A(n9998), .ZN(n9957) );
  INV_X1 U6708 ( .A(n10000), .ZN(n10008) );
  NAND2_X1 U6709 ( .A1(n6984), .A2(n6384), .ZN(n9998) );
  INV_X1 U6710 ( .A(n9703), .ZN(n9656) );
  OR3_X1 U6711 ( .A1(n7785), .A2(n7895), .A3(n7836), .ZN(n7042) );
  NAND2_X1 U6712 ( .A1(n7810), .A2(n7809), .ZN(n7910) );
  AND2_X1 U6713 ( .A1(n7155), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8238) );
  NAND2_X1 U6714 ( .A1(n7022), .A2(n8527), .ZN(n8236) );
  INV_X1 U6715 ( .A(n8382), .ZN(n8342) );
  OR2_X1 U6716 ( .A1(n5844), .A2(n8516), .ZN(n8534) );
  AOI21_X1 U6717 ( .B1(n8574), .B2(n5919), .A(n5918), .ZN(n8560) );
  INV_X1 U6718 ( .A(n8605), .ZN(n8582) );
  INV_X1 U6719 ( .A(n7926), .ZN(n8600) );
  NAND2_X1 U6720 ( .A1(n7374), .A2(n8527), .ZN(n8645) );
  AOI21_X1 U6721 ( .B1(n5958), .B2(n10035), .A(n10036), .ZN(n7367) );
  OR2_X1 U6722 ( .A1(n7018), .A2(n7017), .ZN(n10070) );
  INV_X1 U6723 ( .A(n10066), .ZN(n8767) );
  NAND2_X1 U6724 ( .A1(n8610), .A2(n8759), .ZN(n10066) );
  NAND2_X1 U6725 ( .A1(n5947), .A2(n5948), .ZN(n10030) );
  NAND2_X1 U6726 ( .A1(n5874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5876) );
  INV_X1 U6727 ( .A(n9056), .ZN(n6044) );
  AND2_X1 U6728 ( .A1(n9236), .A2(n9063), .ZN(n9280) );
  INV_X1 U6729 ( .A(n4448), .ZN(n6278) );
  OR2_X1 U6730 ( .A1(n6506), .A2(n9329), .ZN(n9438) );
  NAND2_X1 U6731 ( .A1(n9223), .A2(n9311), .ZN(n9499) );
  INV_X1 U6732 ( .A(n9654), .ZN(n9705) );
  INV_X1 U6733 ( .A(n9557), .ZN(n9708) );
  AND2_X1 U6734 ( .A1(n6417), .A2(n9850), .ZN(n6977) );
  INV_X1 U6735 ( .A(n9731), .ZN(n9732) );
  INV_X1 U6736 ( .A(n9961), .ZN(n10010) );
  INV_X1 U6737 ( .A(n6977), .ZN(n6575) );
  INV_X1 U6738 ( .A(n6411), .ZN(n9848) );
  OR2_X1 U6739 ( .A1(n6416), .A2(n6402), .ZN(n6411) );
  INV_X1 U6740 ( .A(n8395), .ZN(n8366) );
  INV_X1 U6741 ( .A(n8681), .ZN(n8486) );
  NAND2_X1 U6742 ( .A1(n7026), .A2(n7025), .ZN(n8230) );
  INV_X1 U6743 ( .A(n8236), .ZN(n8226) );
  INV_X1 U6744 ( .A(n8388), .ZN(n8372) );
  XNOR2_X1 U6745 ( .A(n8447), .B(n8455), .ZN(n8675) );
  OR2_X1 U6746 ( .A1(n4273), .A2(n7370), .ZN(n8597) );
  INV_X2 U6747 ( .A(n10081), .ZN(n10084) );
  INV_X1 U6748 ( .A(n10076), .ZN(n10074) );
  AND2_X1 U6749 ( .A1(n7040), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10037) );
  XNOR2_X1 U6750 ( .A(n5876), .B(n5875), .ZN(n7785) );
  INV_X1 U6751 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10180) );
  INV_X1 U6752 ( .A(n9500), .ZN(n9339) );
  INV_X1 U6753 ( .A(n9098), .ZN(n9685) );
  INV_X1 U6754 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9874) );
  OR2_X1 U6755 ( .A1(n6506), .A2(n6487), .ZN(n9923) );
  OR2_X1 U6756 ( .A1(n10017), .A2(n6418), .ZN(n6419) );
  OR3_X1 U6757 ( .A1(n9801), .A2(n9800), .A3(n9799), .ZN(n9842) );
  INV_X1 U6758 ( .A(n6577), .ZN(n9849) );
  INV_X1 U6759 ( .A(n6379), .ZN(n7301) );
  INV_X1 U6760 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10197) );
  INV_X1 U6761 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6465) );
  NOR2_X1 U6762 ( .A1(n10280), .A2(n10279), .ZN(n10278) );
  NOR2_X1 U6763 ( .A1(n10112), .A2(n10111), .ZN(n10110) );
  AND2_X1 U6764 ( .A1(n6422), .A2(n10037), .ZN(P2_U3966) );
  NAND2_X1 U6765 ( .A1(n5966), .A2(n5965), .ZN(P2_U3516) );
  NAND2_X1 U6766 ( .A1(n6420), .A2(n6419), .ZN(P1_U3518) );
  INV_X1 U6767 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6430) );
  INV_X1 U6768 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6440) );
  INV_X1 U6769 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U6770 ( .A1(n5067), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5046) );
  INV_X1 U6771 ( .A(SI_2_), .ZN(n5243) );
  OAI211_X1 U6772 ( .C1(n5067), .C2(n6432), .A(n5046), .B(n5243), .ZN(n5057)
         );
  NOR2_X1 U6773 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5048) );
  NAND2_X1 U6774 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6775 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5047) );
  OAI21_X1 U6776 ( .B1(n5048), .B2(n5223), .A(n5047), .ZN(n5049) );
  NAND2_X1 U6777 ( .A1(n5067), .A2(n5049), .ZN(n5056) );
  INV_X1 U6778 ( .A(n5067), .ZN(n5054) );
  NOR2_X1 U6779 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5052) );
  AND2_X1 U6780 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5222) );
  INV_X1 U6781 ( .A(n5222), .ZN(n5051) );
  NAND2_X1 U6782 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5050) );
  OAI21_X1 U6783 ( .B1(n5052), .B2(n5051), .A(n5050), .ZN(n5053) );
  NAND2_X1 U6784 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  INV_X1 U6785 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U6786 ( .A1(n5067), .A2(n6447), .ZN(n5058) );
  OAI211_X1 U6787 ( .C1(n5226), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5058), .B(
        SI_2_), .ZN(n5059) );
  NAND2_X1 U6788 ( .A1(n5060), .A2(n5059), .ZN(n5255) );
  NAND2_X1 U6789 ( .A1(n5256), .A2(n5255), .ZN(n5064) );
  INV_X1 U6790 ( .A(n5061), .ZN(n5062) );
  NAND2_X1 U6791 ( .A1(n5062), .A2(SI_3_), .ZN(n5063) );
  XNOR2_X1 U6792 ( .A(n5066), .B(SI_4_), .ZN(n5275) );
  INV_X1 U6793 ( .A(n5275), .ZN(n5065) );
  INV_X4 U6794 ( .A(n5067), .ZN(n6005) );
  NAND2_X1 U6795 ( .A1(n5293), .A2(SI_5_), .ZN(n5311) );
  NAND2_X1 U6796 ( .A1(n5066), .A2(SI_4_), .ZN(n5291) );
  MUX2_X1 U6797 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5067), .Z(n5070) );
  XNOR2_X1 U6798 ( .A(n5070), .B(SI_6_), .ZN(n5313) );
  NOR2_X1 U6799 ( .A1(n5293), .A2(SI_5_), .ZN(n5068) );
  NOR2_X1 U6800 ( .A1(n5313), .A2(n5068), .ZN(n5069) );
  NAND2_X1 U6801 ( .A1(n5070), .A2(SI_6_), .ZN(n5071) );
  NAND2_X1 U6802 ( .A1(n5074), .A2(SI_7_), .ZN(n5075) );
  INV_X1 U6803 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6449) );
  INV_X4 U6804 ( .A(n6005), .ZN(n5245) );
  INV_X1 U6805 ( .A(SI_8_), .ZN(n5076) );
  INV_X1 U6806 ( .A(n5077), .ZN(n5078) );
  NAND2_X1 U6807 ( .A1(n5078), .A2(SI_8_), .ZN(n5079) );
  NAND2_X1 U6808 ( .A1(n5351), .A2(n5079), .ZN(n5339) );
  INV_X1 U6809 ( .A(SI_10_), .ZN(n5081) );
  INV_X1 U6810 ( .A(n5082), .ZN(n5083) );
  NAND2_X1 U6811 ( .A1(n5083), .A2(SI_10_), .ZN(n5084) );
  INV_X1 U6812 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6463) );
  INV_X1 U6813 ( .A(SI_9_), .ZN(n5087) );
  NAND2_X1 U6814 ( .A1(n5088), .A2(n5087), .ZN(n5364) );
  NAND2_X1 U6815 ( .A1(n5351), .A2(n5364), .ZN(n5384) );
  INV_X1 U6816 ( .A(n5388), .ZN(n5089) );
  NAND2_X1 U6817 ( .A1(n5092), .A2(SI_11_), .ZN(n5093) );
  MUX2_X1 U6818 ( .A(n6459), .B(n6457), .S(n5245), .Z(n5096) );
  INV_X1 U6819 ( .A(SI_12_), .ZN(n5095) );
  INV_X1 U6820 ( .A(n5096), .ZN(n5097) );
  NAND2_X1 U6821 ( .A1(n5097), .A2(SI_12_), .ZN(n5098) );
  MUX2_X1 U6822 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5245), .Z(n5100) );
  INV_X1 U6823 ( .A(n5404), .ZN(n5104) );
  INV_X1 U6824 ( .A(n5100), .ZN(n5102) );
  INV_X1 U6825 ( .A(SI_13_), .ZN(n5101) );
  INV_X1 U6826 ( .A(n5107), .ZN(n5108) );
  MUX2_X1 U6827 ( .A(n6478), .B(n10197), .S(n4410), .Z(n5110) );
  INV_X1 U6828 ( .A(SI_15_), .ZN(n5109) );
  INV_X1 U6829 ( .A(n5110), .ZN(n5111) );
  NAND2_X1 U6830 ( .A1(n5111), .A2(SI_15_), .ZN(n5112) );
  OAI21_X2 U6831 ( .B1(n5465), .B2(n5466), .A(n5113), .ZN(n5480) );
  INV_X1 U6832 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5114) );
  MUX2_X1 U6833 ( .A(n5114), .B(n6556), .S(n5245), .Z(n5116) );
  INV_X1 U6834 ( .A(SI_16_), .ZN(n5115) );
  NAND2_X1 U6835 ( .A1(n5116), .A2(n5115), .ZN(n5119) );
  INV_X1 U6836 ( .A(n5116), .ZN(n5117) );
  NAND2_X1 U6837 ( .A1(n5117), .A2(SI_16_), .ZN(n5118) );
  INV_X1 U6838 ( .A(SI_17_), .ZN(n10188) );
  INV_X1 U6839 ( .A(n5498), .ZN(n5121) );
  NAND2_X1 U6840 ( .A1(n5122), .A2(SI_17_), .ZN(n5123) );
  MUX2_X1 U6841 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5245), .Z(n5125) );
  INV_X1 U6842 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6875) );
  MUX2_X1 U6843 ( .A(n10180), .B(n6875), .S(n5226), .Z(n5127) );
  INV_X1 U6844 ( .A(SI_19_), .ZN(n5126) );
  INV_X1 U6845 ( .A(n5127), .ZN(n5128) );
  NAND2_X1 U6846 ( .A1(n5128), .A2(SI_19_), .ZN(n5129) );
  OAI21_X2 U6847 ( .B1(n5541), .B2(n5540), .A(n5130), .ZN(n5556) );
  INV_X1 U6848 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7121) );
  INV_X1 U6849 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7118) );
  MUX2_X1 U6850 ( .A(n7121), .B(n7118), .S(n4410), .Z(n5132) );
  INV_X1 U6851 ( .A(SI_20_), .ZN(n5131) );
  NAND2_X1 U6852 ( .A1(n5132), .A2(n5131), .ZN(n5135) );
  INV_X1 U6853 ( .A(n5132), .ZN(n5133) );
  NAND2_X1 U6854 ( .A1(n5133), .A2(SI_20_), .ZN(n5134) );
  INV_X1 U6855 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7270) );
  INV_X1 U6856 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7220) );
  MUX2_X1 U6857 ( .A(n7270), .B(n7220), .S(n4410), .Z(n5137) );
  INV_X1 U6858 ( .A(n5137), .ZN(n5138) );
  NAND2_X1 U6859 ( .A1(n5138), .A2(SI_21_), .ZN(n5139) );
  INV_X1 U6860 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7300) );
  INV_X1 U6861 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7303) );
  MUX2_X1 U6862 ( .A(n7300), .B(n7303), .S(n5245), .Z(n5141) );
  INV_X1 U6863 ( .A(SI_22_), .ZN(n5140) );
  NAND2_X1 U6864 ( .A1(n5141), .A2(n5140), .ZN(n5144) );
  INV_X1 U6865 ( .A(n5141), .ZN(n5142) );
  NAND2_X1 U6866 ( .A1(n5142), .A2(SI_22_), .ZN(n5143) );
  NAND2_X1 U6867 ( .A1(n5144), .A2(n5143), .ZN(n5570) );
  INV_X1 U6868 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7632) );
  INV_X1 U6869 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5145) );
  MUX2_X1 U6870 ( .A(n7632), .B(n5145), .S(n5245), .Z(n5147) );
  INV_X1 U6871 ( .A(SI_23_), .ZN(n5146) );
  NAND2_X1 U6872 ( .A1(n5147), .A2(n5146), .ZN(n5150) );
  INV_X1 U6873 ( .A(n5147), .ZN(n5148) );
  NAND2_X1 U6874 ( .A1(n5148), .A2(SI_23_), .ZN(n5149) );
  INV_X1 U6875 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7783) );
  INV_X1 U6876 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7759) );
  MUX2_X1 U6877 ( .A(n7783), .B(n7759), .S(n4410), .Z(n5151) );
  XNOR2_X1 U6878 ( .A(n5151), .B(SI_24_), .ZN(n5599) );
  INV_X1 U6879 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6880 ( .A1(n5152), .A2(SI_24_), .ZN(n5153) );
  INV_X1 U6881 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7838) );
  INV_X1 U6882 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5155) );
  MUX2_X1 U6883 ( .A(n7838), .B(n5155), .S(n4410), .Z(n5157) );
  INV_X1 U6884 ( .A(SI_25_), .ZN(n5156) );
  NAND2_X1 U6885 ( .A1(n5157), .A2(n5156), .ZN(n5160) );
  INV_X1 U6886 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U6887 ( .A1(n5158), .A2(SI_25_), .ZN(n5159) );
  NAND2_X1 U6888 ( .A1(n5160), .A2(n5159), .ZN(n5610) );
  INV_X1 U6889 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7893) );
  INV_X1 U6890 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5161) );
  MUX2_X1 U6891 ( .A(n7893), .B(n5161), .S(n4410), .Z(n5163) );
  INV_X1 U6892 ( .A(SI_26_), .ZN(n5162) );
  NAND2_X1 U6893 ( .A1(n5163), .A2(n5162), .ZN(n5166) );
  INV_X1 U6894 ( .A(n5163), .ZN(n5164) );
  NAND2_X1 U6895 ( .A1(n5164), .A2(SI_26_), .ZN(n5165) );
  INV_X1 U6896 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8801) );
  INV_X1 U6897 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5168) );
  MUX2_X1 U6898 ( .A(n8801), .B(n5168), .S(n4410), .Z(n5169) );
  INV_X1 U6899 ( .A(SI_27_), .ZN(n10211) );
  NAND2_X1 U6900 ( .A1(n5169), .A2(n10211), .ZN(n5172) );
  INV_X1 U6901 ( .A(n5169), .ZN(n5170) );
  NAND2_X1 U6902 ( .A1(n5170), .A2(SI_27_), .ZN(n5171) );
  INV_X1 U6903 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8798) );
  INV_X1 U6904 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5173) );
  MUX2_X1 U6905 ( .A(n8798), .B(n5173), .S(n5245), .Z(n5175) );
  XNOR2_X1 U6906 ( .A(n5175), .B(SI_28_), .ZN(n5648) );
  INV_X1 U6907 ( .A(SI_28_), .ZN(n5174) );
  NAND2_X1 U6908 ( .A1(n5175), .A2(n5174), .ZN(n5176) );
  INV_X1 U6909 ( .A(SI_29_), .ZN(n5664) );
  MUX2_X1 U6910 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4807), .Z(n5665) );
  MUX2_X1 U6911 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n5245), .Z(n5681) );
  XNOR2_X1 U6912 ( .A(n5681), .B(SI_30_), .ZN(n5178) );
  AND4_X2 U6914 ( .A1(n5181), .A2(n5180), .A3(n5179), .A4(n5409), .ZN(n5482)
         );
  NOR2_X2 U6915 ( .A1(n5483), .A2(n5182), .ZN(n5184) );
  NOR2_X2 U6916 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5242) );
  AND2_X2 U6917 ( .A1(n5242), .A2(n5183), .ZN(n5273) );
  NOR2_X1 U6918 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5187) );
  NOR2_X1 U6919 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5186) );
  NOR2_X1 U6920 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5185) );
  NAND4_X1 U6921 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5875), .ZN(n5197)
         );
  INV_X1 U6922 ( .A(n5197), .ZN(n5189) );
  NOR3_X1 U6923 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_26__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6924 ( .A1(n5189), .A2(n5188), .ZN(n5190) );
  OAI21_X2 U6925 ( .B1(n5500), .B2(n5190), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5193) );
  INV_X1 U6926 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6927 ( .A1(n9065), .A2(n4276), .ZN(n5195) );
  INV_X1 U6928 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7935) );
  OR2_X1 U6929 ( .A1(n4468), .A2(n7935), .ZN(n5194) );
  INV_X1 U6930 ( .A(n5877), .ZN(n5200) );
  NAND2_X1 U6931 ( .A1(n5200), .A2(n5199), .ZN(n5204) );
  NOR2_X2 U6932 ( .A1(n5204), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5203) );
  INV_X1 U6933 ( .A(n5203), .ZN(n8791) );
  NAND2_X1 U6934 ( .A1(n5204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5205) );
  MUX2_X1 U6935 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5205), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5206) );
  CLKBUF_X3 U6936 ( .A(n5282), .Z(n5695) );
  NAND2_X1 U6937 ( .A1(n5695), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5210) );
  AND2_X2 U6938 ( .A1(n5216), .A2(n7934), .ZN(n5283) );
  NAND2_X1 U6939 ( .A1(n5670), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6940 ( .A1(n7936), .A2(n7934), .ZN(n5214) );
  NAND2_X1 U6941 ( .A1(n5671), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5208) );
  AND3_X1 U6942 ( .A1(n5210), .A2(n5209), .A3(n5208), .ZN(n5703) );
  NAND2_X1 U6943 ( .A1(n5703), .A2(n7028), .ZN(n5711) );
  NAND2_X1 U6944 ( .A1(n5494), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5220) );
  AND2_X4 U6945 ( .A1(n5216), .A2(n5215), .ZN(n5622) );
  NAND2_X1 U6946 ( .A1(n5250), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U6947 ( .A1(n5283), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5217) );
  INV_X1 U6948 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U6949 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5221) );
  XNOR2_X1 U6950 ( .A(n10174), .B(n5221), .ZN(n6663) );
  NAND2_X1 U6951 ( .A1(n9054), .A2(n5222), .ZN(n5235) );
  OAI21_X1 U6952 ( .B1(n5223), .B2(n9054), .A(n5235), .ZN(n5225) );
  INV_X1 U6953 ( .A(SI_1_), .ZN(n5224) );
  OR2_X1 U6954 ( .A1(n5263), .A2(n6444), .ZN(n5228) );
  NAND2_X1 U6955 ( .A1(n5622), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6956 ( .A1(n5494), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6957 ( .A1(n5250), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6958 ( .A1(n5283), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5229) );
  INV_X1 U6959 ( .A(n7034), .ZN(n5237) );
  NAND2_X1 U6960 ( .A1(n6005), .A2(SI_0_), .ZN(n5234) );
  INV_X1 U6961 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6962 ( .A1(n5234), .A2(n5233), .ZN(n5236) );
  AND2_X1 U6963 ( .A1(n5236), .A2(n5235), .ZN(n8803) );
  MUX2_X1 U6964 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8803), .S(n6650), .Z(n7434) );
  INV_X1 U6965 ( .A(n7531), .ZN(n5249) );
  NAND2_X1 U6966 ( .A1(n5622), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6967 ( .A1(n5494), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6968 ( .A1(n5283), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6969 ( .A1(n5282), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5238) );
  INV_X1 U6970 ( .A(n7157), .ZN(n8262) );
  OR2_X1 U6971 ( .A1(n5242), .A2(n5270), .ZN(n5258) );
  INV_X1 U6972 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5257) );
  XNOR2_X1 U6973 ( .A(n5244), .B(n5243), .ZN(n5247) );
  XNOR2_X1 U6974 ( .A(n5247), .B(n5246), .ZN(n6446) );
  NAND2_X1 U6975 ( .A1(n7157), .A2(n8761), .ZN(n5737) );
  NAND2_X1 U6976 ( .A1(n5282), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6977 ( .A1(n5494), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5253) );
  INV_X1 U6978 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U6979 ( .A1(n5622), .A2(n8640), .ZN(n5252) );
  NAND2_X1 U6980 ( .A1(n5283), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5251) );
  AND4_X2 U6981 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n7535)
         );
  XNOR2_X1 U6982 ( .A(n5255), .B(n5256), .ZN(n6439) );
  NAND2_X1 U6983 ( .A1(n5258), .A2(n5257), .ZN(n5259) );
  NAND2_X1 U6984 ( .A1(n5259), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5261) );
  INV_X1 U6985 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5260) );
  XNOR2_X1 U6986 ( .A(n5261), .B(n5260), .ZN(n8286) );
  OR2_X1 U6987 ( .A1(n6650), .A2(n8286), .ZN(n5262) );
  NAND2_X1 U6988 ( .A1(n8261), .A2(n7156), .ZN(n5723) );
  NAND2_X1 U6989 ( .A1(n7470), .A2(n5723), .ZN(n6933) );
  INV_X1 U6990 ( .A(n6933), .ZN(n6936) );
  NAND2_X1 U6991 ( .A1(n5694), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6992 ( .A1(n5282), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5267) );
  OAI21_X1 U6993 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5285), .ZN(n5264) );
  INV_X1 U6994 ( .A(n5264), .ZN(n7479) );
  NAND2_X1 U6995 ( .A1(n5622), .A2(n7479), .ZN(n5266) );
  NAND2_X1 U6996 ( .A1(n5207), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5265) );
  NAND4_X1 U6997 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n8260)
         );
  NOR2_X1 U6998 ( .A1(n5273), .A2(n5270), .ZN(n5269) );
  MUX2_X1 U6999 ( .A(n5270), .B(n5269), .S(P2_IR_REG_4__SCAN_IN), .Z(n5271) );
  INV_X1 U7000 ( .A(n5271), .ZN(n5274) );
  NAND2_X1 U7001 ( .A1(n5273), .A2(n5272), .ZN(n5485) );
  NAND2_X1 U7002 ( .A1(n5274), .A2(n5485), .ZN(n6837) );
  XNOR2_X1 U7003 ( .A(n4269), .B(n5275), .ZN(n6429) );
  NAND2_X1 U7004 ( .A1(n6429), .A2(n5294), .ZN(n5278) );
  OR2_X1 U7005 ( .A1(n5691), .A2(n4515), .ZN(n5277) );
  NAND2_X1 U7006 ( .A1(n5897), .A2(n5279), .ZN(n5727) );
  NAND2_X1 U7007 ( .A1(n8260), .A2(n10043), .ZN(n5729) );
  NAND2_X2 U7008 ( .A1(n5727), .A2(n5729), .ZN(n5896) );
  INV_X1 U7009 ( .A(n7470), .ZN(n5280) );
  NOR2_X1 U7010 ( .A1(n5896), .A2(n5280), .ZN(n5281) );
  NAND2_X1 U7011 ( .A1(n5282), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U7012 ( .A1(n5494), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U7013 ( .A1(n5207), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5288) );
  INV_X1 U7014 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U7015 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  AND2_X1 U7016 ( .A1(n5302), .A2(n5286), .ZN(n7376) );
  NAND2_X1 U7017 ( .A1(n5647), .A2(n7376), .ZN(n5287) );
  XNOR2_X1 U7018 ( .A(n5293), .B(SI_5_), .ZN(n5308) );
  XNOR2_X1 U7019 ( .A(n5310), .B(n5308), .ZN(n6425) );
  NAND2_X1 U7020 ( .A1(n6425), .A2(n4277), .ZN(n5298) );
  INV_X2 U7021 ( .A(n5691), .ZN(n5545) );
  INV_X2 U7022 ( .A(n6650), .ZN(n6472) );
  NAND2_X1 U7023 ( .A1(n5485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5295) );
  MUX2_X1 U7024 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5295), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5296) );
  AND2_X1 U7025 ( .A1(n5296), .A2(n5315), .ZN(n6856) );
  AOI22_X1 U7026 ( .A1(n5545), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6472), .B2(
        n6856), .ZN(n5297) );
  NAND2_X1 U7027 ( .A1(n5695), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U7028 ( .A1(n5694), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5306) );
  INV_X1 U7029 ( .A(n5622), .ZN(n5300) );
  INV_X2 U7030 ( .A(n5300), .ZN(n5647) );
  INV_X1 U7031 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U7032 ( .A1(n5302), .A2(n5301), .ZN(n5303) );
  AND2_X1 U7033 ( .A1(n5323), .A2(n5303), .ZN(n7445) );
  NAND2_X1 U7034 ( .A1(n5647), .A2(n7445), .ZN(n5305) );
  NAND2_X1 U7035 ( .A1(n5207), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5304) );
  INV_X1 U7036 ( .A(n5308), .ZN(n5309) );
  NAND2_X1 U7037 ( .A1(n5310), .A2(n5309), .ZN(n5312) );
  NAND2_X1 U7038 ( .A1(n6433), .A2(n4276), .ZN(n5320) );
  NAND2_X1 U7039 ( .A1(n5315), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5314) );
  MUX2_X1 U7040 ( .A(n5314), .B(P2_IR_REG_31__SCAN_IN), .S(n5316), .Z(n5318)
         );
  INV_X1 U7041 ( .A(n5315), .ZN(n5317) );
  NAND2_X1 U7042 ( .A1(n5317), .A2(n5316), .ZN(n5332) );
  NAND2_X1 U7043 ( .A1(n5318), .A2(n5332), .ZN(n8302) );
  INV_X1 U7044 ( .A(n8302), .ZN(n8299) );
  AOI22_X1 U7045 ( .A1(n5545), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6472), .B2(
        n8299), .ZN(n5319) );
  INV_X1 U7046 ( .A(n7448), .ZN(n10051) );
  NAND2_X1 U7047 ( .A1(n10051), .A2(n8258), .ZN(n5741) );
  NAND2_X1 U7048 ( .A1(n5694), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U7049 ( .A1(n5207), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U7050 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  AND2_X1 U7051 ( .A1(n5345), .A2(n5324), .ZN(n7555) );
  NAND2_X1 U7052 ( .A1(n5647), .A2(n7555), .ZN(n5326) );
  NAND2_X1 U7053 ( .A1(n5695), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5325) );
  XNOR2_X1 U7054 ( .A(n5330), .B(n5329), .ZN(n6427) );
  NAND2_X1 U7055 ( .A1(n6427), .A2(n4276), .ZN(n5337) );
  NAND2_X1 U7056 ( .A1(n5332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5331) );
  MUX2_X1 U7057 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5331), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5335) );
  INV_X1 U7058 ( .A(n5332), .ZN(n5334) );
  NAND2_X1 U7059 ( .A1(n5334), .A2(n5333), .ZN(n5353) );
  AND2_X1 U7060 ( .A1(n5335), .A2(n5353), .ZN(n6891) );
  AOI22_X1 U7061 ( .A1(n5545), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6472), .B2(
        n6891), .ZN(n5336) );
  NAND2_X1 U7062 ( .A1(n5337), .A2(n5336), .ZN(n7558) );
  NAND2_X1 U7063 ( .A1(n7653), .A2(n7558), .ZN(n5746) );
  INV_X1 U7064 ( .A(n7653), .ZN(n8256) );
  NAND2_X1 U7065 ( .A1(n5746), .A2(n5747), .ZN(n5905) );
  INV_X1 U7066 ( .A(n7547), .ZN(n5338) );
  XNOR2_X1 U7067 ( .A(n5339), .B(n5340), .ZN(n6434) );
  NAND2_X1 U7068 ( .A1(n6434), .A2(n4277), .ZN(n5343) );
  NAND2_X1 U7069 ( .A1(n5353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5341) );
  XNOR2_X1 U7070 ( .A(n5341), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8317) );
  AOI22_X1 U7071 ( .A1(n5545), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6472), .B2(
        n8317), .ZN(n5342) );
  NAND2_X1 U7072 ( .A1(n5343), .A2(n5342), .ZN(n7658) );
  NAND2_X1 U7073 ( .A1(n5694), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U7074 ( .A1(n5695), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U7075 ( .A1(n5345), .A2(n5344), .ZN(n5346) );
  NAND2_X1 U7076 ( .A1(n5647), .A2(n4299), .ZN(n5348) );
  NAND2_X1 U7077 ( .A1(n5207), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5347) );
  OR2_X1 U7078 ( .A1(n7658), .A2(n7694), .ZN(n5749) );
  NAND2_X1 U7079 ( .A1(n7658), .A2(n7694), .ZN(n7689) );
  NAND2_X1 U7080 ( .A1(n5383), .A2(n5351), .ZN(n5363) );
  AND2_X1 U7081 ( .A1(n5352), .A2(n5364), .ZN(n5362) );
  XNOR2_X1 U7082 ( .A(n5363), .B(n5362), .ZN(n6450) );
  NAND2_X1 U7083 ( .A1(n6450), .A2(n4277), .ZN(n5355) );
  NAND2_X1 U7084 ( .A1(n5411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5369) );
  XNOR2_X1 U7085 ( .A(n5369), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8330) );
  AOI22_X1 U7086 ( .A1(n5545), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8330), .B2(
        n6472), .ZN(n5354) );
  NAND2_X1 U7087 ( .A1(n5695), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U7088 ( .A1(n5694), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U7089 ( .A1(n5356), .A2(n10148), .ZN(n5357) );
  AND2_X1 U7090 ( .A1(n5376), .A2(n5357), .ZN(n8626) );
  NAND2_X1 U7091 ( .A1(n5647), .A2(n8626), .ZN(n5359) );
  NAND2_X1 U7092 ( .A1(n5207), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5358) );
  OR2_X1 U7094 ( .A1(n8627), .A2(n7768), .ZN(n5754) );
  NAND2_X1 U7095 ( .A1(n8627), .A2(n7768), .ZN(n5751) );
  INV_X1 U7096 ( .A(n7690), .ZN(n5722) );
  NAND2_X1 U7097 ( .A1(n5363), .A2(n5362), .ZN(n5365) );
  NAND2_X1 U7098 ( .A1(n5365), .A2(n5364), .ZN(n5368) );
  INV_X1 U7099 ( .A(n5366), .ZN(n5367) );
  NAND2_X1 U7100 ( .A1(n6452), .A2(n4276), .ZN(n5374) );
  NAND2_X1 U7101 ( .A1(n5369), .A2(n5409), .ZN(n5370) );
  NAND2_X1 U7102 ( .A1(n5370), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5371) );
  INV_X1 U7103 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U7104 ( .A1(n5371), .A2(n5408), .ZN(n5393) );
  OR2_X1 U7105 ( .A1(n5371), .A2(n5408), .ZN(n5372) );
  AOI22_X1 U7106 ( .A1(n8344), .A2(n6472), .B1(n5545), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U7107 ( .A1(n5695), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U7108 ( .A1(n5694), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5380) );
  INV_X1 U7109 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U7110 ( .A1(n5376), .A2(n5375), .ZN(n5377) );
  AND2_X1 U7111 ( .A1(n5398), .A2(n5377), .ZN(n7777) );
  NAND2_X1 U7112 ( .A1(n5622), .A2(n7777), .ZN(n5379) );
  NAND2_X1 U7113 ( .A1(n5207), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U7114 ( .A1(n7774), .A2(n7816), .ZN(n5758) );
  INV_X1 U7115 ( .A(n5384), .ZN(n5385) );
  NAND2_X1 U7116 ( .A1(n5383), .A2(n5385), .ZN(n5387) );
  NAND2_X1 U7117 ( .A1(n5387), .A2(n5386), .ZN(n5389) );
  NAND2_X1 U7118 ( .A1(n5389), .A2(n5388), .ZN(n5392) );
  INV_X1 U7119 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U7120 ( .A1(n6454), .A2(n4276), .ZN(n5396) );
  NAND2_X1 U7121 ( .A1(n5393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U7122 ( .A(n5394), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6913) );
  AOI22_X1 U7123 ( .A1(n6913), .A2(n6472), .B1(n5545), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U7124 ( .A1(n5695), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U7125 ( .A1(n5694), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5402) );
  INV_X1 U7126 ( .A(n5418), .ZN(n5434) );
  INV_X1 U7127 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U7128 ( .A1(n5398), .A2(n7815), .ZN(n5399) );
  AND2_X1 U7129 ( .A1(n5434), .A2(n5399), .ZN(n7813) );
  NAND2_X1 U7130 ( .A1(n5647), .A2(n7813), .ZN(n5401) );
  NAND4_X1 U7131 ( .A1(n5403), .A2(n5402), .A3(n5401), .A4(n5400), .ZN(n8253)
         );
  INV_X1 U7132 ( .A(n8253), .ZN(n7919) );
  NAND2_X1 U7133 ( .A1(n7819), .A2(n7919), .ZN(n5851) );
  INV_X1 U7134 ( .A(n5851), .ZN(n5763) );
  AND2_X1 U7135 ( .A1(n5406), .A2(n5444), .ZN(n5442) );
  XNOR2_X1 U7136 ( .A(n5443), .B(n5442), .ZN(n6469) );
  NAND2_X1 U7137 ( .A1(n6469), .A2(n4277), .ZN(n5417) );
  INV_X1 U7138 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5407) );
  NAND3_X1 U7139 ( .A1(n5409), .A2(n5408), .A3(n5407), .ZN(n5410) );
  INV_X1 U7140 ( .A(n5426), .ZN(n5413) );
  INV_X1 U7141 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U7142 ( .A1(n5413), .A2(n5412), .ZN(n5428) );
  NAND2_X1 U7143 ( .A1(n5428), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5414) );
  MUX2_X1 U7144 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5414), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n5415) );
  AOI22_X1 U7145 ( .A1(n6919), .A2(n6472), .B1(n5545), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U7146 ( .A1(n5695), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U7147 ( .A1(n5694), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5422) );
  INV_X1 U7148 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6968) );
  NAND2_X1 U7149 ( .A1(n5436), .A2(n6968), .ZN(n5419) );
  AND2_X1 U7150 ( .A1(n5455), .A2(n5419), .ZN(n8175) );
  NAND2_X1 U7151 ( .A1(n5647), .A2(n8175), .ZN(n5421) );
  NAND2_X1 U7152 ( .A1(n5670), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5420) );
  XNOR2_X1 U7153 ( .A(n5424), .B(n5425), .ZN(n6456) );
  NAND2_X1 U7154 ( .A1(n6456), .A2(n4276), .ZN(n5432) );
  NAND2_X1 U7155 ( .A1(n5426), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5427) );
  MUX2_X1 U7156 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5427), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n5429) );
  NAND2_X1 U7157 ( .A1(n5429), .A2(n5428), .ZN(n6917) );
  OAI22_X1 U7158 ( .A1(n6917), .A2(n6650), .B1(n4468), .B2(n6459), .ZN(n5430)
         );
  INV_X1 U7159 ( .A(n5430), .ZN(n5431) );
  NAND2_X1 U7160 ( .A1(n5695), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U7161 ( .A1(n5694), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5439) );
  INV_X1 U7162 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U7163 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  AND2_X1 U7164 ( .A1(n5436), .A2(n5435), .ZN(n7916) );
  NAND2_X1 U7165 ( .A1(n5647), .A2(n7916), .ZN(n5438) );
  NAND2_X1 U7166 ( .A1(n5207), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5437) );
  OR2_X1 U7167 ( .A1(n8743), .A2(n8172), .ZN(n5850) );
  AND2_X1 U7168 ( .A1(n5850), .A2(n7839), .ZN(n7859) );
  NAND2_X1 U7169 ( .A1(n5443), .A2(n5442), .ZN(n5445) );
  NAND2_X1 U7170 ( .A1(n5445), .A2(n5444), .ZN(n5447) );
  NAND2_X1 U7171 ( .A1(n6479), .A2(n4276), .ZN(n5453) );
  NAND2_X1 U7172 ( .A1(n5448), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U7173 ( .A1(n5450), .A2(n10130), .ZN(n5467) );
  OR2_X1 U7174 ( .A1(n5450), .A2(n10130), .ZN(n5451) );
  AOI22_X1 U7175 ( .A1(n7136), .A2(n6472), .B1(n5545), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U7176 ( .A1(n5695), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U7177 ( .A1(n5694), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5459) );
  INV_X1 U7178 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U7179 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  AND2_X1 U7180 ( .A1(n5475), .A2(n5456), .ZN(n8073) );
  NAND2_X1 U7181 ( .A1(n5622), .A2(n8073), .ZN(n5458) );
  NAND2_X1 U7182 ( .A1(n5670), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U7183 ( .A1(n8733), .A2(n8171), .ZN(n5770) );
  NAND2_X1 U7184 ( .A1(n5769), .A2(n5770), .ZN(n7885) );
  NAND2_X1 U7185 ( .A1(n8743), .A2(n8172), .ZN(n7862) );
  INV_X1 U7186 ( .A(n7862), .ZN(n7863) );
  NAND2_X1 U7187 ( .A1(n5765), .A2(n7863), .ZN(n5461) );
  NAND2_X1 U7188 ( .A1(n8737), .A2(n8071), .ZN(n5766) );
  NAND2_X1 U7189 ( .A1(n5461), .A2(n5766), .ZN(n5462) );
  NOR2_X1 U7190 ( .A1(n7885), .A2(n5462), .ZN(n5463) );
  XNOR2_X1 U7191 ( .A(n5465), .B(n5466), .ZN(n6476) );
  NAND2_X1 U7192 ( .A1(n6476), .A2(n4277), .ZN(n5470) );
  NAND2_X1 U7193 ( .A1(n5467), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5468) );
  XNOR2_X1 U7194 ( .A(n5468), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7209) );
  AOI22_X1 U7195 ( .A1(n7209), .A2(n6472), .B1(n5545), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5469) );
  NAND2_X2 U7196 ( .A1(n5470), .A2(n5469), .ZN(n8728) );
  NAND2_X1 U7197 ( .A1(n5694), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U7198 ( .A1(n5695), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5471) );
  AND2_X1 U7199 ( .A1(n5472), .A2(n5471), .ZN(n5479) );
  INV_X1 U7200 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U7201 ( .A1(n5475), .A2(n5474), .ZN(n5476) );
  NAND2_X1 U7202 ( .A1(n5492), .A2(n5476), .ZN(n7902) );
  OR2_X1 U7203 ( .A1(n7902), .A2(n5669), .ZN(n5478) );
  NAND2_X1 U7204 ( .A1(n5670), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U7205 ( .A1(n8728), .A2(n8604), .ZN(n5772) );
  NAND2_X1 U7206 ( .A1(n5773), .A2(n5772), .ZN(n5916) );
  XNOR2_X1 U7207 ( .A(n5480), .B(n5032), .ZN(n6482) );
  NAND2_X1 U7208 ( .A1(n6482), .A2(n4277), .ZN(n5490) );
  NOR2_X1 U7209 ( .A1(n5483), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7210 ( .A1(n5482), .A2(n5484), .ZN(n5486) );
  OAI21_X1 U7211 ( .B1(n5486), .B2(n5485), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5487) );
  MUX2_X1 U7212 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5487), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5488) );
  AND2_X1 U7213 ( .A1(n5500), .A2(n5488), .ZN(n7624) );
  AOI22_X1 U7214 ( .A1(n5545), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6472), .B2(
        n7624), .ZN(n5489) );
  INV_X1 U7215 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U7216 ( .A1(n5492), .A2(n5491), .ZN(n5493) );
  AND2_X1 U7217 ( .A1(n5508), .A2(n5493), .ZN(n8618) );
  NAND2_X1 U7218 ( .A1(n8618), .A2(n5622), .ZN(n5497) );
  AOI22_X1 U7219 ( .A1(n5695), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n5671), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7220 ( .A1(n5670), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7221 ( .A1(n8721), .A2(n8248), .ZN(n5779) );
  NAND2_X1 U7222 ( .A1(n6570), .A2(n4277), .ZN(n5505) );
  NAND2_X1 U7223 ( .A1(n5500), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5501) );
  MUX2_X1 U7224 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5501), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5503) );
  AND2_X1 U7225 ( .A1(n5503), .A2(n5502), .ZN(n8361) );
  AOI22_X1 U7226 ( .A1(n5545), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6472), .B2(
        n8361), .ZN(n5504) );
  NAND2_X2 U7227 ( .A1(n5505), .A2(n5504), .ZN(n8717) );
  INV_X1 U7228 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7229 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  NAND2_X1 U7230 ( .A1(n5520), .A2(n5509), .ZN(n8142) );
  OR2_X1 U7231 ( .A1(n8142), .A2(n5669), .ZN(n5512) );
  AOI22_X1 U7232 ( .A1(n5695), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n5671), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7233 ( .A1(n5670), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5510) );
  OR2_X2 U7234 ( .A1(n8717), .A2(n8606), .ZN(n5783) );
  NAND2_X1 U7235 ( .A1(n8717), .A2(n8606), .ZN(n5782) );
  XNOR2_X1 U7236 ( .A(n5514), .B(n5513), .ZN(n6789) );
  NAND2_X1 U7237 ( .A1(n6789), .A2(n4276), .ZN(n5518) );
  NAND2_X1 U7238 ( .A1(n5502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5515) );
  MUX2_X1 U7239 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5515), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n5516) );
  NAND2_X1 U7240 ( .A1(n5516), .A2(n5542), .ZN(n8368) );
  INV_X1 U7241 ( .A(n8368), .ZN(n8379) );
  AOI22_X1 U7242 ( .A1(n5545), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6472), .B2(
        n8379), .ZN(n5517) );
  INV_X1 U7243 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7244 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  NAND2_X1 U7245 ( .A1(n5548), .A2(n5521), .ZN(n8202) );
  OR2_X1 U7246 ( .A1(n8202), .A2(n5669), .ZN(n5526) );
  INV_X1 U7247 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U7248 ( .A1(n5670), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7249 ( .A1(n5671), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5522) );
  OAI211_X1 U7250 ( .C1(n5674), .C2(n8362), .A(n5523), .B(n5522), .ZN(n5524)
         );
  INV_X1 U7251 ( .A(n5524), .ZN(n5525) );
  NAND2_X1 U7252 ( .A1(n5526), .A2(n5525), .ZN(n8568) );
  INV_X1 U7253 ( .A(n8568), .ZN(n5917) );
  OR2_X1 U7254 ( .A1(n8711), .A2(n5917), .ZN(n5796) );
  NAND2_X1 U7255 ( .A1(n8711), .A2(n5917), .ZN(n5788) );
  NAND2_X1 U7256 ( .A1(n7219), .A2(n4277), .ZN(n5530) );
  OR2_X1 U7257 ( .A1(n4468), .A2(n7270), .ZN(n5529) );
  INV_X1 U7258 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8095) );
  INV_X1 U7259 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7260 ( .A1(n5562), .A2(n5533), .ZN(n5534) );
  NAND2_X1 U7261 ( .A1(n5574), .A2(n5534), .ZN(n8528) );
  INV_X1 U7262 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U7263 ( .A1(n5695), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7264 ( .A1(n5671), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5535) );
  OAI211_X1 U7265 ( .C1(n8529), .C2(n5699), .A(n5536), .B(n5535), .ZN(n5537)
         );
  INV_X1 U7266 ( .A(n5537), .ZN(n5538) );
  INV_X1 U7267 ( .A(n8543), .ZN(n5580) );
  OR2_X1 U7268 ( .A1(n8698), .A2(n5580), .ZN(n5843) );
  XNOR2_X1 U7269 ( .A(n5541), .B(n5540), .ZN(n6873) );
  NAND2_X1 U7270 ( .A1(n6873), .A2(n4277), .ZN(n5547) );
  AOI22_X1 U7271 ( .A1(n5545), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7373), .B2(
        n6472), .ZN(n5546) );
  NAND2_X1 U7272 ( .A1(n5548), .A2(n8095), .ZN(n5549) );
  NAND2_X1 U7273 ( .A1(n5560), .A2(n5549), .ZN(n8096) );
  INV_X1 U7274 ( .A(n8096), .ZN(n8563) );
  NAND2_X1 U7275 ( .A1(n8563), .A2(n5622), .ZN(n5554) );
  INV_X1 U7276 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U7277 ( .A1(n5670), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7278 ( .A1(n5671), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5550) );
  OAI211_X1 U7279 ( .C1(n5674), .C2(n8380), .A(n5551), .B(n5550), .ZN(n5552)
         );
  INV_X1 U7280 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U7281 ( .A1(n8707), .A2(n8203), .ZN(n8540) );
  NAND2_X1 U7282 ( .A1(n5797), .A2(n8540), .ZN(n8559) );
  INV_X1 U7283 ( .A(n8559), .ZN(n8567) );
  XNOR2_X1 U7284 ( .A(n5556), .B(n5555), .ZN(n7117) );
  NAND2_X1 U7285 ( .A1(n7117), .A2(n4276), .ZN(n5558) );
  OR2_X1 U7286 ( .A1(n4468), .A2(n7121), .ZN(n5557) );
  INV_X1 U7287 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7288 ( .A1(n5560), .A2(n5559), .ZN(n5561) );
  AND2_X1 U7289 ( .A1(n5562), .A2(n5561), .ZN(n8550) );
  NAND2_X1 U7290 ( .A1(n8550), .A2(n5622), .ZN(n5568) );
  INV_X1 U7291 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7292 ( .A1(n5695), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7293 ( .A1(n5671), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5563) );
  OAI211_X1 U7294 ( .C1(n5565), .C2(n5699), .A(n5564), .B(n5563), .ZN(n5566)
         );
  INV_X1 U7295 ( .A(n5566), .ZN(n5567) );
  XNOR2_X1 U7296 ( .A(n5571), .B(n5570), .ZN(n7298) );
  NAND2_X1 U7297 ( .A1(n7298), .A2(n4276), .ZN(n5573) );
  OR2_X1 U7298 ( .A1(n4468), .A2(n7300), .ZN(n5572) );
  INV_X1 U7299 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U7300 ( .A1(n5574), .A2(n8190), .ZN(n5575) );
  AND2_X1 U7301 ( .A1(n5591), .A2(n5575), .ZN(n8510) );
  INV_X1 U7302 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7303 ( .A1(n5695), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7304 ( .A1(n5671), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5576) );
  OAI211_X1 U7305 ( .C1(n5578), .C2(n5699), .A(n5577), .B(n5576), .ZN(n5579)
         );
  NAND2_X1 U7306 ( .A1(n8691), .A2(n8537), .ZN(n5793) );
  AND2_X1 U7307 ( .A1(n5843), .A2(n8514), .ZN(n5790) );
  NAND2_X1 U7308 ( .A1(n8701), .A2(n8536), .ZN(n5845) );
  NAND2_X1 U7309 ( .A1(n5845), .A2(n8540), .ZN(n5791) );
  AND2_X1 U7310 ( .A1(n8698), .A2(n5580), .ZN(n8516) );
  AOI21_X1 U7311 ( .B1(n5790), .B2(n5791), .A(n8516), .ZN(n5581) );
  NAND2_X1 U7312 ( .A1(n7629), .A2(n4277), .ZN(n5589) );
  OR2_X1 U7313 ( .A1(n4468), .A2(n7632), .ZN(n5588) );
  INV_X1 U7314 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7315 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  NAND2_X1 U7316 ( .A1(n5602), .A2(n5592), .ZN(n8498) );
  INV_X1 U7317 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U7318 ( .A1(n5695), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7319 ( .A1(n5671), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5593) );
  OAI211_X1 U7320 ( .C1(n8499), .C2(n5699), .A(n5594), .B(n5593), .ZN(n5595)
         );
  INV_X1 U7321 ( .A(n5595), .ZN(n5596) );
  INV_X1 U7322 ( .A(n8502), .ZN(n8494) );
  NAND2_X1 U7323 ( .A1(n7757), .A2(n4277), .ZN(n5601) );
  OR2_X1 U7324 ( .A1(n4468), .A2(n7783), .ZN(n5600) );
  INV_X1 U7325 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U7326 ( .A1(n5602), .A2(n8155), .ZN(n5603) );
  NAND2_X1 U7327 ( .A1(n8484), .A2(n5622), .ZN(n5609) );
  INV_X1 U7328 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7329 ( .A1(n5695), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7330 ( .A1(n5694), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5604) );
  OAI211_X1 U7331 ( .C1(n5606), .C2(n5699), .A(n5605), .B(n5604), .ZN(n5607)
         );
  INV_X1 U7332 ( .A(n5607), .ZN(n5608) );
  XNOR2_X2 U7333 ( .A(n8681), .B(n8246), .ZN(n8487) );
  OR2_X1 U7334 ( .A1(n8681), .A2(n8505), .ZN(n8467) );
  NAND2_X1 U7335 ( .A1(n8466), .A2(n8467), .ZN(n5623) );
  NAND2_X1 U7336 ( .A1(n7798), .A2(n4277), .ZN(n5613) );
  OR2_X1 U7337 ( .A1(n4468), .A2(n7838), .ZN(n5612) );
  NAND2_X2 U7338 ( .A1(n5613), .A2(n5612), .ZN(n8678) );
  INV_X1 U7339 ( .A(n5628), .ZN(n5630) );
  INV_X1 U7340 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7341 ( .A1(n5616), .A2(n5615), .ZN(n5617) );
  INV_X1 U7342 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7343 ( .A1(n5695), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7344 ( .A1(n5671), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5618) );
  OAI211_X1 U7345 ( .C1(n5620), .C2(n5699), .A(n5619), .B(n5618), .ZN(n5621)
         );
  NAND2_X1 U7346 ( .A1(n8678), .A2(n8218), .ZN(n5814) );
  NAND2_X1 U7347 ( .A1(n7875), .A2(n4276), .ZN(n5627) );
  OR2_X1 U7348 ( .A1(n4468), .A2(n7893), .ZN(n5626) );
  INV_X1 U7349 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7350 ( .A1(n5630), .A2(n5629), .ZN(n5631) );
  NAND2_X1 U7351 ( .A1(n5641), .A2(n5631), .ZN(n8451) );
  INV_X1 U7352 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U7353 ( .A1(n5695), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7354 ( .A1(n5671), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5632) );
  OAI211_X1 U7355 ( .C1(n8450), .C2(n5699), .A(n5633), .B(n5632), .ZN(n5634)
         );
  INV_X1 U7356 ( .A(n5634), .ZN(n5635) );
  NAND2_X1 U7357 ( .A1(n8673), .A2(n8437), .ZN(n5818) );
  INV_X2 U7358 ( .A(n5928), .ZN(n8455) );
  NAND2_X1 U7359 ( .A1(n8799), .A2(n4276), .ZN(n5640) );
  OR2_X1 U7360 ( .A1(n4468), .A2(n8801), .ZN(n5639) );
  INV_X1 U7361 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U7362 ( .A1(n5641), .A2(n8065), .ZN(n5642) );
  INV_X1 U7363 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7364 ( .A1(n5695), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7365 ( .A1(n5671), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5643) );
  OAI211_X1 U7366 ( .C1(n5645), .C2(n5699), .A(n5644), .B(n5643), .ZN(n5646)
         );
  INV_X1 U7367 ( .A(n8435), .ZN(n5820) );
  OR2_X1 U7368 ( .A1(n8666), .A2(n8217), .ZN(n5824) );
  NAND2_X1 U7369 ( .A1(n9859), .A2(n4277), .ZN(n5651) );
  OR2_X1 U7370 ( .A1(n4468), .A2(n8798), .ZN(n5650) );
  INV_X1 U7371 ( .A(n5654), .ZN(n5652) );
  NAND2_X1 U7372 ( .A1(n5652), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8419) );
  INV_X1 U7373 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7374 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  NAND2_X1 U7375 ( .A1(n8419), .A2(n5655), .ZN(n8025) );
  INV_X1 U7376 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10223) );
  NAND2_X1 U7377 ( .A1(n5695), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7378 ( .A1(n5670), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5656) );
  OAI211_X1 U7379 ( .C1(n5321), .C2(n10223), .A(n5657), .B(n5656), .ZN(n5658)
         );
  INV_X1 U7380 ( .A(n5658), .ZN(n5659) );
  NAND2_X1 U7381 ( .A1(n8017), .A2(n8438), .ZN(n5661) );
  INV_X1 U7382 ( .A(n5936), .ZN(n5662) );
  XNOR2_X1 U7383 ( .A(n5665), .B(n5664), .ZN(n5666) );
  NAND2_X1 U7384 ( .A1(n8034), .A2(n4276), .ZN(n5668) );
  INV_X1 U7385 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7933) );
  OR2_X1 U7386 ( .A1(n4468), .A2(n7933), .ZN(n5667) );
  OR2_X1 U7387 ( .A1(n8419), .A2(n5669), .ZN(n5678) );
  INV_X1 U7388 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7389 ( .A1(n5670), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7390 ( .A1(n5671), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5672) );
  OAI211_X1 U7391 ( .C1(n5675), .C2(n5674), .A(n5673), .B(n5672), .ZN(n5676)
         );
  INV_X1 U7392 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U7393 ( .A1(n8417), .A2(n7634), .ZN(n5830) );
  INV_X1 U7394 ( .A(n8410), .ZN(n5829) );
  INV_X1 U7395 ( .A(n5830), .ZN(n5679) );
  OAI211_X1 U7396 ( .C1(n8659), .C2(n5711), .A(n5707), .B(n7373), .ZN(n5710)
         );
  INV_X1 U7397 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U7398 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  INV_X1 U7399 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5690) );
  INV_X1 U7400 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5686) );
  MUX2_X1 U7401 ( .A(n5690), .B(n5686), .S(n4807), .Z(n5687) );
  XNOR2_X1 U7402 ( .A(n5687), .B(SI_31_), .ZN(n5688) );
  NOR2_X1 U7403 ( .A1(n4468), .A2(n5690), .ZN(n5692) );
  INV_X1 U7404 ( .A(n5704), .ZN(n5693) );
  INV_X1 U7405 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7406 ( .A1(n5671), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7407 ( .A1(n5695), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5696) );
  OAI211_X1 U7408 ( .C1(n5699), .C2(n5698), .A(n5697), .B(n5696), .ZN(n8412)
         );
  INV_X1 U7409 ( .A(n8412), .ZN(n5702) );
  NAND2_X1 U7410 ( .A1(n8402), .A2(n5702), .ZN(n5833) );
  NAND2_X1 U7411 ( .A1(n5703), .A2(n7373), .ZN(n5701) );
  NAND3_X1 U7412 ( .A1(n8402), .A2(n7028), .A3(n8390), .ZN(n5700) );
  MUX2_X1 U7413 ( .A(n5701), .B(n5700), .S(n8651), .Z(n5709) );
  NOR2_X1 U7414 ( .A1(n8402), .A2(n5702), .ZN(n5834) );
  INV_X1 U7415 ( .A(n5703), .ZN(n8398) );
  AOI211_X1 U7416 ( .C1(n5834), .C2(n5711), .A(n7373), .B(n5835), .ZN(n5705)
         );
  INV_X1 U7417 ( .A(n5705), .ZN(n5706) );
  OAI211_X1 U7418 ( .C1(n5710), .C2(n5842), .A(n5709), .B(n5708), .ZN(n5721)
         );
  NAND3_X1 U7419 ( .A1(n5834), .A2(n7373), .A3(n5711), .ZN(n5713) );
  INV_X1 U7420 ( .A(n5835), .ZN(n5836) );
  NAND3_X1 U7421 ( .A1(n5842), .A2(n8390), .A3(n5836), .ZN(n5712) );
  OAI21_X1 U7422 ( .B1(n5842), .B2(n5713), .A(n5712), .ZN(n5720) );
  NAND2_X1 U7423 ( .A1(n5543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5714) );
  MUX2_X1 U7424 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5714), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5715) );
  NAND2_X1 U7425 ( .A1(n5715), .A2(n5716), .ZN(n7119) );
  INV_X1 U7426 ( .A(n7119), .ZN(n5944) );
  NAND2_X1 U7427 ( .A1(n7028), .A2(n5944), .ZN(n5938) );
  INV_X1 U7428 ( .A(n5938), .ZN(n5719) );
  INV_X1 U7429 ( .A(n7017), .ZN(n5718) );
  INV_X1 U7430 ( .A(n5793), .ZN(n5795) );
  NAND2_X1 U7431 ( .A1(n7765), .A2(n5722), .ZN(n5853) );
  NAND3_X1 U7432 ( .A1(n5756), .A2(n5837), .A3(n5754), .ZN(n5753) );
  NAND2_X1 U7433 ( .A1(n5848), .A2(n5727), .ZN(n5736) );
  AOI21_X1 U7434 ( .B1(n5723), .B2(n5729), .A(n5736), .ZN(n5725) );
  INV_X1 U7435 ( .A(n5741), .ZN(n5724) );
  NOR3_X1 U7436 ( .A1(n5725), .A2(n4849), .A3(n5724), .ZN(n5745) );
  AND2_X1 U7437 ( .A1(n4483), .A2(n7102), .ZN(n7099) );
  NOR2_X1 U7438 ( .A1(n7099), .A2(n7268), .ZN(n5726) );
  OAI211_X1 U7439 ( .C1(n6779), .C2(n5726), .A(n5738), .B(n5889), .ZN(n5728)
         );
  AND2_X1 U7440 ( .A1(n7470), .A2(n5727), .ZN(n5731) );
  NAND4_X1 U7441 ( .A1(n5737), .A2(n5731), .A3(n5728), .A4(n5839), .ZN(n5734)
         );
  NAND3_X1 U7442 ( .A1(n5734), .A2(n5733), .A3(n5732), .ZN(n5735) );
  AOI21_X1 U7443 ( .B1(n5837), .B2(n5736), .A(n5735), .ZN(n5743) );
  AOI21_X1 U7444 ( .B1(n5848), .B2(n7547), .A(n5837), .ZN(n5742) );
  INV_X1 U7445 ( .A(n5889), .ZN(n6778) );
  OAI211_X1 U7446 ( .C1(n6778), .C2(n7099), .A(n5737), .B(n5890), .ZN(n5739)
         );
  NAND3_X1 U7447 ( .A1(n5739), .A2(n5837), .A3(n5738), .ZN(n5740) );
  OAI211_X1 U7448 ( .C1(n5743), .C2(n5742), .A(n5741), .B(n5740), .ZN(n5744)
         );
  INV_X1 U7449 ( .A(n5905), .ZN(n7549) );
  MUX2_X1 U7450 ( .A(n5747), .B(n5746), .S(n5839), .Z(n5748) );
  MUX2_X1 U7451 ( .A(n7689), .B(n5749), .S(n5839), .Z(n5750) );
  AOI21_X1 U7452 ( .B1(n5853), .B2(n5753), .A(n5752), .ZN(n5762) );
  INV_X1 U7453 ( .A(n5754), .ZN(n5755) );
  NAND2_X1 U7454 ( .A1(n5758), .A2(n5755), .ZN(n5757) );
  NAND3_X1 U7455 ( .A1(n5757), .A2(n5756), .A3(n7839), .ZN(n5760) );
  NAND2_X1 U7456 ( .A1(n5758), .A2(n5851), .ZN(n5759) );
  MUX2_X1 U7457 ( .A(n5760), .B(n5759), .S(n5837), .Z(n5761) );
  INV_X1 U7458 ( .A(n5765), .ZN(n5767) );
  INV_X1 U7459 ( .A(n5766), .ZN(n7878) );
  MUX2_X1 U7460 ( .A(n5767), .B(n7878), .S(n5839), .Z(n5768) );
  MUX2_X1 U7461 ( .A(n5770), .B(n5769), .S(n5839), .Z(n5771) );
  NAND2_X1 U7462 ( .A1(n4631), .A2(n5771), .ZN(n5776) );
  NAND2_X1 U7463 ( .A1(n5778), .A2(n5779), .ZN(n8608) );
  INV_X1 U7464 ( .A(n8608), .ZN(n5775) );
  MUX2_X1 U7465 ( .A(n5773), .B(n5772), .S(n5839), .Z(n5774) );
  OAI211_X1 U7466 ( .C1(n5777), .C2(n5776), .A(n5775), .B(n5774), .ZN(n5781)
         );
  MUX2_X1 U7467 ( .A(n5779), .B(n5778), .S(n5839), .Z(n5780) );
  AOI21_X1 U7468 ( .B1(n5781), .B2(n5780), .A(n8595), .ZN(n5787) );
  NAND2_X1 U7469 ( .A1(n5788), .A2(n5782), .ZN(n5785) );
  NAND2_X1 U7470 ( .A1(n5796), .A2(n5783), .ZN(n5784) );
  MUX2_X1 U7471 ( .A(n5785), .B(n5784), .S(n5839), .Z(n5786) );
  INV_X1 U7472 ( .A(n5799), .ZN(n5789) );
  INV_X1 U7473 ( .A(n8516), .ZN(n5792) );
  MUX2_X1 U7474 ( .A(n5795), .B(n5794), .S(n5839), .Z(n5810) );
  NAND2_X1 U7475 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  OAI21_X1 U7476 ( .B1(n5799), .B2(n5798), .A(n8540), .ZN(n5801) );
  INV_X1 U7477 ( .A(n5845), .ZN(n5800) );
  AOI211_X1 U7478 ( .C1(n5801), .C2(n8514), .A(n5800), .B(n8516), .ZN(n5804)
         );
  NAND3_X1 U7479 ( .A1(n5802), .A2(n5837), .A3(n5843), .ZN(n5803) );
  OAI21_X1 U7480 ( .B1(n5804), .B2(n5803), .A(n8502), .ZN(n5809) );
  NAND2_X1 U7481 ( .A1(n8519), .A2(n5837), .ZN(n5806) );
  NAND2_X1 U7482 ( .A1(n5924), .A2(n5839), .ZN(n5805) );
  MUX2_X1 U7483 ( .A(n5806), .B(n5805), .S(n8688), .Z(n5807) );
  NAND2_X1 U7484 ( .A1(n8681), .A2(n8505), .ZN(n5811) );
  MUX2_X1 U7485 ( .A(n5811), .B(n8467), .S(n5839), .Z(n5812) );
  NAND2_X1 U7486 ( .A1(n5817), .A2(n5813), .ZN(n5816) );
  NAND2_X1 U7487 ( .A1(n8455), .A2(n5814), .ZN(n5815) );
  MUX2_X1 U7488 ( .A(n5816), .B(n5815), .S(n5839), .Z(n5821) );
  MUX2_X1 U7489 ( .A(n5818), .B(n5817), .S(n5839), .Z(n5819) );
  OAI211_X1 U7490 ( .C1(n4289), .C2(n5821), .A(n5820), .B(n5819), .ZN(n5823)
         );
  NAND2_X1 U7491 ( .A1(n5823), .A2(n5822), .ZN(n5827) );
  AOI21_X1 U7492 ( .B1(n5826), .B2(n5824), .A(n5839), .ZN(n5825) );
  NAND3_X1 U7493 ( .A1(n8017), .A2(n8438), .A3(n5837), .ZN(n5828) );
  MUX2_X1 U7494 ( .A(n5831), .B(n5830), .S(n5839), .Z(n5832) );
  NAND3_X1 U7495 ( .A1(n5842), .A2(n5837), .A3(n5836), .ZN(n5841) );
  INV_X1 U7496 ( .A(n5838), .ZN(n5840) );
  INV_X1 U7497 ( .A(n5842), .ZN(n5863) );
  INV_X1 U7498 ( .A(n5923), .ZN(n8517) );
  INV_X1 U7499 ( .A(n5843), .ZN(n5844) );
  NAND2_X1 U7500 ( .A1(n8514), .A2(n5845), .ZN(n8546) );
  INV_X1 U7501 ( .A(n8546), .ZN(n8541) );
  INV_X1 U7502 ( .A(n7099), .ZN(n6687) );
  NAND4_X1 U7503 ( .A1(n6936), .A2(n5944), .A3(n5889), .A4(n6687), .ZN(n5846)
         );
  NOR4_X1 U7504 ( .A1(n5846), .A2(n7540), .A3(n5896), .A4(n6779), .ZN(n5849)
         );
  AND2_X2 U7505 ( .A1(n5848), .A2(n5847), .ZN(n7106) );
  NAND4_X1 U7506 ( .A1(n5849), .A2(n7549), .A3(n7106), .A4(n7439), .ZN(n5852)
         );
  NOR4_X1 U7507 ( .A1(n5852), .A2(n7850), .A3(n5908), .A4(n7750), .ZN(n5856)
         );
  INV_X1 U7508 ( .A(n7885), .ZN(n5855) );
  INV_X1 U7509 ( .A(n5853), .ZN(n5854) );
  NAND4_X1 U7510 ( .A1(n5856), .A2(n5855), .A3(n7864), .A4(n5854), .ZN(n5857)
         );
  NAND4_X1 U7511 ( .A1(n8541), .A2(n8567), .A3(n4291), .A4(n5858), .ZN(n5859)
         );
  NOR4_X1 U7512 ( .A1(n8494), .A2(n8517), .A3(n8534), .A4(n5859), .ZN(n5860)
         );
  NAND4_X1 U7513 ( .A1(n8455), .A2(n8465), .A3(n5860), .A4(n8487), .ZN(n5861)
         );
  NAND3_X1 U7514 ( .A1(n5864), .A2(n5863), .A3(n5862), .ZN(n5865) );
  XNOR2_X1 U7515 ( .A(n5865), .B(n8390), .ZN(n5866) );
  OAI22_X1 U7516 ( .A1(n5866), .A2(n7028), .B1(n5944), .B2(n5939), .ZN(n5867)
         );
  NAND2_X1 U7517 ( .A1(n5869), .A2(n5717), .ZN(n5870) );
  INV_X1 U7518 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5872) );
  XNOR2_X1 U7519 ( .A(n5873), .B(n5872), .ZN(n7040) );
  OR2_X1 U7520 ( .A1(n7040), .A2(P2_U3152), .ZN(n7630) );
  NAND2_X1 U7521 ( .A1(n5878), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5879) );
  XNOR2_X1 U7522 ( .A(n5879), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5948) );
  INV_X1 U7523 ( .A(n5948), .ZN(n7895) );
  NOR2_X1 U7524 ( .A1(n5880), .A2(n5270), .ZN(n5881) );
  MUX2_X1 U7525 ( .A(n5270), .B(n5881), .S(P2_IR_REG_25__SCAN_IN), .Z(n5882)
         );
  INV_X1 U7526 ( .A(n5882), .ZN(n5883) );
  AND2_X1 U7527 ( .A1(n5878), .A2(n5883), .ZN(n5949) );
  INV_X1 U7528 ( .A(n5949), .ZN(n7836) );
  NAND2_X1 U7529 ( .A1(n5933), .A2(n7028), .ZN(n7024) );
  OR2_X1 U7530 ( .A1(n7024), .A2(n7017), .ZN(n7041) );
  NAND2_X1 U7531 ( .A1(n10031), .A2(n7041), .ZN(n6694) );
  INV_X1 U7532 ( .A(n7024), .ZN(n6473) );
  INV_X1 U7533 ( .A(n6658), .ZN(n5940) );
  NOR3_X1 U7534 ( .A1(n6694), .A2(n8800), .A3(n8603), .ZN(n5886) );
  OAI21_X1 U7535 ( .B1(n7630), .B2(n5933), .A(P2_B_REG_SCAN_IN), .ZN(n5885) );
  OR2_X1 U7536 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U7537 ( .A1(n5888), .A2(n5887), .ZN(P2_U3244) );
  NAND2_X1 U7538 ( .A1(n5890), .A2(n5889), .ZN(n6774) );
  NAND2_X1 U7539 ( .A1(n5891), .A2(n7580), .ZN(n5892) );
  NAND2_X1 U7540 ( .A1(n6775), .A2(n5892), .ZN(n7539) );
  NAND2_X1 U7541 ( .A1(n4467), .A2(n7541), .ZN(n5893) );
  OAI21_X2 U7542 ( .B1(n5894), .B2(n7539), .A(n5893), .ZN(n6932) );
  AND2_X1 U7543 ( .A1(n6933), .A2(n5896), .ZN(n5895) );
  NOR2_X1 U7544 ( .A1(n8261), .A2(n8636), .ZN(n7482) );
  NAND2_X1 U7545 ( .A1(n5896), .A2(n7482), .ZN(n5899) );
  NAND2_X1 U7546 ( .A1(n7176), .A2(n10043), .ZN(n5898) );
  NAND2_X1 U7547 ( .A1(n5899), .A2(n5898), .ZN(n7104) );
  NOR2_X1 U7548 ( .A1(n8259), .A2(n5900), .ZN(n5901) );
  NAND2_X1 U7549 ( .A1(n8258), .A2(n7448), .ZN(n5903) );
  NAND2_X1 U7550 ( .A1(n7308), .A2(n10051), .ZN(n5904) );
  NAND2_X1 U7551 ( .A1(n7545), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U7552 ( .A1(n7653), .A2(n10061), .ZN(n5906) );
  INV_X1 U7553 ( .A(n7694), .ZN(n8255) );
  NAND2_X1 U7554 ( .A1(n7658), .A2(n8255), .ZN(n5910) );
  INV_X1 U7555 ( .A(n7768), .ZN(n8254) );
  INV_X1 U7556 ( .A(n7774), .ZN(n8754) );
  NAND2_X1 U7557 ( .A1(n7819), .A2(n8253), .ZN(n7848) );
  NAND2_X1 U7558 ( .A1(n7850), .A2(n7848), .ZN(n5914) );
  INV_X1 U7559 ( .A(n7848), .ZN(n5911) );
  NOR2_X1 U7560 ( .A1(n7750), .A2(n5911), .ZN(n5912) );
  AOI22_X1 U7561 ( .A1(n5912), .A2(n7850), .B1(n8172), .B2(n7847), .ZN(n5913)
         );
  INV_X1 U7562 ( .A(n8071), .ZN(n8251) );
  INV_X1 U7563 ( .A(n8171), .ZN(n8250) );
  INV_X1 U7564 ( .A(n8728), .ZN(n7905) );
  INV_X1 U7565 ( .A(n8606), .ZN(n8581) );
  NAND2_X1 U7566 ( .A1(n8711), .A2(n8568), .ZN(n5919) );
  INV_X1 U7567 ( .A(n8711), .ZN(n8578) );
  NAND2_X1 U7568 ( .A1(n8560), .A2(n8559), .ZN(n8558) );
  NAND2_X1 U7569 ( .A1(n8558), .A2(n5034), .ZN(n8547) );
  NAND2_X1 U7570 ( .A1(n8547), .A2(n8546), .ZN(n8545) );
  NAND2_X1 U7571 ( .A1(n8545), .A2(n5035), .ZN(n8524) );
  NAND2_X1 U7572 ( .A1(n8524), .A2(n5920), .ZN(n5922) );
  NAND2_X1 U7573 ( .A1(n8698), .A2(n8543), .ZN(n5921) );
  INV_X1 U7574 ( .A(n8537), .ZN(n8247) );
  NAND2_X1 U7575 ( .A1(n8486), .A2(n8505), .ZN(n5927) );
  INV_X1 U7576 ( .A(n8678), .ZN(n8478) );
  AND2_X1 U7577 ( .A1(n8478), .A2(n8218), .ZN(n8445) );
  INV_X1 U7578 ( .A(n8673), .ZN(n8449) );
  AOI22_X1 U7579 ( .A1(n5928), .A2(n8445), .B1(n8437), .B2(n8449), .ZN(n5929)
         );
  NAND2_X1 U7580 ( .A1(n5930), .A2(n5929), .ZN(n8427) );
  NAND2_X1 U7581 ( .A1(n8433), .A2(n8217), .ZN(n5931) );
  OAI21_X1 U7582 ( .B1(n5932), .B2(n5936), .A(n8408), .ZN(n7924) );
  NAND2_X1 U7583 ( .A1(n7028), .A2(n7119), .ZN(n7369) );
  XNOR2_X1 U7584 ( .A(n5933), .B(n7369), .ZN(n5934) );
  NAND2_X1 U7585 ( .A1(n5934), .A2(n8390), .ZN(n8610) );
  AND2_X1 U7586 ( .A1(n7119), .A2(n7373), .ZN(n5935) );
  NAND2_X1 U7587 ( .A1(n7299), .A2(n5935), .ZN(n8759) );
  XNOR2_X1 U7588 ( .A(n5937), .B(n5936), .ZN(n5942) );
  AND2_X1 U7589 ( .A1(n5939), .A2(n5938), .ZN(n8535) );
  INV_X2 U7590 ( .A(n8535), .ZN(n8614) );
  OR2_X1 U7591 ( .A1(n8217), .A2(n8603), .ZN(n5941) );
  OAI21_X1 U7592 ( .B1(n7634), .B2(n8605), .A(n5941), .ZN(n7937) );
  NAND2_X1 U7593 ( .A1(n5943), .A2(n7102), .ZN(n7530) );
  AND2_X2 U7594 ( .A1(n7554), .A2(n10061), .ZN(n7654) );
  INV_X1 U7595 ( .A(n7658), .ZN(n10071) );
  INV_X1 U7596 ( .A(n7819), .ZN(n8748) );
  AND2_X2 U7597 ( .A1(n8448), .A2(n8433), .ZN(n8429) );
  OAI211_X1 U7598 ( .C1(n8429), .C2(n8406), .A(n8763), .B(n8416), .ZN(n7927)
         );
  INV_X1 U7599 ( .A(P2_B_REG_SCAN_IN), .ZN(n8396) );
  XNOR2_X1 U7600 ( .A(n7785), .B(n8396), .ZN(n5946) );
  INV_X1 U7601 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U7602 ( .A1(n5949), .A2(n5948), .ZN(n10036) );
  INV_X1 U7603 ( .A(n7367), .ZN(n5964) );
  NOR4_X1 U7604 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5953) );
  NOR4_X1 U7605 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5952) );
  NOR4_X1 U7606 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5951) );
  NOR4_X1 U7607 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5950) );
  NAND4_X1 U7608 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n5960)
         );
  NOR2_X1 U7609 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .ZN(
        n5957) );
  NOR4_X1 U7610 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5956) );
  NOR4_X1 U7611 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5955) );
  NOR4_X1 U7612 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5954) );
  NAND4_X1 U7613 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n5959)
         );
  OAI21_X1 U7614 ( .B1(n5960), .B2(n5959), .A(n5958), .ZN(n7014) );
  AND2_X1 U7615 ( .A1(n7785), .A2(n7895), .ZN(n10033) );
  NOR2_X1 U7616 ( .A1(n10030), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5961) );
  NOR2_X1 U7617 ( .A1(n6694), .A2(n7013), .ZN(n5962) );
  NAND2_X1 U7618 ( .A1(n7014), .A2(n5962), .ZN(n7366) );
  NOR2_X1 U7619 ( .A1(n7366), .A2(n7037), .ZN(n5963) );
  OR2_X1 U7620 ( .A1(n10076), .A2(n10223), .ZN(n5965) );
  NOR2_X2 U7621 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5969) );
  NOR2_X2 U7622 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5968) );
  NOR2_X2 U7623 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5967) );
  NAND3_X1 U7624 ( .A1(n5972), .A2(n5971), .A3(n6305), .ZN(n5973) );
  NAND2_X1 U7625 ( .A1(n6214), .A2(n6309), .ZN(n6302) );
  NOR2_X1 U7626 ( .A1(n5973), .A2(n6302), .ZN(n5974) );
  NAND2_X1 U7627 ( .A1(n6171), .A2(n5974), .ZN(n6387) );
  NOR2_X1 U7628 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5975) );
  NOR2_X1 U7629 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5979) );
  NOR2_X1 U7630 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5978) );
  XNOR2_X2 U7631 ( .A(n5983), .B(n5982), .ZN(n5986) );
  AND2_X2 U7632 ( .A1(n9854), .A2(n5987), .ZN(n6061) );
  NAND2_X1 U7633 ( .A1(n6061), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5991) );
  BUF_X2 U7634 ( .A(n5986), .Z(n5988) );
  NAND2_X1 U7635 ( .A1(n6057), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5990) );
  AND2_X2 U7636 ( .A1(n5988), .A2(n5987), .ZN(n6056) );
  NAND2_X1 U7637 ( .A1(n6056), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5989) );
  XNOR2_X1 U7638 ( .A(n5992), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9868) );
  INV_X1 U7639 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5993) );
  INV_X1 U7640 ( .A(n5994), .ZN(n5996) );
  NOR2_X1 U7641 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  MUX2_X1 U7642 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9868), .S(n9056), .Z(n7092) );
  NAND2_X1 U7643 ( .A1(n7004), .A2(n7092), .ZN(n6634) );
  NAND2_X1 U7644 ( .A1(n6057), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7645 ( .A1(n6056), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7646 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6006) );
  NAND2_X1 U7647 ( .A1(n6044), .A2(n6518), .ZN(n6007) );
  NAND2_X1 U7648 ( .A1(n6633), .A2(n9956), .ZN(n6997) );
  NAND2_X1 U7649 ( .A1(n6634), .A2(n6997), .ZN(n9288) );
  INV_X1 U7650 ( .A(n9956), .ZN(n6716) );
  NAND2_X1 U7651 ( .A1(n6057), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7652 ( .A1(n6061), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7653 ( .A1(n6056), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7654 ( .A1(n9066), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7655 ( .A1(n6044), .A2(n6519), .ZN(n6013) );
  NAND2_X1 U7656 ( .A1(n6335), .A2(n6993), .ZN(n9290) );
  NAND2_X1 U7657 ( .A1(n9356), .A2(n6755), .ZN(n9286) );
  NAND2_X1 U7658 ( .A1(n6057), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7659 ( .A1(n6056), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7660 ( .A1(n6061), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6017) );
  INV_X1 U7661 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7662 ( .A1(n6060), .A2(n6015), .ZN(n6016) );
  AND4_X2 U7663 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n6339)
         );
  INV_X1 U7664 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7665 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  NAND2_X1 U7666 ( .A1(n6022), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7667 ( .A1(n6044), .A2(n6520), .ZN(n6024) );
  NAND2_X1 U7668 ( .A1(n9355), .A2(n4860), .ZN(n9202) );
  NAND2_X1 U7669 ( .A1(n6056), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7670 ( .A1(n6057), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7671 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6038), .ZN(n7067) );
  INV_X1 U7672 ( .A(n7067), .ZN(n6025) );
  NAND2_X1 U7673 ( .A1(n6060), .A2(n6025), .ZN(n6027) );
  INV_X2 U7674 ( .A(n6061), .ZN(n6070) );
  INV_X2 U7675 ( .A(n6070), .ZN(n8046) );
  NAND2_X1 U7676 ( .A1(n6061), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6026) );
  INV_X1 U7677 ( .A(n6030), .ZN(n6032) );
  NOR2_X1 U7678 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6031) );
  NAND2_X1 U7679 ( .A1(n6032), .A2(n6031), .ZN(n6045) );
  NAND2_X1 U7680 ( .A1(n6045), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6034) );
  INV_X1 U7681 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6033) );
  XNOR2_X1 U7682 ( .A(n6034), .B(n6033), .ZN(n6521) );
  NAND2_X1 U7683 ( .A1(n6429), .A2(n6091), .ZN(n6037) );
  NAND2_X1 U7684 ( .A1(n9066), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6036) );
  OAI211_X1 U7685 ( .C1(n9056), .C2(n6521), .A(n6037), .B(n6036), .ZN(n7073)
         );
  NAND2_X1 U7686 ( .A1(n7284), .A2(n7073), .ZN(n9295) );
  INV_X1 U7687 ( .A(n7284), .ZN(n9354) );
  AND2_X1 U7688 ( .A1(n6038), .A2(n6698), .ZN(n6039) );
  NOR2_X1 U7689 ( .A1(n6058), .A2(n6039), .ZN(n7288) );
  NAND2_X1 U7690 ( .A1(n6060), .A2(n7288), .ZN(n6043) );
  NAND2_X1 U7691 ( .A1(n6057), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7692 ( .A1(n8046), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7693 ( .A1(n6056), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6040) );
  AND4_X2 U7694 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n6800)
         );
  NAND2_X1 U7695 ( .A1(n6425), .A2(n6091), .ZN(n6052) );
  NAND2_X1 U7696 ( .A1(n6047), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6046) );
  MUX2_X1 U7697 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6046), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n6050) );
  INV_X1 U7698 ( .A(n6047), .ZN(n6049) );
  INV_X1 U7699 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7700 ( .A1(n6049), .A2(n6048), .ZN(n6066) );
  NAND2_X1 U7701 ( .A1(n6050), .A2(n6066), .ZN(n6522) );
  INV_X1 U7702 ( .A(n6522), .ZN(n6707) );
  AOI22_X1 U7703 ( .A1(n9066), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6424), .B2(
        n6707), .ZN(n6051) );
  NAND2_X1 U7704 ( .A1(n6433), .A2(n6091), .ZN(n6055) );
  NAND2_X1 U7705 ( .A1(n6066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6053) );
  XNOR2_X1 U7706 ( .A(n6053), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6684) );
  AOI22_X1 U7707 ( .A1(n9066), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6044), .B2(
        n6684), .ZN(n6054) );
  NAND2_X1 U7708 ( .A1(n6056), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7709 ( .A1(n6057), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6064) );
  OR2_X1 U7710 ( .A1(n6058), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6059) );
  AND2_X1 U7711 ( .A1(n6072), .A2(n6059), .ZN(n7084) );
  NAND2_X1 U7712 ( .A1(n6060), .A2(n7084), .ZN(n6063) );
  NAND2_X1 U7713 ( .A1(n6061), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7714 ( .A1(n6427), .A2(n6091), .ZN(n6069) );
  OAI21_X1 U7715 ( .B1(n6066), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U7716 ( .A(n6067), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6524) );
  AOI22_X1 U7717 ( .A1(n6286), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6424), .B2(
        n6524), .ZN(n6068) );
  NAND2_X1 U7718 ( .A1(n9057), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7719 ( .A1(n8046), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7720 ( .A1(n6072), .A2(n6071), .ZN(n6073) );
  AND2_X1 U7721 ( .A1(n6084), .A2(n6073), .ZN(n7320) );
  NAND2_X1 U7722 ( .A1(n6060), .A2(n7320), .ZN(n6075) );
  NAND2_X1 U7723 ( .A1(n9059), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7724 ( .A1(n7561), .A2(n7423), .ZN(n9070) );
  NAND2_X1 U7725 ( .A1(n6434), .A2(n6091), .ZN(n6082) );
  INV_X1 U7726 ( .A(n6171), .ZN(n6078) );
  NAND2_X1 U7727 ( .A1(n6078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6079) );
  MUX2_X1 U7728 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6079), .S(n10238), .Z(n6080)
         );
  OR2_X1 U7729 ( .A1(n6078), .A2(n10238), .ZN(n6102) );
  NAND2_X1 U7730 ( .A1(n6080), .A2(n6102), .ZN(n6541) );
  INV_X1 U7731 ( .A(n6541), .ZN(n6546) );
  AOI22_X1 U7732 ( .A1(n9066), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6424), .B2(
        n6546), .ZN(n6081) );
  NAND2_X1 U7733 ( .A1(n9057), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7734 ( .A1(n8046), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7735 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  NAND2_X1 U7736 ( .A1(n6110), .A2(n6085), .ZN(n7422) );
  INV_X1 U7737 ( .A(n7422), .ZN(n7229) );
  NAND2_X1 U7738 ( .A1(n6060), .A2(n7229), .ZN(n6088) );
  INV_X4 U7739 ( .A(n6086), .ZN(n9059) );
  NAND2_X1 U7740 ( .A1(n6056), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7741 ( .A1(n7414), .A2(n7570), .ZN(n9077) );
  INV_X1 U7742 ( .A(n6102), .ZN(n6093) );
  INV_X1 U7743 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7744 ( .A1(n6093), .A2(n6092), .ZN(n6105) );
  NAND2_X1 U7745 ( .A1(n6105), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6094) );
  XNOR2_X1 U7746 ( .A(n6094), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6816) );
  AOI22_X1 U7747 ( .A1(n9066), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6424), .B2(
        n6816), .ZN(n6095) );
  NAND2_X2 U7748 ( .A1(n6096), .A2(n6095), .ZN(n6327) );
  NAND2_X1 U7749 ( .A1(n9057), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7750 ( .A1(n9059), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6100) );
  OR2_X1 U7751 ( .A1(n6112), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6097) );
  AND2_X1 U7752 ( .A1(n6097), .A2(n6124), .ZN(n7710) );
  NAND2_X1 U7753 ( .A1(n6060), .A2(n7710), .ZN(n6099) );
  NAND2_X1 U7754 ( .A1(n9058), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7755 ( .A1(n6327), .A2(n7644), .ZN(n9081) );
  NAND2_X1 U7756 ( .A1(n6450), .A2(n6091), .ZN(n6108) );
  NAND2_X1 U7757 ( .A1(n6102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6103) );
  MUX2_X1 U7758 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6103), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n6104) );
  INV_X1 U7759 ( .A(n6104), .ZN(n6106) );
  INV_X1 U7760 ( .A(n6105), .ZN(n6120) );
  NOR2_X1 U7761 ( .A1(n6106), .A2(n6120), .ZN(n6767) );
  AOI22_X1 U7762 ( .A1(n9066), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6424), .B2(
        n6767), .ZN(n6107) );
  NAND2_X1 U7763 ( .A1(n9059), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7764 ( .A1(n9057), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6115) );
  AND2_X1 U7765 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  NOR2_X1 U7766 ( .A1(n6112), .A2(n6111), .ZN(n7641) );
  NAND2_X1 U7767 ( .A1(n6060), .A2(n7641), .ZN(n6114) );
  NAND2_X1 U7768 ( .A1(n9058), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7769 ( .A1(n7640), .A2(n7712), .ZN(n9078) );
  OR2_X1 U7770 ( .A1(n7640), .A2(n7712), .ZN(n9080) );
  NAND2_X1 U7771 ( .A1(n9080), .A2(n9076), .ZN(n7329) );
  NAND2_X1 U7772 ( .A1(n9192), .A2(n7329), .ZN(n6117) );
  OAI21_X2 U7773 ( .B1(n7236), .B2(n6118), .A(n9172), .ZN(n7357) );
  NAND2_X1 U7774 ( .A1(n6454), .A2(n6091), .ZN(n6123) );
  INV_X1 U7775 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7776 ( .A1(n6120), .A2(n6119), .ZN(n6130) );
  NAND2_X1 U7777 ( .A1(n6130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6121) );
  XNOR2_X1 U7778 ( .A(n6121), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7275) );
  AOI22_X1 U7779 ( .A1(n9066), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6424), .B2(
        n7275), .ZN(n6122) );
  NAND2_X1 U7780 ( .A1(n9057), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7781 ( .A1(n8046), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7782 ( .A1(n6124), .A2(n6820), .ZN(n6125) );
  AND2_X1 U7783 ( .A1(n6135), .A2(n6125), .ZN(n7522) );
  NAND2_X1 U7784 ( .A1(n6060), .A2(n7522), .ZN(n6127) );
  NAND2_X1 U7785 ( .A1(n9059), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7786 ( .A1(n6456), .A2(n6091), .ZN(n6133) );
  NAND2_X1 U7787 ( .A1(n6144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6131) );
  XNOR2_X1 U7788 ( .A(n6131), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7387) );
  AOI22_X1 U7789 ( .A1(n9066), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6424), .B2(
        n7387), .ZN(n6132) );
  NAND2_X1 U7790 ( .A1(n9057), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6140) );
  AND2_X1 U7791 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  NOR2_X1 U7792 ( .A1(n6150), .A2(n6136), .ZN(n7678) );
  NAND2_X1 U7793 ( .A1(n4448), .A2(n7678), .ZN(n6139) );
  NAND2_X1 U7794 ( .A1(n9059), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7795 ( .A1(n9058), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7796 ( .A1(n9824), .A2(n7666), .ZN(n9109) );
  NAND2_X1 U7797 ( .A1(n9112), .A2(n9109), .ZN(n9248) );
  NAND3_X1 U7798 ( .A1(n9109), .A2(n9902), .A3(n9347), .ZN(n6143) );
  NAND2_X1 U7799 ( .A1(n6469), .A2(n6091), .ZN(n6149) );
  OAI21_X1 U7800 ( .B1(n6144), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6146) );
  INV_X1 U7801 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7802 ( .A1(n6146), .A2(n6145), .ZN(n6156) );
  OR2_X1 U7803 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  AOI22_X1 U7804 ( .A1(n9066), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9365), .B2(
        n6424), .ZN(n6148) );
  OR2_X1 U7805 ( .A1(n6150), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6151) );
  AND2_X1 U7806 ( .A1(n6160), .A2(n6151), .ZN(n7790) );
  NAND2_X1 U7807 ( .A1(n7790), .A2(n4448), .ZN(n6155) );
  NAND2_X1 U7808 ( .A1(n9057), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7809 ( .A1(n9058), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7810 ( .A1(n9059), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6152) );
  OR2_X1 U7811 ( .A1(n9818), .A2(n9095), .ZN(n9174) );
  NAND2_X1 U7812 ( .A1(n6156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6157) );
  XNOR2_X1 U7813 ( .A(n6157), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9378) );
  AOI22_X1 U7814 ( .A1(n9378), .A2(n6424), .B1(n9066), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n6158) );
  INV_X1 U7815 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7816 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  AND2_X1 U7817 ( .A1(n4297), .A2(n6161), .ZN(n9711) );
  NAND2_X1 U7818 ( .A1(n9711), .A2(n4448), .ZN(n6166) );
  NAND2_X1 U7819 ( .A1(n9059), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7820 ( .A1(n9057), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6162) );
  AND2_X1 U7821 ( .A1(n6163), .A2(n6162), .ZN(n6165) );
  NAND2_X1 U7822 ( .A1(n9058), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7823 ( .A1(n9814), .A2(n9098), .ZN(n9177) );
  NAND2_X1 U7824 ( .A1(n6476), .A2(n6091), .ZN(n6176) );
  NAND2_X1 U7825 ( .A1(n6173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6172) );
  MUX2_X1 U7826 ( .A(n6172), .B(P1_IR_REG_31__SCAN_IN), .S(n6181), .Z(n6174)
         );
  INV_X1 U7827 ( .A(n6173), .ZN(n6184) );
  NAND2_X1 U7828 ( .A1(n6174), .A2(n4365), .ZN(n9393) );
  INV_X1 U7829 ( .A(n9393), .ZN(n9389) );
  AOI22_X1 U7830 ( .A1(n9066), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6424), .B2(
        n9389), .ZN(n6175) );
  INV_X1 U7831 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10234) );
  AND2_X1 U7832 ( .A1(n4297), .A2(n10234), .ZN(n6177) );
  OR2_X1 U7833 ( .A1(n6177), .A2(n6188), .ZN(n9692) );
  AOI22_X1 U7834 ( .A1(n9057), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n9059), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7835 ( .A1(n9058), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6178) );
  OAI211_X1 U7836 ( .C1(n9692), .C2(n6278), .A(n6179), .B(n6178), .ZN(n9704)
         );
  INV_X1 U7837 ( .A(n9704), .ZN(n9655) );
  NAND2_X1 U7838 ( .A1(n9807), .A2(n9655), .ZN(n9178) );
  NAND2_X1 U7839 ( .A1(n9683), .A2(n9684), .ZN(n9682) );
  NAND2_X1 U7840 ( .A1(n6482), .A2(n6091), .ZN(n6187) );
  NAND2_X1 U7841 ( .A1(n4365), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6180) );
  MUX2_X1 U7842 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6180), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n6185) );
  INV_X1 U7843 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7844 ( .A1(n6184), .A2(n6183), .ZN(n6192) );
  NAND2_X1 U7845 ( .A1(n6185), .A2(n6192), .ZN(n9415) );
  INV_X1 U7846 ( .A(n9415), .ZN(n9400) );
  AOI22_X1 U7847 ( .A1(n9066), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6424), .B2(
        n9400), .ZN(n6186) );
  NOR2_X1 U7848 ( .A1(n6188), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6189) );
  OR2_X1 U7849 ( .A1(n6195), .A2(n6189), .ZN(n9668) );
  AOI22_X1 U7850 ( .A1(n9057), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8046), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7851 ( .A1(n9059), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6190) );
  OAI211_X1 U7852 ( .C1(n9668), .C2(n6278), .A(n6191), .B(n6190), .ZN(n9686)
         );
  INV_X1 U7853 ( .A(n9686), .ZN(n9631) );
  OR2_X1 U7854 ( .A1(n9673), .A2(n9631), .ZN(n9182) );
  NAND2_X1 U7855 ( .A1(n9673), .A2(n9631), .ZN(n9168) );
  NAND2_X1 U7856 ( .A1(n9182), .A2(n9168), .ZN(n9650) );
  NAND2_X1 U7857 ( .A1(n6570), .A2(n6091), .ZN(n6194) );
  XNOR2_X1 U7858 ( .A(n6204), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9429) );
  AOI22_X1 U7859 ( .A1(n9066), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6424), .B2(
        n9429), .ZN(n6193) );
  OR2_X1 U7860 ( .A1(n6195), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6196) );
  AND2_X1 U7861 ( .A1(n6222), .A2(n6196), .ZN(n9641) );
  NAND2_X1 U7862 ( .A1(n9641), .A2(n4448), .ZN(n6201) );
  INV_X1 U7863 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U7864 ( .A1(n8046), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7865 ( .A1(n9059), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6197) );
  OAI211_X1 U7866 ( .C1(n6282), .C2(n9406), .A(n6198), .B(n6197), .ZN(n6199)
         );
  INV_X1 U7867 ( .A(n6199), .ZN(n6200) );
  NAND2_X1 U7868 ( .A1(n6789), .A2(n6091), .ZN(n6206) );
  NAND2_X1 U7869 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n6203) );
  XNOR2_X1 U7870 ( .A(n6213), .B(n4939), .ZN(n9911) );
  AOI22_X1 U7871 ( .A1(n9066), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6424), .B2(
        n9911), .ZN(n6205) );
  XNOR2_X1 U7872 ( .A(n6222), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U7873 ( .A1(n9623), .A2(n4448), .ZN(n6212) );
  INV_X1 U7874 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7875 ( .A1(n9059), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7876 ( .A1(n8046), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6207) );
  OAI211_X1 U7877 ( .C1(n6282), .C2(n6209), .A(n6208), .B(n6207), .ZN(n6210)
         );
  INV_X1 U7878 ( .A(n6210), .ZN(n6211) );
  OR2_X1 U7879 ( .A1(n9642), .A2(n9657), .ZN(n9611) );
  NAND2_X1 U7880 ( .A1(n9612), .A2(n9187), .ZN(n9595) );
  NAND2_X1 U7881 ( .A1(n9595), .A2(n9594), .ZN(n6230) );
  NAND2_X1 U7882 ( .A1(n6873), .A2(n6091), .ZN(n6218) );
  INV_X1 U7883 ( .A(n6304), .ZN(n6215) );
  NAND2_X1 U7884 ( .A1(n6215), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n6216) );
  AOI22_X1 U7885 ( .A1(n9164), .A2(n6424), .B1(n9066), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n6217) );
  INV_X1 U7886 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6220) );
  INV_X1 U7887 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6219) );
  OAI21_X1 U7888 ( .B1(n6222), .B2(n6220), .A(n6219), .ZN(n6223) );
  NAND2_X1 U7889 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6221) );
  OR2_X2 U7890 ( .A1(n6222), .A2(n6221), .ZN(n6233) );
  NAND2_X1 U7891 ( .A1(n6223), .A2(n6233), .ZN(n9601) );
  OR2_X1 U7892 ( .A1(n9601), .A2(n6278), .ZN(n6229) );
  INV_X1 U7893 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7894 ( .A1(n9059), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7895 ( .A1(n9058), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6224) );
  OAI211_X1 U7896 ( .C1(n6282), .C2(n6226), .A(n6225), .B(n6224), .ZN(n6227)
         );
  INV_X1 U7897 ( .A(n6227), .ZN(n6228) );
  OR2_X1 U7898 ( .A1(n9785), .A2(n9615), .ZN(n9124) );
  NAND2_X1 U7899 ( .A1(n9785), .A2(n9615), .ZN(n9201) );
  NAND2_X1 U7900 ( .A1(n7117), .A2(n6091), .ZN(n6232) );
  NAND2_X1 U7901 ( .A1(n6286), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6231) );
  INV_X1 U7902 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U7903 ( .A1(n6233), .A2(n8999), .ZN(n6234) );
  NAND2_X1 U7904 ( .A1(n4296), .A2(n6234), .ZN(n9000) );
  INV_X1 U7905 ( .A(n9000), .ZN(n9586) );
  NAND2_X1 U7906 ( .A1(n9586), .A2(n4448), .ZN(n6239) );
  INV_X1 U7907 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10191) );
  NAND2_X1 U7908 ( .A1(n9057), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7909 ( .A1(n9058), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6235) );
  OAI211_X1 U7910 ( .C1(n10191), .C2(n6086), .A(n6236), .B(n6235), .ZN(n6237)
         );
  INV_X1 U7911 ( .A(n6237), .ZN(n6238) );
  OR2_X1 U7912 ( .A1(n9587), .A2(n9562), .ZN(n9245) );
  INV_X1 U7913 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8944) );
  AND2_X2 U7914 ( .A1(n6251), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6257) );
  NOR2_X1 U7915 ( .A1(n6251), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6242) );
  OR2_X1 U7916 ( .A1(n6257), .A2(n6242), .ZN(n9550) );
  INV_X1 U7917 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7918 ( .A1(n9059), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7919 ( .A1(n8046), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6243) );
  OAI211_X1 U7920 ( .C1(n6282), .C2(n6245), .A(n6244), .B(n6243), .ZN(n6246)
         );
  INV_X1 U7921 ( .A(n6246), .ZN(n6247) );
  INV_X1 U7922 ( .A(n9244), .ZN(n9217) );
  NAND2_X1 U7923 ( .A1(n7219), .A2(n6091), .ZN(n6249) );
  NAND2_X1 U7924 ( .A1(n6286), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6248) );
  AND2_X1 U7925 ( .A1(n4296), .A2(n8944), .ZN(n6250) );
  NOR2_X1 U7926 ( .A1(n6251), .A2(n6250), .ZN(n9570) );
  INV_X1 U7927 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U7928 ( .A1(n9059), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7929 ( .A1(n9058), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6252) );
  OAI211_X1 U7930 ( .C1(n6282), .C2(n9777), .A(n6253), .B(n6252), .ZN(n6254)
         );
  AOI21_X2 U7931 ( .B1(n9570), .B2(n4448), .A(n6254), .ZN(n9578) );
  OR2_X2 U7932 ( .A1(n9571), .A2(n9578), .ZN(n9545) );
  NAND2_X1 U7933 ( .A1(n9571), .A2(n9578), .ZN(n9142) );
  NAND2_X1 U7934 ( .A1(n6286), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6255) );
  AND2_X2 U7935 ( .A1(n6257), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6267) );
  NOR2_X1 U7936 ( .A1(n6257), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6258) );
  NOR2_X1 U7937 ( .A1(n6267), .A2(n6258), .ZN(n9527) );
  NAND2_X1 U7938 ( .A1(n9527), .A2(n4448), .ZN(n6264) );
  INV_X1 U7939 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U7940 ( .A1(n9057), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7941 ( .A1(n9059), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6259) );
  OAI211_X1 U7942 ( .C1(n6261), .C2(n6070), .A(n6260), .B(n6259), .ZN(n6262)
         );
  INV_X1 U7943 ( .A(n6262), .ZN(n6263) );
  NAND2_X1 U7944 ( .A1(n9761), .A2(n9548), .ZN(n9145) );
  NAND2_X1 U7945 ( .A1(n6286), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6265) );
  OR2_X1 U7946 ( .A1(n6267), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7947 ( .A1(n9520), .A2(n4448), .ZN(n6273) );
  INV_X1 U7948 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10189) );
  NAND2_X1 U7949 ( .A1(n9057), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7950 ( .A1(n9059), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6269) );
  OAI211_X1 U7951 ( .C1(n10189), .C2(n6070), .A(n6270), .B(n6269), .ZN(n6271)
         );
  INV_X1 U7952 ( .A(n6271), .ZN(n6272) );
  NAND2_X1 U7953 ( .A1(n7798), .A2(n6091), .ZN(n6275) );
  NAND2_X1 U7954 ( .A1(n6286), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6274) );
  INV_X1 U7955 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U7956 ( .A1(n6276), .A2(n8954), .ZN(n6277) );
  NAND2_X1 U7957 ( .A1(n6277), .A2(n4298), .ZN(n9505) );
  INV_X1 U7958 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7959 ( .A1(n9058), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7960 ( .A1(n9059), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6279) );
  OAI211_X1 U7961 ( .C1(n6282), .C2(n6281), .A(n6280), .B(n6279), .ZN(n6283)
         );
  INV_X1 U7962 ( .A(n6283), .ZN(n6284) );
  AND2_X2 U7963 ( .A1(n9501), .A2(n9340), .ZN(n9147) );
  NAND2_X1 U7964 ( .A1(n6286), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7965 ( .A1(n9059), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U7966 ( .A1(n9057), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6291) );
  INV_X1 U7967 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9031) );
  NOR2_X2 U7968 ( .A1(n4298), .A2(n9031), .ZN(n6295) );
  AOI21_X1 U7969 ( .B1(n9031), .B2(n4298), .A(n6295), .ZN(n9491) );
  NAND2_X1 U7970 ( .A1(n4448), .A2(n9491), .ZN(n6290) );
  NAND2_X1 U7971 ( .A1(n9058), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7972 ( .A1(n9066), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7973 ( .A1(n9059), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7974 ( .A1(n9057), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7975 ( .A1(n6295), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U7976 ( .A1(n4448), .A2(n6296), .ZN(n6298) );
  NAND2_X1 U7977 ( .A1(n9058), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6297) );
  OR2_X2 U7978 ( .A1(n9474), .A2(n9488), .ZN(n9457) );
  XNOR2_X1 U7979 ( .A(n8043), .B(n6301), .ZN(n6315) );
  NAND2_X1 U7980 ( .A1(n6302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6303) );
  INV_X1 U7981 ( .A(n6311), .ZN(n6306) );
  INV_X1 U7982 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7983 ( .A1(n6306), .A2(n6305), .ZN(n6312) );
  NAND2_X1 U7984 ( .A1(n6312), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6307) );
  XNOR2_X1 U7985 ( .A(n6307), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U7986 ( .A1(n6379), .A2(n9164), .ZN(n6314) );
  XNOR2_X2 U7987 ( .A(n6310), .B(n6309), .ZN(n9276) );
  INV_X1 U7988 ( .A(n9276), .ZN(n6983) );
  NAND2_X1 U7989 ( .A1(n6311), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U7990 ( .A1(n6983), .A2(n9284), .ZN(n6313) );
  NAND2_X1 U7991 ( .A1(n6315), .A2(n9708), .ZN(n6326) );
  NAND2_X1 U7992 ( .A1(n9057), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U7993 ( .A1(n9059), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6321) );
  INV_X1 U7994 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U7995 ( .A1(n8932), .A2(n6316), .ZN(n6318) );
  INV_X1 U7996 ( .A(n6316), .ZN(n6317) );
  AND2_X2 U7997 ( .A1(n6318), .A2(n8037), .ZN(n9469) );
  NAND2_X1 U7998 ( .A1(n4448), .A2(n9469), .ZN(n6320) );
  NAND2_X1 U7999 ( .A1(n9058), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6319) );
  AND4_X2 U8000 ( .A1(n6322), .A2(n6321), .A3(n6320), .A4(n6319), .ZN(n8903)
         );
  AND2_X1 U8001 ( .A1(n6595), .A2(n6729), .ZN(n9703) );
  INV_X1 U8002 ( .A(n6729), .ZN(n6579) );
  NOR2_X1 U8003 ( .A1(n9500), .A2(n9654), .ZN(n6324) );
  NAND2_X1 U8004 ( .A1(n6326), .A2(n6325), .ZN(n9480) );
  INV_X1 U8005 ( .A(n7414), .ZN(n9999) );
  INV_X1 U8006 ( .A(n7640), .ZN(n7248) );
  INV_X1 U8007 ( .A(n9824), .ZN(n7608) );
  INV_X1 U8008 ( .A(n9818), .ZN(n7792) );
  INV_X1 U8009 ( .A(n9642), .ZN(n9797) );
  INV_X1 U8010 ( .A(n9587), .ZN(n9779) );
  AND2_X2 U8011 ( .A1(n9526), .A2(n9517), .ZN(n9518) );
  OR2_X2 U8012 ( .A1(n9503), .A2(n9742), .ZN(n9489) );
  NAND2_X1 U8013 ( .A1(n6984), .A2(n9276), .ZN(n10000) );
  AOI21_X1 U8014 ( .B1(n9489), .B2(n9474), .A(n10000), .ZN(n6328) );
  AND2_X1 U8015 ( .A1(n9465), .A2(n6328), .ZN(n9479) );
  NAND2_X1 U8016 ( .A1(n9276), .A2(n9440), .ZN(n6384) );
  INV_X1 U8017 ( .A(n7008), .ZN(n6332) );
  NAND2_X1 U8018 ( .A1(n6754), .A2(n9249), .ZN(n6337) );
  NAND2_X1 U8019 ( .A1(n6335), .A2(n6755), .ZN(n6336) );
  NAND2_X1 U8020 ( .A1(n6337), .A2(n6336), .ZN(n7048) );
  NAND2_X1 U8021 ( .A1(n7048), .A2(n6338), .ZN(n6341) );
  NAND2_X1 U8022 ( .A1(n6339), .A2(n4860), .ZN(n6340) );
  NAND2_X1 U8023 ( .A1(n7061), .A2(n7062), .ZN(n6343) );
  NAND2_X1 U8024 ( .A1(n7284), .A2(n9972), .ZN(n6342) );
  NAND2_X1 U8025 ( .A1(n7292), .A2(n9353), .ZN(n7078) );
  AND2_X2 U8026 ( .A1(n9205), .A2(n9207), .ZN(n7287) );
  OR2_X1 U8027 ( .A1(n9352), .A2(n7089), .ZN(n6345) );
  NAND2_X1 U8028 ( .A1(n6346), .A2(n6345), .ZN(n7313) );
  INV_X1 U8029 ( .A(n7423), .ZN(n9351) );
  INV_X1 U8030 ( .A(n7712), .ZN(n9349) );
  NAND2_X1 U8031 ( .A1(n9087), .A2(n9081), .ZN(n7334) );
  INV_X1 U8032 ( .A(n7570), .ZN(n9350) );
  NAND2_X1 U8033 ( .A1(n7414), .A2(n9350), .ZN(n7241) );
  NAND2_X1 U8034 ( .A1(n7241), .A2(n7712), .ZN(n6350) );
  INV_X1 U8035 ( .A(n7241), .ZN(n6349) );
  AOI22_X1 U8036 ( .A1(n7640), .A2(n6350), .B1(n6349), .B2(n9349), .ZN(n6351)
         );
  INV_X1 U8037 ( .A(n7644), .ZN(n9348) );
  OR2_X1 U8038 ( .A1(n6327), .A2(n9348), .ZN(n6353) );
  NAND2_X1 U8039 ( .A1(n7361), .A2(n9347), .ZN(n7354) );
  NOR2_X1 U8040 ( .A1(n7361), .A2(n9347), .ZN(n7356) );
  NAND2_X1 U8041 ( .A1(n7610), .A2(n9248), .ZN(n7609) );
  NAND2_X1 U8042 ( .A1(n9824), .A2(n9346), .ZN(n6354) );
  AND2_X1 U8043 ( .A1(n9818), .A2(n9706), .ZN(n6355) );
  OR2_X1 U8044 ( .A1(n9818), .A2(n9706), .ZN(n6356) );
  OR2_X1 U8045 ( .A1(n9807), .A2(n9704), .ZN(n6357) );
  NAND2_X1 U8046 ( .A1(n9807), .A2(n9704), .ZN(n6358) );
  NAND2_X1 U8047 ( .A1(n6359), .A2(n6358), .ZN(n9661) );
  NAND2_X1 U8048 ( .A1(n9661), .A2(n9650), .ZN(n6361) );
  NAND2_X1 U8049 ( .A1(n9673), .A2(n9686), .ZN(n6360) );
  AND2_X1 U8050 ( .A1(n9642), .A2(n9345), .ZN(n6362) );
  INV_X1 U8051 ( .A(n6362), .ZN(n6363) );
  OR2_X1 U8052 ( .A1(n9642), .A2(n9345), .ZN(n6365) );
  OR2_X1 U8053 ( .A1(n9785), .A2(n9344), .ZN(n6366) );
  NAND2_X1 U8054 ( .A1(n9605), .A2(n6366), .ZN(n6368) );
  NAND2_X1 U8055 ( .A1(n9785), .A2(n9344), .ZN(n6367) );
  NAND2_X1 U8056 ( .A1(n6368), .A2(n6367), .ZN(n9581) );
  AND2_X1 U8057 ( .A1(n9587), .A2(n9598), .ZN(n6369) );
  NAND2_X1 U8058 ( .A1(n9554), .A2(n9534), .ZN(n6370) );
  OAI21_X1 U8059 ( .B1(n9535), .B2(n9517), .A(n9512), .ZN(n6375) );
  NAND2_X1 U8060 ( .A1(n6375), .A2(n6374), .ZN(n9497) );
  NAND2_X1 U8061 ( .A1(n9484), .A2(n6376), .ZN(n6377) );
  NAND2_X1 U8062 ( .A1(n6377), .A2(n5037), .ZN(n8033) );
  XOR2_X1 U8063 ( .A(n9316), .B(n6378), .Z(n9483) );
  NAND2_X1 U8064 ( .A1(n6379), .A2(n9440), .ZN(n6380) );
  NAND2_X2 U8065 ( .A1(n9276), .A2(n9284), .ZN(n6586) );
  CLKBUF_X3 U8066 ( .A(n6710), .Z(n8927) );
  AND2_X1 U8067 ( .A1(n8927), .A2(n9440), .ZN(n6381) );
  INV_X1 U8068 ( .A(n6384), .ZN(n9324) );
  NAND2_X1 U8069 ( .A1(n6595), .A2(n9324), .ZN(n9331) );
  NAND2_X1 U8070 ( .A1(n6381), .A2(n9331), .ZN(n9689) );
  AND2_X1 U8071 ( .A1(n9276), .A2(n9164), .ZN(n9323) );
  NAND2_X1 U8072 ( .A1(n9323), .A2(n7301), .ZN(n9811) );
  NAND2_X1 U8073 ( .A1(n6595), .A2(n6384), .ZN(n6733) );
  INV_X1 U8074 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6398) );
  INV_X1 U8075 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6394) );
  INV_X1 U8076 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6390) );
  XNOR2_X2 U8077 ( .A(n6389), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7876) );
  OR2_X1 U8078 ( .A1(n6391), .A2(n6390), .ZN(n6392) );
  NAND2_X1 U8079 ( .A1(n6393), .A2(n6392), .ZN(n6403) );
  XNOR2_X1 U8080 ( .A(n6395), .B(n6394), .ZN(n7760) );
  NOR2_X1 U8081 ( .A1(n6403), .A2(n7760), .ZN(n6396) );
  NAND2_X1 U8082 ( .A1(n6397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6399) );
  XNOR2_X1 U8083 ( .A(n6399), .B(n6398), .ZN(n7598) );
  AND2_X1 U8084 ( .A1(n7598), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6400) );
  NAND2_X1 U8085 ( .A1(n6984), .A2(n9323), .ZN(n6981) );
  INV_X1 U8086 ( .A(n7876), .ZN(n6416) );
  NAND3_X1 U8087 ( .A1(n6403), .A2(P1_B_REG_SCAN_IN), .A3(n7760), .ZN(n6401)
         );
  OAI21_X1 U8088 ( .B1(P1_B_REG_SCAN_IN), .B2(n7760), .A(n6401), .ZN(n6402) );
  INV_X1 U8089 ( .A(n6403), .ZN(n7799) );
  OAI22_X1 U8090 ( .A1(n6411), .A2(P1_D_REG_1__SCAN_IN), .B1(n7876), .B2(n7799), .ZN(n6573) );
  NOR4_X1 U8091 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6407) );
  NOR4_X1 U8092 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6406) );
  NOR4_X1 U8093 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6405) );
  NOR4_X1 U8094 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6404) );
  NAND4_X1 U8095 ( .A1(n6407), .A2(n6406), .A3(n6405), .A4(n6404), .ZN(n6413)
         );
  NOR4_X1 U8096 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10134) );
  NOR2_X1 U8097 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n6410) );
  NOR4_X1 U8098 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6409) );
  NOR4_X1 U8099 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6408) );
  NAND4_X1 U8100 ( .A1(n10134), .A2(n6410), .A3(n6409), .A4(n6408), .ZN(n6412)
         );
  OAI21_X1 U8101 ( .B1(n6413), .B2(n6412), .A(n9848), .ZN(n6572) );
  AND2_X1 U8102 ( .A1(n6573), .A2(n6572), .ZN(n6414) );
  INV_X1 U8103 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8104 ( .A1(n9848), .A2(n6415), .ZN(n6417) );
  NAND2_X1 U8105 ( .A1(n6416), .A2(n7760), .ZN(n9850) );
  AND3_X2 U8106 ( .A1(n6980), .A2(n6638), .A3(n6575), .ZN(n10017) );
  NAND2_X1 U8107 ( .A1(n9740), .A2(n10017), .ZN(n6420) );
  INV_X1 U8108 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6418) );
  INV_X1 U8109 ( .A(n7598), .ZN(n6421) );
  OR2_X1 U8110 ( .A1(n6731), .A2(n6421), .ZN(n6484) );
  INV_X1 U8111 ( .A(n9336), .ZN(P1_U4006) );
  INV_X1 U8112 ( .A(n7042), .ZN(n6422) );
  NAND2_X1 U8113 ( .A1(n6595), .A2(n7598), .ZN(n6423) );
  NAND2_X1 U8114 ( .A1(n6423), .A2(n6484), .ZN(n6506) );
  OAI21_X1 U8115 ( .B1(n6506), .B2(n6424), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  INV_X1 U8116 ( .A(n6425), .ZN(n6441) );
  AND2_X1 U8117 ( .A1(n9054), .A2(P2_U3152), .ZN(n8795) );
  AND2_X1 U8118 ( .A1(n4807), .A2(P2_U3152), .ZN(n8793) );
  AOI22_X1 U8119 ( .A1(n6856), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8793), .ZN(n6426) );
  OAI21_X1 U8120 ( .B1(n6441), .B2(n4275), .A(n6426), .ZN(P2_U3353) );
  INV_X1 U8121 ( .A(n6427), .ZN(n6442) );
  AOI22_X1 U8122 ( .A1(n6891), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8793), .ZN(n6428) );
  OAI21_X1 U8123 ( .B1(n6442), .B2(n4275), .A(n6428), .ZN(P2_U3351) );
  INV_X1 U8124 ( .A(n8793), .ZN(n8802) );
  INV_X1 U8125 ( .A(n6429), .ZN(n6438) );
  OAI222_X1 U8126 ( .A1(n8802), .A2(n4515), .B1(n4275), .B2(n6438), .C1(
        P2_U3152), .C2(n6837), .ZN(P2_U3354) );
  OAI222_X1 U8127 ( .A1(n8802), .A2(n6430), .B1(n4275), .B2(n6439), .C1(
        P2_U3152), .C2(n8286), .ZN(P2_U3355) );
  NAND2_X1 U8128 ( .A1(n9849), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6431) );
  OAI21_X1 U8129 ( .B1(n9849), .B2(n6573), .A(n6431), .ZN(P1_U3441) );
  OAI222_X1 U8130 ( .A1(n6663), .A2(P2_U3152), .B1(n4275), .B2(n6444), .C1(
        n4413), .C2(n8802), .ZN(P2_U3357) );
  OAI222_X1 U8131 ( .A1(n6661), .A2(P2_U3152), .B1(n4275), .B2(n6446), .C1(
        n6432), .C2(n8802), .ZN(P2_U3356) );
  INV_X1 U8132 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10236) );
  INV_X1 U8133 ( .A(n6433), .ZN(n6436) );
  OAI222_X1 U8134 ( .A1(n8802), .A2(n10236), .B1(n4275), .B2(n6436), .C1(
        P2_U3152), .C2(n8302), .ZN(P2_U3352) );
  INV_X1 U8135 ( .A(n6434), .ZN(n6448) );
  AOI22_X1 U8136 ( .A1(n8317), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n8793), .ZN(n6435) );
  OAI21_X1 U8137 ( .B1(n6448), .B2(n4275), .A(n6435), .ZN(P2_U3350) );
  NOR2_X1 U8138 ( .A1(n5245), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9864) );
  INV_X1 U8139 ( .A(n9864), .ZN(n7758) );
  INV_X1 U8140 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6437) );
  OAI222_X1 U8141 ( .A1(n7758), .A2(n6437), .B1(n9866), .B2(n6436), .C1(
        P1_U3084), .C2(n6523), .ZN(P1_U3347) );
  INV_X1 U8142 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10120) );
  OAI222_X1 U8143 ( .A1(n7758), .A2(n10120), .B1(n9866), .B2(n6438), .C1(
        P1_U3084), .C2(n6521), .ZN(P1_U3349) );
  INV_X1 U8144 ( .A(n6520), .ZN(n6564) );
  OAI222_X1 U8145 ( .A1(n7758), .A2(n6440), .B1(n9866), .B2(n6439), .C1(
        P1_U3084), .C2(n6564), .ZN(P1_U3350) );
  OAI222_X1 U8146 ( .A1(n7758), .A2(n4485), .B1(n9866), .B2(n6441), .C1(
        P1_U3084), .C2(n6522), .ZN(P1_U3348) );
  INV_X1 U8147 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6443) );
  INV_X1 U8148 ( .A(n6524), .ZN(n6532) );
  OAI222_X1 U8149 ( .A1(n7758), .A2(n6443), .B1(n9866), .B2(n6442), .C1(
        P1_U3084), .C2(n6532), .ZN(P1_U3346) );
  INV_X1 U8150 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6445) );
  INV_X1 U8151 ( .A(n6518), .ZN(n6512) );
  OAI222_X1 U8152 ( .A1(n7758), .A2(n6445), .B1(n9866), .B2(n6444), .C1(
        P1_U3084), .C2(n6512), .ZN(P1_U3352) );
  INV_X1 U8153 ( .A(n6519), .ZN(n6626) );
  OAI222_X1 U8154 ( .A1(n7758), .A2(n6447), .B1(n9866), .B2(n6446), .C1(
        P1_U3084), .C2(n6626), .ZN(P1_U3351) );
  OAI222_X1 U8155 ( .A1(n7758), .A2(n6449), .B1(n9866), .B2(n6448), .C1(
        P1_U3084), .C2(n6541), .ZN(P1_U3345) );
  INV_X1 U8156 ( .A(n6450), .ZN(n6462) );
  AOI22_X1 U8157 ( .A1(n8330), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8793), .ZN(n6451) );
  OAI21_X1 U8158 ( .B1(n6462), .B2(n4275), .A(n6451), .ZN(P2_U3349) );
  INV_X1 U8159 ( .A(n6452), .ZN(n6464) );
  AOI22_X1 U8160 ( .A1(n8344), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8793), .ZN(n6453) );
  OAI21_X1 U8161 ( .B1(n6464), .B2(n4275), .A(n6453), .ZN(P2_U3348) );
  INV_X1 U8162 ( .A(n6454), .ZN(n6460) );
  INV_X1 U8163 ( .A(n7275), .ZN(n7272) );
  INV_X1 U8164 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6455) );
  OAI222_X1 U8165 ( .A1(n9866), .A2(n6460), .B1(n7272), .B2(P1_U3084), .C1(
        n6455), .C2(n7758), .ZN(P1_U3342) );
  INV_X1 U8166 ( .A(n6456), .ZN(n6458) );
  INV_X1 U8167 ( .A(n7387), .ZN(n7273) );
  OAI222_X1 U8168 ( .A1(n7758), .A2(n6457), .B1(n9866), .B2(n6458), .C1(
        P1_U3084), .C2(n7273), .ZN(P1_U3341) );
  OAI222_X1 U8169 ( .A1(n8802), .A2(n6459), .B1(n4275), .B2(n6458), .C1(
        P2_U3152), .C2(n6917), .ZN(P2_U3346) );
  INV_X1 U8170 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6461) );
  INV_X1 U8171 ( .A(n6913), .ZN(n6888) );
  OAI222_X1 U8172 ( .A1(n8802), .A2(n6461), .B1(n4275), .B2(n6460), .C1(n6888), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8173 ( .A(n6767), .ZN(n6545) );
  OAI222_X1 U8174 ( .A1(n7758), .A2(n6463), .B1(n6545), .B2(P1_U3084), .C1(
        n9866), .C2(n6462), .ZN(P1_U3344) );
  INV_X1 U8175 ( .A(n6816), .ZN(n6809) );
  OAI222_X1 U8176 ( .A1(n7758), .A2(n6465), .B1(n6809), .B2(P1_U3084), .C1(
        n9866), .C2(n6464), .ZN(P1_U3343) );
  NAND2_X1 U8177 ( .A1(n8398), .A2(P2_U3966), .ZN(n6466) );
  OAI21_X1 U8178 ( .B1(n5686), .B2(P2_U3966), .A(n6466), .ZN(P2_U3583) );
  INV_X1 U8179 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8180 ( .A1(n4483), .A2(P2_U3966), .ZN(n6467) );
  OAI21_X1 U8181 ( .B1(n6468), .B2(P2_U3966), .A(n6467), .ZN(P2_U3552) );
  INV_X1 U8182 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6470) );
  INV_X1 U8183 ( .A(n6469), .ZN(n6471) );
  INV_X1 U8184 ( .A(n6919), .ZN(n6969) );
  OAI222_X1 U8185 ( .A1(n8802), .A2(n6470), .B1(n4275), .B2(n6471), .C1(n6969), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8186 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10194) );
  INV_X1 U8187 ( .A(n9365), .ZN(n9359) );
  OAI222_X1 U8188 ( .A1(n7758), .A2(n10194), .B1(n9359), .B2(P1_U3084), .C1(
        n9866), .C2(n6471), .ZN(P1_U3340) );
  OAI21_X1 U8189 ( .B1(n10031), .B2(n5871), .A(n6472), .ZN(n6475) );
  NAND2_X1 U8190 ( .A1(n10031), .A2(n6473), .ZN(n6474) );
  NOR2_X1 U8191 ( .A1(n8366), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8192 ( .A(n6476), .ZN(n6477) );
  OAI222_X1 U8193 ( .A1(n7758), .A2(n10197), .B1(n9866), .B2(n6477), .C1(
        P1_U3084), .C2(n9393), .ZN(P1_U3338) );
  INV_X1 U8194 ( .A(n7209), .ZN(n7142) );
  OAI222_X1 U8195 ( .A1(n8802), .A2(n6478), .B1(n4275), .B2(n6477), .C1(
        P2_U3152), .C2(n7142), .ZN(P2_U3343) );
  INV_X1 U8196 ( .A(n6479), .ZN(n6480) );
  INV_X1 U8197 ( .A(n7136), .ZN(n7130) );
  OAI222_X1 U8198 ( .A1(n8802), .A2(n10183), .B1(n4275), .B2(n6480), .C1(n7130), .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8199 ( .A(n9378), .ZN(n9366) );
  OAI222_X1 U8200 ( .A1(n7758), .A2(n6481), .B1(n9366), .B2(P1_U3084), .C1(
        n9866), .C2(n6480), .ZN(P1_U3339) );
  INV_X1 U8201 ( .A(n6482), .ZN(n6555) );
  AOI22_X1 U8202 ( .A1(n7624), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8793), .ZN(n6483) );
  OAI21_X1 U8203 ( .B1(n6555), .B2(n4275), .A(n6483), .ZN(P2_U3342) );
  INV_X1 U8204 ( .A(P1_U3083), .ZN(n6485) );
  NAND2_X1 U8205 ( .A1(n6485), .A2(n6484), .ZN(n9442) );
  INV_X1 U8206 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U8207 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6490) );
  XOR2_X1 U8208 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6518), .Z(n6486) );
  INV_X1 U8209 ( .A(n6486), .ZN(n6489) );
  INV_X1 U8210 ( .A(n6510), .ZN(n6488) );
  NOR2_X1 U8211 ( .A1(n6729), .A2(P1_U3084), .ZN(n9860) );
  NAND2_X1 U8212 ( .A1(n9860), .A2(n6613), .ZN(n6487) );
  AOI211_X1 U8213 ( .C1(n6490), .C2(n6489), .A(n6488), .B(n9923), .ZN(n6496)
         );
  NAND2_X1 U8214 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6615) );
  XNOR2_X1 U8215 ( .A(n6518), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6491) );
  NOR2_X1 U8216 ( .A1(n6491), .A2(n6615), .ZN(n6517) );
  INV_X1 U8217 ( .A(n6613), .ZN(n8044) );
  NAND2_X1 U8218 ( .A1(n9860), .A2(n8044), .ZN(n9329) );
  AOI211_X1 U8219 ( .C1(n6615), .C2(n6491), .A(n6517), .B(n9438), .ZN(n6495)
         );
  NOR2_X1 U8220 ( .A1(n6613), .A2(P1_U3084), .ZN(n9863) );
  NAND2_X1 U8221 ( .A1(n9863), .A2(n6729), .ZN(n6492) );
  INV_X1 U8222 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6493) );
  OAI22_X1 U8223 ( .A1(n9918), .A2(n6512), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6493), .ZN(n6494) );
  NOR3_X1 U8224 ( .A1(n6496), .A2(n6495), .A3(n6494), .ZN(n6497) );
  OAI21_X1 U8225 ( .B1(n9442), .B2(n6498), .A(n6497), .ZN(P1_U3242) );
  INV_X1 U8226 ( .A(n9442), .ZN(n9927) );
  INV_X1 U8227 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7096) );
  NAND2_X1 U8228 ( .A1(n8044), .A2(n7096), .ZN(n6499) );
  NAND2_X1 U8229 ( .A1(n6579), .A2(n6499), .ZN(n6503) );
  INV_X1 U8230 ( .A(n9860), .ZN(n6501) );
  INV_X1 U8231 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6591) );
  INV_X1 U8232 ( .A(n9863), .ZN(n6500) );
  OAI21_X1 U8233 ( .B1(n6501), .B2(n6591), .A(n6500), .ZN(n6502) );
  NAND2_X1 U8234 ( .A1(n6503), .A2(n6587), .ZN(n6616) );
  OAI211_X1 U8235 ( .C1(n6503), .C2(n6587), .A(n6502), .B(n6616), .ZN(n6505)
         );
  INV_X1 U8236 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6504) );
  OAI22_X1 U8237 ( .A1(n6506), .A2(n6505), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6504), .ZN(n6508) );
  NOR3_X1 U8238 ( .A1(n9923), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6587), .ZN(
        n6507) );
  AOI211_X1 U8239 ( .C1(n9927), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n6508), .B(
        n6507), .ZN(n6509) );
  INV_X1 U8240 ( .A(n6509), .ZN(P1_U3241) );
  XNOR2_X1 U8241 ( .A(n6541), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6543) );
  INV_X1 U8242 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10116) );
  INV_X1 U8243 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6516) );
  INV_X1 U8244 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6515) );
  INV_X1 U8245 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6514) );
  INV_X1 U8246 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6513) );
  INV_X1 U8247 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6511) );
  XOR2_X1 U8248 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6519), .Z(n6624) );
  NAND2_X1 U8249 ( .A1(n6623), .A2(n6624), .ZN(n6622) );
  OAI21_X1 U8250 ( .B1(n6626), .B2(n6513), .A(n6622), .ZN(n6561) );
  XOR2_X1 U8251 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6520), .Z(n6562) );
  XOR2_X1 U8252 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6521), .Z(n6607) );
  NOR2_X1 U8253 ( .A1(n6606), .A2(n6607), .ZN(n6605) );
  XNOR2_X1 U8254 ( .A(n6522), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6703) );
  OAI21_X1 U8255 ( .B1(n6522), .B2(n6516), .A(n6701), .ZN(n6676) );
  XNOR2_X1 U8256 ( .A(n6684), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6677) );
  NOR2_X1 U8257 ( .A1(n6676), .A2(n6677), .ZN(n6675) );
  XNOR2_X1 U8258 ( .A(n6524), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6531) );
  OAI22_X1 U8259 ( .A1(n6530), .A2(n6531), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n6524), .ZN(n6544) );
  XOR2_X1 U8260 ( .A(n6544), .B(n6543), .Z(n6529) );
  INV_X1 U8261 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7321) );
  INV_X1 U8262 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7085) );
  INV_X1 U8263 ( .A(n6521), .ZN(n6612) );
  XNOR2_X1 U8264 ( .A(n6519), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6620) );
  XNOR2_X1 U8265 ( .A(n6520), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6558) );
  NOR2_X1 U8266 ( .A1(n6559), .A2(n6558), .ZN(n6557) );
  XNOR2_X1 U8267 ( .A(n6521), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6603) );
  XNOR2_X1 U8268 ( .A(n6522), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6700) );
  INV_X1 U8269 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7290) );
  XNOR2_X1 U8270 ( .A(n6523), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U8271 ( .A1(n6680), .A2(n6679), .ZN(n6678) );
  OAI21_X1 U8272 ( .B1(n6523), .B2(n7085), .A(n6678), .ZN(n6534) );
  XNOR2_X1 U8273 ( .A(n6524), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6535) );
  XNOR2_X1 U8274 ( .A(n6546), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6547) );
  XNOR2_X1 U8275 ( .A(n6548), .B(n6547), .ZN(n6525) );
  INV_X1 U8276 ( .A(n9438), .ZN(n9913) );
  NAND2_X1 U8277 ( .A1(n6525), .A2(n9913), .ZN(n6528) );
  AND2_X1 U8278 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3084), .ZN(n7425) );
  NOR2_X1 U8279 ( .A1(n9918), .A2(n6541), .ZN(n6526) );
  AOI211_X1 U8280 ( .C1(n9927), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n7425), .B(
        n6526), .ZN(n6527) );
  OAI211_X1 U8281 ( .C1(n6529), .C2(n9923), .A(n6528), .B(n6527), .ZN(P1_U3249) );
  XOR2_X1 U8282 ( .A(n6530), .B(n6531), .Z(n6540) );
  NAND2_X1 U8283 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7569) );
  OAI21_X1 U8284 ( .B1(n9918), .B2(n6532), .A(n7569), .ZN(n6538) );
  AOI21_X1 U8285 ( .B1(n6535), .B2(n6534), .A(n6533), .ZN(n6536) );
  NOR2_X1 U8286 ( .A1(n6536), .A2(n9438), .ZN(n6537) );
  AOI211_X1 U8287 ( .C1(n9927), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n6538), .B(
        n6537), .ZN(n6539) );
  OAI21_X1 U8288 ( .B1(n9923), .B2(n6540), .A(n6539), .ZN(P1_U3248) );
  XNOR2_X1 U8289 ( .A(n6767), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n6763) );
  INV_X1 U8290 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6542) );
  AOI22_X1 U8291 ( .A1(n6544), .A2(n6543), .B1(n6542), .B2(n6541), .ZN(n6764)
         );
  XOR2_X1 U8292 ( .A(n6764), .B(n6763), .Z(n6554) );
  NAND2_X1 U8293 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7642) );
  OAI21_X1 U8294 ( .B1(n9918), .B2(n6545), .A(n7642), .ZN(n6552) );
  XNOR2_X1 U8295 ( .A(n6767), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6550) );
  OAI22_X1 U8296 ( .A1(n6548), .A2(n6547), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6546), .ZN(n6549) );
  AOI211_X1 U8297 ( .C1(n6550), .C2(n6549), .A(n9438), .B(n6766), .ZN(n6551)
         );
  AOI211_X1 U8298 ( .C1(n9927), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n6552), .B(
        n6551), .ZN(n6553) );
  OAI21_X1 U8299 ( .B1(n9923), .B2(n6554), .A(n6553), .ZN(P1_U3250) );
  OAI222_X1 U8300 ( .A1(n7758), .A2(n6556), .B1(n9415), .B2(P1_U3084), .C1(
        n9866), .C2(n6555), .ZN(P1_U3337) );
  INV_X1 U8301 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6569) );
  AOI211_X1 U8302 ( .C1(n6559), .C2(n6558), .A(n6557), .B(n9438), .ZN(n6567)
         );
  INV_X1 U8303 ( .A(n9923), .ZN(n9410) );
  OAI211_X1 U8304 ( .C1(n6562), .C2(n6561), .A(n9410), .B(n6560), .ZN(n6563)
         );
  INV_X1 U8305 ( .A(n6563), .ZN(n6566) );
  NAND2_X1 U8306 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3084), .ZN(n6728) );
  OAI21_X1 U8307 ( .B1(n9918), .B2(n6564), .A(n6728), .ZN(n6565) );
  NOR3_X1 U8308 ( .A1(n6567), .A2(n6566), .A3(n6565), .ZN(n6568) );
  OAI21_X1 U8309 ( .B1(n9442), .B2(n6569), .A(n6568), .ZN(P1_U3244) );
  INV_X1 U8310 ( .A(n6570), .ZN(n6641) );
  AOI22_X1 U8311 ( .A1(n9429), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9864), .ZN(n6571) );
  OAI21_X1 U8312 ( .B1(n6641), .B2(n9866), .A(n6571), .ZN(P1_U3336) );
  INV_X1 U8313 ( .A(n6572), .ZN(n6574) );
  OR2_X1 U8314 ( .A1(n6574), .A2(n6573), .ZN(n6978) );
  NOR2_X1 U8315 ( .A1(n6978), .A2(n6575), .ZN(n6597) );
  INV_X1 U8316 ( .A(n6597), .ZN(n6576) );
  NAND2_X1 U8317 ( .A1(n6576), .A2(n6981), .ZN(n6735) );
  AND2_X1 U8318 ( .A1(n6735), .A2(n6577), .ZN(n7646) );
  INV_X1 U8319 ( .A(n7092), .ZN(n6998) );
  NOR2_X1 U8320 ( .A1(n9331), .A2(n9849), .ZN(n6578) );
  NAND2_X1 U8321 ( .A1(n6597), .A2(n6578), .ZN(n6730) );
  INV_X1 U8322 ( .A(n9048), .ZN(n9019) );
  NAND2_X1 U8323 ( .A1(n6735), .A2(n6980), .ZN(n6750) );
  AOI22_X1 U8324 ( .A1(n9019), .A2(n9357), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6750), .ZN(n6600) );
  INV_X1 U8325 ( .A(n6312), .ZN(n6580) );
  NAND2_X1 U8326 ( .A1(n6580), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6584) );
  INV_X1 U8327 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6581) );
  OAI21_X1 U8328 ( .B1(n6582), .B2(n6581), .A(n6312), .ZN(n6583) );
  NAND2_X1 U8329 ( .A1(n6797), .A2(n6334), .ZN(n6590) );
  OR2_X2 U8330 ( .A1(n6586), .A2(n6585), .ZN(n6715) );
  OAI22_X1 U8331 ( .A1(n8892), .A2(n6998), .B1(n6731), .B2(n6587), .ZN(n6588)
         );
  INV_X1 U8332 ( .A(n6588), .ZN(n6589) );
  AND2_X1 U8333 ( .A1(n6590), .A2(n6589), .ZN(n6594) );
  OR2_X1 U8334 ( .A1(n6731), .A2(n6591), .ZN(n6593) );
  OAI211_X2 U8335 ( .C1(n7004), .C2(n8892), .A(n6593), .B(n6592), .ZN(n6711)
         );
  OAI21_X1 U8336 ( .B1(n6594), .B2(n6711), .A(n6712), .ZN(n6614) );
  NOR2_X1 U8337 ( .A1(n6595), .A2(n9849), .ZN(n6596) );
  AND2_X1 U8338 ( .A1(n6596), .A2(n9998), .ZN(n6598) );
  NAND2_X1 U8339 ( .A1(n6614), .A2(n9043), .ZN(n6599) );
  OAI211_X1 U8340 ( .C1(n9053), .C2(n6998), .A(n6600), .B(n6599), .ZN(P1_U3230) );
  INV_X1 U8341 ( .A(n9918), .ZN(n9418) );
  NAND2_X1 U8342 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n6801) );
  INV_X1 U8343 ( .A(n6801), .ZN(n6611) );
  OAI21_X1 U8344 ( .B1(n6603), .B2(n6602), .A(n6601), .ZN(n6604) );
  INV_X1 U8345 ( .A(n6604), .ZN(n6609) );
  AOI21_X1 U8346 ( .B1(n6607), .B2(n6606), .A(n6605), .ZN(n6608) );
  OAI22_X1 U8347 ( .A1(n6609), .A2(n9438), .B1(n6608), .B2(n9923), .ZN(n6610)
         );
  AOI211_X1 U8348 ( .C1(n9418), .C2(n6612), .A(n6611), .B(n6610), .ZN(n6618)
         );
  MUX2_X1 U8349 ( .A(n6615), .B(n6614), .S(n6613), .Z(n6617) );
  OAI211_X1 U8350 ( .C1(n6617), .C2(n6729), .A(P1_U4006), .B(n6616), .ZN(n6631) );
  OAI211_X1 U8351 ( .C1(n9874), .C2(n9442), .A(n6618), .B(n6631), .ZN(P1_U3245) );
  INV_X1 U8352 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6632) );
  AOI211_X1 U8353 ( .C1(n6621), .C2(n6620), .A(n6619), .B(n9438), .ZN(n6629)
         );
  OAI211_X1 U8354 ( .C1(n6624), .C2(n6623), .A(n9410), .B(n6622), .ZN(n6625)
         );
  INV_X1 U8355 ( .A(n6625), .ZN(n6628) );
  OAI22_X1 U8356 ( .A1(n9918), .A2(n6626), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n4669), .ZN(n6627) );
  NOR3_X1 U8357 ( .A1(n6629), .A2(n6628), .A3(n6627), .ZN(n6630) );
  OAI211_X1 U8358 ( .C1(n6632), .C2(n9442), .A(n6631), .B(n6630), .ZN(P1_U3243) );
  NOR2_X1 U8359 ( .A1(n7004), .A2(n7092), .ZN(n9283) );
  INV_X1 U8360 ( .A(n6634), .ZN(n7003) );
  INV_X1 U8361 ( .A(n6984), .ZN(n6635) );
  OAI211_X1 U8362 ( .C1(n9283), .C2(n7003), .A(n9331), .B(n6635), .ZN(n6636)
         );
  OAI21_X1 U8363 ( .B1(n6633), .B2(n9656), .A(n6636), .ZN(n7093) );
  AOI21_X1 U8364 ( .B1(n7092), .B2(n6984), .A(n7093), .ZN(n6640) );
  INV_X1 U8365 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10149) );
  NAND2_X1 U8366 ( .A1(n10015), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6637) );
  OAI21_X1 U8367 ( .B1(n6640), .B2(n10015), .A(n6637), .ZN(P1_U3454) );
  AND3_X2 U8368 ( .A1(n6980), .A2(n6638), .A3(n6977), .ZN(n10029) );
  NAND2_X1 U8369 ( .A1(n10026), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6639) );
  OAI21_X1 U8370 ( .B1(n6640), .B2(n10026), .A(n6639), .ZN(P1_U3523) );
  INV_X1 U8371 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6642) );
  INV_X1 U8372 ( .A(n8361), .ZN(n7622) );
  OAI222_X1 U8373 ( .A1(n8802), .A2(n6642), .B1(n4275), .B2(n6641), .C1(n7622), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U8374 ( .A1(n10031), .A2(n7024), .ZN(n6645) );
  OR2_X1 U8375 ( .A1(n6658), .A2(P2_U3152), .ZN(n8796) );
  OAI21_X1 U8376 ( .B1(n7042), .B2(n8796), .A(n7630), .ZN(n6643) );
  INV_X1 U8377 ( .A(n6643), .ZN(n6644) );
  NAND2_X1 U8378 ( .A1(n6645), .A2(n6644), .ZN(n6652) );
  NAND2_X1 U8379 ( .A1(n6652), .A2(n6650), .ZN(n6646) );
  NAND2_X1 U8380 ( .A1(n6646), .A2(n8257), .ZN(n6660) );
  NAND2_X1 U8381 ( .A1(n6660), .A2(n6658), .ZN(n8382) );
  NAND2_X1 U8382 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7185) );
  INV_X1 U8383 ( .A(n7185), .ZN(n6657) );
  XNOR2_X1 U8384 ( .A(n6837), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6654) );
  XNOR2_X1 U8385 ( .A(n6661), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n8279) );
  XNOR2_X1 U8386 ( .A(n6663), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n8269) );
  AND2_X1 U8387 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8268) );
  NAND2_X1 U8388 ( .A1(n8269), .A2(n8268), .ZN(n8267) );
  INV_X1 U8389 ( .A(n6663), .ZN(n8263) );
  NAND2_X1 U8390 ( .A1(n8263), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U8391 ( .A1(n8267), .A2(n6647), .ZN(n8278) );
  NAND2_X1 U8392 ( .A1(n8279), .A2(n8278), .ZN(n8277) );
  INV_X1 U8393 ( .A(n6661), .ZN(n8274) );
  NAND2_X1 U8394 ( .A1(n8274), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U8395 ( .A1(n8277), .A2(n6648), .ZN(n8293) );
  XNOR2_X1 U8396 ( .A(n8286), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n8294) );
  NAND2_X1 U8397 ( .A1(n8293), .A2(n8294), .ZN(n8292) );
  INV_X1 U8398 ( .A(n8286), .ZN(n8284) );
  NAND2_X1 U8399 ( .A1(n8284), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U8400 ( .A1(n8292), .A2(n6649), .ZN(n6653) );
  AND2_X1 U8401 ( .A1(n6650), .A2(n8800), .ZN(n6651) );
  NAND2_X1 U8402 ( .A1(n6652), .A2(n6651), .ZN(n8383) );
  NAND2_X1 U8403 ( .A1(n6653), .A2(n6654), .ZN(n6829) );
  OAI211_X1 U8404 ( .C1(n6654), .C2(n6653), .A(n8386), .B(n6829), .ZN(n6655)
         );
  INV_X1 U8405 ( .A(n6655), .ZN(n6656) );
  AOI211_X1 U8406 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n8366), .A(n6657), .B(
        n6656), .ZN(n6674) );
  NOR2_X1 U8407 ( .A1(n6658), .A2(n8800), .ZN(n6659) );
  INV_X1 U8408 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6662) );
  MUX2_X1 U8409 ( .A(n6662), .B(P2_REG2_REG_2__SCAN_IN), .S(n6661), .Z(n8276)
         );
  XNOR2_X1 U8410 ( .A(n6663), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n8266) );
  AND2_X1 U8411 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n8265) );
  NAND2_X1 U8412 ( .A1(n8266), .A2(n8265), .ZN(n8264) );
  NAND2_X1 U8413 ( .A1(n8263), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U8414 ( .A1(n8264), .A2(n6664), .ZN(n8275) );
  NAND2_X1 U8415 ( .A1(n8274), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U8416 ( .A1(n8288), .A2(n8287), .ZN(n6667) );
  INV_X1 U8417 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6665) );
  MUX2_X1 U8418 ( .A(n6665), .B(P2_REG2_REG_3__SCAN_IN), .S(n8286), .Z(n6666)
         );
  NAND2_X1 U8419 ( .A1(n6667), .A2(n6666), .ZN(n8291) );
  NAND2_X1 U8420 ( .A1(n8284), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8421 ( .A1(n8291), .A2(n6671), .ZN(n6669) );
  INV_X1 U8422 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6836) );
  MUX2_X1 U8423 ( .A(n6836), .B(P2_REG2_REG_4__SCAN_IN), .S(n6837), .Z(n6668)
         );
  MUX2_X1 U8424 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6836), .S(n6837), .Z(n6670)
         );
  NAND3_X1 U8425 ( .A1(n8291), .A2(n6671), .A3(n6670), .ZN(n6672) );
  NAND3_X1 U8426 ( .A1(n8388), .A2(n6841), .A3(n6672), .ZN(n6673) );
  OAI211_X1 U8427 ( .C1(n8382), .C2(n6837), .A(n6674), .B(n6673), .ZN(P2_U3249) );
  INV_X1 U8428 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6686) );
  AND2_X1 U8429 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7351) );
  AOI21_X1 U8430 ( .B1(n6677), .B2(n6676), .A(n6675), .ZN(n6682) );
  OAI211_X1 U8431 ( .C1(n6680), .C2(n6679), .A(n6678), .B(n9913), .ZN(n6681)
         );
  OAI21_X1 U8432 ( .B1(n6682), .B2(n9923), .A(n6681), .ZN(n6683) );
  AOI211_X1 U8433 ( .C1(n9418), .C2(n6684), .A(n7351), .B(n6683), .ZN(n6685)
         );
  OAI21_X1 U8434 ( .B1(n9442), .B2(n6686), .A(n6685), .ZN(P1_U3247) );
  AND2_X1 U8435 ( .A1(n6777), .A2(n6687), .ZN(n7431) );
  INV_X1 U8436 ( .A(n7431), .ZN(n6689) );
  NOR2_X1 U8437 ( .A1(n7534), .A2(n8605), .ZN(n7098) );
  AOI21_X1 U8438 ( .B1(n8614), .B2(n6689), .A(n7098), .ZN(n7430) );
  INV_X1 U8439 ( .A(n7430), .ZN(n6691) );
  OAI22_X1 U8440 ( .A1(n7431), .A2(n8767), .B1(n7018), .B2(n7102), .ZN(n6690)
         );
  NOR2_X1 U8441 ( .A1(n6691), .A2(n6690), .ZN(n10039) );
  OR2_X1 U8442 ( .A1(n6692), .A2(n7037), .ZN(n6693) );
  NOR2_X1 U8443 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  NAND2_X1 U8444 ( .A1(n7014), .A2(n6695), .ZN(n6696) );
  NAND2_X1 U8445 ( .A1(n10081), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6697) );
  OAI21_X1 U8446 ( .B1(n10039), .B2(n10081), .A(n6697), .ZN(P2_U3520) );
  INV_X1 U8447 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6709) );
  NOR2_X1 U8448 ( .A1(n6698), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7262) );
  XOR2_X1 U8449 ( .A(n6700), .B(n6699), .Z(n6705) );
  OAI211_X1 U8450 ( .C1(n6703), .C2(n6702), .A(n9410), .B(n6701), .ZN(n6704)
         );
  OAI21_X1 U8451 ( .B1(n6705), .B2(n9438), .A(n6704), .ZN(n6706) );
  AOI211_X1 U8452 ( .C1(n9418), .C2(n6707), .A(n7262), .B(n6706), .ZN(n6708)
         );
  OAI21_X1 U8453 ( .B1(n9442), .B2(n6709), .A(n6708), .ZN(P1_U3246) );
  OR2_X2 U8454 ( .A1(n6711), .A2(n8880), .ZN(n6713) );
  NAND2_X1 U8455 ( .A1(n6713), .A2(n6712), .ZN(n6742) );
  XNOR2_X1 U8456 ( .A(n6714), .B(n8927), .ZN(n6744) );
  BUF_X2 U8457 ( .A(n6715), .Z(n8832) );
  OAI22_X1 U8458 ( .A1(n6727), .A2(n6633), .B1(n6716), .B2(n8832), .ZN(n6741)
         );
  NAND2_X1 U8459 ( .A1(n6744), .A2(n6741), .ZN(n6717) );
  NAND2_X1 U8460 ( .A1(n6742), .A2(n6717), .ZN(n6719) );
  OR2_X1 U8461 ( .A1(n6741), .A2(n6744), .ZN(n6718) );
  XNOR2_X1 U8462 ( .A(n6720), .B(n8880), .ZN(n6723) );
  OAI22_X1 U8463 ( .A1(n6727), .A2(n6335), .B1(n6755), .B2(n8832), .ZN(n6721)
         );
  INV_X1 U8464 ( .A(n6721), .ZN(n6722) );
  NAND2_X1 U8465 ( .A1(n6723), .A2(n6722), .ZN(n6724) );
  XNOR2_X1 U8466 ( .A(n6726), .B(n8880), .ZN(n6795) );
  OAI22_X1 U8467 ( .A1(n6727), .A2(n6339), .B1(n4860), .B2(n8832), .ZN(n6793)
         );
  XOR2_X1 U8468 ( .A(n6792), .B(n6791), .Z(n6740) );
  OAI21_X1 U8469 ( .B1(n9048), .B2(n7284), .A(n6728), .ZN(n6738) );
  NAND2_X1 U8470 ( .A1(n6731), .A2(n7598), .ZN(n9330) );
  INV_X1 U8471 ( .A(n9330), .ZN(n6732) );
  AND2_X1 U8472 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  NAND2_X1 U8473 ( .A1(n6735), .A2(n6734), .ZN(n6736) );
  NAND2_X1 U8474 ( .A1(n6736), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9047) );
  OAI22_X1 U8475 ( .A1(n6335), .A2(n9032), .B1(n9047), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n6737) );
  AOI211_X1 U8476 ( .C1(n9022), .C2(n7053), .A(n6738), .B(n6737), .ZN(n6739)
         );
  OAI21_X1 U8477 ( .B1(n6740), .B2(n9024), .A(n6739), .ZN(P1_U3216) );
  XNOR2_X1 U8478 ( .A(n6742), .B(n6741), .ZN(n6743) );
  XNOR2_X1 U8479 ( .A(n6744), .B(n6743), .ZN(n6747) );
  AOI22_X1 U8480 ( .A1(n9019), .A2(n9356), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6750), .ZN(n6746) );
  AOI22_X1 U8481 ( .A1(n9022), .A2(n9956), .B1(n9050), .B2(n6334), .ZN(n6745)
         );
  OAI211_X1 U8482 ( .C1(n6747), .C2(n9024), .A(n6746), .B(n6745), .ZN(P1_U3220) );
  XOR2_X1 U8483 ( .A(n6748), .B(n6749), .Z(n6753) );
  AOI22_X1 U8484 ( .A1(n9019), .A2(n9355), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6750), .ZN(n6752) );
  AOI22_X1 U8485 ( .A1(n9022), .A2(n6993), .B1(n9050), .B2(n9357), .ZN(n6751)
         );
  OAI211_X1 U8486 ( .C1(n6753), .C2(n9024), .A(n6752), .B(n6751), .ZN(P1_U3235) );
  INV_X1 U8487 ( .A(n9811), .ZN(n10005) );
  XOR2_X1 U8488 ( .A(n6754), .B(n9249), .Z(n6989) );
  INV_X1 U8489 ( .A(n6989), .ZN(n6761) );
  OAI211_X1 U8490 ( .C1(n6755), .C2(n7008), .A(n10008), .B(n7049), .ZN(n6990)
         );
  OAI21_X1 U8491 ( .B1(n6755), .B2(n9998), .A(n6990), .ZN(n6760) );
  XNOR2_X1 U8492 ( .A(n6756), .B(n9249), .ZN(n6758) );
  OAI22_X1 U8493 ( .A1(n9656), .A2(n6339), .B1(n6633), .B2(n9654), .ZN(n6757)
         );
  AOI21_X1 U8494 ( .B1(n6758), .B2(n9708), .A(n6757), .ZN(n6759) );
  OAI21_X1 U8495 ( .B1(n6989), .B2(n9689), .A(n6759), .ZN(n6982) );
  AOI211_X1 U8496 ( .C1(n10005), .C2(n6761), .A(n6760), .B(n6982), .ZN(n9964)
         );
  NAND2_X1 U8497 ( .A1(n10026), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6762) );
  OAI21_X1 U8498 ( .B1(n9964), .B2(n10026), .A(n6762), .ZN(P1_U3525) );
  XOR2_X1 U8499 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6816), .Z(n6811) );
  OAI22_X1 U8500 ( .A1(n6764), .A2(n6763), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6767), .ZN(n6812) );
  XOR2_X1 U8501 ( .A(n6812), .B(n6811), .Z(n6773) );
  AND2_X1 U8502 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7714) );
  INV_X1 U8503 ( .A(n7714), .ZN(n6765) );
  OAI21_X1 U8504 ( .B1(n9918), .B2(n6809), .A(n6765), .ZN(n6771) );
  XNOR2_X1 U8505 ( .A(n6816), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6768) );
  AOI211_X1 U8506 ( .C1(n6769), .C2(n6768), .A(n9438), .B(n6815), .ZN(n6770)
         );
  AOI211_X1 U8507 ( .C1(n9927), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n6771), .B(
        n6770), .ZN(n6772) );
  OAI21_X1 U8508 ( .B1(n9923), .B2(n6773), .A(n6772), .ZN(P1_U3251) );
  INV_X1 U8509 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6788) );
  OAI21_X1 U8510 ( .B1(n6774), .B2(n6776), .A(n6775), .ZN(n7583) );
  INV_X1 U8511 ( .A(n6777), .ZN(n6781) );
  NOR2_X1 U8512 ( .A1(n6779), .A2(n6778), .ZN(n6780) );
  AOI211_X1 U8513 ( .C1(n6781), .C2(n6774), .A(n8535), .B(n6780), .ZN(n6784)
         );
  OR2_X1 U8514 ( .A1(n4467), .A2(n8605), .ZN(n6783) );
  NAND2_X1 U8515 ( .A1(n4483), .A2(n8580), .ZN(n6782) );
  NAND2_X1 U8516 ( .A1(n6783), .A2(n6782), .ZN(n7023) );
  NOR2_X1 U8517 ( .A1(n6784), .A2(n7023), .ZN(n7577) );
  INV_X1 U8518 ( .A(n7576), .ZN(n6785) );
  AOI21_X1 U8519 ( .B1(n8762), .B2(n7580), .A(n6785), .ZN(n6786) );
  OAI211_X1 U8520 ( .C1(n8767), .C2(n7583), .A(n7577), .B(n6786), .ZN(n6930)
         );
  NAND2_X1 U8521 ( .A1(n6930), .A2(n10076), .ZN(n6787) );
  OAI21_X1 U8522 ( .B1(n10076), .B2(n6788), .A(n6787), .ZN(P2_U3454) );
  INV_X1 U8523 ( .A(n6789), .ZN(n6807) );
  AOI22_X1 U8524 ( .A1(n9911), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9864), .ZN(n6790) );
  OAI21_X1 U8525 ( .B1(n6807), .B2(n9866), .A(n6790), .ZN(P1_U3335) );
  INV_X1 U8526 ( .A(n6793), .ZN(n6794) );
  NAND2_X1 U8527 ( .A1(n6795), .A2(n6794), .ZN(n6796) );
  OAI22_X1 U8528 ( .A1(n6727), .A2(n7284), .B1(n9972), .B2(n8832), .ZN(n7253)
         );
  OAI22_X1 U8529 ( .A1(n7284), .A2(n8832), .B1(n6725), .B2(n9972), .ZN(n6798)
         );
  XNOR2_X1 U8530 ( .A(n6798), .B(n8927), .ZN(n7254) );
  XOR2_X1 U8531 ( .A(n7253), .B(n7254), .Z(n6799) );
  XNOR2_X1 U8532 ( .A(n7256), .B(n6799), .ZN(n6805) );
  OAI22_X1 U8533 ( .A1(n6339), .A2(n9032), .B1(n9047), .B2(n7067), .ZN(n6804)
         );
  NAND2_X1 U8534 ( .A1(n9022), .A2(n7073), .ZN(n6802) );
  OAI211_X1 U8535 ( .C1(n6800), .C2(n9048), .A(n6802), .B(n6801), .ZN(n6803)
         );
  AOI211_X1 U8536 ( .C1(n6805), .C2(n9043), .A(n6804), .B(n6803), .ZN(n6806)
         );
  INV_X1 U8537 ( .A(n6806), .ZN(P1_U3228) );
  INV_X1 U8538 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6808) );
  OAI222_X1 U8539 ( .A1(n8802), .A2(n6808), .B1(n4275), .B2(n6807), .C1(
        P2_U3152), .C2(n8368), .ZN(P2_U3340) );
  INV_X1 U8540 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9908) );
  MUX2_X1 U8541 ( .A(n9908), .B(P1_REG1_REG_11__SCAN_IN), .S(n7275), .Z(n6814)
         );
  INV_X1 U8542 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6810) );
  NOR2_X1 U8543 ( .A1(n6813), .A2(n6814), .ZN(n7271) );
  AOI21_X1 U8544 ( .B1(n6814), .B2(n6813), .A(n7271), .ZN(n6825) );
  XNOR2_X1 U8545 ( .A(n7272), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n6818) );
  NAND2_X1 U8546 ( .A1(n6817), .A2(n6818), .ZN(n7274) );
  OAI21_X1 U8547 ( .B1(n6818), .B2(n6817), .A(n7274), .ZN(n6819) );
  NAND2_X1 U8548 ( .A1(n6819), .A2(n9913), .ZN(n6824) );
  NOR2_X1 U8549 ( .A1(n6820), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7525) );
  INV_X1 U8550 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6821) );
  NOR2_X1 U8551 ( .A1(n9442), .A2(n6821), .ZN(n6822) );
  AOI211_X1 U8552 ( .C1(n9418), .C2(n7275), .A(n7525), .B(n6822), .ZN(n6823)
         );
  OAI211_X1 U8553 ( .C1(n6825), .C2(n9923), .A(n6824), .B(n6823), .ZN(P1_U3252) );
  INV_X1 U8554 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6826) );
  XNOR2_X1 U8555 ( .A(n6856), .B(n6826), .ZN(n6831) );
  INV_X1 U8556 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6827) );
  OR2_X1 U8557 ( .A1(n6837), .A2(n6827), .ZN(n6828) );
  NAND2_X1 U8558 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  NAND2_X1 U8559 ( .A1(n6830), .A2(n6831), .ZN(n6848) );
  OAI21_X1 U8560 ( .B1(n6831), .B2(n6830), .A(n6848), .ZN(n6832) );
  NOR2_X1 U8561 ( .A1(n8383), .A2(n6832), .ZN(n6835) );
  INV_X1 U8562 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U8563 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7175) );
  OAI21_X1 U8564 ( .B1(n8395), .B2(n6833), .A(n7175), .ZN(n6834) );
  AOI211_X1 U8565 ( .C1(n8342), .C2(n6856), .A(n6835), .B(n6834), .ZN(n6845)
         );
  OR2_X1 U8566 ( .A1(n6837), .A2(n6836), .ZN(n6840) );
  NAND2_X1 U8567 ( .A1(n6841), .A2(n6840), .ZN(n6839) );
  INV_X1 U8568 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7372) );
  MUX2_X1 U8569 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7372), .S(n6856), .Z(n6838)
         );
  NAND2_X1 U8570 ( .A1(n6839), .A2(n6838), .ZN(n8304) );
  MUX2_X1 U8571 ( .A(n7372), .B(P2_REG2_REG_5__SCAN_IN), .S(n6856), .Z(n6842)
         );
  NAND3_X1 U8572 ( .A1(n6842), .A2(n6841), .A3(n6840), .ZN(n6843) );
  NAND3_X1 U8573 ( .A1(n8388), .A2(n8304), .A3(n6843), .ZN(n6844) );
  NAND2_X1 U8574 ( .A1(n6845), .A2(n6844), .ZN(P2_U3250) );
  INV_X1 U8575 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6846) );
  XNOR2_X1 U8576 ( .A(n6891), .B(n6846), .ZN(n6851) );
  NAND2_X1 U8577 ( .A1(n6856), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6847) );
  NAND2_X1 U8578 ( .A1(n6848), .A2(n6847), .ZN(n8309) );
  XNOR2_X1 U8579 ( .A(n8302), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U8580 ( .A1(n8309), .A2(n8310), .ZN(n8308) );
  NAND2_X1 U8581 ( .A1(n8299), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U8582 ( .A1(n8308), .A2(n6849), .ZN(n6850) );
  NAND2_X1 U8583 ( .A1(n6850), .A2(n6851), .ZN(n6893) );
  OAI21_X1 U8584 ( .B1(n6851), .B2(n6850), .A(n6893), .ZN(n6852) );
  NOR2_X1 U8585 ( .A1(n8383), .A2(n6852), .ZN(n6855) );
  INV_X1 U8586 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U8587 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7307) );
  OAI21_X1 U8588 ( .B1(n8395), .B2(n6853), .A(n7307), .ZN(n6854) );
  AOI211_X1 U8589 ( .C1(n8342), .C2(n6891), .A(n6855), .B(n6854), .ZN(n6865)
         );
  NAND2_X1 U8590 ( .A1(n6856), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U8591 ( .A1(n8304), .A2(n8303), .ZN(n6858) );
  INV_X1 U8592 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7441) );
  MUX2_X1 U8593 ( .A(n7441), .B(P2_REG2_REG_6__SCAN_IN), .S(n8302), .Z(n6857)
         );
  NAND2_X1 U8594 ( .A1(n6858), .A2(n6857), .ZN(n8307) );
  NAND2_X1 U8595 ( .A1(n8299), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6862) );
  NAND2_X1 U8596 ( .A1(n8307), .A2(n6862), .ZN(n6860) );
  INV_X1 U8597 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7552) );
  MUX2_X1 U8598 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7552), .S(n6891), .Z(n6859)
         );
  MUX2_X1 U8599 ( .A(n7552), .B(P2_REG2_REG_7__SCAN_IN), .S(n6891), .Z(n6861)
         );
  NAND3_X1 U8600 ( .A1(n8307), .A2(n6862), .A3(n6861), .ZN(n6863) );
  NAND3_X1 U8601 ( .A1(n8388), .A2(n8320), .A3(n6863), .ZN(n6864) );
  NAND2_X1 U8602 ( .A1(n6865), .A2(n6864), .ZN(P2_U3252) );
  AOI22_X1 U8603 ( .A1(n8388), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n8386), .ZN(n6870) );
  INV_X1 U8604 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U8605 ( .A1(n8388), .A2(n6866), .ZN(n6867) );
  OAI211_X1 U8606 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n8383), .A(n6867), .B(
        n8382), .ZN(n6868) );
  INV_X1 U8607 ( .A(n6868), .ZN(n6869) );
  MUX2_X1 U8608 ( .A(n6870), .B(n6869), .S(P2_IR_REG_0__SCAN_IN), .Z(n6872) );
  AOI22_X1 U8609 ( .A1(n8366), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n6871) );
  NAND2_X1 U8610 ( .A1(n6872), .A2(n6871), .ZN(P2_U3245) );
  INV_X1 U8611 ( .A(n6873), .ZN(n6874) );
  OAI222_X1 U8612 ( .A1(n8802), .A2(n10180), .B1(n4275), .B2(n6874), .C1(
        P2_U3152), .C2(n8390), .ZN(P2_U3339) );
  OAI222_X1 U8613 ( .A1(n7758), .A2(n6875), .B1(n9866), .B2(n6874), .C1(n9440), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  MUX2_X1 U8614 ( .A(n4418), .B(P2_REG2_REG_11__SCAN_IN), .S(n6913), .Z(n6887)
         );
  NAND2_X1 U8615 ( .A1(n6891), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U8616 ( .A1(n8320), .A2(n8319), .ZN(n6878) );
  INV_X1 U8617 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6876) );
  MUX2_X1 U8618 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6876), .S(n8317), .Z(n6877)
         );
  NAND2_X1 U8619 ( .A1(n6878), .A2(n6877), .ZN(n8333) );
  NAND2_X1 U8620 ( .A1(n8317), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U8621 ( .A1(n8333), .A2(n8332), .ZN(n6881) );
  INV_X1 U8622 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6879) );
  MUX2_X1 U8623 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6879), .S(n8330), .Z(n6880)
         );
  NAND2_X1 U8624 ( .A1(n8330), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U8625 ( .A1(n8347), .A2(n8346), .ZN(n6883) );
  INV_X1 U8626 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7773) );
  MUX2_X1 U8627 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7773), .S(n8344), .Z(n6882)
         );
  NAND2_X1 U8628 ( .A1(n6883), .A2(n6882), .ZN(n8349) );
  NAND2_X1 U8629 ( .A1(n8344), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U8630 ( .A1(n8349), .A2(n6884), .ZN(n6886) );
  INV_X1 U8631 ( .A(n6915), .ZN(n6885) );
  AOI21_X1 U8632 ( .B1(n6887), .B2(n6886), .A(n6885), .ZN(n6904) );
  NOR2_X1 U8633 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7815), .ZN(n6890) );
  NOR2_X1 U8634 ( .A1(n8382), .A2(n6888), .ZN(n6889) );
  AOI211_X1 U8635 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n8366), .A(n6890), .B(
        n6889), .ZN(n6903) );
  NAND2_X1 U8636 ( .A1(n6891), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8637 ( .A1(n6893), .A2(n6892), .ZN(n8323) );
  XNOR2_X1 U8638 ( .A(n8317), .B(n10082), .ZN(n8324) );
  NAND2_X1 U8639 ( .A1(n8323), .A2(n8324), .ZN(n8322) );
  NAND2_X1 U8640 ( .A1(n8317), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U8641 ( .A1(n8322), .A2(n6894), .ZN(n8336) );
  INV_X1 U8642 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6895) );
  XNOR2_X1 U8643 ( .A(n8330), .B(n6895), .ZN(n8337) );
  NAND2_X1 U8644 ( .A1(n8336), .A2(n8337), .ZN(n8335) );
  NAND2_X1 U8645 ( .A1(n8330), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8646 ( .A1(n8335), .A2(n6896), .ZN(n8351) );
  INV_X1 U8647 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6897) );
  XNOR2_X1 U8648 ( .A(n8344), .B(n6897), .ZN(n8352) );
  NAND2_X1 U8649 ( .A1(n8351), .A2(n8352), .ZN(n8350) );
  NAND2_X1 U8650 ( .A1(n8344), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U8651 ( .A1(n8350), .A2(n6898), .ZN(n6901) );
  INV_X1 U8652 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6899) );
  XNOR2_X1 U8653 ( .A(n6913), .B(n6899), .ZN(n6900) );
  NAND2_X1 U8654 ( .A1(n6901), .A2(n6900), .ZN(n6906) );
  OAI211_X1 U8655 ( .C1(n6901), .C2(n6900), .A(n6906), .B(n8386), .ZN(n6902)
         );
  OAI211_X1 U8656 ( .C1(n6904), .C2(n8372), .A(n6903), .B(n6902), .ZN(P2_U3256) );
  INV_X1 U8657 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10182) );
  XNOR2_X1 U8658 ( .A(n7136), .B(n10182), .ZN(n7138) );
  NAND2_X1 U8659 ( .A1(n6913), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U8660 ( .A1(n6906), .A2(n6905), .ZN(n6952) );
  INV_X1 U8661 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6907) );
  XNOR2_X1 U8662 ( .A(n6917), .B(n6907), .ZN(n6953) );
  NAND2_X1 U8663 ( .A1(n6917), .A2(n6907), .ZN(n6908) );
  NAND2_X1 U8664 ( .A1(n6950), .A2(n6908), .ZN(n6972) );
  INV_X1 U8665 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6909) );
  XNOR2_X1 U8666 ( .A(n6919), .B(n6909), .ZN(n6971) );
  NAND2_X1 U8667 ( .A1(n6972), .A2(n6971), .ZN(n6911) );
  OR2_X1 U8668 ( .A1(n6919), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8669 ( .A1(n6911), .A2(n6910), .ZN(n7139) );
  XOR2_X1 U8670 ( .A(n7138), .B(n7139), .Z(n6929) );
  INV_X1 U8671 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8672 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8074) );
  OAI21_X1 U8673 ( .B1(n8395), .B2(n6912), .A(n8074), .ZN(n6927) );
  OR2_X1 U8674 ( .A1(n6913), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6914) );
  INV_X1 U8675 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6916) );
  MUX2_X1 U8676 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6916), .S(n6917), .Z(n6957)
         );
  INV_X1 U8677 ( .A(n6917), .ZN(n6961) );
  NAND2_X1 U8678 ( .A1(n6961), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U8679 ( .A1(n6955), .A2(n6918), .ZN(n6966) );
  OR2_X1 U8680 ( .A1(n6919), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8681 ( .A1(n6919), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U8682 ( .A1(n6923), .A2(n6920), .ZN(n6967) );
  NAND2_X1 U8683 ( .A1(n6964), .A2(n6923), .ZN(n6921) );
  INV_X1 U8684 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7129) );
  MUX2_X1 U8685 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n7129), .S(n7136), .Z(n6922)
         );
  NAND2_X1 U8686 ( .A1(n6921), .A2(n6922), .ZN(n7132) );
  INV_X1 U8687 ( .A(n6922), .ZN(n6924) );
  NAND3_X1 U8688 ( .A1(n6964), .A2(n6924), .A3(n6923), .ZN(n6925) );
  AOI21_X1 U8689 ( .B1(n7132), .B2(n6925), .A(n8372), .ZN(n6926) );
  AOI211_X1 U8690 ( .C1(n8342), .C2(n7136), .A(n6927), .B(n6926), .ZN(n6928)
         );
  OAI21_X1 U8691 ( .B1(n8383), .B2(n6929), .A(n6928), .ZN(P2_U3259) );
  INV_X1 U8692 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U8693 ( .A1(n6930), .A2(n10084), .ZN(n6931) );
  OAI21_X1 U8694 ( .B1(n10084), .B2(n10144), .A(n6931), .ZN(P2_U3521) );
  INV_X1 U8695 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U8696 ( .A1(n6932), .A2(n6933), .ZN(n7484) );
  OR2_X1 U8697 ( .A1(n6932), .A2(n6933), .ZN(n6934) );
  NAND2_X1 U8698 ( .A1(n7484), .A2(n6934), .ZN(n8638) );
  INV_X1 U8699 ( .A(n8638), .ZN(n6944) );
  OAI21_X1 U8700 ( .B1(n6936), .B2(n6935), .A(n7471), .ZN(n6938) );
  OAI22_X1 U8701 ( .A1(n7176), .A2(n8605), .B1(n4467), .B2(n8603), .ZN(n6937)
         );
  AOI21_X1 U8702 ( .B1(n6938), .B2(n8614), .A(n6937), .ZN(n6940) );
  INV_X1 U8703 ( .A(n8610), .ZN(n7763) );
  NAND2_X1 U8704 ( .A1(n8638), .A2(n7763), .ZN(n6939) );
  NAND2_X1 U8705 ( .A1(n6940), .A2(n6939), .ZN(n8644) );
  INV_X1 U8706 ( .A(n8644), .ZN(n6943) );
  AND2_X1 U8707 ( .A1(n7528), .A2(n8636), .ZN(n6941) );
  NOR2_X1 U8708 ( .A1(n7477), .A2(n6941), .ZN(n8642) );
  AOI22_X1 U8709 ( .A1(n8642), .A2(n8763), .B1(n8762), .B2(n8636), .ZN(n6942)
         );
  OAI211_X1 U8710 ( .C1(n6944), .C2(n8759), .A(n6943), .B(n6942), .ZN(n6947)
         );
  NAND2_X1 U8711 ( .A1(n6947), .A2(n10084), .ZN(n6945) );
  OAI21_X1 U8712 ( .B1(n10084), .B2(n6946), .A(n6945), .ZN(P2_U3523) );
  INV_X1 U8713 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8714 ( .A1(n6947), .A2(n10076), .ZN(n6948) );
  OAI21_X1 U8715 ( .B1(n10076), .B2(n6949), .A(n6948), .ZN(P2_U3460) );
  INV_X1 U8716 ( .A(n6950), .ZN(n6951) );
  AOI21_X1 U8717 ( .B1(n6953), .B2(n6952), .A(n6951), .ZN(n6963) );
  INV_X1 U8718 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8719 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7917) );
  OAI21_X1 U8720 ( .B1(n8395), .B2(n6954), .A(n7917), .ZN(n6960) );
  INV_X1 U8721 ( .A(n6955), .ZN(n6956) );
  AOI211_X1 U8722 ( .C1(n6958), .C2(n6957), .A(n8372), .B(n6956), .ZN(n6959)
         );
  AOI211_X1 U8723 ( .C1(n8342), .C2(n6961), .A(n6960), .B(n6959), .ZN(n6962)
         );
  OAI21_X1 U8724 ( .B1(n6963), .B2(n8383), .A(n6962), .ZN(P2_U3257) );
  INV_X1 U8725 ( .A(n6964), .ZN(n6965) );
  AOI21_X1 U8726 ( .B1(n6967), .B2(n6966), .A(n6965), .ZN(n6976) );
  NOR2_X1 U8727 ( .A1(n6968), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8174) );
  NOR2_X1 U8728 ( .A1(n8382), .A2(n6969), .ZN(n6970) );
  AOI211_X1 U8729 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n8366), .A(n8174), .B(
        n6970), .ZN(n6975) );
  XNOR2_X1 U8730 ( .A(n6972), .B(n6971), .ZN(n6973) );
  NAND2_X1 U8731 ( .A1(n6973), .A2(n8386), .ZN(n6974) );
  OAI211_X1 U8732 ( .C1(n6976), .C2(n8372), .A(n6975), .B(n6974), .ZN(P2_U3258) );
  NOR2_X1 U8733 ( .A1(n6978), .A2(n6977), .ZN(n6979) );
  NAND2_X1 U8734 ( .A1(n6980), .A2(n6979), .ZN(n6987) );
  NAND2_X2 U8735 ( .A1(n6987), .A2(n9667), .ZN(n9670) );
  INV_X1 U8736 ( .A(n6982), .ZN(n6995) );
  AND2_X1 U8737 ( .A1(n6984), .A2(n6983), .ZN(n6985) );
  NAND2_X1 U8738 ( .A1(n9670), .A2(n6985), .ZN(n9714) );
  INV_X1 U8739 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6986) );
  OAI22_X1 U8740 ( .A1(n9670), .A2(n6986), .B1(n4669), .B2(n9667), .ZN(n6992)
         );
  OR2_X1 U8741 ( .A1(n6987), .A2(n9164), .ZN(n9675) );
  AND2_X1 U8742 ( .A1(n9323), .A2(n9284), .ZN(n6988) );
  NAND2_X1 U8743 ( .A1(n9670), .A2(n6988), .ZN(n9697) );
  OAI22_X1 U8744 ( .A1(n9675), .A2(n6990), .B1(n6989), .B2(n9697), .ZN(n6991)
         );
  AOI211_X1 U8745 ( .C1(n9672), .C2(n6993), .A(n6992), .B(n6991), .ZN(n6994)
         );
  OAI21_X1 U8746 ( .B1(n9694), .B2(n6995), .A(n6994), .ZN(P1_U3289) );
  AND2_X1 U8747 ( .A1(n9331), .A2(n8927), .ZN(n6996) );
  NAND2_X1 U8748 ( .A1(n9670), .A2(n6996), .ZN(n9716) );
  NAND2_X1 U8749 ( .A1(n6997), .A2(n9287), .ZN(n7002) );
  NOR2_X1 U8750 ( .A1(n7004), .A2(n6998), .ZN(n6999) );
  XNOR2_X1 U8751 ( .A(n7002), .B(n6999), .ZN(n9960) );
  INV_X1 U8752 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7000) );
  NOR2_X1 U8753 ( .A1(n9670), .A2(n7000), .ZN(n7011) );
  INV_X1 U8754 ( .A(n9287), .ZN(n7001) );
  NOR2_X1 U8755 ( .A1(n9288), .A2(n7001), .ZN(n9252) );
  AOI211_X1 U8756 ( .C1(n7003), .C2(n7002), .A(n9557), .B(n9252), .ZN(n7006)
         );
  OAI22_X1 U8757 ( .A1(n9656), .A2(n6335), .B1(n7004), .B2(n9654), .ZN(n7005)
         );
  NOR2_X1 U8758 ( .A1(n7006), .A2(n7005), .ZN(n9959) );
  NOR3_X1 U8759 ( .A1(n10000), .A2(n7008), .A3(n7007), .ZN(n9955) );
  AOI22_X1 U8760 ( .A1(n9955), .A2(n9440), .B1(n9710), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7009) );
  INV_X1 U8761 ( .A(n9670), .ZN(n9694) );
  AOI21_X1 U8762 ( .B1(n9959), .B2(n7009), .A(n9694), .ZN(n7010) );
  AOI211_X1 U8763 ( .C1(n9672), .C2(n9956), .A(n7011), .B(n7010), .ZN(n7012)
         );
  OAI21_X1 U8764 ( .B1(n9716), .B2(n9960), .A(n7012), .ZN(P1_U3290) );
  AND2_X1 U8765 ( .A1(n7014), .A2(n7013), .ZN(n7015) );
  INV_X1 U8766 ( .A(n10031), .ZN(n7016) );
  NAND2_X1 U8767 ( .A1(n7026), .A2(n7017), .ZN(n8221) );
  INV_X1 U8768 ( .A(n8221), .ZN(n8235) );
  OR2_X1 U8769 ( .A1(n7018), .A2(n7119), .ZN(n7375) );
  INV_X1 U8770 ( .A(n7375), .ZN(n7019) );
  AND2_X1 U8771 ( .A1(n10031), .A2(n7019), .ZN(n7020) );
  NAND2_X1 U8772 ( .A1(n7021), .A2(n7020), .ZN(n7022) );
  AOI22_X1 U8773 ( .A1(n8235), .A2(n7023), .B1(n7580), .B2(n8236), .ZN(n7047)
         );
  AND2_X1 U8774 ( .A1(n10070), .A2(n7024), .ZN(n7025) );
  NOR2_X1 U8775 ( .A1(n7534), .A2(n8012), .ZN(n7030) );
  XNOR2_X1 U8776 ( .A(n7124), .B(n7580), .ZN(n7029) );
  NAND2_X1 U8777 ( .A1(n7030), .A2(n7029), .ZN(n7033) );
  INV_X1 U8778 ( .A(n7029), .ZN(n7032) );
  INV_X1 U8779 ( .A(n7030), .ZN(n7031) );
  NAND2_X1 U8780 ( .A1(n7032), .A2(n7031), .ZN(n7122) );
  NAND2_X1 U8781 ( .A1(n4483), .A2(n7991), .ZN(n7097) );
  OAI21_X1 U8782 ( .B1(n7036), .B2(n7035), .A(n7123), .ZN(n7045) );
  INV_X1 U8783 ( .A(n7037), .ZN(n7038) );
  NAND2_X1 U8784 ( .A1(n7039), .A2(n7038), .ZN(n7044) );
  AND3_X1 U8785 ( .A1(n7042), .A2(n7041), .A3(n7040), .ZN(n7043) );
  NAND2_X1 U8786 ( .A1(n7044), .A2(n7043), .ZN(n7155) );
  OR2_X1 U8787 ( .A1(n7155), .A2(P2_U3152), .ZN(n7125) );
  AOI22_X1 U8788 ( .A1(n8184), .A2(n7045), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n7125), .ZN(n7046) );
  NAND2_X1 U8789 ( .A1(n7047), .A2(n7046), .ZN(P2_U3224) );
  XNOR2_X1 U8790 ( .A(n7048), .B(n9251), .ZN(n9965) );
  NAND2_X1 U8791 ( .A1(n9670), .A2(n4373), .ZN(n9645) );
  OAI21_X1 U8792 ( .B1(n7050), .B2(n4860), .A(n7069), .ZN(n9966) );
  INV_X1 U8793 ( .A(n9670), .ZN(n9712) );
  AOI22_X1 U8794 ( .A1(n9712), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9710), .B2(
        n6015), .ZN(n7051) );
  OAI21_X1 U8795 ( .B1(n9645), .B2(n9966), .A(n7051), .ZN(n7052) );
  AOI21_X1 U8796 ( .B1(n9672), .B2(n7053), .A(n7052), .ZN(n7060) );
  OAI21_X1 U8797 ( .B1(n9251), .B2(n7054), .A(n7055), .ZN(n7057) );
  OAI22_X1 U8798 ( .A1(n9656), .A2(n7284), .B1(n6335), .B2(n9654), .ZN(n7056)
         );
  AOI21_X1 U8799 ( .B1(n7057), .B2(n9708), .A(n7056), .ZN(n7058) );
  OAI21_X1 U8800 ( .B1(n9965), .B2(n9689), .A(n7058), .ZN(n9967) );
  NAND2_X1 U8801 ( .A1(n9967), .A2(n9670), .ZN(n7059) );
  OAI211_X1 U8802 ( .C1(n9965), .C2(n9697), .A(n7060), .B(n7059), .ZN(P1_U3288) );
  XNOR2_X1 U8803 ( .A(n7061), .B(n4897), .ZN(n9971) );
  XNOR2_X1 U8804 ( .A(n7063), .B(n4897), .ZN(n7065) );
  OAI22_X1 U8805 ( .A1(n9656), .A2(n6800), .B1(n6339), .B2(n9654), .ZN(n7064)
         );
  AOI21_X1 U8806 ( .B1(n7065), .B2(n9708), .A(n7064), .ZN(n7066) );
  OAI21_X1 U8807 ( .B1(n9971), .B2(n9689), .A(n7066), .ZN(n9974) );
  NAND2_X1 U8808 ( .A1(n9974), .A2(n9670), .ZN(n7075) );
  INV_X1 U8809 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7068) );
  OAI22_X1 U8810 ( .A1(n9670), .A2(n7068), .B1(n7067), .B2(n9667), .ZN(n7072)
         );
  AND2_X1 U8811 ( .A1(n7069), .A2(n7073), .ZN(n7070) );
  OR2_X1 U8812 ( .A1(n7070), .A2(n7286), .ZN(n9973) );
  NOR2_X1 U8813 ( .A1(n9645), .A2(n9973), .ZN(n7071) );
  AOI211_X1 U8814 ( .C1(n9672), .C2(n7073), .A(n7072), .B(n7071), .ZN(n7074)
         );
  OAI211_X1 U8815 ( .C1(n9971), .C2(n9697), .A(n7075), .B(n7074), .ZN(P1_U3287) );
  INV_X1 U8816 ( .A(n7076), .ZN(n7077) );
  INV_X1 U8817 ( .A(n7287), .ZN(n9253) );
  NAND2_X1 U8818 ( .A1(n7077), .A2(n9253), .ZN(n9979) );
  NAND2_X1 U8819 ( .A1(n9979), .A2(n7078), .ZN(n7079) );
  XNOR2_X1 U8820 ( .A(n9073), .B(n7079), .ZN(n9986) );
  XNOR2_X1 U8821 ( .A(n9073), .B(n7080), .ZN(n7082) );
  OAI22_X1 U8822 ( .A1(n9656), .A2(n7423), .B1(n6800), .B2(n9654), .ZN(n7081)
         );
  AOI21_X1 U8823 ( .B1(n7082), .B2(n9708), .A(n7081), .ZN(n7083) );
  OAI21_X1 U8824 ( .B1(n9689), .B2(n9986), .A(n7083), .ZN(n9988) );
  NAND2_X1 U8825 ( .A1(n9988), .A2(n9670), .ZN(n7091) );
  INV_X1 U8826 ( .A(n7084), .ZN(n7349) );
  OAI22_X1 U8827 ( .A1(n9670), .A2(n7085), .B1(n7349), .B2(n9667), .ZN(n7088)
         );
  NAND2_X1 U8828 ( .A1(n7285), .A2(n7089), .ZN(n7086) );
  NAND2_X1 U8829 ( .A1(n7316), .A2(n7086), .ZN(n9987) );
  NOR2_X1 U8830 ( .A1(n9987), .A2(n9645), .ZN(n7087) );
  AOI211_X1 U8831 ( .C1(n9672), .C2(n7089), .A(n7088), .B(n7087), .ZN(n7090)
         );
  OAI211_X1 U8832 ( .C1(n9986), .C2(n9697), .A(n7091), .B(n7090), .ZN(P1_U3285) );
  INV_X1 U8833 ( .A(n9645), .ZN(n9700) );
  OAI21_X1 U8834 ( .B1(n9700), .B2(n9672), .A(n7092), .ZN(n7095) );
  AOI22_X1 U8835 ( .A1(n7093), .A2(n9670), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9710), .ZN(n7094) );
  OAI211_X1 U8836 ( .C1(n9670), .C2(n7096), .A(n7095), .B(n7094), .ZN(P1_U3291) );
  AOI21_X1 U8837 ( .B1(n8184), .B2(n7097), .A(n8236), .ZN(n7103) );
  AOI22_X1 U8838 ( .A1(n8235), .A2(n7098), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n7125), .ZN(n7101) );
  INV_X1 U8839 ( .A(n8209), .ZN(n8185) );
  NAND2_X1 U8840 ( .A1(n8185), .A2(n7099), .ZN(n7100) );
  OAI211_X1 U8841 ( .C1(n7103), .C2(n7102), .A(n7101), .B(n7100), .ZN(P2_U3234) );
  INV_X1 U8842 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7114) );
  INV_X1 U8843 ( .A(n7104), .ZN(n7105) );
  XNOR2_X1 U8844 ( .A(n7107), .B(n7106), .ZN(n7383) );
  XNOR2_X1 U8845 ( .A(n7108), .B(n4274), .ZN(n7109) );
  AOI222_X1 U8846 ( .A1(n8614), .A2(n7109), .B1(n8260), .B2(n8580), .C1(n8258), 
        .C2(n8582), .ZN(n7371) );
  INV_X1 U8847 ( .A(n7442), .ZN(n7111) );
  AOI211_X1 U8848 ( .C1(n5900), .C2(n7110), .A(n10052), .B(n7111), .ZN(n7380)
         );
  AOI21_X1 U8849 ( .B1(n8762), .B2(n5900), .A(n7380), .ZN(n7112) );
  OAI211_X1 U8850 ( .C1(n8767), .C2(n7383), .A(n7371), .B(n7112), .ZN(n7115)
         );
  NAND2_X1 U8851 ( .A1(n7115), .A2(n10076), .ZN(n7113) );
  OAI21_X1 U8852 ( .B1(n10076), .B2(n7114), .A(n7113), .ZN(P2_U3466) );
  NAND2_X1 U8853 ( .A1(n7115), .A2(n10084), .ZN(n7116) );
  OAI21_X1 U8854 ( .B1(n10084), .B2(n6826), .A(n7116), .ZN(P2_U3525) );
  INV_X1 U8855 ( .A(n7117), .ZN(n7120) );
  OAI222_X1 U8856 ( .A1(n9866), .A2(n7120), .B1(P1_U3084), .B2(n9276), .C1(
        n7118), .C2(n7758), .ZN(P1_U3333) );
  OAI222_X1 U8857 ( .A1(n8802), .A2(n7121), .B1(n4275), .B2(n7120), .C1(n7119), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OR2_X1 U8858 ( .A1(n4467), .A2(n8012), .ZN(n7148) );
  XNOR2_X1 U8859 ( .A(n7154), .B(n7153), .ZN(n7128) );
  INV_X1 U8860 ( .A(n8204), .ZN(n8186) );
  INV_X1 U8861 ( .A(n8205), .ZN(n8187) );
  AOI22_X1 U8862 ( .A1(n8186), .A2(n8261), .B1(n8187), .B2(n5891), .ZN(n7127)
         );
  AOI22_X1 U8863 ( .A1(n7125), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8236), .B2(
        n8761), .ZN(n7126) );
  OAI211_X1 U8864 ( .C1(n7128), .C2(n8230), .A(n7127), .B(n7126), .ZN(P2_U3239) );
  NAND2_X1 U8865 ( .A1(n7130), .A2(n7129), .ZN(n7131) );
  NAND2_X1 U8866 ( .A1(n7132), .A2(n7131), .ZN(n7133) );
  NAND2_X1 U8867 ( .A1(n7133), .A2(n7142), .ZN(n7206) );
  OAI21_X1 U8868 ( .B1(n7133), .B2(n7142), .A(n7206), .ZN(n7135) );
  OR2_X1 U8869 ( .A1(n7135), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7207) );
  INV_X1 U8870 ( .A(n7207), .ZN(n7134) );
  AOI21_X1 U8871 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7135), .A(n7134), .ZN(
        n7147) );
  NOR2_X1 U8872 ( .A1(n7136), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7137) );
  AOI21_X1 U8873 ( .B1(n7139), .B2(n7138), .A(n7137), .ZN(n7210) );
  XOR2_X1 U8874 ( .A(n7209), .B(n7210), .Z(n7141) );
  INV_X1 U8875 ( .A(n7208), .ZN(n7140) );
  OAI211_X1 U8876 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n7141), .A(n7140), .B(
        n8386), .ZN(n7146) );
  AND2_X1 U8877 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7144) );
  NOR2_X1 U8878 ( .A1(n8382), .A2(n7142), .ZN(n7143) );
  AOI211_X1 U8879 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n8366), .A(n7144), .B(
        n7143), .ZN(n7145) );
  OAI211_X1 U8880 ( .C1(n7147), .C2(n8372), .A(n7146), .B(n7145), .ZN(P2_U3260) );
  INV_X1 U8881 ( .A(n7148), .ZN(n7151) );
  INV_X1 U8882 ( .A(n7149), .ZN(n7150) );
  NAND2_X1 U8883 ( .A1(n7151), .A2(n7150), .ZN(n7152) );
  XNOR2_X1 U8884 ( .A(n7124), .B(n8636), .ZN(n7162) );
  OR2_X1 U8885 ( .A1(n7535), .A2(n8012), .ZN(n7163) );
  XNOR2_X1 U8886 ( .A(n7162), .B(n7163), .ZN(n7166) );
  XNOR2_X1 U8887 ( .A(n7167), .B(n7166), .ZN(n7161) );
  OAI22_X1 U8888 ( .A1(n8226), .A2(n7156), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8640), .ZN(n7159) );
  OAI22_X1 U8889 ( .A1(n7176), .A2(n8204), .B1(n8205), .B2(n4467), .ZN(n7158)
         );
  AOI211_X1 U8890 ( .C1(n8238), .C2(n8640), .A(n7159), .B(n7158), .ZN(n7160)
         );
  OAI21_X1 U8891 ( .B1(n8230), .B2(n7161), .A(n7160), .ZN(P2_U3220) );
  INV_X1 U8892 ( .A(n7162), .ZN(n7164) );
  NOR2_X1 U8893 ( .A1(n7164), .A2(n7163), .ZN(n7165) );
  NOR2_X1 U8894 ( .A1(n7176), .A2(n8012), .ZN(n7169) );
  XNOR2_X1 U8895 ( .A(n7124), .B(n5279), .ZN(n7168) );
  NAND2_X1 U8896 ( .A1(n7169), .A2(n7168), .ZN(n7172) );
  INV_X1 U8897 ( .A(n7168), .ZN(n7171) );
  INV_X1 U8898 ( .A(n7169), .ZN(n7170) );
  NAND2_X1 U8899 ( .A1(n7171), .A2(n7170), .ZN(n7173) );
  AND2_X1 U8900 ( .A1(n7172), .A2(n7173), .ZN(n7182) );
  XNOR2_X1 U8901 ( .A(n7124), .B(n7378), .ZN(n7196) );
  OR2_X1 U8902 ( .A1(n7474), .A2(n8012), .ZN(n7195) );
  XNOR2_X1 U8903 ( .A(n7196), .B(n7195), .ZN(n7194) );
  XOR2_X1 U8904 ( .A(n7193), .B(n7194), .Z(n7179) );
  NAND2_X1 U8905 ( .A1(n8238), .A2(n7376), .ZN(n7174) );
  OAI211_X1 U8906 ( .C1(n8226), .C2(n7378), .A(n7175), .B(n7174), .ZN(n7178)
         );
  OAI22_X1 U8907 ( .A1(n7308), .A2(n8204), .B1(n8205), .B2(n7176), .ZN(n7177)
         );
  AOI211_X1 U8908 ( .C1(n7179), .C2(n8184), .A(n7178), .B(n7177), .ZN(n7180)
         );
  INV_X1 U8909 ( .A(n7180), .ZN(P2_U3229) );
  OAI21_X1 U8910 ( .B1(n7183), .B2(n7182), .A(n7181), .ZN(n7188) );
  NAND2_X1 U8911 ( .A1(n8238), .A2(n7479), .ZN(n7184) );
  OAI211_X1 U8912 ( .C1(n8226), .C2(n10043), .A(n7185), .B(n7184), .ZN(n7187)
         );
  OAI22_X1 U8913 ( .A1(n7535), .A2(n8205), .B1(n8204), .B2(n7474), .ZN(n7186)
         );
  AOI211_X1 U8914 ( .C1(n8184), .C2(n7188), .A(n7187), .B(n7186), .ZN(n7189)
         );
  INV_X1 U8915 ( .A(n7189), .ZN(P2_U3232) );
  AND2_X1 U8916 ( .A1(n8258), .A2(n7991), .ZN(n7190) );
  XNOR2_X1 U8917 ( .A(n7124), .B(n7448), .ZN(n7191) );
  NAND2_X1 U8918 ( .A1(n7191), .A2(n7190), .ZN(n7192) );
  AND2_X1 U8919 ( .A1(n7304), .A2(n7192), .ZN(n7200) );
  INV_X1 U8920 ( .A(n7195), .ZN(n7198) );
  INV_X1 U8921 ( .A(n7196), .ZN(n7197) );
  NAND2_X1 U8922 ( .A1(n7199), .A2(n7200), .ZN(n7305) );
  OAI21_X1 U8923 ( .B1(n7200), .B2(n7199), .A(n7305), .ZN(n7204) );
  NAND2_X1 U8924 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8300) );
  NAND2_X1 U8925 ( .A1(n8238), .A2(n7445), .ZN(n7201) );
  OAI211_X1 U8926 ( .C1(n8226), .C2(n10051), .A(n8300), .B(n7201), .ZN(n7203)
         );
  OAI22_X1 U8927 ( .A1(n7474), .A2(n8205), .B1(n8204), .B2(n7653), .ZN(n7202)
         );
  AOI211_X1 U8928 ( .C1(n7204), .C2(n8184), .A(n7203), .B(n7202), .ZN(n7205)
         );
  INV_X1 U8929 ( .A(n7205), .ZN(P2_U3241) );
  NAND2_X1 U8930 ( .A1(n7207), .A2(n7206), .ZN(n7615) );
  XNOR2_X1 U8931 ( .A(n7624), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n7614) );
  XNOR2_X1 U8932 ( .A(n7615), .B(n7614), .ZN(n7218) );
  XOR2_X1 U8933 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n7624), .Z(n7212) );
  AOI21_X1 U8934 ( .B1(n7210), .B2(n7209), .A(n7208), .ZN(n7211) );
  NAND2_X1 U8935 ( .A1(n7211), .A2(n7212), .ZN(n7623) );
  OAI21_X1 U8936 ( .B1(n7212), .B2(n7211), .A(n7623), .ZN(n7213) );
  NAND2_X1 U8937 ( .A1(n7213), .A2(n8386), .ZN(n7217) );
  INV_X1 U8938 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U8939 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8130) );
  OAI21_X1 U8940 ( .B1(n8395), .B2(n7214), .A(n8130), .ZN(n7215) );
  AOI21_X1 U8941 ( .B1(n8342), .B2(n7624), .A(n7215), .ZN(n7216) );
  OAI211_X1 U8942 ( .C1(n8372), .C2(n7218), .A(n7217), .B(n7216), .ZN(P2_U3261) );
  INV_X1 U8943 ( .A(n7219), .ZN(n7269) );
  OAI222_X1 U8944 ( .A1(n9866), .A2(n7269), .B1(P1_U3084), .B2(n9165), .C1(
        n7220), .C2(n7758), .ZN(P1_U3332) );
  NAND2_X1 U8945 ( .A1(n7324), .A2(n9070), .ZN(n7221) );
  XOR2_X1 U8946 ( .A(n9256), .B(n7221), .Z(n7227) );
  INV_X1 U8947 ( .A(n7242), .ZN(n7223) );
  AOI21_X1 U8948 ( .B1(n9256), .B2(n7222), .A(n7223), .ZN(n10004) );
  INV_X1 U8949 ( .A(n9689), .ZN(n7225) );
  OAI22_X1 U8950 ( .A1(n9656), .A2(n7712), .B1(n7423), .B2(n9654), .ZN(n7224)
         );
  AOI21_X1 U8951 ( .B1(n10004), .B2(n7225), .A(n7224), .ZN(n7226) );
  OAI21_X1 U8952 ( .B1(n7227), .B2(n9557), .A(n7226), .ZN(n10002) );
  INV_X1 U8953 ( .A(n10002), .ZN(n7235) );
  INV_X1 U8954 ( .A(n9697), .ZN(n7233) );
  NOR2_X1 U8955 ( .A1(n7318), .A2(n9999), .ZN(n7228) );
  OR2_X1 U8956 ( .A1(n7244), .A2(n7228), .ZN(n10001) );
  AOI22_X1 U8957 ( .A1(n9712), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7229), .B2(
        n9710), .ZN(n7231) );
  NAND2_X1 U8958 ( .A1(n9672), .A2(n7414), .ZN(n7230) );
  OAI211_X1 U8959 ( .C1(n10001), .C2(n9645), .A(n7231), .B(n7230), .ZN(n7232)
         );
  AOI21_X1 U8960 ( .B1(n10004), .B2(n7233), .A(n7232), .ZN(n7234) );
  OAI21_X1 U8961 ( .B1(n7235), .B2(n9694), .A(n7234), .ZN(P1_U3283) );
  NAND2_X1 U8962 ( .A1(n7236), .A2(n9076), .ZN(n7237) );
  NAND2_X1 U8963 ( .A1(n9080), .A2(n9078), .ZN(n9259) );
  XNOR2_X1 U8964 ( .A(n7237), .B(n9259), .ZN(n7240) );
  NAND2_X1 U8965 ( .A1(n9703), .A2(n9348), .ZN(n7238) );
  OAI21_X1 U8966 ( .B1(n7570), .B2(n9654), .A(n7238), .ZN(n7239) );
  AOI21_X1 U8967 ( .B1(n7240), .B2(n9708), .A(n7239), .ZN(n10014) );
  NAND2_X1 U8968 ( .A1(n7242), .A2(n7241), .ZN(n7332) );
  INV_X1 U8969 ( .A(n9259), .ZN(n7243) );
  XNOR2_X1 U8970 ( .A(n7332), .B(n7243), .ZN(n10011) );
  OR2_X1 U8971 ( .A1(n7244), .A2(n7248), .ZN(n7245) );
  AND2_X1 U8972 ( .A1(n7336), .A2(n7245), .ZN(n10009) );
  NAND2_X1 U8973 ( .A1(n10009), .A2(n9700), .ZN(n7247) );
  AOI22_X1 U8974 ( .A1(n9712), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7641), .B2(
        n9710), .ZN(n7246) );
  OAI211_X1 U8975 ( .C1(n7248), .C2(n9714), .A(n7247), .B(n7246), .ZN(n7249)
         );
  AOI21_X1 U8976 ( .B1(n10011), .B2(n9677), .A(n7249), .ZN(n7250) );
  OAI21_X1 U8977 ( .B1(n10014), .B2(n9694), .A(n7250), .ZN(P1_U3282) );
  NAND2_X1 U8978 ( .A1(n8924), .A2(n9353), .ZN(n7252) );
  NAND2_X1 U8979 ( .A1(n8883), .A2(n7292), .ZN(n7251) );
  AND2_X1 U8980 ( .A1(n7252), .A2(n7251), .ZN(n7402) );
  NAND2_X1 U8981 ( .A1(n7254), .A2(n7253), .ZN(n7255) );
  OAI21_X1 U8982 ( .B1(n6800), .B2(n8892), .A(n7257), .ZN(n7258) );
  XNOR2_X1 U8983 ( .A(n7258), .B(n8927), .ZN(n7259) );
  AND2_X1 U8984 ( .A1(n7407), .A2(n7403), .ZN(n7261) );
  NAND2_X1 U8985 ( .A1(n7261), .A2(n7402), .ZN(n7345) );
  OAI21_X1 U8986 ( .B1(n7402), .B2(n7261), .A(n7345), .ZN(n7266) );
  INV_X1 U8987 ( .A(n9047), .ZN(n9035) );
  AOI22_X1 U8988 ( .A1(n9050), .A2(n9354), .B1(n9035), .B2(n7288), .ZN(n7264)
         );
  AOI21_X1 U8989 ( .B1(n9019), .B2(n9352), .A(n7262), .ZN(n7263) );
  OAI211_X1 U8990 ( .C1(n9982), .C2(n9053), .A(n7264), .B(n7263), .ZN(n7265)
         );
  AOI21_X1 U8991 ( .B1(n7266), .B2(n9043), .A(n7265), .ZN(n7267) );
  INV_X1 U8992 ( .A(n7267), .ZN(P1_U3225) );
  OAI222_X1 U8993 ( .A1(n8802), .A2(n7270), .B1(n4275), .B2(n7269), .C1(n7268), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  XNOR2_X1 U8994 ( .A(n7387), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7384) );
  AOI21_X1 U8995 ( .B1(n9908), .B2(n7272), .A(n7271), .ZN(n7385) );
  XOR2_X1 U8996 ( .A(n7385), .B(n7384), .Z(n7281) );
  NAND2_X1 U8997 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7679) );
  OAI21_X1 U8998 ( .B1(n9918), .B2(n7273), .A(n7679), .ZN(n7279) );
  XNOR2_X1 U8999 ( .A(n7387), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7277) );
  AOI211_X1 U9000 ( .C1(n7277), .C2(n7276), .A(n9438), .B(n7386), .ZN(n7278)
         );
  AOI211_X1 U9001 ( .C1(n9927), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7279), .B(
        n7278), .ZN(n7280) );
  OAI21_X1 U9002 ( .B1(n9923), .B2(n7281), .A(n7280), .ZN(P1_U3253) );
  XNOR2_X1 U9003 ( .A(n7287), .B(n7282), .ZN(n7283) );
  OAI222_X1 U9004 ( .A1(n9656), .A2(n7568), .B1(n9654), .B2(n7284), .C1(n9557), 
        .C2(n7283), .ZN(n9984) );
  OAI211_X1 U9005 ( .C1(n7286), .C2(n9982), .A(n10008), .B(n7285), .ZN(n9980)
         );
  NAND2_X1 U9006 ( .A1(n7076), .A2(n7287), .ZN(n9978) );
  NAND3_X1 U9007 ( .A1(n9979), .A2(n9677), .A3(n9978), .ZN(n7294) );
  INV_X1 U9008 ( .A(n7288), .ZN(n7289) );
  OAI22_X1 U9009 ( .A1(n9670), .A2(n7290), .B1(n7289), .B2(n9667), .ZN(n7291)
         );
  AOI21_X1 U9010 ( .B1(n9672), .B2(n7292), .A(n7291), .ZN(n7293) );
  OAI211_X1 U9011 ( .C1(n9675), .C2(n9980), .A(n7294), .B(n7293), .ZN(n7295)
         );
  AOI21_X1 U9012 ( .B1(n9984), .B2(n9670), .A(n7295), .ZN(n7296) );
  INV_X1 U9013 ( .A(n7296), .ZN(P1_U3286) );
  NAND2_X1 U9014 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n8257), .ZN(n7297) );
  OAI21_X1 U9015 ( .B1(n8218), .B2(n8257), .A(n7297), .ZN(P2_U3577) );
  INV_X1 U9016 ( .A(n7298), .ZN(n7302) );
  OAI222_X1 U9017 ( .A1(n8802), .A2(n7300), .B1(n4275), .B2(n7302), .C1(
        P2_U3152), .C2(n7299), .ZN(P2_U3336) );
  OAI222_X1 U9018 ( .A1(n7758), .A2(n7303), .B1(n9866), .B2(n7302), .C1(n7301), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  NOR2_X1 U9019 ( .A1(n7653), .A2(n8012), .ZN(n7454) );
  XNOR2_X1 U9020 ( .A(n7124), .B(n7558), .ZN(n7453) );
  XNOR2_X1 U9021 ( .A(n7454), .B(n7453), .ZN(n7451) );
  XOR2_X1 U9022 ( .A(n7451), .B(n7452), .Z(n7311) );
  NAND2_X1 U9023 ( .A1(n8238), .A2(n7555), .ZN(n7306) );
  OAI211_X1 U9024 ( .C1(n8226), .C2(n10061), .A(n7307), .B(n7306), .ZN(n7310)
         );
  OAI22_X1 U9025 ( .A1(n7308), .A2(n8205), .B1(n8204), .B2(n7694), .ZN(n7309)
         );
  AOI211_X1 U9026 ( .C1(n7311), .C2(n8184), .A(n7310), .B(n7309), .ZN(n7312)
         );
  INV_X1 U9027 ( .A(n7312), .ZN(P2_U3215) );
  AOI21_X1 U9028 ( .B1(n7076), .B2(n7314), .A(n7313), .ZN(n7315) );
  XNOR2_X1 U9029 ( .A(n7315), .B(n9255), .ZN(n9996) );
  NAND2_X1 U9030 ( .A1(n7316), .A2(n7561), .ZN(n7317) );
  NAND2_X1 U9031 ( .A1(n7317), .A2(n10008), .ZN(n7319) );
  OR2_X1 U9032 ( .A1(n7319), .A2(n7318), .ZN(n9992) );
  INV_X1 U9033 ( .A(n7320), .ZN(n7567) );
  OAI22_X1 U9034 ( .A1(n9670), .A2(n7321), .B1(n7567), .B2(n9667), .ZN(n7322)
         );
  AOI21_X1 U9035 ( .B1(n9672), .B2(n7561), .A(n7322), .ZN(n7323) );
  OAI21_X1 U9036 ( .B1(n9992), .B2(n9675), .A(n7323), .ZN(n7327) );
  OAI21_X1 U9037 ( .B1(n9255), .B2(n9072), .A(n7324), .ZN(n7325) );
  AOI222_X1 U9038 ( .A1(n9708), .A2(n7325), .B1(n9350), .B2(n9703), .C1(n9352), 
        .C2(n9705), .ZN(n9993) );
  NOR2_X1 U9039 ( .A1(n9993), .A2(n9694), .ZN(n7326) );
  AOI211_X1 U9040 ( .C1(n9677), .C2(n9996), .A(n7327), .B(n7326), .ZN(n7328)
         );
  INV_X1 U9041 ( .A(n7328), .ZN(P1_U3284) );
  INV_X1 U9042 ( .A(n7329), .ZN(n9085) );
  AOI21_X1 U9043 ( .B1(n7236), .B2(n9085), .A(n4690), .ZN(n7330) );
  INV_X1 U9044 ( .A(n7334), .ZN(n9263) );
  XNOR2_X1 U9045 ( .A(n7330), .B(n9263), .ZN(n7331) );
  OAI222_X1 U9046 ( .A1(n9656), .A2(n7681), .B1(n9654), .B2(n7712), .C1(n7331), 
        .C2(n9557), .ZN(n7585) );
  INV_X1 U9047 ( .A(n7585), .ZN(n7342) );
  AOI22_X1 U9048 ( .A1(n7332), .A2(n4374), .B1(n9349), .B2(n7640), .ZN(n7335)
         );
  OAI21_X1 U9049 ( .B1(n7335), .B2(n7334), .A(n7333), .ZN(n7587) );
  INV_X1 U9050 ( .A(n7336), .ZN(n7337) );
  INV_X1 U9051 ( .A(n6327), .ZN(n7717) );
  OAI211_X1 U9052 ( .C1(n7337), .C2(n7717), .A(n10008), .B(n7360), .ZN(n7584)
         );
  AOI22_X1 U9053 ( .A1(n9712), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7710), .B2(
        n9710), .ZN(n7339) );
  NAND2_X1 U9054 ( .A1(n9672), .A2(n6327), .ZN(n7338) );
  OAI211_X1 U9055 ( .C1(n7584), .C2(n9675), .A(n7339), .B(n7338), .ZN(n7340)
         );
  AOI21_X1 U9056 ( .B1(n9677), .B2(n7587), .A(n7340), .ZN(n7341) );
  OAI21_X1 U9057 ( .B1(n7342), .B2(n9694), .A(n7341), .ZN(P1_U3281) );
  OAI22_X1 U9058 ( .A1(n4520), .A2(n6725), .B1(n7568), .B2(n8892), .ZN(n7343)
         );
  XNOR2_X1 U9059 ( .A(n7343), .B(n8927), .ZN(n7398) );
  NAND2_X1 U9060 ( .A1(n8924), .A2(n9352), .ZN(n7344) );
  OAI21_X1 U9061 ( .B1(n4520), .B2(n8892), .A(n7344), .ZN(n7394) );
  INV_X1 U9062 ( .A(n7394), .ZN(n7399) );
  XNOR2_X1 U9063 ( .A(n7398), .B(n7399), .ZN(n7347) );
  NAND2_X1 U9064 ( .A1(n7345), .A2(n7407), .ZN(n7346) );
  NAND2_X1 U9065 ( .A1(n7346), .A2(n7347), .ZN(n7563) );
  OAI21_X1 U9066 ( .B1(n7347), .B2(n7346), .A(n7563), .ZN(n7348) );
  NAND2_X1 U9067 ( .A1(n7348), .A2(n9043), .ZN(n7353) );
  OAI22_X1 U9068 ( .A1(n6800), .A2(n9032), .B1(n9047), .B2(n7349), .ZN(n7350)
         );
  AOI211_X1 U9069 ( .C1(n9019), .C2(n9351), .A(n7351), .B(n7350), .ZN(n7352)
         );
  OAI211_X1 U9070 ( .C1(n4520), .C2(n9053), .A(n7353), .B(n7352), .ZN(P1_U3237) );
  INV_X1 U9071 ( .A(n7354), .ZN(n7355) );
  OR2_X1 U9072 ( .A1(n7356), .A2(n7355), .ZN(n9261) );
  XOR2_X1 U9073 ( .A(n7357), .B(n9261), .Z(n7358) );
  AOI222_X1 U9074 ( .A1(n9708), .A2(n7358), .B1(n9346), .B2(n9703), .C1(n9348), 
        .C2(n9705), .ZN(n9904) );
  XOR2_X1 U9075 ( .A(n7359), .B(n9261), .Z(n9907) );
  AOI21_X1 U9076 ( .B1(n7361), .B2(n7360), .A(n7605), .ZN(n9901) );
  NAND2_X1 U9077 ( .A1(n9901), .A2(n9700), .ZN(n7363) );
  AOI22_X1 U9078 ( .A1(n9712), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7522), .B2(
        n9710), .ZN(n7362) );
  OAI211_X1 U9079 ( .C1(n9902), .C2(n9714), .A(n7363), .B(n7362), .ZN(n7364)
         );
  AOI21_X1 U9080 ( .B1(n9677), .B2(n9907), .A(n7364), .ZN(n7365) );
  OAI21_X1 U9081 ( .B1(n9904), .B2(n9694), .A(n7365), .ZN(P1_U3280) );
  INV_X1 U9082 ( .A(n7366), .ZN(n7368) );
  NAND2_X1 U9083 ( .A1(n7368), .A2(n7367), .ZN(n7374) );
  OR2_X1 U9084 ( .A1(n7369), .A2(n8390), .ZN(n7762) );
  AND2_X1 U9085 ( .A1(n8610), .A2(n7762), .ZN(n7370) );
  MUX2_X1 U9086 ( .A(n7372), .B(n7371), .S(n8645), .Z(n7382) );
  OR2_X1 U9087 ( .A1(n7374), .A2(n7373), .ZN(n7926) );
  INV_X1 U9088 ( .A(n7376), .ZN(n7377) );
  OAI22_X1 U9089 ( .A1(n8620), .A2(n7378), .B1(n8527), .B2(n7377), .ZN(n7379)
         );
  AOI21_X1 U9090 ( .B1(n8600), .B2(n7380), .A(n7379), .ZN(n7381) );
  OAI211_X1 U9091 ( .C1(n7383), .C2(n8597), .A(n7382), .B(n7381), .ZN(P2_U3291) );
  XOR2_X1 U9092 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9365), .Z(n9360) );
  OAI22_X1 U9093 ( .A1(n7385), .A2(n7384), .B1(n7387), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n9361) );
  XOR2_X1 U9094 ( .A(n9361), .B(n9360), .Z(n7393) );
  NAND2_X1 U9095 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7727) );
  OAI21_X1 U9096 ( .B1(n9918), .B2(n9359), .A(n7727), .ZN(n7391) );
  XNOR2_X1 U9097 ( .A(n9365), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7388) );
  AOI211_X1 U9098 ( .C1(n7389), .C2(n7388), .A(n9438), .B(n9364), .ZN(n7390)
         );
  AOI211_X1 U9099 ( .C1(n9927), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7391), .B(
        n7390), .ZN(n7392) );
  OAI21_X1 U9100 ( .B1(n9923), .B2(n7393), .A(n7392), .ZN(P1_U3254) );
  NAND2_X1 U9101 ( .A1(n7398), .A2(n7394), .ZN(n7401) );
  INV_X1 U9102 ( .A(n7401), .ZN(n7406) );
  INV_X2 U9103 ( .A(n8832), .ZN(n8923) );
  NAND2_X1 U9104 ( .A1(n9351), .A2(n8923), .ZN(n7396) );
  NAND2_X1 U9105 ( .A1(n7396), .A2(n7395), .ZN(n7397) );
  XNOR2_X1 U9106 ( .A(n7397), .B(n8927), .ZN(n7410) );
  AOI22_X1 U9107 ( .A1(n8924), .A2(n9351), .B1(n7561), .B2(n8883), .ZN(n7408)
         );
  XNOR2_X1 U9108 ( .A(n7410), .B(n7408), .ZN(n7565) );
  INV_X1 U9109 ( .A(n7398), .ZN(n7400) );
  NAND2_X1 U9110 ( .A1(n7400), .A2(n7399), .ZN(n7562) );
  AND2_X1 U9111 ( .A1(n7565), .A2(n7562), .ZN(n7405) );
  NAND3_X1 U9112 ( .A1(n7403), .A2(n7402), .A3(n7401), .ZN(n7404) );
  OAI211_X2 U9113 ( .C1(n7407), .C2(n7406), .A(n7405), .B(n7404), .ZN(n7564)
         );
  INV_X1 U9114 ( .A(n7408), .ZN(n7409) );
  NAND2_X1 U9115 ( .A1(n7410), .A2(n7409), .ZN(n7418) );
  NAND2_X1 U9116 ( .A1(n7414), .A2(n8883), .ZN(n7412) );
  NAND2_X1 U9117 ( .A1(n8924), .A2(n9350), .ZN(n7411) );
  NAND2_X1 U9118 ( .A1(n7412), .A2(n7411), .ZN(n7492) );
  INV_X1 U9119 ( .A(n7492), .ZN(n7413) );
  AND2_X1 U9120 ( .A1(n7418), .A2(n7413), .ZN(n7503) );
  AND2_X1 U9121 ( .A1(n7564), .A2(n7503), .ZN(n7419) );
  NAND2_X1 U9122 ( .A1(n9350), .A2(n8883), .ZN(n7415) );
  NAND2_X1 U9123 ( .A1(n7416), .A2(n7415), .ZN(n7417) );
  XNOR2_X1 U9124 ( .A(n7417), .B(n8880), .ZN(n7506) );
  NOR2_X1 U9125 ( .A1(n7419), .A2(n7506), .ZN(n7637) );
  INV_X1 U9126 ( .A(n7637), .ZN(n7421) );
  NAND2_X1 U9127 ( .A1(n7564), .A2(n7418), .ZN(n7494) );
  AND2_X1 U9128 ( .A1(n7494), .A2(n7492), .ZN(n7636) );
  OAI21_X1 U9129 ( .B1(n7636), .B2(n7419), .A(n7506), .ZN(n7420) );
  OAI211_X1 U9130 ( .C1(n7421), .C2(n7636), .A(n9043), .B(n7420), .ZN(n7427)
         );
  OAI22_X1 U9131 ( .A1(n7423), .A2(n9032), .B1(n9047), .B2(n7422), .ZN(n7424)
         );
  AOI211_X1 U9132 ( .C1(n9019), .C2(n9349), .A(n7425), .B(n7424), .ZN(n7426)
         );
  OAI211_X1 U9133 ( .C1(n9999), .C2(n9053), .A(n7427), .B(n7426), .ZN(P1_U3219) );
  NAND2_X1 U9134 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n8257), .ZN(n7428) );
  OAI21_X1 U9135 ( .B1(n8217), .B2(n8257), .A(n7428), .ZN(P2_U3579) );
  INV_X1 U9136 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7429) );
  OAI22_X1 U9137 ( .A1(n4273), .A2(n7430), .B1(n7429), .B2(n8527), .ZN(n7433)
         );
  NOR2_X1 U9138 ( .A1(n8597), .A2(n7431), .ZN(n7432) );
  AOI211_X1 U9139 ( .C1(n4273), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7433), .B(
        n7432), .ZN(n7436) );
  NAND2_X1 U9140 ( .A1(n8600), .A2(n8763), .ZN(n8630) );
  OAI21_X1 U9141 ( .B1(n8643), .B2(n8637), .A(n7434), .ZN(n7435) );
  NAND2_X1 U9142 ( .A1(n7436), .A2(n7435), .ZN(P2_U3296) );
  XNOR2_X1 U9143 ( .A(n7437), .B(n7439), .ZN(n10050) );
  OAI21_X1 U9144 ( .B1(n7439), .B2(n7438), .A(n7548), .ZN(n7440) );
  AOI222_X1 U9145 ( .A1(n8614), .A2(n7440), .B1(n8256), .B2(n8582), .C1(n8259), 
        .C2(n8580), .ZN(n10054) );
  MUX2_X1 U9146 ( .A(n7441), .B(n10054), .S(n8645), .Z(n7450) );
  INV_X1 U9147 ( .A(n7554), .ZN(n7444) );
  NAND2_X1 U9148 ( .A1(n7442), .A2(n7448), .ZN(n7443) );
  NAND2_X1 U9149 ( .A1(n7444), .A2(n7443), .ZN(n10053) );
  INV_X1 U9150 ( .A(n7445), .ZN(n7446) );
  OAI22_X1 U9151 ( .A1(n8630), .A2(n10053), .B1(n7446), .B2(n8527), .ZN(n7447)
         );
  AOI21_X1 U9152 ( .B1(n8637), .B2(n7448), .A(n7447), .ZN(n7449) );
  OAI211_X1 U9153 ( .C1(n10050), .C2(n8597), .A(n7450), .B(n7449), .ZN(
        P2_U3290) );
  NAND2_X1 U9154 ( .A1(n7454), .A2(n7453), .ZN(n7455) );
  XNOR2_X1 U9155 ( .A(n7658), .B(n7998), .ZN(n7456) );
  NOR2_X1 U9156 ( .A1(n7694), .A2(n8012), .ZN(n7457) );
  XNOR2_X1 U9157 ( .A(n7456), .B(n7457), .ZN(n7592) );
  INV_X1 U9158 ( .A(n7456), .ZN(n7458) );
  AND2_X1 U9159 ( .A1(n7458), .A2(n7457), .ZN(n7459) );
  XNOR2_X1 U9160 ( .A(n8627), .B(n7124), .ZN(n7463) );
  INV_X1 U9161 ( .A(n7463), .ZN(n7461) );
  NOR2_X1 U9162 ( .A1(n7768), .A2(n8012), .ZN(n7462) );
  INV_X1 U9163 ( .A(n7462), .ZN(n7460) );
  NAND2_X1 U9164 ( .A1(n7461), .A2(n7460), .ZN(n7734) );
  NAND2_X1 U9165 ( .A1(n7463), .A2(n7462), .ZN(n7732) );
  NAND2_X1 U9166 ( .A1(n7734), .A2(n7732), .ZN(n7464) );
  XNOR2_X1 U9167 ( .A(n7733), .B(n7464), .ZN(n7469) );
  AOI22_X1 U9168 ( .A1(n8186), .A2(n4626), .B1(n8238), .B2(n8626), .ZN(n7468)
         );
  INV_X1 U9169 ( .A(n8627), .ZN(n7688) );
  NOR2_X1 U9170 ( .A1(n10148), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8329) );
  INV_X1 U9171 ( .A(n8329), .ZN(n7465) );
  OAI21_X1 U9172 ( .B1(n8226), .B2(n7688), .A(n7465), .ZN(n7466) );
  AOI21_X1 U9173 ( .B1(n8187), .B2(n8255), .A(n7466), .ZN(n7467) );
  OAI211_X1 U9174 ( .C1(n7469), .C2(n8230), .A(n7468), .B(n7467), .ZN(P2_U3233) );
  NAND2_X1 U9175 ( .A1(n7471), .A2(n7470), .ZN(n7473) );
  INV_X1 U9176 ( .A(n5896), .ZN(n7472) );
  XNOR2_X1 U9177 ( .A(n7473), .B(n7472), .ZN(n7476) );
  OAI22_X1 U9178 ( .A1(n7535), .A2(n8603), .B1(n7474), .B2(n8605), .ZN(n7475)
         );
  AOI21_X1 U9179 ( .B1(n7476), .B2(n8614), .A(n7475), .ZN(n10049) );
  OR2_X1 U9180 ( .A1(n7477), .A2(n10043), .ZN(n7478) );
  NAND2_X1 U9181 ( .A1(n7110), .A2(n7478), .ZN(n10044) );
  AOI22_X1 U9182 ( .A1(n4273), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n7479), .B2(
        n8641), .ZN(n7480) );
  OAI21_X1 U9183 ( .B1(n8630), .B2(n10044), .A(n7480), .ZN(n7481) );
  AOI21_X1 U9184 ( .B1(n8637), .B2(n5279), .A(n7481), .ZN(n7487) );
  INV_X1 U9185 ( .A(n7482), .ZN(n7483) );
  NAND2_X1 U9186 ( .A1(n7484), .A2(n7483), .ZN(n7485) );
  XNOR2_X1 U9187 ( .A(n7485), .B(n5896), .ZN(n10046) );
  NAND2_X1 U9188 ( .A1(n8555), .A2(n10046), .ZN(n7486) );
  OAI211_X1 U9189 ( .C1(n4273), .C2(n10049), .A(n7487), .B(n7486), .ZN(
        P2_U3292) );
  NAND2_X1 U9190 ( .A1(n9349), .A2(n8923), .ZN(n7488) );
  NAND2_X1 U9191 ( .A1(n7489), .A2(n7488), .ZN(n7490) );
  XNOR2_X1 U9192 ( .A(n7490), .B(n8880), .ZN(n7499) );
  NOR2_X1 U9193 ( .A1(n6727), .A2(n7712), .ZN(n7491) );
  AOI21_X1 U9194 ( .B1(n7640), .B2(n8883), .A(n7491), .ZN(n7500) );
  NAND2_X1 U9195 ( .A1(n7499), .A2(n7500), .ZN(n7704) );
  AND2_X1 U9196 ( .A1(n7704), .A2(n7492), .ZN(n7493) );
  NAND2_X1 U9197 ( .A1(n9348), .A2(n8883), .ZN(n7495) );
  NAND2_X1 U9198 ( .A1(n7496), .A2(n7495), .ZN(n7497) );
  XNOR2_X1 U9199 ( .A(n7497), .B(n8927), .ZN(n7511) );
  NOR2_X1 U9200 ( .A1(n6727), .A2(n7644), .ZN(n7498) );
  AOI21_X1 U9201 ( .B1(n6327), .B2(n8883), .A(n7498), .ZN(n7512) );
  XNOR2_X1 U9202 ( .A(n7511), .B(n7512), .ZN(n7705) );
  INV_X1 U9203 ( .A(n7499), .ZN(n7502) );
  INV_X1 U9204 ( .A(n7500), .ZN(n7501) );
  NAND2_X1 U9205 ( .A1(n7502), .A2(n7501), .ZN(n7635) );
  AND2_X1 U9206 ( .A1(n7503), .A2(n7635), .ZN(n7504) );
  NAND2_X1 U9207 ( .A1(n7564), .A2(n7505), .ZN(n7510) );
  NAND2_X1 U9208 ( .A1(n7635), .A2(n7506), .ZN(n7507) );
  NAND2_X1 U9209 ( .A1(n7507), .A2(n7704), .ZN(n7508) );
  NAND2_X1 U9210 ( .A1(n7705), .A2(n7508), .ZN(n7509) );
  INV_X1 U9211 ( .A(n7511), .ZN(n7513) );
  NAND2_X1 U9212 ( .A1(n7513), .A2(n7512), .ZN(n7517) );
  AND2_X1 U9213 ( .A1(n7519), .A2(n7517), .ZN(n7521) );
  XNOR2_X1 U9214 ( .A(n7514), .B(n8880), .ZN(n7672) );
  OR2_X1 U9215 ( .A1(n9902), .A2(n8892), .ZN(n7516) );
  NAND2_X1 U9216 ( .A1(n8924), .A2(n9347), .ZN(n7515) );
  NAND2_X1 U9217 ( .A1(n7516), .A2(n7515), .ZN(n7673) );
  XNOR2_X1 U9218 ( .A(n7672), .B(n7673), .ZN(n7520) );
  AND2_X1 U9219 ( .A1(n7520), .A2(n7517), .ZN(n7518) );
  OAI211_X1 U9220 ( .C1(n7521), .C2(n7520), .A(n9043), .B(n7676), .ZN(n7527)
         );
  INV_X1 U9221 ( .A(n7522), .ZN(n7523) );
  OAI22_X1 U9222 ( .A1(n7644), .A2(n9032), .B1(n9047), .B2(n7523), .ZN(n7524)
         );
  AOI211_X1 U9223 ( .C1(n9019), .C2(n9346), .A(n7525), .B(n7524), .ZN(n7526)
         );
  OAI211_X1 U9224 ( .C1(n9902), .C2(n9053), .A(n7527), .B(n7526), .ZN(P1_U3234) );
  INV_X1 U9225 ( .A(n7528), .ZN(n7529) );
  AOI21_X1 U9226 ( .B1(n8761), .B2(n7530), .A(n7529), .ZN(n8764) );
  NAND2_X1 U9227 ( .A1(n7540), .A2(n7531), .ZN(n7532) );
  NAND2_X1 U9228 ( .A1(n7533), .A2(n7532), .ZN(n7537) );
  OAI22_X1 U9229 ( .A1(n7535), .A2(n8605), .B1(n7534), .B2(n8603), .ZN(n7536)
         );
  AOI21_X1 U9230 ( .B1(n7537), .B2(n8614), .A(n7536), .ZN(n8766) );
  AOI22_X1 U9231 ( .A1(n8641), .A2(P2_REG3_REG_2__SCAN_IN), .B1(
        P2_REG2_REG_2__SCAN_IN), .B2(n4273), .ZN(n7538) );
  OAI21_X1 U9232 ( .B1(n4273), .B2(n8766), .A(n7538), .ZN(n7543) );
  XNOR2_X1 U9233 ( .A(n7539), .B(n7540), .ZN(n8768) );
  OAI22_X1 U9234 ( .A1(n7541), .A2(n8620), .B1(n8597), .B2(n8768), .ZN(n7542)
         );
  AOI211_X1 U9235 ( .C1(n8643), .C2(n8764), .A(n7543), .B(n7542), .ZN(n7544)
         );
  INV_X1 U9236 ( .A(n7544), .ZN(P2_U3294) );
  XNOR2_X1 U9237 ( .A(n7546), .B(n7549), .ZN(n10059) );
  NAND2_X1 U9238 ( .A1(n7548), .A2(n7547), .ZN(n7550) );
  XNOR2_X1 U9239 ( .A(n7550), .B(n7549), .ZN(n7551) );
  AOI222_X1 U9240 ( .A1(n8614), .A2(n7551), .B1(n8255), .B2(n8582), .C1(n8258), 
        .C2(n8580), .ZN(n10062) );
  MUX2_X1 U9241 ( .A(n7552), .B(n10062), .S(n8645), .Z(n7560) );
  INV_X1 U9242 ( .A(n7654), .ZN(n7553) );
  OAI211_X1 U9243 ( .C1(n10061), .C2(n7554), .A(n7553), .B(n8763), .ZN(n10060)
         );
  INV_X1 U9244 ( .A(n7555), .ZN(n7556) );
  OAI22_X1 U9245 ( .A1(n7926), .A2(n10060), .B1(n7556), .B2(n8527), .ZN(n7557)
         );
  AOI21_X1 U9246 ( .B1(n8637), .B2(n7558), .A(n7557), .ZN(n7559) );
  OAI211_X1 U9247 ( .C1(n10059), .C2(n8597), .A(n7560), .B(n7559), .ZN(
        P2_U3289) );
  INV_X1 U9248 ( .A(n7561), .ZN(n9994) );
  AND2_X1 U9249 ( .A1(n7563), .A2(n7562), .ZN(n7566) );
  OAI211_X1 U9250 ( .C1(n7566), .C2(n7565), .A(n9043), .B(n7564), .ZN(n7574)
         );
  OAI22_X1 U9251 ( .A1(n7568), .A2(n9032), .B1(n9047), .B2(n7567), .ZN(n7572)
         );
  OAI21_X1 U9252 ( .B1(n9048), .B2(n7570), .A(n7569), .ZN(n7571) );
  NOR2_X1 U9253 ( .A1(n7572), .A2(n7571), .ZN(n7573) );
  OAI211_X1 U9254 ( .C1(n9994), .C2(n9053), .A(n7574), .B(n7573), .ZN(P1_U3211) );
  INV_X1 U9255 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7575) );
  OAI22_X1 U9256 ( .A1(n7926), .A2(n7576), .B1(n7575), .B2(n8527), .ZN(n7579)
         );
  NOR2_X1 U9257 ( .A1(n7577), .A2(n4273), .ZN(n7578) );
  AOI211_X1 U9258 ( .C1(n4273), .C2(P2_REG2_REG_1__SCAN_IN), .A(n7579), .B(
        n7578), .ZN(n7582) );
  NAND2_X1 U9259 ( .A1(n8637), .A2(n7580), .ZN(n7581) );
  OAI211_X1 U9260 ( .C1(n8597), .C2(n7583), .A(n7582), .B(n7581), .ZN(P2_U3295) );
  OAI21_X1 U9261 ( .B1(n7717), .B2(n9998), .A(n7584), .ZN(n7586) );
  AOI211_X1 U9262 ( .C1(n10010), .C2(n7587), .A(n7586), .B(n7585), .ZN(n7590)
         );
  NAND2_X1 U9263 ( .A1(n10015), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7588) );
  OAI21_X1 U9264 ( .B1(n7590), .B2(n10015), .A(n7588), .ZN(P1_U3484) );
  NAND2_X1 U9265 ( .A1(n10026), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7589) );
  OAI21_X1 U9266 ( .B1(n7590), .B2(n10026), .A(n7589), .ZN(P1_U3533) );
  XOR2_X1 U9267 ( .A(n7592), .B(n7591), .Z(n7596) );
  NAND2_X1 U9268 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8315) );
  NAND2_X1 U9269 ( .A1(n8238), .A2(n4299), .ZN(n7593) );
  OAI211_X1 U9270 ( .C1(n8226), .C2(n10071), .A(n8315), .B(n7593), .ZN(n7595)
         );
  OAI22_X1 U9271 ( .A1(n7653), .A2(n8205), .B1(n8204), .B2(n7768), .ZN(n7594)
         );
  AOI211_X1 U9272 ( .C1(n7596), .C2(n8184), .A(n7595), .B(n7594), .ZN(n7597)
         );
  INV_X1 U9273 ( .A(n7597), .ZN(P2_U3223) );
  INV_X1 U9274 ( .A(n7629), .ZN(n7600) );
  OR2_X1 U9275 ( .A1(n7598), .A2(P1_U3084), .ZN(n9332) );
  INV_X1 U9276 ( .A(n9332), .ZN(n9325) );
  AOI21_X1 U9277 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9864), .A(n9325), .ZN(
        n7599) );
  OAI21_X1 U9278 ( .B1(n7600), .B2(n9866), .A(n7599), .ZN(P1_U3330) );
  AOI21_X1 U9279 ( .B1(n7601), .B2(n9248), .A(n9557), .ZN(n7604) );
  OAI22_X1 U9280 ( .A1(n9656), .A2(n9095), .B1(n7681), .B2(n9654), .ZN(n7602)
         );
  AOI21_X1 U9281 ( .B1(n7604), .B2(n7603), .A(n7602), .ZN(n9826) );
  INV_X1 U9282 ( .A(n7605), .ZN(n7606) );
  AOI211_X1 U9283 ( .C1(n9824), .C2(n7606), .A(n10000), .B(n7788), .ZN(n9823)
         );
  INV_X1 U9284 ( .A(n9675), .ZN(n9719) );
  AOI22_X1 U9285 ( .A1(n9712), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7678), .B2(
        n9710), .ZN(n7607) );
  OAI21_X1 U9286 ( .B1(n7608), .B2(n9714), .A(n7607), .ZN(n7612) );
  OAI21_X1 U9287 ( .B1(n7610), .B2(n9248), .A(n7609), .ZN(n9827) );
  NOR2_X1 U9288 ( .A1(n9827), .A2(n9716), .ZN(n7611) );
  AOI211_X1 U9289 ( .C1(n9823), .C2(n9719), .A(n7612), .B(n7611), .ZN(n7613)
         );
  OAI21_X1 U9290 ( .B1(n9826), .B2(n9694), .A(n7613), .ZN(P1_U3279) );
  NAND2_X1 U9291 ( .A1(n7624), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7616) );
  XOR2_X1 U9292 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8361), .Z(n7617) );
  NAND2_X1 U9293 ( .A1(n7617), .A2(n7618), .ZN(n8357) );
  OAI211_X1 U9294 ( .C1(n7618), .C2(n7617), .A(n8388), .B(n8357), .ZN(n7621)
         );
  AND2_X1 U9295 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7619) );
  AOI21_X1 U9296 ( .B1(n8366), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7619), .ZN(
        n7620) );
  OAI211_X1 U9297 ( .C1(n8382), .C2(n7622), .A(n7621), .B(n7620), .ZN(n7628)
         );
  OAI21_X1 U9298 ( .B1(n7624), .B2(P2_REG1_REG_16__SCAN_IN), .A(n7623), .ZN(
        n7626) );
  XNOR2_X1 U9299 ( .A(n8361), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7625) );
  NOR2_X1 U9300 ( .A1(n7625), .A2(n7626), .ZN(n8360) );
  AOI211_X1 U9301 ( .C1(n7626), .C2(n7625), .A(n8360), .B(n8383), .ZN(n7627)
         );
  OR2_X1 U9302 ( .A1(n7628), .A2(n7627), .ZN(P2_U3262) );
  NAND2_X1 U9303 ( .A1(n7629), .A2(n8795), .ZN(n7631) );
  OAI211_X1 U9304 ( .C1(n7632), .C2(n8802), .A(n7631), .B(n7630), .ZN(P2_U3335) );
  NAND2_X1 U9305 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8257), .ZN(n7633) );
  OAI21_X1 U9306 ( .B1(n7634), .B2(n8257), .A(n7633), .ZN(P2_U3581) );
  NAND2_X1 U9307 ( .A1(n7704), .A2(n7635), .ZN(n7639) );
  OR2_X1 U9308 ( .A1(n7637), .A2(n7636), .ZN(n7638) );
  NOR3_X1 U9309 ( .A1(n7637), .A2(n7636), .A3(n7639), .ZN(n7707) );
  AOI21_X1 U9310 ( .B1(n7639), .B2(n7638), .A(n7707), .ZN(n7648) );
  AND2_X1 U9311 ( .A1(n7640), .A2(n9957), .ZN(n10007) );
  AOI22_X1 U9312 ( .A1(n9050), .A2(n9350), .B1(n9035), .B2(n7641), .ZN(n7643)
         );
  OAI211_X1 U9313 ( .C1(n7644), .C2(n9048), .A(n7643), .B(n7642), .ZN(n7645)
         );
  AOI21_X1 U9314 ( .B1(n7646), .B2(n10007), .A(n7645), .ZN(n7647) );
  OAI21_X1 U9315 ( .B1(n7648), .B2(n9024), .A(n7647), .ZN(P1_U3229) );
  INV_X1 U9316 ( .A(n7691), .ZN(n7650) );
  AOI21_X1 U9317 ( .B1(n5908), .B2(n7651), .A(n7650), .ZN(n7652) );
  OAI222_X1 U9318 ( .A1(n8605), .A2(n7768), .B1(n8603), .B2(n7653), .C1(n8535), 
        .C2(n7652), .ZN(n10073) );
  MUX2_X1 U9319 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10073), .S(n8645), .Z(n7662)
         );
  OAI211_X1 U9320 ( .C1(n7654), .C2(n10071), .A(n8763), .B(n7686), .ZN(n10068)
         );
  NAND2_X1 U9321 ( .A1(n7657), .A2(n7656), .ZN(n10067) );
  NAND3_X1 U9322 ( .A1(n7655), .A2(n10067), .A3(n8555), .ZN(n7660) );
  AOI22_X1 U9323 ( .A1(n8637), .A2(n7658), .B1(n8641), .B2(n4299), .ZN(n7659)
         );
  OAI211_X1 U9324 ( .C1(n7926), .C2(n10068), .A(n7660), .B(n7659), .ZN(n7661)
         );
  OR2_X1 U9325 ( .A1(n7662), .A2(n7661), .ZN(P2_U3288) );
  NAND2_X1 U9326 ( .A1(n9346), .A2(n8883), .ZN(n7663) );
  NAND2_X1 U9327 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  XNOR2_X1 U9328 ( .A(n7665), .B(n8880), .ZN(n7671) );
  INV_X1 U9329 ( .A(n7671), .ZN(n7669) );
  NOR2_X1 U9330 ( .A1(n6727), .A2(n7666), .ZN(n7667) );
  AOI21_X1 U9331 ( .B1(n9824), .B2(n8883), .A(n7667), .ZN(n7670) );
  INV_X1 U9332 ( .A(n7670), .ZN(n7668) );
  NAND2_X1 U9333 ( .A1(n7669), .A2(n7668), .ZN(n7720) );
  NAND2_X1 U9334 ( .A1(n7671), .A2(n7670), .ZN(n7718) );
  NAND2_X1 U9335 ( .A1(n7720), .A2(n7718), .ZN(n7677) );
  INV_X1 U9336 ( .A(n7672), .ZN(n7674) );
  NAND2_X1 U9337 ( .A1(n7674), .A2(n7673), .ZN(n7675) );
  XOR2_X1 U9338 ( .A(n7677), .B(n7719), .Z(n7684) );
  AOI22_X1 U9339 ( .A1(n9019), .A2(n9706), .B1(n9035), .B2(n7678), .ZN(n7680)
         );
  OAI211_X1 U9340 ( .C1(n7681), .C2(n9032), .A(n7680), .B(n7679), .ZN(n7682)
         );
  AOI21_X1 U9341 ( .B1(n9022), .B2(n9824), .A(n7682), .ZN(n7683) );
  OAI21_X1 U9342 ( .B1(n7684), .B2(n9024), .A(n7683), .ZN(P1_U3222) );
  INV_X1 U9343 ( .A(n8759), .ZN(n7700) );
  OAI21_X1 U9344 ( .B1(n4371), .B2(n7690), .A(n7685), .ZN(n8634) );
  NAND2_X1 U9345 ( .A1(n7686), .A2(n8627), .ZN(n7687) );
  NAND2_X1 U9346 ( .A1(n7775), .A2(n7687), .ZN(n8629) );
  OAI22_X1 U9347 ( .A1(n8629), .A2(n10052), .B1(n7688), .B2(n10070), .ZN(n7699) );
  NAND2_X1 U9348 ( .A1(n8634), .A2(n7763), .ZN(n7698) );
  NAND3_X1 U9349 ( .A1(n7691), .A2(n7690), .A3(n7689), .ZN(n7692) );
  NAND2_X1 U9350 ( .A1(n7693), .A2(n7692), .ZN(n7696) );
  OAI22_X1 U9351 ( .A1(n7694), .A2(n8603), .B1(n7816), .B2(n8605), .ZN(n7695)
         );
  AOI21_X1 U9352 ( .B1(n7696), .B2(n8614), .A(n7695), .ZN(n7697) );
  NAND2_X1 U9353 ( .A1(n7698), .A2(n7697), .ZN(n8631) );
  AOI211_X1 U9354 ( .C1(n7700), .C2(n8634), .A(n7699), .B(n8631), .ZN(n7703)
         );
  NAND2_X1 U9355 ( .A1(n10081), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7701) );
  OAI21_X1 U9356 ( .B1(n7703), .B2(n10081), .A(n7701), .ZN(P2_U3529) );
  NAND2_X1 U9357 ( .A1(n10074), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7702) );
  OAI21_X1 U9358 ( .B1(n7703), .B2(n10074), .A(n7702), .ZN(P2_U3478) );
  INV_X1 U9359 ( .A(n7704), .ZN(n7706) );
  NOR3_X1 U9360 ( .A1(n7707), .A2(n7706), .A3(n7705), .ZN(n7709) );
  INV_X1 U9361 ( .A(n7519), .ZN(n7708) );
  OAI21_X1 U9362 ( .B1(n7709), .B2(n7708), .A(n9043), .ZN(n7716) );
  INV_X1 U9363 ( .A(n7710), .ZN(n7711) );
  OAI22_X1 U9364 ( .A1(n7712), .A2(n9032), .B1(n9047), .B2(n7711), .ZN(n7713)
         );
  AOI211_X1 U9365 ( .C1(n9019), .C2(n9347), .A(n7714), .B(n7713), .ZN(n7715)
         );
  OAI211_X1 U9366 ( .C1(n7717), .C2(n9053), .A(n7716), .B(n7715), .ZN(P1_U3215) );
  NAND2_X1 U9367 ( .A1(n9818), .A2(n8923), .ZN(n7722) );
  NAND2_X1 U9368 ( .A1(n8924), .A2(n9706), .ZN(n7721) );
  NAND2_X1 U9369 ( .A1(n7722), .A2(n7721), .ZN(n7822) );
  NAND2_X1 U9370 ( .A1(n9706), .A2(n8923), .ZN(n7723) );
  NAND2_X1 U9371 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  XNOR2_X1 U9372 ( .A(n7725), .B(n8927), .ZN(n7823) );
  XOR2_X1 U9373 ( .A(n7822), .B(n7823), .Z(n7726) );
  XNOR2_X1 U9374 ( .A(n7824), .B(n7726), .ZN(n7731) );
  AOI22_X1 U9375 ( .A1(n9050), .A2(n9346), .B1(n9035), .B2(n7790), .ZN(n7728)
         );
  OAI211_X1 U9376 ( .C1(n9098), .C2(n9048), .A(n7728), .B(n7727), .ZN(n7729)
         );
  AOI21_X1 U9377 ( .B1(n9022), .B2(n9818), .A(n7729), .ZN(n7730) );
  OAI21_X1 U9378 ( .B1(n7731), .B2(n9024), .A(n7730), .ZN(P1_U3232) );
  XNOR2_X1 U9379 ( .A(n7774), .B(n7124), .ZN(n7736) );
  NOR2_X1 U9380 ( .A1(n7816), .A2(n8012), .ZN(n7737) );
  NAND2_X1 U9381 ( .A1(n7736), .A2(n7737), .ZN(n7807) );
  INV_X1 U9382 ( .A(n7736), .ZN(n7806) );
  INV_X1 U9383 ( .A(n7737), .ZN(n7738) );
  NAND2_X1 U9384 ( .A1(n7806), .A2(n7738), .ZN(n7739) );
  NAND2_X1 U9385 ( .A1(n7807), .A2(n7739), .ZN(n7741) );
  AOI21_X1 U9386 ( .B1(n7740), .B2(n7741), .A(n8230), .ZN(n7743) );
  INV_X1 U9387 ( .A(n7741), .ZN(n7742) );
  NAND2_X1 U9388 ( .A1(n7743), .A2(n7808), .ZN(n7746) );
  AND2_X1 U9389 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8343) );
  OAI22_X1 U9390 ( .A1(n7919), .A2(n8204), .B1(n8205), .B2(n7768), .ZN(n7744)
         );
  AOI211_X1 U9391 ( .C1(n8238), .C2(n7777), .A(n8343), .B(n7744), .ZN(n7745)
         );
  OAI211_X1 U9392 ( .C1(n8754), .C2(n8226), .A(n7746), .B(n7745), .ZN(P2_U3219) );
  XOR2_X1 U9393 ( .A(n7747), .B(n7750), .Z(n7748) );
  INV_X1 U9394 ( .A(n8172), .ZN(n8252) );
  AOI222_X1 U9395 ( .A1(n8614), .A2(n7748), .B1(n4626), .B2(n8580), .C1(n8252), 
        .C2(n8582), .ZN(n8752) );
  NAND2_X1 U9396 ( .A1(n7749), .A2(n7750), .ZN(n7849) );
  OAI21_X1 U9397 ( .B1(n7749), .B2(n7750), .A(n7849), .ZN(n8753) );
  INV_X1 U9398 ( .A(n8753), .ZN(n7755) );
  NOR2_X1 U9399 ( .A1(n4366), .A2(n8748), .ZN(n7751) );
  OR2_X1 U9400 ( .A1(n7842), .A2(n7751), .ZN(n8749) );
  AOI22_X1 U9401 ( .A1(n4273), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7813), .B2(
        n8641), .ZN(n7753) );
  NAND2_X1 U9402 ( .A1(n8637), .A2(n7819), .ZN(n7752) );
  OAI211_X1 U9403 ( .C1(n8749), .C2(n8630), .A(n7753), .B(n7752), .ZN(n7754)
         );
  AOI21_X1 U9404 ( .B1(n7755), .B2(n8555), .A(n7754), .ZN(n7756) );
  OAI21_X1 U9405 ( .B1(n8752), .B2(n4273), .A(n7756), .ZN(P2_U3285) );
  INV_X1 U9406 ( .A(n7757), .ZN(n7784) );
  OAI222_X1 U9407 ( .A1(n9866), .A2(n7784), .B1(P1_U3084), .B2(n7760), .C1(
        n7759), .C2(n7758), .ZN(P1_U3329) );
  XNOR2_X1 U9408 ( .A(n7761), .B(n4623), .ZN(n7764) );
  INV_X1 U9409 ( .A(n7764), .ZN(n8760) );
  NOR2_X1 U9410 ( .A1(n4273), .A2(n7762), .ZN(n8639) );
  INV_X1 U9411 ( .A(n8639), .ZN(n8622) );
  NAND2_X1 U9412 ( .A1(n7764), .A2(n7763), .ZN(n7772) );
  XNOR2_X1 U9413 ( .A(n7766), .B(n7765), .ZN(n7770) );
  NAND2_X1 U9414 ( .A1(n8253), .A2(n8582), .ZN(n7767) );
  OAI21_X1 U9415 ( .B1(n7768), .B2(n8603), .A(n7767), .ZN(n7769) );
  AOI21_X1 U9416 ( .B1(n7770), .B2(n8614), .A(n7769), .ZN(n7771) );
  AND2_X1 U9417 ( .A1(n7772), .A2(n7771), .ZN(n8758) );
  MUX2_X1 U9418 ( .A(n8758), .B(n7773), .S(n4273), .Z(n7782) );
  AND2_X1 U9419 ( .A1(n7775), .A2(n7774), .ZN(n7776) );
  OR2_X1 U9420 ( .A1(n7776), .A2(n4366), .ZN(n8755) );
  INV_X1 U9421 ( .A(n8755), .ZN(n7780) );
  INV_X1 U9422 ( .A(n7777), .ZN(n7778) );
  OAI22_X1 U9423 ( .A1(n8620), .A2(n8754), .B1(n8527), .B2(n7778), .ZN(n7779)
         );
  AOI21_X1 U9424 ( .B1(n7780), .B2(n8643), .A(n7779), .ZN(n7781) );
  OAI211_X1 U9425 ( .C1(n8760), .C2(n8622), .A(n7782), .B(n7781), .ZN(P2_U3286) );
  OAI222_X1 U9426 ( .A1(P2_U3152), .A2(n7785), .B1(n4275), .B2(n7784), .C1(
        n7783), .C2(n8802), .ZN(P2_U3334) );
  OAI21_X1 U9427 ( .B1(n9265), .B2(n4370), .A(n7786), .ZN(n7787) );
  AOI222_X1 U9428 ( .A1(n9708), .A2(n7787), .B1(n9346), .B2(n9705), .C1(n9685), 
        .C2(n9703), .ZN(n9821) );
  OR2_X1 U9429 ( .A1(n7788), .A2(n7792), .ZN(n7789) );
  AND2_X1 U9430 ( .A1(n4369), .A2(n7789), .ZN(n9819) );
  AOI22_X1 U9431 ( .A1(n9712), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7790), .B2(
        n9710), .ZN(n7791) );
  OAI21_X1 U9432 ( .B1(n7792), .B2(n9714), .A(n7791), .ZN(n7796) );
  INV_X1 U9433 ( .A(n9265), .ZN(n7793) );
  XNOR2_X1 U9434 ( .A(n4491), .B(n7793), .ZN(n9822) );
  NOR2_X1 U9435 ( .A1(n9822), .A2(n9716), .ZN(n7795) );
  AOI211_X1 U9436 ( .C1(n9819), .C2(n9700), .A(n7796), .B(n7795), .ZN(n7797)
         );
  OAI21_X1 U9437 ( .B1(n9821), .B2(n9712), .A(n7797), .ZN(P1_U3278) );
  INV_X1 U9438 ( .A(n7798), .ZN(n7837) );
  AOI22_X1 U9439 ( .A1(n7799), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n9864), .ZN(n7800) );
  OAI21_X1 U9440 ( .B1(n7837), .B2(n9866), .A(n7800), .ZN(P1_U3328) );
  XNOR2_X1 U9441 ( .A(n7819), .B(n7124), .ZN(n7911) );
  AND2_X1 U9442 ( .A1(n8253), .A2(n7991), .ZN(n7801) );
  NAND2_X1 U9443 ( .A1(n7911), .A2(n7801), .ZN(n7908) );
  INV_X1 U9444 ( .A(n7911), .ZN(n7803) );
  INV_X1 U9445 ( .A(n7801), .ZN(n7802) );
  NAND2_X1 U9446 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  AND2_X1 U9447 ( .A1(n7908), .A2(n7804), .ZN(n7809) );
  INV_X1 U9448 ( .A(n7809), .ZN(n7805) );
  AOI21_X1 U9449 ( .B1(n7808), .B2(n7805), .A(n8230), .ZN(n7812) );
  NOR3_X1 U9450 ( .A1(n8209), .A2(n7816), .A3(n7806), .ZN(n7811) );
  OAI21_X1 U9451 ( .B1(n7812), .B2(n7811), .A(n7910), .ZN(n7821) );
  NAND2_X1 U9452 ( .A1(n8238), .A2(n7813), .ZN(n7814) );
  OAI21_X1 U9453 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7815), .A(n7814), .ZN(n7818) );
  OAI22_X1 U9454 ( .A1(n8172), .A2(n8204), .B1(n8205), .B2(n7816), .ZN(n7817)
         );
  AOI211_X1 U9455 ( .C1(n7819), .C2(n8236), .A(n7818), .B(n7817), .ZN(n7820)
         );
  NAND2_X1 U9456 ( .A1(n7821), .A2(n7820), .ZN(P2_U3238) );
  NAND2_X1 U9457 ( .A1(n7824), .A2(n7823), .ZN(n7825) );
  NAND2_X1 U9458 ( .A1(n9685), .A2(n8923), .ZN(n7826) );
  NAND2_X1 U9459 ( .A1(n7827), .A2(n7826), .ZN(n7828) );
  XNOR2_X1 U9460 ( .A(n7828), .B(n8880), .ZN(n8827) );
  NAND2_X1 U9461 ( .A1(n4411), .A2(n8883), .ZN(n7830) );
  NAND2_X1 U9462 ( .A1(n9685), .A2(n8924), .ZN(n7829) );
  NAND2_X1 U9463 ( .A1(n7830), .A2(n7829), .ZN(n8812) );
  XNOR2_X1 U9464 ( .A(n8827), .B(n8812), .ZN(n7831) );
  XNOR2_X1 U9465 ( .A(n8813), .B(n7831), .ZN(n7835) );
  AOI22_X1 U9466 ( .A1(n9019), .A2(n9704), .B1(n9035), .B2(n9711), .ZN(n7832)
         );
  NAND2_X1 U9467 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9362) );
  OAI211_X1 U9468 ( .C1(n9095), .C2(n9032), .A(n7832), .B(n9362), .ZN(n7833)
         );
  AOI21_X1 U9469 ( .B1(n9022), .B2(n4411), .A(n7833), .ZN(n7834) );
  OAI21_X1 U9470 ( .B1(n7835), .B2(n9024), .A(n7834), .ZN(P1_U3213) );
  OAI222_X1 U9471 ( .A1(n8802), .A2(n7838), .B1(n4275), .B2(n7837), .C1(
        P2_U3152), .C2(n7836), .ZN(P2_U3333) );
  NAND2_X1 U9472 ( .A1(n7860), .A2(n7839), .ZN(n7840) );
  XNOR2_X1 U9473 ( .A(n7840), .B(n7850), .ZN(n7841) );
  AOI222_X1 U9474 ( .A1(n8614), .A2(n7841), .B1(n8251), .B2(n8582), .C1(n8253), 
        .C2(n8580), .ZN(n8746) );
  INV_X1 U9475 ( .A(n7842), .ZN(n7845) );
  INV_X1 U9476 ( .A(n7843), .ZN(n7844) );
  AOI21_X1 U9477 ( .B1(n8743), .B2(n7845), .A(n7844), .ZN(n8744) );
  AOI22_X1 U9478 ( .A1(n4273), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7916), .B2(
        n8641), .ZN(n7846) );
  OAI21_X1 U9479 ( .B1(n8620), .B2(n7847), .A(n7846), .ZN(n7853) );
  NAND2_X1 U9480 ( .A1(n7849), .A2(n7848), .ZN(n7851) );
  XNOR2_X1 U9481 ( .A(n7851), .B(n7850), .ZN(n8747) );
  NOR2_X1 U9482 ( .A1(n8747), .A2(n8597), .ZN(n7852) );
  AOI211_X1 U9483 ( .C1(n8744), .C2(n8643), .A(n7853), .B(n7852), .ZN(n7854)
         );
  OAI21_X1 U9484 ( .B1(n4273), .B2(n8746), .A(n7854), .ZN(P2_U3284) );
  AND2_X1 U9485 ( .A1(n7855), .A2(n7864), .ZN(n7857) );
  OR2_X1 U9486 ( .A1(n7857), .A2(n7856), .ZN(n8740) );
  OAI22_X1 U9487 ( .A1(n8172), .A2(n8603), .B1(n8171), .B2(n8605), .ZN(n7858)
         );
  INV_X1 U9488 ( .A(n7858), .ZN(n7869) );
  NAND2_X1 U9489 ( .A1(n7860), .A2(n7859), .ZN(n7866) );
  INV_X1 U9490 ( .A(n7864), .ZN(n7861) );
  AOI21_X1 U9491 ( .B1(n7866), .B2(n7862), .A(n7861), .ZN(n7879) );
  NOR2_X1 U9492 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  AND2_X1 U9493 ( .A1(n7866), .A2(n7865), .ZN(n7867) );
  OAI21_X1 U9494 ( .B1(n7879), .B2(n7867), .A(n8614), .ZN(n7868) );
  OAI211_X1 U9495 ( .C1(n8740), .C2(n8610), .A(n7869), .B(n7868), .ZN(n8742)
         );
  NAND2_X1 U9496 ( .A1(n8742), .A2(n8645), .ZN(n7874) );
  NAND2_X1 U9497 ( .A1(n7843), .A2(n8737), .ZN(n7870) );
  AND2_X1 U9498 ( .A1(n7887), .A2(n7870), .ZN(n8738) );
  INV_X1 U9499 ( .A(n8737), .ZN(n8178) );
  AOI22_X1 U9500 ( .A1(n4273), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8175), .B2(
        n8641), .ZN(n7871) );
  OAI21_X1 U9501 ( .B1(n8620), .B2(n8178), .A(n7871), .ZN(n7872) );
  AOI21_X1 U9502 ( .B1(n8738), .B2(n8643), .A(n7872), .ZN(n7873) );
  OAI211_X1 U9503 ( .C1(n8740), .C2(n8622), .A(n7874), .B(n7873), .ZN(P2_U3283) );
  INV_X1 U9504 ( .A(n7875), .ZN(n7894) );
  AOI22_X1 U9505 ( .A1(n7876), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9864), .ZN(n7877) );
  OAI21_X1 U9506 ( .B1(n7894), .B2(n9866), .A(n7877), .ZN(P1_U3327) );
  OAI21_X1 U9507 ( .B1(n7879), .B2(n7878), .A(n7885), .ZN(n7881) );
  NAND3_X1 U9508 ( .A1(n7881), .A2(n8614), .A3(n7880), .ZN(n7883) );
  OAI22_X1 U9509 ( .A1(n8604), .A2(n8605), .B1(n8071), .B2(n8603), .ZN(n7882)
         );
  INV_X1 U9510 ( .A(n7882), .ZN(n8076) );
  AND2_X1 U9511 ( .A1(n7883), .A2(n8076), .ZN(n8735) );
  OAI21_X1 U9512 ( .B1(n7886), .B2(n7885), .A(n7884), .ZN(n8731) );
  AOI21_X1 U9513 ( .B1(n7887), .B2(n8733), .A(n10052), .ZN(n7888) );
  AND2_X1 U9514 ( .A1(n7901), .A2(n7888), .ZN(n8732) );
  NAND2_X1 U9515 ( .A1(n8732), .A2(n8600), .ZN(n7890) );
  AOI22_X1 U9516 ( .A1(n4273), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8073), .B2(
        n8641), .ZN(n7889) );
  OAI211_X1 U9517 ( .C1(n4969), .C2(n8620), .A(n7890), .B(n7889), .ZN(n7891)
         );
  AOI21_X1 U9518 ( .B1(n8731), .B2(n8555), .A(n7891), .ZN(n7892) );
  OAI21_X1 U9519 ( .B1(n4273), .B2(n8735), .A(n7892), .ZN(P2_U3282) );
  OAI222_X1 U9520 ( .A1(P2_U3152), .A2(n7895), .B1(n4275), .B2(n7894), .C1(
        n7893), .C2(n8802), .ZN(P2_U3332) );
  XNOR2_X1 U9521 ( .A(n7896), .B(n4631), .ZN(n8730) );
  OAI211_X1 U9522 ( .C1(n7898), .C2(n4631), .A(n4386), .B(n8614), .ZN(n7900)
         );
  OAI22_X1 U9523 ( .A1(n8248), .A2(n8605), .B1(n8171), .B2(n8603), .ZN(n8234)
         );
  INV_X1 U9524 ( .A(n8234), .ZN(n7899) );
  NAND2_X1 U9525 ( .A1(n7900), .A2(n7899), .ZN(n8726) );
  AOI211_X1 U9526 ( .C1(n8728), .C2(n7901), .A(n10052), .B(n8615), .ZN(n8727)
         );
  NAND2_X1 U9527 ( .A1(n8727), .A2(n8600), .ZN(n7904) );
  INV_X1 U9528 ( .A(n7902), .ZN(n8237) );
  AOI22_X1 U9529 ( .A1(n4273), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8237), .B2(
        n8641), .ZN(n7903) );
  OAI211_X1 U9530 ( .C1(n7905), .C2(n8620), .A(n7904), .B(n7903), .ZN(n7906)
         );
  AOI21_X1 U9531 ( .B1(n8726), .B2(n8645), .A(n7906), .ZN(n7907) );
  OAI21_X1 U9532 ( .B1(n8730), .B2(n8597), .A(n7907), .ZN(P2_U3281) );
  XNOR2_X1 U9533 ( .A(n8743), .B(n7998), .ZN(n7940) );
  NOR2_X1 U9534 ( .A1(n8172), .A2(n8012), .ZN(n7938) );
  XNOR2_X1 U9535 ( .A(n7940), .B(n7938), .ZN(n7913) );
  AND2_X1 U9536 ( .A1(n7913), .A2(n7908), .ZN(n7909) );
  NAND3_X1 U9537 ( .A1(n8185), .A2(n8253), .A3(n7911), .ZN(n7912) );
  OAI21_X1 U9538 ( .B1(n7910), .B2(n8230), .A(n7912), .ZN(n7915) );
  INV_X1 U9539 ( .A(n7913), .ZN(n7914) );
  NAND2_X1 U9540 ( .A1(n7915), .A2(n7914), .ZN(n7923) );
  NAND2_X1 U9541 ( .A1(n8238), .A2(n7916), .ZN(n7918) );
  NAND2_X1 U9542 ( .A1(n7918), .A2(n7917), .ZN(n7921) );
  OAI22_X1 U9543 ( .A1(n7919), .A2(n8205), .B1(n8204), .B2(n8071), .ZN(n7920)
         );
  AOI211_X1 U9544 ( .C1(n8743), .C2(n8236), .A(n7921), .B(n7920), .ZN(n7922)
         );
  OAI211_X1 U9545 ( .C1(n8230), .C2(n7942), .A(n7923), .B(n7922), .ZN(P2_U3226) );
  NAND2_X1 U9546 ( .A1(n7924), .A2(n8555), .ZN(n7931) );
  INV_X1 U9547 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7925) );
  OAI22_X1 U9548 ( .A1(n8025), .A2(n8527), .B1(n7925), .B2(n8645), .ZN(n7929)
         );
  NOR2_X1 U9549 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  AOI211_X1 U9550 ( .C1(n8637), .C2(n8017), .A(n7929), .B(n7928), .ZN(n7930)
         );
  OAI211_X1 U9551 ( .C1(n4273), .C2(n7932), .A(n7931), .B(n7930), .ZN(P2_U3268) );
  INV_X1 U9552 ( .A(n8034), .ZN(n9858) );
  OAI222_X1 U9553 ( .A1(P2_U3152), .A2(n7934), .B1(n4275), .B2(n9858), .C1(
        n7933), .C2(n8802), .ZN(P2_U3329) );
  INV_X1 U9554 ( .A(n9065), .ZN(n9856) );
  OAI222_X1 U9555 ( .A1(P2_U3152), .A2(n7936), .B1(n4275), .B2(n9856), .C1(
        n7935), .C2(n8802), .ZN(P2_U3328) );
  INV_X1 U9556 ( .A(n7937), .ZN(n8029) );
  INV_X1 U9557 ( .A(n7938), .ZN(n7939) );
  NAND2_X1 U9558 ( .A1(n7940), .A2(n7939), .ZN(n7941) );
  XNOR2_X1 U9559 ( .A(n8737), .B(n7124), .ZN(n7943) );
  NOR2_X1 U9560 ( .A1(n8071), .A2(n8012), .ZN(n7944) );
  NAND2_X1 U9561 ( .A1(n7943), .A2(n7944), .ZN(n7947) );
  INV_X1 U9562 ( .A(n7943), .ZN(n8070) );
  INV_X1 U9563 ( .A(n7944), .ZN(n7945) );
  NAND2_X1 U9564 ( .A1(n8070), .A2(n7945), .ZN(n7946) );
  NAND2_X1 U9565 ( .A1(n7947), .A2(n7946), .ZN(n8168) );
  XNOR2_X1 U9566 ( .A(n8733), .B(n7998), .ZN(n7951) );
  NOR2_X1 U9567 ( .A1(n8171), .A2(n8012), .ZN(n7949) );
  XNOR2_X1 U9568 ( .A(n7951), .B(n7949), .ZN(n8081) );
  AND2_X1 U9569 ( .A1(n8081), .A2(n7947), .ZN(n7948) );
  XNOR2_X1 U9570 ( .A(n8721), .B(n7998), .ZN(n8126) );
  OR2_X1 U9571 ( .A1(n8248), .A2(n8012), .ZN(n8124) );
  XNOR2_X1 U9572 ( .A(n8728), .B(n7124), .ZN(n7955) );
  NOR2_X1 U9573 ( .A1(n8604), .A2(n8012), .ZN(n8231) );
  INV_X1 U9574 ( .A(n7949), .ZN(n7950) );
  NAND2_X1 U9575 ( .A1(n7951), .A2(n7950), .ZN(n8121) );
  OAI21_X1 U9576 ( .B1(n7955), .B2(n8231), .A(n8121), .ZN(n7952) );
  AOI21_X1 U9577 ( .B1(n8126), .B2(n8124), .A(n7952), .ZN(n7953) );
  INV_X1 U9578 ( .A(n8126), .ZN(n7958) );
  INV_X1 U9579 ( .A(n7955), .ZN(n8122) );
  INV_X1 U9580 ( .A(n8231), .ZN(n7954) );
  OAI21_X1 U9581 ( .B1(n8122), .B2(n7954), .A(n8124), .ZN(n7957) );
  NOR2_X1 U9582 ( .A1(n8124), .A2(n7954), .ZN(n7956) );
  AOI22_X1 U9583 ( .A1(n7958), .A2(n7957), .B1(n7956), .B2(n7955), .ZN(n7959)
         );
  NAND2_X1 U9584 ( .A1(n7960), .A2(n7959), .ZN(n8138) );
  XNOR2_X1 U9585 ( .A(n8717), .B(n7124), .ZN(n7961) );
  NOR2_X1 U9586 ( .A1(n8606), .A2(n8012), .ZN(n7962) );
  NAND2_X1 U9587 ( .A1(n7961), .A2(n7962), .ZN(n7965) );
  INV_X1 U9588 ( .A(n7961), .ZN(n8199) );
  INV_X1 U9589 ( .A(n7962), .ZN(n7963) );
  NAND2_X1 U9590 ( .A1(n8199), .A2(n7963), .ZN(n7964) );
  AND2_X1 U9591 ( .A1(n7965), .A2(n7964), .ZN(n8139) );
  XNOR2_X1 U9592 ( .A(n8711), .B(n7124), .ZN(n7966) );
  AND2_X1 U9593 ( .A1(n8568), .A2(n7991), .ZN(n7967) );
  NAND2_X1 U9594 ( .A1(n7966), .A2(n7967), .ZN(n7970) );
  INV_X1 U9595 ( .A(n7966), .ZN(n8092) );
  INV_X1 U9596 ( .A(n7967), .ZN(n7968) );
  NAND2_X1 U9597 ( .A1(n8092), .A2(n7968), .ZN(n7969) );
  XNOR2_X1 U9598 ( .A(n8707), .B(n7998), .ZN(n7974) );
  NOR2_X1 U9599 ( .A1(n8203), .A2(n8012), .ZN(n7972) );
  XNOR2_X1 U9600 ( .A(n7974), .B(n7972), .ZN(n8093) );
  AND2_X1 U9601 ( .A1(n8093), .A2(n7970), .ZN(n7971) );
  INV_X1 U9602 ( .A(n7972), .ZN(n7973) );
  NAND2_X1 U9603 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  XNOR2_X1 U9604 ( .A(n8701), .B(n7124), .ZN(n7976) );
  NOR2_X1 U9605 ( .A1(n8536), .A2(n8012), .ZN(n7977) );
  NAND2_X1 U9606 ( .A1(n7976), .A2(n7977), .ZN(n8105) );
  INV_X1 U9607 ( .A(n7976), .ZN(n8104) );
  INV_X1 U9608 ( .A(n7977), .ZN(n7978) );
  NAND2_X1 U9609 ( .A1(n8104), .A2(n7978), .ZN(n7979) );
  NAND2_X1 U9610 ( .A1(n8105), .A2(n7979), .ZN(n8163) );
  XNOR2_X1 U9611 ( .A(n8691), .B(n7124), .ZN(n8181) );
  OR2_X1 U9612 ( .A1(n8537), .A2(n8012), .ZN(n8183) );
  INV_X1 U9613 ( .A(n8183), .ZN(n7985) );
  NAND2_X1 U9614 ( .A1(n8181), .A2(n7985), .ZN(n7980) );
  XNOR2_X1 U9615 ( .A(n8698), .B(n7124), .ZN(n7984) );
  AND2_X1 U9616 ( .A1(n8543), .A2(n7991), .ZN(n7982) );
  NAND2_X1 U9617 ( .A1(n7984), .A2(n7982), .ZN(n8179) );
  NAND2_X1 U9618 ( .A1(n7980), .A2(n8179), .ZN(n7986) );
  INV_X1 U9619 ( .A(n8105), .ZN(n7981) );
  INV_X1 U9620 ( .A(n7982), .ZN(n7983) );
  XNOR2_X1 U9621 ( .A(n7984), .B(n7983), .ZN(n8106) );
  OAI22_X1 U9622 ( .A1(n7986), .A2(n8106), .B1(n7985), .B2(n8181), .ZN(n7987)
         );
  XNOR2_X1 U9623 ( .A(n8688), .B(n7124), .ZN(n7992) );
  XNOR2_X1 U9624 ( .A(n8681), .B(n7124), .ZN(n7994) );
  AND2_X1 U9625 ( .A1(n8519), .A2(n7991), .ZN(n8083) );
  INV_X1 U9626 ( .A(n7989), .ZN(n7990) );
  AND2_X1 U9627 ( .A1(n8246), .A2(n7991), .ZN(n7995) );
  INV_X1 U9628 ( .A(n7994), .ZN(n8148) );
  INV_X1 U9629 ( .A(n7995), .ZN(n8151) );
  XNOR2_X1 U9630 ( .A(n8678), .B(n7998), .ZN(n8210) );
  OR2_X1 U9631 ( .A1(n8218), .A2(n8012), .ZN(n7999) );
  NOR2_X1 U9632 ( .A1(n8210), .A2(n7999), .ZN(n8000) );
  AOI21_X1 U9633 ( .B1(n8210), .B2(n7999), .A(n8000), .ZN(n8115) );
  XNOR2_X1 U9634 ( .A(n8673), .B(n7124), .ZN(n8001) );
  NOR2_X1 U9635 ( .A1(n8437), .A2(n8012), .ZN(n8002) );
  NAND2_X1 U9636 ( .A1(n8001), .A2(n8002), .ZN(n8005) );
  INV_X1 U9637 ( .A(n8001), .ZN(n8061) );
  INV_X1 U9638 ( .A(n8002), .ZN(n8003) );
  NAND2_X1 U9639 ( .A1(n8061), .A2(n8003), .ZN(n8004) );
  NAND2_X1 U9640 ( .A1(n8005), .A2(n8004), .ZN(n8211) );
  XNOR2_X1 U9641 ( .A(n8666), .B(n7124), .ZN(n8006) );
  NOR2_X1 U9642 ( .A1(n8217), .A2(n8012), .ZN(n8007) );
  NAND2_X1 U9643 ( .A1(n8006), .A2(n8007), .ZN(n8011) );
  INV_X1 U9644 ( .A(n8006), .ZN(n8009) );
  INV_X1 U9645 ( .A(n8007), .ZN(n8008) );
  NAND2_X1 U9646 ( .A1(n8009), .A2(n8008), .ZN(n8010) );
  NAND2_X1 U9647 ( .A1(n8062), .A2(n8011), .ZN(n8024) );
  NOR2_X1 U9648 ( .A1(n8438), .A2(n8012), .ZN(n8013) );
  XNOR2_X1 U9649 ( .A(n8013), .B(n7124), .ZN(n8015) );
  INV_X1 U9650 ( .A(n8015), .ZN(n8016) );
  NOR3_X1 U9651 ( .A1(n8406), .A2(n8236), .A3(n8016), .ZN(n8014) );
  AOI21_X1 U9652 ( .B1(n8406), .B2(n8016), .A(n8014), .ZN(n8023) );
  OAI21_X1 U9653 ( .B1(n8406), .B2(n8226), .A(n8230), .ZN(n8022) );
  NOR3_X1 U9654 ( .A1(n8406), .A2(n8015), .A3(n8236), .ZN(n8019) );
  NOR2_X1 U9655 ( .A1(n8017), .A2(n8016), .ZN(n8018) );
  NAND2_X1 U9656 ( .A1(n8024), .A2(n8020), .ZN(n8021) );
  OAI211_X1 U9657 ( .C1(n8024), .C2(n8023), .A(n8022), .B(n8021), .ZN(n8028)
         );
  INV_X1 U9658 ( .A(n8025), .ZN(n8026) );
  AOI22_X1 U9659 ( .A1(n8026), .A2(n8238), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8027) );
  OAI211_X1 U9660 ( .C1(n8029), .C2(n8221), .A(n8028), .B(n8027), .ZN(P2_U3222) );
  NAND2_X1 U9661 ( .A1(n9066), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8030) );
  INV_X1 U9662 ( .A(n9488), .ZN(n9463) );
  OR2_X2 U9663 ( .A1(n9736), .A2(n8903), .ZN(n9166) );
  AND2_X2 U9664 ( .A1(n9166), .A2(n9226), .ZN(n9459) );
  NAND2_X1 U9665 ( .A1(n8034), .A2(n6091), .ZN(n8036) );
  NAND2_X1 U9666 ( .A1(n9066), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U9667 ( .A1(n9059), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8041) );
  NAND2_X1 U9668 ( .A1(n9057), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8040) );
  NAND2_X1 U9669 ( .A1(n4448), .A2(n8054), .ZN(n8039) );
  NAND2_X1 U9670 ( .A1(n8046), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U9671 ( .A1(n8044), .A2(P1_B_REG_SCAN_IN), .ZN(n8045) );
  NAND2_X1 U9672 ( .A1(n9703), .A2(n8045), .ZN(n9445) );
  NAND2_X1 U9673 ( .A1(n9057), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U9674 ( .A1(n9058), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U9675 ( .A1(n9059), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8047) );
  AND3_X1 U9676 ( .A1(n8049), .A2(n8048), .A3(n8047), .ZN(n9241) );
  NOR2_X1 U9677 ( .A1(n9445), .A2(n9241), .ZN(n8050) );
  NOR2_X1 U9678 ( .A1(n9730), .A2(n9645), .ZN(n8057) );
  AOI22_X1 U9679 ( .A1(n9712), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8054), .B2(
        n9710), .ZN(n8055) );
  OAI21_X1 U9680 ( .B1(n9729), .B2(n9714), .A(n8055), .ZN(n8056) );
  AOI211_X1 U9681 ( .C1(n9728), .C2(n9670), .A(n8057), .B(n8056), .ZN(n8058)
         );
  OAI21_X1 U9682 ( .B1(n9734), .B2(n9716), .A(n8058), .ZN(P1_U3355) );
  INV_X1 U9683 ( .A(n8059), .ZN(n8060) );
  NOR3_X1 U9684 ( .A1(n8061), .A2(n8437), .A3(n8209), .ZN(n8063) );
  OAI21_X1 U9685 ( .B1(n8064), .B2(n8063), .A(n8062), .ZN(n8069) );
  NOR2_X1 U9686 ( .A1(n8065), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8067) );
  OAI22_X1 U9687 ( .A1(n8438), .A2(n8204), .B1(n8437), .B2(n8205), .ZN(n8066)
         );
  AOI211_X1 U9688 ( .C1(n8238), .C2(n8431), .A(n8067), .B(n8066), .ZN(n8068)
         );
  OAI211_X1 U9689 ( .C1(n8433), .C2(n8226), .A(n8069), .B(n8068), .ZN(P2_U3216) );
  NOR3_X1 U9690 ( .A1(n8209), .A2(n8071), .A3(n8070), .ZN(n8072) );
  AOI21_X1 U9691 ( .B1(n4364), .B2(n8184), .A(n8072), .ZN(n8082) );
  NAND2_X1 U9692 ( .A1(n8238), .A2(n8073), .ZN(n8075) );
  OAI211_X1 U9693 ( .C1(n8221), .C2(n8076), .A(n8075), .B(n8074), .ZN(n8079)
         );
  NOR2_X1 U9694 ( .A1(n8077), .A2(n8230), .ZN(n8078) );
  AOI211_X1 U9695 ( .C1(n8733), .C2(n8236), .A(n8079), .B(n8078), .ZN(n8080)
         );
  OAI21_X1 U9696 ( .B1(n8082), .B2(n8081), .A(n8080), .ZN(P2_U3217) );
  AOI22_X1 U9697 ( .A1(n8084), .A2(n8184), .B1(n8185), .B2(n8519), .ZN(n8089)
         );
  INV_X1 U9698 ( .A(n8238), .ZN(n8216) );
  AOI22_X1 U9699 ( .A1(n8187), .A2(n8247), .B1(n8186), .B2(n8246), .ZN(n8086)
         );
  NAND2_X1 U9700 ( .A1(P2_U3152), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8085) );
  OAI211_X1 U9701 ( .C1(n8216), .C2(n8498), .A(n8086), .B(n8085), .ZN(n8087)
         );
  AOI21_X1 U9702 ( .B1(n8688), .B2(n8236), .A(n8087), .ZN(n8088) );
  OAI21_X1 U9703 ( .B1(n8089), .B2(n8147), .A(n8088), .ZN(P2_U3218) );
  OAI21_X1 U9704 ( .B1(n8093), .B2(n8090), .A(n8091), .ZN(n8101) );
  NOR3_X1 U9705 ( .A1(n8093), .A2(n8092), .A3(n8209), .ZN(n8094) );
  OAI21_X1 U9706 ( .B1(n8094), .B2(n8187), .A(n8568), .ZN(n8099) );
  INV_X1 U9707 ( .A(n8536), .ZN(n8569) );
  OAI22_X1 U9708 ( .A1(n8216), .A2(n8096), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8095), .ZN(n8097) );
  AOI21_X1 U9709 ( .B1(n8186), .B2(n8569), .A(n8097), .ZN(n8098) );
  OAI211_X1 U9710 ( .C1(n8565), .C2(n8226), .A(n8099), .B(n8098), .ZN(n8100)
         );
  AOI21_X1 U9711 ( .B1(n8101), .B2(n8184), .A(n8100), .ZN(n8102) );
  INV_X1 U9712 ( .A(n8102), .ZN(P2_U3221) );
  INV_X1 U9713 ( .A(n8106), .ZN(n8103) );
  AOI21_X1 U9714 ( .B1(n8160), .B2(n8103), .A(n8230), .ZN(n8109) );
  NOR3_X1 U9715 ( .A1(n8104), .A2(n8536), .A3(n8209), .ZN(n8108) );
  NAND2_X1 U9716 ( .A1(n8160), .A2(n8105), .ZN(n8107) );
  NAND2_X1 U9717 ( .A1(n8107), .A2(n8106), .ZN(n8180) );
  OAI21_X1 U9718 ( .B1(n8109), .B2(n8108), .A(n8180), .ZN(n8114) );
  INV_X1 U9719 ( .A(n8528), .ZN(n8110) );
  AOI22_X1 U9720 ( .A1(n8238), .A2(n8110), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8113) );
  AOI22_X1 U9721 ( .A1(n8187), .A2(n8569), .B1(n8186), .B2(n8247), .ZN(n8112)
         );
  NAND2_X1 U9722 ( .A1(n8698), .A2(n8236), .ZN(n8111) );
  NAND4_X1 U9723 ( .A1(n8114), .A2(n8113), .A3(n8112), .A4(n8111), .ZN(
        P2_U3225) );
  OAI211_X1 U9724 ( .C1(n8116), .C2(n8115), .A(n8212), .B(n8184), .ZN(n8120)
         );
  INV_X1 U9725 ( .A(n8437), .ZN(n8245) );
  AOI22_X1 U9726 ( .A1(n8245), .A2(n8582), .B1(n8580), .B2(n8246), .ZN(n8471)
         );
  AOI22_X1 U9727 ( .A1(n8475), .A2(n8238), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8117) );
  OAI21_X1 U9728 ( .B1(n8471), .B2(n8221), .A(n8117), .ZN(n8118) );
  AOI21_X1 U9729 ( .B1(n8678), .B2(n8236), .A(n8118), .ZN(n8119) );
  NAND2_X1 U9730 ( .A1(n8120), .A2(n8119), .ZN(P2_U3227) );
  NAND2_X1 U9731 ( .A1(n8077), .A2(n8121), .ZN(n8123) );
  NOR2_X1 U9732 ( .A1(n8123), .A2(n8122), .ZN(n8227) );
  NOR2_X1 U9733 ( .A1(n8209), .A2(n8604), .ZN(n8232) );
  AOI21_X1 U9734 ( .B1(n8227), .B2(n8184), .A(n8232), .ZN(n8137) );
  NAND2_X1 U9735 ( .A1(n8123), .A2(n8122), .ZN(n8228) );
  INV_X1 U9736 ( .A(n8124), .ZN(n8125) );
  XNOR2_X1 U9737 ( .A(n8126), .B(n8125), .ZN(n8128) );
  INV_X1 U9738 ( .A(n8128), .ZN(n8127) );
  NAND2_X1 U9739 ( .A1(n8228), .A2(n8127), .ZN(n8136) );
  OAI21_X1 U9740 ( .B1(n8227), .B2(n8231), .A(n8228), .ZN(n8129) );
  NAND3_X1 U9741 ( .A1(n8129), .A2(n8184), .A3(n8128), .ZN(n8135) );
  NAND2_X1 U9742 ( .A1(n8238), .A2(n8618), .ZN(n8131) );
  NAND2_X1 U9743 ( .A1(n8131), .A2(n8130), .ZN(n8133) );
  OAI22_X1 U9744 ( .A1(n8604), .A2(n8205), .B1(n8204), .B2(n8606), .ZN(n8132)
         );
  AOI211_X1 U9745 ( .C1(n8721), .C2(n8236), .A(n8133), .B(n8132), .ZN(n8134)
         );
  OAI211_X1 U9746 ( .C1(n8137), .C2(n8136), .A(n8135), .B(n8134), .ZN(P2_U3228) );
  OAI211_X1 U9747 ( .C1(n8139), .C2(n8138), .A(n8198), .B(n8184), .ZN(n8146)
         );
  NAND2_X1 U9748 ( .A1(n8568), .A2(n8582), .ZN(n8141) );
  OR2_X1 U9749 ( .A1(n8248), .A2(n8603), .ZN(n8140) );
  NAND2_X1 U9750 ( .A1(n8141), .A2(n8140), .ZN(n8589) );
  AOI22_X1 U9751 ( .A1(n8235), .A2(n8589), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8145) );
  NAND2_X1 U9752 ( .A1(n8717), .A2(n8236), .ZN(n8144) );
  INV_X1 U9753 ( .A(n8142), .ZN(n8592) );
  NAND2_X1 U9754 ( .A1(n8238), .A2(n8592), .ZN(n8143) );
  NAND4_X1 U9755 ( .A1(n8146), .A2(n8145), .A3(n8144), .A4(n8143), .ZN(
        P2_U3230) );
  NOR2_X1 U9756 ( .A1(n8147), .A2(n4307), .ZN(n8149) );
  XNOR2_X1 U9757 ( .A(n8149), .B(n8148), .ZN(n8152) );
  OAI22_X1 U9758 ( .A1(n8152), .A2(n8230), .B1(n8505), .B2(n8209), .ZN(n8150)
         );
  OAI21_X1 U9759 ( .B1(n8152), .B2(n8151), .A(n8150), .ZN(n8159) );
  OR2_X1 U9760 ( .A1(n8218), .A2(n8605), .ZN(n8154) );
  NAND2_X1 U9761 ( .A1(n8519), .A2(n8580), .ZN(n8153) );
  NAND2_X1 U9762 ( .A1(n8154), .A2(n8153), .ZN(n8488) );
  INV_X1 U9763 ( .A(n8488), .ZN(n8156) );
  OAI22_X1 U9764 ( .A1(n8156), .A2(n8221), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8155), .ZN(n8157) );
  AOI21_X1 U9765 ( .B1(n8484), .B2(n8238), .A(n8157), .ZN(n8158) );
  OAI211_X1 U9766 ( .C1(n8486), .C2(n8226), .A(n8159), .B(n8158), .ZN(P2_U3231) );
  INV_X1 U9767 ( .A(n8160), .ZN(n8161) );
  AOI211_X1 U9768 ( .C1(n8163), .C2(n8162), .A(n8230), .B(n8161), .ZN(n8167)
         );
  AOI22_X1 U9769 ( .A1(n8238), .A2(n8550), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8165) );
  INV_X1 U9770 ( .A(n8203), .ZN(n8583) );
  AOI22_X1 U9771 ( .A1(n8186), .A2(n8543), .B1(n8187), .B2(n8583), .ZN(n8164)
         );
  OAI211_X1 U9772 ( .C1(n8553), .C2(n8226), .A(n8165), .B(n8164), .ZN(n8166)
         );
  OR2_X1 U9773 ( .A1(n8167), .A2(n8166), .ZN(P2_U3235) );
  AOI211_X1 U9774 ( .C1(n8169), .C2(n8168), .A(n8230), .B(n4364), .ZN(n8170)
         );
  INV_X1 U9775 ( .A(n8170), .ZN(n8177) );
  OAI22_X1 U9776 ( .A1(n8172), .A2(n8205), .B1(n8204), .B2(n8171), .ZN(n8173)
         );
  AOI211_X1 U9777 ( .C1(n8238), .C2(n8175), .A(n8174), .B(n8173), .ZN(n8176)
         );
  OAI211_X1 U9778 ( .C1(n8178), .C2(n8226), .A(n8177), .B(n8176), .ZN(P2_U3236) );
  NAND2_X1 U9779 ( .A1(n8180), .A2(n8179), .ZN(n8182) );
  XNOR2_X1 U9780 ( .A(n8182), .B(n8181), .ZN(n8195) );
  NAND2_X1 U9781 ( .A1(n8184), .A2(n8183), .ZN(n8194) );
  NAND3_X1 U9782 ( .A1(n8195), .A2(n8185), .A3(n8247), .ZN(n8193) );
  AOI22_X1 U9783 ( .A1(n8187), .A2(n8543), .B1(n8186), .B2(n8519), .ZN(n8189)
         );
  NAND2_X1 U9784 ( .A1(n8238), .A2(n8510), .ZN(n8188) );
  OAI211_X1 U9785 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n8190), .A(n8189), .B(n8188), .ZN(n8191) );
  AOI21_X1 U9786 ( .B1(n4433), .B2(n8236), .A(n8191), .ZN(n8192) );
  OAI211_X1 U9787 ( .C1(n8195), .C2(n8194), .A(n8193), .B(n8192), .ZN(P2_U3237) );
  INV_X1 U9788 ( .A(n8196), .ZN(n8197) );
  AOI21_X1 U9789 ( .B1(n8198), .B2(n8197), .A(n8230), .ZN(n8201) );
  NOR3_X1 U9790 ( .A1(n8199), .A2(n8606), .A3(n8209), .ZN(n8200) );
  OAI21_X1 U9791 ( .B1(n8201), .B2(n8200), .A(n8090), .ZN(n8208) );
  INV_X1 U9792 ( .A(n8202), .ZN(n8576) );
  AND2_X1 U9793 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8365) );
  OAI22_X1 U9794 ( .A1(n8606), .A2(n8205), .B1(n8204), .B2(n8203), .ZN(n8206)
         );
  AOI211_X1 U9795 ( .C1(n8238), .C2(n8576), .A(n8365), .B(n8206), .ZN(n8207)
         );
  OAI211_X1 U9796 ( .C1(n8578), .C2(n8226), .A(n8208), .B(n8207), .ZN(P2_U3240) );
  NOR3_X1 U9797 ( .A1(n8210), .A2(n8218), .A3(n8209), .ZN(n8215) );
  AOI21_X1 U9798 ( .B1(n8212), .B2(n8211), .A(n8230), .ZN(n8214) );
  OAI21_X1 U9799 ( .B1(n8215), .B2(n8214), .A(n8213), .ZN(n8225) );
  NOR2_X1 U9800 ( .A1(n8451), .A2(n8216), .ZN(n8223) );
  OR2_X1 U9801 ( .A1(n8217), .A2(n8605), .ZN(n8220) );
  OR2_X1 U9802 ( .A1(n8218), .A2(n8603), .ZN(n8219) );
  NOR2_X1 U9803 ( .A1(n8457), .A2(n8221), .ZN(n8222) );
  AOI211_X1 U9804 ( .C1(P2_REG3_REG_26__SCAN_IN), .C2(P2_U3152), .A(n8223), 
        .B(n8222), .ZN(n8224) );
  OAI211_X1 U9805 ( .C1(n8449), .C2(n8226), .A(n8225), .B(n8224), .ZN(P2_U3242) );
  INV_X1 U9806 ( .A(n8227), .ZN(n8229) );
  NAND2_X1 U9807 ( .A1(n8229), .A2(n8228), .ZN(n8233) );
  NOR3_X1 U9808 ( .A1(n8233), .A2(n8231), .A3(n8230), .ZN(n8244) );
  NAND2_X1 U9809 ( .A1(n8233), .A2(n8232), .ZN(n8242) );
  AOI22_X1 U9810 ( .A1(n8235), .A2(n8234), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n8241) );
  NAND2_X1 U9811 ( .A1(n8236), .A2(n8728), .ZN(n8240) );
  NAND2_X1 U9812 ( .A1(n8238), .A2(n8237), .ZN(n8239) );
  NAND4_X1 U9813 ( .A1(n8242), .A2(n8241), .A3(n8240), .A4(n8239), .ZN(n8243)
         );
  OR2_X1 U9814 ( .A1(n8244), .A2(n8243), .ZN(P2_U3243) );
  MUX2_X1 U9815 ( .A(n8412), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8257), .Z(
        P2_U3582) );
  INV_X1 U9816 ( .A(n8438), .ZN(n8414) );
  INV_X2 U9817 ( .A(P2_U3966), .ZN(n8257) );
  MUX2_X1 U9818 ( .A(n8414), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8257), .Z(
        P2_U3580) );
  MUX2_X1 U9819 ( .A(n8245), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8257), .Z(
        P2_U3578) );
  MUX2_X1 U9820 ( .A(n8246), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8257), .Z(
        P2_U3576) );
  MUX2_X1 U9821 ( .A(n8519), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8257), .Z(
        P2_U3575) );
  MUX2_X1 U9822 ( .A(n8247), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8257), .Z(
        P2_U3574) );
  MUX2_X1 U9823 ( .A(n8543), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8257), .Z(
        P2_U3573) );
  MUX2_X1 U9824 ( .A(n8569), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8257), .Z(
        P2_U3572) );
  MUX2_X1 U9825 ( .A(n8583), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8257), .Z(
        P2_U3571) );
  MUX2_X1 U9826 ( .A(n8568), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8257), .Z(
        P2_U3570) );
  MUX2_X1 U9827 ( .A(n8581), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8257), .Z(
        P2_U3569) );
  INV_X1 U9828 ( .A(n8248), .ZN(n8249) );
  MUX2_X1 U9829 ( .A(n8249), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8257), .Z(
        P2_U3568) );
  MUX2_X1 U9830 ( .A(n5915), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8257), .Z(
        P2_U3567) );
  MUX2_X1 U9831 ( .A(n8250), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8257), .Z(
        P2_U3566) );
  MUX2_X1 U9832 ( .A(n8251), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8257), .Z(
        P2_U3565) );
  MUX2_X1 U9833 ( .A(n8252), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8257), .Z(
        P2_U3564) );
  MUX2_X1 U9834 ( .A(n8253), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8257), .Z(
        P2_U3563) );
  MUX2_X1 U9835 ( .A(n4626), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8257), .Z(
        P2_U3562) );
  MUX2_X1 U9836 ( .A(n8254), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8257), .Z(
        P2_U3561) );
  MUX2_X1 U9837 ( .A(n8255), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8257), .Z(
        P2_U3560) );
  MUX2_X1 U9838 ( .A(n8256), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8257), .Z(
        P2_U3559) );
  MUX2_X1 U9839 ( .A(n8258), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8257), .Z(
        P2_U3558) );
  MUX2_X1 U9840 ( .A(n8259), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8257), .Z(
        P2_U3557) );
  MUX2_X1 U9841 ( .A(n8260), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8257), .Z(
        P2_U3556) );
  MUX2_X1 U9842 ( .A(n8261), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8257), .Z(
        P2_U3555) );
  MUX2_X1 U9843 ( .A(n8262), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8257), .Z(
        P2_U3554) );
  MUX2_X1 U9844 ( .A(n5891), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8257), .Z(
        P2_U3553) );
  NAND2_X1 U9845 ( .A1(n8342), .A2(n8263), .ZN(n8273) );
  OAI211_X1 U9846 ( .C1(n8266), .C2(n8265), .A(n8388), .B(n8264), .ZN(n8272)
         );
  AOI22_X1 U9847 ( .A1(n8366), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8271) );
  OAI211_X1 U9848 ( .C1(n8269), .C2(n8268), .A(n8386), .B(n8267), .ZN(n8270)
         );
  NAND4_X1 U9849 ( .A1(n8273), .A2(n8272), .A3(n8271), .A4(n8270), .ZN(
        P2_U3246) );
  NAND2_X1 U9850 ( .A1(n8342), .A2(n8274), .ZN(n8283) );
  OAI211_X1 U9851 ( .C1(n8276), .C2(n8275), .A(n8388), .B(n8288), .ZN(n8282)
         );
  AOI22_X1 U9852 ( .A1(n8366), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n8281) );
  OAI211_X1 U9853 ( .C1(n8279), .C2(n8278), .A(n8386), .B(n8277), .ZN(n8280)
         );
  NAND4_X1 U9854 ( .A1(n8283), .A2(n8282), .A3(n8281), .A4(n8280), .ZN(
        P2_U3247) );
  NAND2_X1 U9855 ( .A1(n8342), .A2(n8284), .ZN(n8298) );
  NOR2_X1 U9856 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8640), .ZN(n8285) );
  AOI21_X1 U9857 ( .B1(n8366), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8285), .ZN(
        n8297) );
  MUX2_X1 U9858 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6665), .S(n8286), .Z(n8289)
         );
  NAND3_X1 U9859 ( .A1(n8289), .A2(n8288), .A3(n8287), .ZN(n8290) );
  NAND3_X1 U9860 ( .A1(n8388), .A2(n8291), .A3(n8290), .ZN(n8296) );
  OAI211_X1 U9861 ( .C1(n8294), .C2(n8293), .A(n8386), .B(n8292), .ZN(n8295)
         );
  NAND4_X1 U9862 ( .A1(n8298), .A2(n8297), .A3(n8296), .A4(n8295), .ZN(
        P2_U3248) );
  NAND2_X1 U9863 ( .A1(n8342), .A2(n8299), .ZN(n8314) );
  INV_X1 U9864 ( .A(n8300), .ZN(n8301) );
  AOI21_X1 U9865 ( .B1(n8366), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8301), .ZN(
        n8313) );
  MUX2_X1 U9866 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7441), .S(n8302), .Z(n8305)
         );
  NAND3_X1 U9867 ( .A1(n8305), .A2(n8304), .A3(n8303), .ZN(n8306) );
  NAND3_X1 U9868 ( .A1(n8388), .A2(n8307), .A3(n8306), .ZN(n8312) );
  OAI211_X1 U9869 ( .C1(n8310), .C2(n8309), .A(n8386), .B(n8308), .ZN(n8311)
         );
  NAND4_X1 U9870 ( .A1(n8314), .A2(n8313), .A3(n8312), .A4(n8311), .ZN(
        P2_U3251) );
  NAND2_X1 U9871 ( .A1(n8342), .A2(n8317), .ZN(n8328) );
  INV_X1 U9872 ( .A(n8315), .ZN(n8316) );
  AOI21_X1 U9873 ( .B1(n8366), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8316), .ZN(
        n8327) );
  MUX2_X1 U9874 ( .A(n6876), .B(P2_REG2_REG_8__SCAN_IN), .S(n8317), .Z(n8318)
         );
  NAND3_X1 U9875 ( .A1(n8320), .A2(n8319), .A3(n8318), .ZN(n8321) );
  NAND3_X1 U9876 ( .A1(n8388), .A2(n8333), .A3(n8321), .ZN(n8326) );
  OAI211_X1 U9877 ( .C1(n8324), .C2(n8323), .A(n8386), .B(n8322), .ZN(n8325)
         );
  NAND4_X1 U9878 ( .A1(n8328), .A2(n8327), .A3(n8326), .A4(n8325), .ZN(
        P2_U3253) );
  NAND2_X1 U9879 ( .A1(n8342), .A2(n8330), .ZN(n8341) );
  AOI21_X1 U9880 ( .B1(n8366), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8329), .ZN(
        n8340) );
  MUX2_X1 U9881 ( .A(n6879), .B(P2_REG2_REG_9__SCAN_IN), .S(n8330), .Z(n8331)
         );
  NAND3_X1 U9882 ( .A1(n8333), .A2(n8332), .A3(n8331), .ZN(n8334) );
  NAND3_X1 U9883 ( .A1(n8388), .A2(n8347), .A3(n8334), .ZN(n8339) );
  OAI211_X1 U9884 ( .C1(n8337), .C2(n8336), .A(n8386), .B(n8335), .ZN(n8338)
         );
  NAND4_X1 U9885 ( .A1(n8341), .A2(n8340), .A3(n8339), .A4(n8338), .ZN(
        P2_U3254) );
  NAND2_X1 U9886 ( .A1(n8342), .A2(n8344), .ZN(n8356) );
  AOI21_X1 U9887 ( .B1(n8366), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8343), .ZN(
        n8355) );
  MUX2_X1 U9888 ( .A(n7773), .B(P2_REG2_REG_10__SCAN_IN), .S(n8344), .Z(n8345)
         );
  NAND3_X1 U9889 ( .A1(n8347), .A2(n8346), .A3(n8345), .ZN(n8348) );
  NAND3_X1 U9890 ( .A1(n8388), .A2(n8349), .A3(n8348), .ZN(n8354) );
  OAI211_X1 U9891 ( .C1(n8352), .C2(n8351), .A(n8386), .B(n8350), .ZN(n8353)
         );
  NAND4_X1 U9892 ( .A1(n8356), .A2(n8355), .A3(n8354), .A4(n8353), .ZN(
        P2_U3255) );
  NAND2_X1 U9893 ( .A1(n8361), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8358) );
  XNOR2_X1 U9894 ( .A(n8379), .B(n8374), .ZN(n8359) );
  NOR2_X1 U9895 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8359), .ZN(n8376) );
  AOI21_X1 U9896 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8359), .A(n8376), .ZN(
        n8373) );
  AOI21_X1 U9897 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8361), .A(n8360), .ZN(
        n8364) );
  AOI22_X1 U9898 ( .A1(n8379), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8362), .B2(
        n8368), .ZN(n8363) );
  NAND2_X1 U9899 ( .A1(n8364), .A2(n8363), .ZN(n8378) );
  OAI21_X1 U9900 ( .B1(n8364), .B2(n8363), .A(n8378), .ZN(n8370) );
  AOI21_X1 U9901 ( .B1(n8366), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8365), .ZN(
        n8367) );
  OAI21_X1 U9902 ( .B1(n8368), .B2(n8382), .A(n8367), .ZN(n8369) );
  AOI21_X1 U9903 ( .B1(n8370), .B2(n8386), .A(n8369), .ZN(n8371) );
  OAI21_X1 U9904 ( .B1(n8373), .B2(n8372), .A(n8371), .ZN(P2_U3263) );
  NOR2_X1 U9905 ( .A1(n8379), .A2(n8374), .ZN(n8375) );
  NOR2_X1 U9906 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  XOR2_X1 U9907 ( .A(n8377), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8389) );
  INV_X1 U9908 ( .A(n8389), .ZN(n8385) );
  OAI21_X1 U9909 ( .B1(n8379), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8378), .ZN(
        n8381) );
  XOR2_X1 U9910 ( .A(n8381), .B(n8380), .Z(n8387) );
  OAI21_X1 U9911 ( .B1(n8387), .B2(n8383), .A(n8382), .ZN(n8384) );
  AOI21_X1 U9912 ( .B1(n8388), .B2(n8385), .A(n8384), .ZN(n8392) );
  AOI22_X1 U9913 ( .A1(n8389), .A2(n8388), .B1(n8387), .B2(n8386), .ZN(n8391)
         );
  NAND2_X1 U9914 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8393) );
  XNOR2_X1 U9915 ( .A(n8651), .B(n8655), .ZN(n8650) );
  NAND2_X1 U9916 ( .A1(n8650), .A2(n8643), .ZN(n8400) );
  NOR2_X1 U9917 ( .A1(n8800), .A2(n8396), .ZN(n8397) );
  NOR2_X1 U9918 ( .A1(n8605), .A2(n8397), .ZN(n8413) );
  NAND2_X1 U9919 ( .A1(n8398), .A2(n8413), .ZN(n8657) );
  NOR2_X1 U9920 ( .A1(n4273), .A2(n8657), .ZN(n8403) );
  AOI21_X1 U9921 ( .B1(n4273), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8403), .ZN(
        n8399) );
  OAI211_X1 U9922 ( .C1(n8651), .C2(n8620), .A(n8400), .B(n8399), .ZN(P2_U3265) );
  NAND2_X1 U9923 ( .A1(n8402), .A2(n8418), .ZN(n8656) );
  NAND3_X1 U9924 ( .A1(n8656), .A2(n8643), .A3(n8655), .ZN(n8405) );
  AOI21_X1 U9925 ( .B1(n4273), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8403), .ZN(
        n8404) );
  OAI211_X1 U9926 ( .C1(n8659), .C2(n8620), .A(n8405), .B(n8404), .ZN(P2_U3266) );
  NAND2_X1 U9927 ( .A1(n8406), .A2(n8438), .ZN(n8407) );
  XNOR2_X1 U9928 ( .A(n8409), .B(n8410), .ZN(n8660) );
  INV_X1 U9929 ( .A(n8660), .ZN(n8425) );
  AOI22_X1 U9930 ( .A1(n8414), .A2(n8580), .B1(n8413), .B2(n8412), .ZN(n8415)
         );
  INV_X1 U9931 ( .A(n8417), .ZN(n8661) );
  NOR2_X1 U9932 ( .A1(n8662), .A2(n8630), .ZN(n8423) );
  INV_X1 U9933 ( .A(n8419), .ZN(n8420) );
  AOI22_X1 U9934 ( .A1(n8420), .A2(n8641), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n4273), .ZN(n8421) );
  OAI21_X1 U9935 ( .B1(n8661), .B2(n8620), .A(n8421), .ZN(n8422) );
  AOI211_X1 U9936 ( .C1(n8664), .C2(n8645), .A(n8423), .B(n8422), .ZN(n8424)
         );
  OAI21_X1 U9937 ( .B1(n8425), .B2(n8597), .A(n8424), .ZN(P2_U3267) );
  OAI21_X1 U9938 ( .B1(n8427), .B2(n8435), .A(n8426), .ZN(n8428) );
  INV_X1 U9939 ( .A(n8428), .ZN(n8670) );
  INV_X1 U9940 ( .A(n8448), .ZN(n8430) );
  AOI21_X1 U9941 ( .B1(n8666), .B2(n8430), .A(n8429), .ZN(n8667) );
  AOI22_X1 U9942 ( .A1(n8431), .A2(n8641), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n4273), .ZN(n8432) );
  OAI21_X1 U9943 ( .B1(n8433), .B2(n8620), .A(n8432), .ZN(n8443) );
  INV_X1 U9944 ( .A(n8434), .ZN(n8436) );
  AOI21_X1 U9945 ( .B1(n8436), .B2(n8435), .A(n8535), .ZN(n8441) );
  OAI22_X1 U9946 ( .A1(n8438), .A2(n8605), .B1(n8437), .B2(n8603), .ZN(n8439)
         );
  AOI21_X1 U9947 ( .B1(n8441), .B2(n8440), .A(n8439), .ZN(n8669) );
  NOR2_X1 U9948 ( .A1(n8669), .A2(n4273), .ZN(n8442) );
  AOI211_X1 U9949 ( .C1(n8667), .C2(n8643), .A(n8443), .B(n8442), .ZN(n8444)
         );
  OAI21_X1 U9950 ( .B1(n8670), .B2(n8597), .A(n8444), .ZN(P2_U3269) );
  NAND2_X1 U9951 ( .A1(n8461), .A2(n8468), .ZN(n8462) );
  INV_X1 U9952 ( .A(n8445), .ZN(n8446) );
  NAND2_X1 U9953 ( .A1(n8462), .A2(n8446), .ZN(n8447) );
  AOI211_X1 U9954 ( .C1(n8673), .C2(n8473), .A(n10052), .B(n8448), .ZN(n8672)
         );
  NOR2_X1 U9955 ( .A1(n8449), .A2(n8620), .ZN(n8453) );
  OAI22_X1 U9956 ( .A1(n8451), .A2(n8527), .B1(n8450), .B2(n8645), .ZN(n8452)
         );
  AOI211_X1 U9957 ( .C1(n8672), .C2(n8600), .A(n8453), .B(n8452), .ZN(n8460)
         );
  OAI211_X1 U9958 ( .C1(n8456), .C2(n8455), .A(n8454), .B(n8614), .ZN(n8458)
         );
  NAND2_X1 U9959 ( .A1(n8458), .A2(n8457), .ZN(n8671) );
  NAND2_X1 U9960 ( .A1(n8671), .A2(n8645), .ZN(n8459) );
  OAI211_X1 U9961 ( .C1(n8675), .C2(n8597), .A(n8460), .B(n8459), .ZN(P2_U3270) );
  INV_X1 U9962 ( .A(n8461), .ZN(n8464) );
  INV_X1 U9963 ( .A(n8462), .ZN(n8463) );
  NAND3_X1 U9964 ( .A1(n8466), .A2(n8468), .A3(n8467), .ZN(n8469) );
  NAND3_X1 U9965 ( .A1(n8470), .A2(n8614), .A3(n8469), .ZN(n8472) );
  NAND2_X1 U9966 ( .A1(n8472), .A2(n8471), .ZN(n8676) );
  INV_X1 U9967 ( .A(n8473), .ZN(n8474) );
  AOI211_X1 U9968 ( .C1(n8678), .C2(n8482), .A(n10052), .B(n8474), .ZN(n8677)
         );
  NAND2_X1 U9969 ( .A1(n8677), .A2(n8600), .ZN(n8477) );
  AOI22_X1 U9970 ( .A1(n8475), .A2(n8641), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n4273), .ZN(n8476) );
  OAI211_X1 U9971 ( .C1(n8478), .C2(n8620), .A(n8477), .B(n8476), .ZN(n8479)
         );
  AOI21_X1 U9972 ( .B1(n8676), .B2(n8645), .A(n8479), .ZN(n8480) );
  OAI21_X1 U9973 ( .B1(n8680), .B2(n8597), .A(n8480), .ZN(P2_U3271) );
  AOI21_X1 U9974 ( .B1(n8487), .B2(n8481), .A(n5926), .ZN(n8685) );
  INV_X1 U9975 ( .A(n8495), .ZN(n8483) );
  AOI21_X1 U9976 ( .B1(n8681), .B2(n8483), .A(n4973), .ZN(n8682) );
  AOI22_X1 U9977 ( .A1(n8484), .A2(n8641), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n4273), .ZN(n8485) );
  OAI21_X1 U9978 ( .B1(n8486), .B2(n8620), .A(n8485), .ZN(n8491) );
  AOI21_X1 U9979 ( .B1(n4329), .B2(n5925), .A(n8535), .ZN(n8489) );
  AOI21_X1 U9980 ( .B1(n8489), .B2(n8466), .A(n8488), .ZN(n8684) );
  NOR2_X1 U9981 ( .A1(n8684), .A2(n4273), .ZN(n8490) );
  AOI211_X1 U9982 ( .C1(n8682), .C2(n8643), .A(n8491), .B(n8490), .ZN(n8492)
         );
  OAI21_X1 U9983 ( .B1(n8685), .B2(n8597), .A(n8492), .ZN(P2_U3272) );
  OAI21_X1 U9984 ( .B1(n4320), .B2(n8494), .A(n8493), .ZN(n8690) );
  INV_X1 U9985 ( .A(n8509), .ZN(n8496) );
  AOI211_X1 U9986 ( .C1(n8688), .C2(n8496), .A(n10052), .B(n8495), .ZN(n8687)
         );
  NOR2_X1 U9987 ( .A1(n8497), .A2(n8620), .ZN(n8501) );
  OAI22_X1 U9988 ( .A1(n8645), .A2(n8499), .B1(n8498), .B2(n8527), .ZN(n8500)
         );
  AOI211_X1 U9989 ( .C1(n8687), .C2(n8600), .A(n8501), .B(n8500), .ZN(n8507)
         );
  XNOR2_X1 U9990 ( .A(n8503), .B(n8502), .ZN(n8504) );
  OAI222_X1 U9991 ( .A1(n8605), .A2(n8505), .B1(n8603), .B2(n8537), .C1(n8504), 
        .C2(n8535), .ZN(n8686) );
  NAND2_X1 U9992 ( .A1(n8686), .A2(n8645), .ZN(n8506) );
  OAI211_X1 U9993 ( .C1(n8690), .C2(n8597), .A(n8507), .B(n8506), .ZN(P2_U3273) );
  XNOR2_X1 U9994 ( .A(n8508), .B(n8517), .ZN(n8695) );
  AOI21_X1 U9995 ( .B1(n4433), .B2(n8525), .A(n8509), .ZN(n8692) );
  INV_X1 U9996 ( .A(n4433), .ZN(n8512) );
  AOI22_X1 U9997 ( .A1(n4273), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8510), .B2(
        n8641), .ZN(n8511) );
  OAI21_X1 U9998 ( .B1(n8512), .B2(n8620), .A(n8511), .ZN(n8522) );
  NAND2_X1 U9999 ( .A1(n8513), .A2(n8567), .ZN(n8566) );
  NAND3_X1 U10000 ( .A1(n8566), .A2(n8541), .A3(n8540), .ZN(n8515) );
  NAND2_X1 U10001 ( .A1(n8515), .A2(n8514), .ZN(n8533) );
  NOR2_X1 U10002 ( .A1(n8532), .A2(n8516), .ZN(n8518) );
  XNOR2_X1 U10003 ( .A(n8518), .B(n8517), .ZN(n8520) );
  AOI211_X1 U10004 ( .C1(n8692), .C2(n8643), .A(n8522), .B(n8521), .ZN(n8523)
         );
  OAI21_X1 U10005 ( .B1(n8597), .B2(n8695), .A(n8523), .ZN(P2_U3274) );
  XNOR2_X1 U10006 ( .A(n8524), .B(n8534), .ZN(n8700) );
  AOI211_X1 U10007 ( .C1(n8698), .C2(n8549), .A(n10052), .B(n4429), .ZN(n8697)
         );
  INV_X1 U10008 ( .A(n8698), .ZN(n8526) );
  NOR2_X1 U10009 ( .A1(n8526), .A2(n8620), .ZN(n8531) );
  OAI22_X1 U10010 ( .A1(n8645), .A2(n8529), .B1(n8528), .B2(n8527), .ZN(n8530)
         );
  AOI211_X1 U10011 ( .C1(n8697), .C2(n8600), .A(n8531), .B(n8530), .ZN(n8539)
         );
  NAND2_X1 U10012 ( .A1(n8696), .A2(n8645), .ZN(n8538) );
  OAI211_X1 U10013 ( .C1(n8700), .C2(n8597), .A(n8539), .B(n8538), .ZN(
        P2_U3275) );
  NAND2_X1 U10014 ( .A1(n8566), .A2(n8540), .ZN(n8542) );
  XNOR2_X1 U10015 ( .A(n8542), .B(n8541), .ZN(n8544) );
  AOI222_X1 U10016 ( .A1(n8614), .A2(n8544), .B1(n8583), .B2(n8580), .C1(n8543), .C2(n8582), .ZN(n8704) );
  OAI21_X1 U10017 ( .B1(n8547), .B2(n8546), .A(n8545), .ZN(n8705) );
  INV_X1 U10018 ( .A(n8705), .ZN(n8556) );
  OR2_X1 U10019 ( .A1(n8561), .A2(n8553), .ZN(n8548) );
  AND2_X1 U10020 ( .A1(n8549), .A2(n8548), .ZN(n8702) );
  NAND2_X1 U10021 ( .A1(n8702), .A2(n8643), .ZN(n8552) );
  AOI22_X1 U10022 ( .A1(n4273), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8550), .B2(
        n8641), .ZN(n8551) );
  OAI211_X1 U10023 ( .C1(n8553), .C2(n8620), .A(n8552), .B(n8551), .ZN(n8554)
         );
  AOI21_X1 U10024 ( .B1(n8556), .B2(n8555), .A(n8554), .ZN(n8557) );
  OAI21_X1 U10025 ( .B1(n4273), .B2(n8704), .A(n8557), .ZN(P2_U3276) );
  OAI21_X1 U10026 ( .B1(n8560), .B2(n8559), .A(n8558), .ZN(n8710) );
  INV_X1 U10027 ( .A(n8575), .ZN(n8562) );
  AOI211_X1 U10028 ( .C1(n8707), .C2(n8562), .A(n10052), .B(n8561), .ZN(n8706)
         );
  AOI22_X1 U10029 ( .A1(n4273), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8563), .B2(
        n8641), .ZN(n8564) );
  OAI21_X1 U10030 ( .B1(n8565), .B2(n8620), .A(n8564), .ZN(n8572) );
  OAI21_X1 U10031 ( .B1(n8567), .B2(n8513), .A(n8566), .ZN(n8570) );
  AOI222_X1 U10032 ( .A1(n8614), .A2(n8570), .B1(n8569), .B2(n8582), .C1(n8568), .C2(n8580), .ZN(n8709) );
  NOR2_X1 U10033 ( .A1(n8709), .A2(n4273), .ZN(n8571) );
  AOI211_X1 U10034 ( .C1(n8706), .C2(n8600), .A(n8572), .B(n8571), .ZN(n8573)
         );
  OAI21_X1 U10035 ( .B1(n8597), .B2(n8710), .A(n8573), .ZN(P2_U3277) );
  XNOR2_X1 U10036 ( .A(n8574), .B(n4291), .ZN(n8715) );
  AOI21_X1 U10037 ( .B1(n8711), .B2(n5031), .A(n8575), .ZN(n8712) );
  AOI22_X1 U10038 ( .A1(n4273), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8576), .B2(
        n8641), .ZN(n8577) );
  OAI21_X1 U10039 ( .B1(n8578), .B2(n8620), .A(n8577), .ZN(n8586) );
  OAI21_X1 U10040 ( .B1(n4317), .B2(n4291), .A(n8579), .ZN(n8584) );
  AOI222_X1 U10041 ( .A1(n8614), .A2(n8584), .B1(n8583), .B2(n8582), .C1(n8581), .C2(n8580), .ZN(n8714) );
  NOR2_X1 U10042 ( .A1(n8714), .A2(n4273), .ZN(n8585) );
  AOI211_X1 U10043 ( .C1(n8712), .C2(n8643), .A(n8586), .B(n8585), .ZN(n8587)
         );
  OAI21_X1 U10044 ( .B1(n8715), .B2(n8597), .A(n8587), .ZN(P2_U3278) );
  XOR2_X1 U10045 ( .A(n4425), .B(n8595), .Z(n8590) );
  AOI21_X1 U10046 ( .B1(n8590), .B2(n8614), .A(n8589), .ZN(n8719) );
  AOI21_X1 U10047 ( .B1(n8616), .B2(n8717), .A(n10052), .ZN(n8591) );
  AND2_X1 U10048 ( .A1(n8591), .A2(n5031), .ZN(n8716) );
  NAND2_X1 U10049 ( .A1(n8717), .A2(n8637), .ZN(n8594) );
  AOI22_X1 U10050 ( .A1(n4273), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8592), .B2(
        n8641), .ZN(n8593) );
  NAND2_X1 U10051 ( .A1(n8594), .A2(n8593), .ZN(n8599) );
  AOI21_X1 U10052 ( .B1(n4843), .B2(n8596), .A(n4334), .ZN(n8720) );
  NOR2_X1 U10053 ( .A1(n8720), .A2(n8597), .ZN(n8598) );
  AOI211_X1 U10054 ( .C1(n8716), .C2(n8600), .A(n8599), .B(n8598), .ZN(n8601)
         );
  OAI21_X1 U10055 ( .B1(n4273), .B2(n8719), .A(n8601), .ZN(P2_U3279) );
  XNOR2_X1 U10056 ( .A(n8602), .B(n8608), .ZN(n8613) );
  OAI22_X1 U10057 ( .A1(n8606), .A2(n8605), .B1(n8604), .B2(n8603), .ZN(n8612)
         );
  OAI21_X1 U10058 ( .B1(n8609), .B2(n8608), .A(n8607), .ZN(n8725) );
  NOR2_X1 U10059 ( .A1(n8725), .A2(n8610), .ZN(n8611) );
  AOI211_X1 U10060 ( .C1(n8614), .C2(n8613), .A(n8612), .B(n8611), .ZN(n8724)
         );
  INV_X1 U10061 ( .A(n8615), .ZN(n8617) );
  AOI21_X1 U10062 ( .B1(n8721), .B2(n8617), .A(n4385), .ZN(n8722) );
  AOI22_X1 U10063 ( .A1(n4273), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8618), .B2(
        n8641), .ZN(n8619) );
  OAI21_X1 U10064 ( .B1(n8621), .B2(n8620), .A(n8619), .ZN(n8624) );
  NOR2_X1 U10065 ( .A1(n8725), .A2(n8622), .ZN(n8623) );
  AOI211_X1 U10066 ( .C1(n8722), .C2(n8643), .A(n8624), .B(n8623), .ZN(n8625)
         );
  OAI21_X1 U10067 ( .B1(n8724), .B2(n4273), .A(n8625), .ZN(P2_U3280) );
  AOI22_X1 U10068 ( .A1(n8637), .A2(n8627), .B1(n8641), .B2(n8626), .ZN(n8628)
         );
  OAI21_X1 U10069 ( .B1(n8630), .B2(n8629), .A(n8628), .ZN(n8633) );
  MUX2_X1 U10070 ( .A(n8631), .B(P2_REG2_REG_9__SCAN_IN), .S(n4273), .Z(n8632)
         );
  AOI211_X1 U10071 ( .C1(n8639), .C2(n8634), .A(n8633), .B(n8632), .ZN(n8635)
         );
  INV_X1 U10072 ( .A(n8635), .ZN(P2_U3287) );
  AOI22_X1 U10073 ( .A1(n8639), .A2(n8638), .B1(n8637), .B2(n8636), .ZN(n8649)
         );
  AOI22_X1 U10074 ( .A1(n4273), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n8641), .B2(
        n8640), .ZN(n8648) );
  NAND2_X1 U10075 ( .A1(n8643), .A2(n8642), .ZN(n8647) );
  NAND2_X1 U10076 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND4_X1 U10077 ( .A1(n8649), .A2(n8648), .A3(n8647), .A4(n8646), .ZN(
        P2_U3293) );
  INV_X1 U10078 ( .A(n8652), .ZN(n8653) );
  MUX2_X1 U10079 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8769), .S(n10084), .Z(
        P2_U3551) );
  NAND3_X1 U10080 ( .A1(n8656), .A2(n8763), .A3(n8655), .ZN(n8658) );
  OAI211_X1 U10081 ( .C1(n8659), .C2(n10070), .A(n8658), .B(n8657), .ZN(n8770)
         );
  MUX2_X1 U10082 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8770), .S(n10084), .Z(
        P2_U3550) );
  OAI22_X1 U10083 ( .A1(n8662), .A2(n10052), .B1(n8661), .B2(n10070), .ZN(
        n8663) );
  MUX2_X1 U10084 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8771), .S(n10084), .Z(
        P2_U3549) );
  MUX2_X1 U10085 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8665), .S(n10084), .Z(
        P2_U3548) );
  AOI22_X1 U10086 ( .A1(n8667), .A2(n8763), .B1(n8762), .B2(n8666), .ZN(n8668)
         );
  OAI211_X1 U10087 ( .C1(n8670), .C2(n8767), .A(n8669), .B(n8668), .ZN(n8772)
         );
  MUX2_X1 U10088 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8772), .S(n10084), .Z(
        P2_U3547) );
  OAI21_X1 U10089 ( .B1(n8675), .B2(n8767), .A(n8674), .ZN(n8773) );
  MUX2_X1 U10090 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8773), .S(n10084), .Z(
        P2_U3546) );
  AOI211_X1 U10091 ( .C1(n8762), .C2(n8678), .A(n8677), .B(n8676), .ZN(n8679)
         );
  OAI21_X1 U10092 ( .B1(n8680), .B2(n8767), .A(n8679), .ZN(n8774) );
  MUX2_X1 U10093 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8774), .S(n10084), .Z(
        P2_U3545) );
  AOI22_X1 U10094 ( .A1(n8682), .A2(n8763), .B1(n8762), .B2(n8681), .ZN(n8683)
         );
  OAI211_X1 U10095 ( .C1(n8685), .C2(n8767), .A(n8684), .B(n8683), .ZN(n8775)
         );
  MUX2_X1 U10096 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8775), .S(n10084), .Z(
        P2_U3544) );
  AOI211_X1 U10097 ( .C1(n8762), .C2(n8688), .A(n8687), .B(n8686), .ZN(n8689)
         );
  OAI21_X1 U10098 ( .B1(n8690), .B2(n8767), .A(n8689), .ZN(n8776) );
  MUX2_X1 U10099 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8776), .S(n10084), .Z(
        P2_U3543) );
  AOI22_X1 U10100 ( .A1(n8692), .A2(n8763), .B1(n8762), .B2(n4433), .ZN(n8693)
         );
  OAI211_X1 U10101 ( .C1(n8695), .C2(n8767), .A(n8694), .B(n8693), .ZN(n8777)
         );
  MUX2_X1 U10102 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8777), .S(n10084), .Z(
        P2_U3542) );
  AOI211_X1 U10103 ( .C1(n8762), .C2(n8698), .A(n8697), .B(n8696), .ZN(n8699)
         );
  OAI21_X1 U10104 ( .B1(n8700), .B2(n8767), .A(n8699), .ZN(n8778) );
  MUX2_X1 U10105 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8778), .S(n10084), .Z(
        P2_U3541) );
  AOI22_X1 U10106 ( .A1(n8702), .A2(n8763), .B1(n8762), .B2(n8701), .ZN(n8703)
         );
  OAI211_X1 U10107 ( .C1(n8705), .C2(n8767), .A(n8704), .B(n8703), .ZN(n8779)
         );
  MUX2_X1 U10108 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8779), .S(n10084), .Z(
        P2_U3540) );
  AOI21_X1 U10109 ( .B1(n8762), .B2(n8707), .A(n8706), .ZN(n8708) );
  OAI211_X1 U10110 ( .C1(n8710), .C2(n8767), .A(n8709), .B(n8708), .ZN(n8780)
         );
  MUX2_X1 U10111 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8780), .S(n10084), .Z(
        P2_U3539) );
  AOI22_X1 U10112 ( .A1(n8712), .A2(n8763), .B1(n8762), .B2(n8711), .ZN(n8713)
         );
  OAI211_X1 U10113 ( .C1(n8715), .C2(n8767), .A(n8714), .B(n8713), .ZN(n8781)
         );
  MUX2_X1 U10114 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8781), .S(n10084), .Z(
        P2_U3538) );
  AOI21_X1 U10115 ( .B1(n8762), .B2(n8717), .A(n8716), .ZN(n8718) );
  OAI211_X1 U10116 ( .C1(n8720), .C2(n8767), .A(n8719), .B(n8718), .ZN(n8782)
         );
  MUX2_X1 U10117 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8782), .S(n10084), .Z(
        P2_U3537) );
  AOI22_X1 U10118 ( .A1(n8722), .A2(n8763), .B1(n8762), .B2(n8721), .ZN(n8723)
         );
  OAI211_X1 U10119 ( .C1(n8759), .C2(n8725), .A(n8724), .B(n8723), .ZN(n8783)
         );
  MUX2_X1 U10120 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8783), .S(n10084), .Z(
        P2_U3536) );
  AOI211_X1 U10121 ( .C1(n8762), .C2(n8728), .A(n8727), .B(n8726), .ZN(n8729)
         );
  OAI21_X1 U10122 ( .B1(n8730), .B2(n8767), .A(n8729), .ZN(n8784) );
  MUX2_X1 U10123 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8784), .S(n10084), .Z(
        P2_U3535) );
  INV_X1 U10124 ( .A(n8731), .ZN(n8736) );
  AOI21_X1 U10125 ( .B1(n8762), .B2(n8733), .A(n8732), .ZN(n8734) );
  OAI211_X1 U10126 ( .C1(n8736), .C2(n8767), .A(n8735), .B(n8734), .ZN(n8785)
         );
  MUX2_X1 U10127 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8785), .S(n10084), .Z(
        P2_U3534) );
  AOI22_X1 U10128 ( .A1(n8738), .A2(n8763), .B1(n8762), .B2(n8737), .ZN(n8739)
         );
  OAI21_X1 U10129 ( .B1(n8740), .B2(n8759), .A(n8739), .ZN(n8741) );
  OR2_X1 U10130 ( .A1(n8742), .A2(n8741), .ZN(n8786) );
  MUX2_X1 U10131 ( .A(n8786), .B(P2_REG1_REG_13__SCAN_IN), .S(n10081), .Z(
        P2_U3533) );
  AOI22_X1 U10132 ( .A1(n8744), .A2(n8763), .B1(n8762), .B2(n8743), .ZN(n8745)
         );
  OAI211_X1 U10133 ( .C1(n8767), .C2(n8747), .A(n8746), .B(n8745), .ZN(n8787)
         );
  MUX2_X1 U10134 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8787), .S(n10084), .Z(
        P2_U3532) );
  OAI22_X1 U10135 ( .A1(n8749), .A2(n10052), .B1(n8748), .B2(n10070), .ZN(
        n8750) );
  INV_X1 U10136 ( .A(n8750), .ZN(n8751) );
  OAI211_X1 U10137 ( .C1(n8767), .C2(n8753), .A(n8752), .B(n8751), .ZN(n8788)
         );
  MUX2_X1 U10138 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8788), .S(n10084), .Z(
        P2_U3531) );
  OAI22_X1 U10139 ( .A1(n8755), .A2(n10052), .B1(n8754), .B2(n10070), .ZN(
        n8756) );
  INV_X1 U10140 ( .A(n8756), .ZN(n8757) );
  OAI211_X1 U10141 ( .C1(n8760), .C2(n8759), .A(n8758), .B(n8757), .ZN(n8789)
         );
  MUX2_X1 U10142 ( .A(n8789), .B(P2_REG1_REG_10__SCAN_IN), .S(n10081), .Z(
        P2_U3530) );
  AOI22_X1 U10143 ( .A1(n8764), .A2(n8763), .B1(n8762), .B2(n8761), .ZN(n8765)
         );
  OAI211_X1 U10144 ( .C1(n8768), .C2(n8767), .A(n8766), .B(n8765), .ZN(n10040)
         );
  MUX2_X1 U10145 ( .A(n10040), .B(P2_REG1_REG_2__SCAN_IN), .S(n10081), .Z(
        P2_U3522) );
  MUX2_X1 U10146 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8769), .S(n10076), .Z(
        P2_U3519) );
  MUX2_X1 U10147 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8770), .S(n10076), .Z(
        P2_U3518) );
  MUX2_X1 U10148 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8771), .S(n10076), .Z(
        P2_U3517) );
  MUX2_X1 U10149 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8772), .S(n10076), .Z(
        P2_U3515) );
  MUX2_X1 U10150 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8773), .S(n10076), .Z(
        P2_U3514) );
  MUX2_X1 U10151 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8774), .S(n10076), .Z(
        P2_U3513) );
  MUX2_X1 U10152 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8775), .S(n10076), .Z(
        P2_U3512) );
  MUX2_X1 U10153 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8776), .S(n10076), .Z(
        P2_U3511) );
  MUX2_X1 U10154 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8777), .S(n10076), .Z(
        P2_U3510) );
  MUX2_X1 U10155 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8778), .S(n10076), .Z(
        P2_U3509) );
  MUX2_X1 U10156 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8779), .S(n10076), .Z(
        P2_U3508) );
  MUX2_X1 U10157 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8780), .S(n10076), .Z(
        P2_U3507) );
  MUX2_X1 U10158 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8781), .S(n10076), .Z(
        P2_U3505) );
  MUX2_X1 U10159 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8782), .S(n10076), .Z(
        P2_U3502) );
  MUX2_X1 U10160 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8783), .S(n10076), .Z(
        P2_U3499) );
  MUX2_X1 U10161 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8784), .S(n10076), .Z(
        P2_U3496) );
  MUX2_X1 U10162 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8785), .S(n10076), .Z(
        P2_U3493) );
  MUX2_X1 U10163 ( .A(n8786), .B(P2_REG0_REG_13__SCAN_IN), .S(n10074), .Z(
        P2_U3490) );
  MUX2_X1 U10164 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8787), .S(n10076), .Z(
        P2_U3487) );
  MUX2_X1 U10165 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8788), .S(n10076), .Z(
        P2_U3484) );
  MUX2_X1 U10166 ( .A(n8789), .B(P2_REG0_REG_10__SCAN_IN), .S(n10074), .Z(
        P2_U3481) );
  INV_X1 U10167 ( .A(n9055), .ZN(n9853) );
  NOR4_X1 U10168 ( .A1(n8791), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5270), .A4(
        P2_U3152), .ZN(n8792) );
  AOI21_X1 U10169 ( .B1(n8793), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8792), .ZN(
        n8794) );
  OAI21_X1 U10170 ( .B1(n9853), .B2(n4275), .A(n8794), .ZN(P2_U3327) );
  NAND2_X1 U10171 ( .A1(n9859), .A2(n8795), .ZN(n8797) );
  OAI211_X1 U10172 ( .C1(n8802), .C2(n8798), .A(n8797), .B(n8796), .ZN(
        P2_U3330) );
  INV_X1 U10173 ( .A(n8799), .ZN(n9867) );
  OAI222_X1 U10174 ( .A1(n8802), .A2(n8801), .B1(n4275), .B2(n9867), .C1(n8800), .C2(P2_U3152), .ZN(P2_U3331) );
  MUX2_X1 U10175 ( .A(n8803), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10176 ( .A(n8827), .ZN(n8804) );
  NAND2_X1 U10177 ( .A1(n9686), .A2(n8883), .ZN(n8805) );
  NAND2_X1 U10178 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  XNOR2_X1 U10179 ( .A(n8807), .B(n8880), .ZN(n8962) );
  NAND2_X1 U10180 ( .A1(n9673), .A2(n8923), .ZN(n8809) );
  NAND2_X1 U10181 ( .A1(n9686), .A2(n8924), .ZN(n8808) );
  AND2_X1 U10182 ( .A1(n8809), .A2(n8808), .ZN(n8821) );
  NAND2_X1 U10183 ( .A1(n8962), .A2(n8821), .ZN(n8972) );
  NAND2_X1 U10184 ( .A1(n9807), .A2(n8883), .ZN(n8811) );
  NAND2_X1 U10185 ( .A1(n9704), .A2(n8924), .ZN(n8810) );
  NAND2_X1 U10186 ( .A1(n8811), .A2(n8810), .ZN(n9040) );
  NAND2_X1 U10187 ( .A1(n9345), .A2(n8923), .ZN(n8814) );
  NAND2_X1 U10188 ( .A1(n8815), .A2(n8814), .ZN(n8816) );
  XNOR2_X1 U10189 ( .A(n8816), .B(n8880), .ZN(n8830) );
  NOR2_X1 U10190 ( .A1(n9657), .A2(n6727), .ZN(n8817) );
  AOI21_X1 U10191 ( .B1(n9642), .B2(n8883), .A(n8817), .ZN(n8829) );
  NOR2_X1 U10192 ( .A1(n8830), .A2(n8829), .ZN(n8974) );
  NAND2_X1 U10193 ( .A1(n9704), .A2(n8923), .ZN(n8818) );
  NAND2_X1 U10194 ( .A1(n8819), .A2(n8818), .ZN(n8820) );
  XNOR2_X1 U10195 ( .A(n8820), .B(n8927), .ZN(n8963) );
  INV_X1 U10196 ( .A(n8821), .ZN(n8961) );
  AOI21_X1 U10197 ( .B1(n9040), .B2(n8963), .A(n8961), .ZN(n8823) );
  NAND3_X1 U10198 ( .A1(n8963), .A2(n8961), .A3(n9040), .ZN(n8822) );
  OAI21_X1 U10199 ( .B1(n8823), .B2(n8962), .A(n8822), .ZN(n8824) );
  NAND2_X1 U10200 ( .A1(n8972), .A2(n8963), .ZN(n8825) );
  NOR2_X1 U10201 ( .A1(n8826), .A2(n8825), .ZN(n8828) );
  NAND2_X1 U10202 ( .A1(n8959), .A2(n8827), .ZN(n8964) );
  NAND2_X1 U10203 ( .A1(n8830), .A2(n8829), .ZN(n8975) );
  XNOR2_X1 U10204 ( .A(n8831), .B(n8927), .ZN(n8833) );
  INV_X1 U10205 ( .A(n9624), .ZN(n9791) );
  OAI22_X1 U10206 ( .A1(n9791), .A2(n8832), .B1(n9632), .B2(n6727), .ZN(n9017)
         );
  NAND2_X1 U10207 ( .A1(n9598), .A2(n8923), .ZN(n8835) );
  NAND2_X1 U10208 ( .A1(n8836), .A2(n8835), .ZN(n8837) );
  XNOR2_X1 U10209 ( .A(n8837), .B(n8927), .ZN(n8996) );
  NAND2_X1 U10210 ( .A1(n9587), .A2(n8923), .ZN(n8839) );
  NAND2_X1 U10211 ( .A1(n9598), .A2(n8924), .ZN(n8838) );
  NAND2_X1 U10212 ( .A1(n8839), .A2(n8838), .ZN(n8995) );
  NOR2_X1 U10213 ( .A1(n8996), .A2(n8995), .ZN(n8994) );
  INV_X1 U10214 ( .A(n8994), .ZN(n8845) );
  NAND2_X1 U10215 ( .A1(n9344), .A2(n8923), .ZN(n8840) );
  NOR2_X1 U10216 ( .A1(n9615), .A2(n6727), .ZN(n8843) );
  NAND2_X1 U10217 ( .A1(n8991), .A2(n8992), .ZN(n8844) );
  INV_X1 U10218 ( .A(n8995), .ZN(n8846) );
  NOR3_X1 U10219 ( .A1(n8846), .A2(n8991), .A3(n8992), .ZN(n8848) );
  OAI21_X1 U10220 ( .B1(n8991), .B2(n8992), .A(n8846), .ZN(n8847) );
  OR2_X1 U10221 ( .A1(n9578), .A2(n8892), .ZN(n8850) );
  NAND2_X1 U10222 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  XNOR2_X1 U10223 ( .A(n8852), .B(n8880), .ZN(n8855) );
  NOR2_X1 U10224 ( .A1(n9578), .A2(n6727), .ZN(n8853) );
  AOI21_X1 U10225 ( .B1(n9571), .B2(n8923), .A(n8853), .ZN(n8854) );
  NOR2_X1 U10226 ( .A1(n8855), .A2(n8854), .ZN(n8941) );
  NAND2_X1 U10227 ( .A1(n9560), .A2(n8924), .ZN(n8856) );
  OAI22_X1 U10228 ( .A1(n9554), .A2(n6725), .B1(n9534), .B2(n8832), .ZN(n8858)
         );
  XNOR2_X1 U10229 ( .A(n8858), .B(n8927), .ZN(n9008) );
  INV_X1 U10230 ( .A(n8868), .ZN(n8866) );
  INV_X1 U10231 ( .A(n9005), .ZN(n8865) );
  NAND2_X1 U10232 ( .A1(n9342), .A2(n8923), .ZN(n8861) );
  NAND2_X1 U10233 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  XNOR2_X1 U10234 ( .A(n8863), .B(n8880), .ZN(n8867) );
  INV_X1 U10235 ( .A(n8867), .ZN(n8864) );
  OAI22_X1 U10236 ( .A1(n4421), .A2(n6715), .B1(n9548), .B2(n6727), .ZN(n8911)
         );
  NAND2_X1 U10237 ( .A1(n9341), .A2(n8923), .ZN(n8869) );
  NAND2_X1 U10238 ( .A1(n8870), .A2(n8869), .ZN(n8871) );
  XNOR2_X1 U10239 ( .A(n8871), .B(n8880), .ZN(n8874) );
  NOR2_X1 U10240 ( .A1(n9535), .A2(n6727), .ZN(n8872) );
  AOI21_X1 U10241 ( .B1(n9758), .B2(n8883), .A(n8872), .ZN(n8873) );
  NAND2_X1 U10242 ( .A1(n8874), .A2(n8873), .ZN(n8876) );
  OAI21_X1 U10243 ( .B1(n8874), .B2(n8873), .A(n8876), .ZN(n8984) );
  OAI22_X1 U10244 ( .A1(n9501), .A2(n8892), .B1(n9516), .B2(n6727), .ZN(n8884)
         );
  OAI22_X1 U10245 ( .A1(n9501), .A2(n6725), .B1(n9516), .B2(n8892), .ZN(n8877)
         );
  XNOR2_X1 U10246 ( .A(n8877), .B(n8927), .ZN(n8885) );
  XOR2_X1 U10247 ( .A(n8884), .B(n8885), .Z(n8952) );
  NAND2_X1 U10248 ( .A1(n9339), .A2(n8923), .ZN(n8878) );
  NAND2_X1 U10249 ( .A1(n8879), .A2(n8878), .ZN(n8881) );
  XNOR2_X1 U10250 ( .A(n8881), .B(n8880), .ZN(n8887) );
  NOR2_X1 U10251 ( .A1(n6727), .A2(n9500), .ZN(n8882) );
  AOI21_X1 U10252 ( .B1(n9742), .B2(n8883), .A(n8882), .ZN(n8888) );
  XNOR2_X1 U10253 ( .A(n8887), .B(n8888), .ZN(n9026) );
  NOR2_X1 U10254 ( .A1(n8885), .A2(n8884), .ZN(n9027) );
  NOR2_X1 U10255 ( .A1(n9026), .A2(n9027), .ZN(n8886) );
  INV_X1 U10256 ( .A(n8887), .ZN(n8890) );
  INV_X1 U10257 ( .A(n8888), .ZN(n8889) );
  NAND2_X1 U10258 ( .A1(n8890), .A2(n8889), .ZN(n8897) );
  XOR2_X1 U10259 ( .A(n8927), .B(n8891), .Z(n8895) );
  INV_X1 U10260 ( .A(n9474), .ZN(n8893) );
  OAI22_X1 U10261 ( .A1(n8893), .A2(n8892), .B1(n9488), .B2(n6727), .ZN(n8894)
         );
  NOR2_X1 U10262 ( .A1(n8895), .A2(n8894), .ZN(n8937) );
  AOI21_X1 U10263 ( .B1(n8895), .B2(n8894), .A(n8937), .ZN(n8896) );
  AOI21_X1 U10264 ( .B1(n9029), .B2(n8897), .A(n8896), .ZN(n8901) );
  INV_X1 U10265 ( .A(n8896), .ZN(n8899) );
  INV_X1 U10266 ( .A(n8897), .ZN(n8898) );
  OAI21_X1 U10267 ( .B1(n8901), .B2(n8931), .A(n9043), .ZN(n8907) );
  INV_X1 U10268 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8902) );
  OAI22_X1 U10269 ( .A1(n9032), .A2(n9500), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8902), .ZN(n8905) );
  OAI22_X1 U10270 ( .A1(n8903), .A2(n9048), .B1(n9047), .B2(n9477), .ZN(n8904)
         );
  AOI211_X1 U10271 ( .C1(n9474), .C2(n9022), .A(n8905), .B(n8904), .ZN(n8906)
         );
  NAND2_X1 U10272 ( .A1(n8907), .A2(n8906), .ZN(P1_U3212) );
  NAND2_X1 U10273 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  XOR2_X1 U10274 ( .A(n8911), .B(n8910), .Z(n8916) );
  AOI22_X1 U10275 ( .A1(n9560), .A2(n9050), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8913) );
  NAND2_X1 U10276 ( .A1(n9527), .A2(n9035), .ZN(n8912) );
  OAI211_X1 U10277 ( .C1(n9535), .C2(n9048), .A(n8913), .B(n8912), .ZN(n8914)
         );
  AOI21_X1 U10278 ( .B1(n9761), .B2(n9022), .A(n8914), .ZN(n8915) );
  OAI21_X1 U10279 ( .B1(n8916), .B2(n9024), .A(n8915), .ZN(P1_U3214) );
  XNOR2_X1 U10280 ( .A(n8991), .B(n8992), .ZN(n8918) );
  XNOR2_X1 U10281 ( .A(n8917), .B(n8918), .ZN(n8922) );
  NAND2_X1 U10282 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9441) );
  OAI21_X1 U10283 ( .B1(n9632), .B2(n9032), .A(n9441), .ZN(n8920) );
  OAI22_X1 U10284 ( .A1(n9562), .A2(n9048), .B1(n9047), .B2(n9601), .ZN(n8919)
         );
  AOI211_X1 U10285 ( .C1(n9785), .C2(n9022), .A(n8920), .B(n8919), .ZN(n8921)
         );
  OAI21_X1 U10286 ( .B1(n8922), .B2(n9024), .A(n8921), .ZN(P1_U3217) );
  NAND2_X1 U10287 ( .A1(n9736), .A2(n8923), .ZN(n8926) );
  NAND2_X1 U10288 ( .A1(n8924), .A2(n8051), .ZN(n8925) );
  NAND2_X1 U10289 ( .A1(n8926), .A2(n8925), .ZN(n8928) );
  XNOR2_X1 U10290 ( .A(n8928), .B(n8927), .ZN(n8930) );
  XNOR2_X1 U10291 ( .A(n8930), .B(n8929), .ZN(n8936) );
  OAI22_X1 U10292 ( .A1(n9032), .A2(n9488), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8932), .ZN(n8935) );
  INV_X1 U10293 ( .A(n9462), .ZN(n9227) );
  INV_X1 U10294 ( .A(n9469), .ZN(n8933) );
  OAI22_X1 U10295 ( .A1(n9227), .A2(n9048), .B1(n9047), .B2(n8933), .ZN(n8934)
         );
  AOI211_X1 U10296 ( .C1(n9736), .C2(n9022), .A(n8935), .B(n8934), .ZN(n8939)
         );
  NAND3_X1 U10297 ( .A1(n8937), .A2(n9043), .A3(n8936), .ZN(n8938) );
  NOR2_X1 U10298 ( .A1(n8941), .A2(n8940), .ZN(n8942) );
  XNOR2_X1 U10299 ( .A(n8943), .B(n8942), .ZN(n8949) );
  OAI22_X1 U10300 ( .A1(n9562), .A2(n9032), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8944), .ZN(n8947) );
  INV_X1 U10301 ( .A(n9570), .ZN(n8945) );
  OAI22_X1 U10302 ( .A1(n9534), .A2(n9048), .B1(n9047), .B2(n8945), .ZN(n8946)
         );
  AOI211_X1 U10303 ( .C1(n9571), .C2(n9022), .A(n8947), .B(n8946), .ZN(n8948)
         );
  OAI21_X1 U10304 ( .B1(n8949), .B2(n9024), .A(n8948), .ZN(P1_U3221) );
  OAI21_X1 U10305 ( .B1(n8952), .B2(n8951), .A(n8950), .ZN(n8953) );
  NAND2_X1 U10306 ( .A1(n8953), .A2(n9043), .ZN(n8958) );
  OAI22_X1 U10307 ( .A1(n9048), .A2(n9500), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8954), .ZN(n8956) );
  NOR2_X1 U10308 ( .A1(n9505), .A2(n9047), .ZN(n8955) );
  AOI211_X1 U10309 ( .C1(n9341), .C2(n9050), .A(n8956), .B(n8955), .ZN(n8957)
         );
  OAI211_X1 U10310 ( .C1(n9501), .C2(n9053), .A(n8958), .B(n8957), .ZN(
        P1_U3223) );
  INV_X1 U10311 ( .A(n8963), .ZN(n8960) );
  NAND2_X1 U10312 ( .A1(n9039), .A2(n9040), .ZN(n9045) );
  XNOR2_X1 U10313 ( .A(n8962), .B(n8961), .ZN(n8966) );
  AND2_X1 U10314 ( .A1(n4500), .A2(n8963), .ZN(n8965) );
  NAND2_X1 U10315 ( .A1(n8965), .A2(n8964), .ZN(n9038) );
  NAND3_X1 U10316 ( .A1(n9045), .A2(n8966), .A3(n9038), .ZN(n8973) );
  INV_X1 U10317 ( .A(n8973), .ZN(n8968) );
  AOI21_X1 U10318 ( .B1(n9045), .B2(n9038), .A(n8966), .ZN(n8967) );
  OAI21_X1 U10319 ( .B1(n8968), .B2(n8967), .A(n9043), .ZN(n8971) );
  AND2_X1 U10320 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9399) );
  OAI22_X1 U10321 ( .A1(n9655), .A2(n9032), .B1(n9047), .B2(n9668), .ZN(n8969)
         );
  AOI211_X1 U10322 ( .C1(n9019), .C2(n9345), .A(n9399), .B(n8969), .ZN(n8970)
         );
  OAI211_X1 U10323 ( .C1(n4442), .C2(n9053), .A(n8971), .B(n8970), .ZN(
        P1_U3224) );
  NAND2_X1 U10324 ( .A1(n8973), .A2(n8972), .ZN(n8978) );
  INV_X1 U10325 ( .A(n8974), .ZN(n8976) );
  NAND2_X1 U10326 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  XNOR2_X1 U10327 ( .A(n8978), .B(n8977), .ZN(n8982) );
  AOI22_X1 U10328 ( .A1(n9050), .A2(n9686), .B1(n9035), .B2(n9641), .ZN(n8979)
         );
  NAND2_X1 U10329 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9420) );
  OAI211_X1 U10330 ( .C1(n9632), .C2(n9048), .A(n8979), .B(n9420), .ZN(n8980)
         );
  AOI21_X1 U10331 ( .B1(n9642), .B2(n9022), .A(n8980), .ZN(n8981) );
  OAI21_X1 U10332 ( .B1(n8982), .B2(n9024), .A(n8981), .ZN(P1_U3226) );
  AOI21_X1 U10333 ( .B1(n8984), .B2(n8983), .A(n8875), .ZN(n8989) );
  AOI22_X1 U10334 ( .A1(n9520), .A2(n9035), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8986) );
  NAND2_X1 U10335 ( .A1(n9342), .A2(n9050), .ZN(n8985) );
  OAI211_X1 U10336 ( .C1(n9516), .C2(n9048), .A(n8986), .B(n8985), .ZN(n8987)
         );
  AOI21_X1 U10337 ( .B1(n9758), .B2(n9022), .A(n8987), .ZN(n8988) );
  OAI21_X1 U10338 ( .B1(n8989), .B2(n9024), .A(n8988), .ZN(P1_U3227) );
  INV_X1 U10339 ( .A(n8991), .ZN(n8990) );
  NOR2_X1 U10340 ( .A1(n4926), .A2(n8990), .ZN(n8993) );
  OAI22_X1 U10341 ( .A1(n8993), .A2(n8992), .B1(n8917), .B2(n8991), .ZN(n8998)
         );
  AOI21_X1 U10342 ( .B1(n8996), .B2(n8995), .A(n8994), .ZN(n8997) );
  XNOR2_X1 U10343 ( .A(n8998), .B(n8997), .ZN(n9004) );
  OAI22_X1 U10344 ( .A1(n9615), .A2(n9032), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8999), .ZN(n9002) );
  OAI22_X1 U10345 ( .A1(n9578), .A2(n9048), .B1(n9047), .B2(n9000), .ZN(n9001)
         );
  AOI211_X1 U10346 ( .C1(n9587), .C2(n9022), .A(n9002), .B(n9001), .ZN(n9003)
         );
  OAI21_X1 U10347 ( .B1(n9004), .B2(n9024), .A(n9003), .ZN(P1_U3231) );
  NAND2_X1 U10348 ( .A1(n9006), .A2(n9005), .ZN(n9007) );
  XOR2_X1 U10349 ( .A(n9008), .B(n9007), .Z(n9013) );
  NOR2_X1 U10350 ( .A1(n9548), .A2(n9048), .ZN(n9011) );
  INV_X1 U10351 ( .A(n9578), .ZN(n9343) );
  AOI22_X1 U10352 ( .A1(n9343), .A2(n9050), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9009) );
  OAI21_X1 U10353 ( .B1(n9550), .B2(n9047), .A(n9009), .ZN(n9010) );
  AOI211_X1 U10354 ( .C1(n9768), .C2(n9022), .A(n9011), .B(n9010), .ZN(n9012)
         );
  OAI21_X1 U10355 ( .B1(n9013), .B2(n9024), .A(n9012), .ZN(P1_U3233) );
  INV_X1 U10356 ( .A(n9014), .ZN(n9015) );
  NOR2_X1 U10357 ( .A1(n9016), .A2(n9015), .ZN(n9018) );
  XNOR2_X1 U10358 ( .A(n9018), .B(n9017), .ZN(n9025) );
  AOI22_X1 U10359 ( .A1(n9344), .A2(n9019), .B1(n9035), .B2(n9623), .ZN(n9020)
         );
  NAND2_X1 U10360 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9916) );
  OAI211_X1 U10361 ( .C1(n9657), .C2(n9032), .A(n9020), .B(n9916), .ZN(n9021)
         );
  AOI21_X1 U10362 ( .B1(n9624), .B2(n9022), .A(n9021), .ZN(n9023) );
  OAI21_X1 U10363 ( .B1(n9025), .B2(n9024), .A(n9023), .ZN(P1_U3236) );
  INV_X1 U10364 ( .A(n8950), .ZN(n9028) );
  OAI21_X1 U10365 ( .B1(n9028), .B2(n9027), .A(n9026), .ZN(n9030) );
  NAND3_X1 U10366 ( .A1(n9030), .A2(n9043), .A3(n9029), .ZN(n9037) );
  OAI22_X1 U10367 ( .A1(n9048), .A2(n9488), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9031), .ZN(n9034) );
  NOR2_X1 U10368 ( .A1(n9516), .A2(n9032), .ZN(n9033) );
  AOI211_X1 U10369 ( .C1(n9035), .C2(n9491), .A(n9034), .B(n9033), .ZN(n9036)
         );
  OAI211_X1 U10370 ( .C1(n9494), .C2(n9053), .A(n9037), .B(n9036), .ZN(
        P1_U3238) );
  INV_X1 U10371 ( .A(n9807), .ZN(n9696) );
  INV_X1 U10372 ( .A(n9038), .ZN(n9046) );
  INV_X1 U10373 ( .A(n9039), .ZN(n9042) );
  INV_X1 U10374 ( .A(n9040), .ZN(n9041) );
  OAI21_X1 U10375 ( .B1(n9042), .B2(n9046), .A(n9041), .ZN(n9044) );
  OAI211_X1 U10376 ( .C1(n9046), .C2(n9045), .A(n9044), .B(n9043), .ZN(n9052)
         );
  NOR2_X1 U10377 ( .A1(n10234), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9383) );
  OAI22_X1 U10378 ( .A1(n9631), .A2(n9048), .B1(n9047), .B2(n9692), .ZN(n9049)
         );
  AOI211_X1 U10379 ( .C1(n9050), .C2(n9685), .A(n9383), .B(n9049), .ZN(n9051)
         );
  OAI211_X1 U10380 ( .C1(n9696), .C2(n9053), .A(n9052), .B(n9051), .ZN(
        P1_U3239) );
  NAND2_X1 U10381 ( .A1(n9057), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U10382 ( .A1(n9058), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U10383 ( .A1(n9059), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9060) );
  AND3_X1 U10384 ( .A1(n9062), .A2(n9061), .A3(n9060), .ZN(n9444) );
  INV_X1 U10385 ( .A(n9444), .ZN(n9337) );
  NOR2_X1 U10386 ( .A1(n6379), .A2(n9165), .ZN(n9063) );
  NAND2_X1 U10387 ( .A1(n9065), .A2(n6091), .ZN(n9068) );
  NAND2_X1 U10388 ( .A1(n9066), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9067) );
  OR2_X1 U10389 ( .A1(n9725), .A2(n9241), .ZN(n9239) );
  NAND2_X1 U10390 ( .A1(n9239), .A2(n9337), .ZN(n9069) );
  NAND2_X1 U10391 ( .A1(n9721), .A2(n9069), .ZN(n9235) );
  INV_X1 U10392 ( .A(n9070), .ZN(n9071) );
  OAI21_X1 U10393 ( .B1(n9072), .B2(n9071), .A(n9299), .ZN(n9075) );
  INV_X1 U10394 ( .A(n9073), .ZN(n9257) );
  INV_X1 U10395 ( .A(n9076), .ZN(n9079) );
  AND2_X1 U10396 ( .A1(n9087), .A2(n9080), .ZN(n9083) );
  INV_X1 U10397 ( .A(n9081), .ZN(n9082) );
  AOI21_X1 U10398 ( .B1(n9084), .B2(n9083), .A(n9082), .ZN(n9091) );
  NAND2_X1 U10399 ( .A1(n9086), .A2(n9085), .ZN(n9089) );
  INV_X1 U10400 ( .A(n9087), .ZN(n9088) );
  AOI21_X1 U10401 ( .B1(n9089), .B2(n9192), .A(n9088), .ZN(n9090) );
  MUX2_X1 U10402 ( .A(n9091), .B(n9090), .S(n9160), .Z(n9092) );
  NAND2_X1 U10403 ( .A1(n9092), .A2(n9261), .ZN(n9110) );
  INV_X1 U10404 ( .A(n9109), .ZN(n9094) );
  AND4_X1 U10405 ( .A1(n9173), .A2(n9175), .A3(n4569), .A4(n9174), .ZN(n9093)
         );
  NAND3_X1 U10406 ( .A1(n9818), .A2(n9095), .A3(n4569), .ZN(n9096) );
  NAND2_X1 U10407 ( .A1(n9098), .A2(n4569), .ZN(n9097) );
  NAND2_X1 U10408 ( .A1(n9096), .A2(n9097), .ZN(n9102) );
  OAI21_X1 U10409 ( .B1(n9706), .B2(n9097), .A(n9818), .ZN(n9101) );
  NOR2_X1 U10410 ( .A1(n9098), .A2(n4569), .ZN(n9103) );
  AND2_X1 U10411 ( .A1(n9103), .A2(n9706), .ZN(n9099) );
  OR2_X1 U10412 ( .A1(n9818), .A2(n9099), .ZN(n9100) );
  AOI22_X1 U10413 ( .A1(n9102), .A2(n4411), .B1(n9101), .B2(n9100), .ZN(n9107)
         );
  INV_X1 U10414 ( .A(n9103), .ZN(n9104) );
  OAI21_X1 U10415 ( .B1(n9174), .B2(n4569), .A(n9104), .ZN(n9105) );
  NAND2_X1 U10416 ( .A1(n9105), .A2(n4873), .ZN(n9106) );
  OR2_X1 U10417 ( .A1(n9902), .A2(n9347), .ZN(n9108) );
  AND2_X1 U10418 ( .A1(n9109), .A2(n9108), .ZN(n9193) );
  NAND2_X1 U10419 ( .A1(n9110), .A2(n9193), .ZN(n9113) );
  NAND3_X1 U10420 ( .A1(n9177), .A2(n9160), .A3(n9195), .ZN(n9111) );
  AOI21_X1 U10421 ( .B1(n9113), .B2(n9112), .A(n9111), .ZN(n9115) );
  MUX2_X1 U10422 ( .A(n9181), .B(n9178), .S(n9160), .Z(n9114) );
  INV_X1 U10423 ( .A(n9650), .ZN(n9663) );
  MUX2_X1 U10424 ( .A(n9182), .B(n9168), .S(n9160), .Z(n9116) );
  AND2_X1 U10425 ( .A1(n9594), .A2(n6202), .ZN(n9117) );
  MUX2_X1 U10426 ( .A(n9117), .B(n9187), .S(n4569), .Z(n9118) );
  NAND2_X1 U10427 ( .A1(n9119), .A2(n9118), .ZN(n9123) );
  NAND3_X1 U10428 ( .A1(n9123), .A2(n9124), .A3(n9120), .ZN(n9122) );
  INV_X1 U10429 ( .A(n9246), .ZN(n9121) );
  NAND3_X1 U10430 ( .A1(n9123), .A2(n9594), .A3(n9201), .ZN(n9125) );
  AND2_X1 U10431 ( .A1(n9245), .A2(n9124), .ZN(n9189) );
  INV_X1 U10432 ( .A(n9126), .ZN(n9127) );
  INV_X1 U10433 ( .A(n9148), .ZN(n9128) );
  NAND2_X1 U10434 ( .A1(n9128), .A2(n9218), .ZN(n9513) );
  INV_X1 U10435 ( .A(n9513), .ZN(n9511) );
  NAND3_X1 U10436 ( .A1(n9129), .A2(n9511), .A3(n9216), .ZN(n9132) );
  INV_X1 U10437 ( .A(n9145), .ZN(n9130) );
  OR2_X1 U10438 ( .A1(n9148), .A2(n9130), .ZN(n9310) );
  NAND2_X1 U10439 ( .A1(n9310), .A2(n9218), .ZN(n9131) );
  AND2_X1 U10440 ( .A1(n9311), .A2(n9131), .ZN(n9221) );
  NAND2_X1 U10441 ( .A1(n9494), .A2(n9147), .ZN(n9133) );
  NAND2_X1 U10442 ( .A1(n9133), .A2(n9500), .ZN(n9135) );
  OAI21_X1 U10443 ( .B1(n9494), .B2(n9147), .A(n9135), .ZN(n9134) );
  OR2_X1 U10444 ( .A1(n9457), .A2(n9160), .ZN(n9141) );
  INV_X1 U10445 ( .A(n9135), .ZN(n9136) );
  NAND4_X1 U10446 ( .A1(n9136), .A2(n9457), .A3(n9160), .A4(n9742), .ZN(n9140)
         );
  OR2_X1 U10447 ( .A1(n9225), .A2(n4569), .ZN(n9139) );
  INV_X1 U10448 ( .A(n9150), .ZN(n9137) );
  NAND4_X1 U10449 ( .A1(n9225), .A2(n9137), .A3(n4569), .A4(n9339), .ZN(n9138)
         );
  NAND2_X1 U10450 ( .A1(n9545), .A2(n9246), .ZN(n9143) );
  AND2_X1 U10451 ( .A1(n9143), .A2(n9142), .ZN(n9144) );
  NAND2_X1 U10452 ( .A1(n9144), .A2(n9531), .ZN(n9306) );
  INV_X1 U10453 ( .A(n9218), .ZN(n9146) );
  NOR2_X1 U10454 ( .A1(n9147), .A2(n9146), .ZN(n9281) );
  NAND2_X1 U10455 ( .A1(n9311), .A2(n9339), .ZN(n9149) );
  AOI21_X1 U10456 ( .B1(n9150), .B2(n9149), .A(n9160), .ZN(n9151) );
  NAND3_X1 U10457 ( .A1(n9152), .A2(n9151), .A3(n9225), .ZN(n9153) );
  MUX2_X1 U10458 ( .A(n9226), .B(n9166), .S(n9160), .Z(n9154) );
  INV_X1 U10459 ( .A(n9241), .ZN(n9338) );
  NAND2_X1 U10460 ( .A1(n9338), .A2(n9337), .ZN(n9155) );
  NAND2_X1 U10461 ( .A1(n9725), .A2(n9155), .ZN(n9232) );
  NAND3_X1 U10462 ( .A1(n9157), .A2(n9232), .A3(n9462), .ZN(n9156) );
  INV_X1 U10463 ( .A(n9240), .ZN(n9158) );
  MUX2_X1 U10464 ( .A(n9462), .B(n9228), .S(n9160), .Z(n9161) );
  INV_X1 U10465 ( .A(n9161), .ZN(n9162) );
  NAND2_X1 U10466 ( .A1(n9232), .A2(n9162), .ZN(n9163) );
  NAND2_X1 U10467 ( .A1(n9165), .A2(n9164), .ZN(n9275) );
  AND2_X1 U10468 ( .A1(n9167), .A2(n9166), .ZN(n9231) );
  INV_X1 U10469 ( .A(n9231), .ZN(n9320) );
  INV_X1 U10470 ( .A(n9168), .ZN(n9169) );
  NOR2_X1 U10471 ( .A1(n9170), .A2(n9169), .ZN(n9199) );
  NAND2_X1 U10472 ( .A1(n9195), .A2(n9193), .ZN(n9171) );
  NOR2_X1 U10473 ( .A1(n9172), .A2(n9171), .ZN(n9180) );
  INV_X1 U10474 ( .A(n9195), .ZN(n9176) );
  OAI211_X1 U10475 ( .C1(n9176), .C2(n9175), .A(n9174), .B(n9173), .ZN(n9179)
         );
  AND2_X1 U10476 ( .A1(n9178), .A2(n9177), .ZN(n9191) );
  OAI21_X1 U10477 ( .B1(n9180), .B2(n9179), .A(n9191), .ZN(n9183) );
  NAND3_X1 U10478 ( .A1(n9183), .A2(n9182), .A3(n9181), .ZN(n9184) );
  NAND2_X1 U10479 ( .A1(n9199), .A2(n9184), .ZN(n9186) );
  INV_X1 U10480 ( .A(n9594), .ZN(n9185) );
  AOI21_X1 U10481 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(n9188) );
  INV_X1 U10482 ( .A(n9188), .ZN(n9190) );
  OAI211_X1 U10483 ( .C1(n4686), .C2(n9190), .A(n9545), .B(n9189), .ZN(n9304)
         );
  INV_X1 U10484 ( .A(n9191), .ZN(n9197) );
  NAND4_X1 U10485 ( .A1(n9195), .A2(n9194), .A3(n9193), .A4(n9192), .ZN(n9196)
         );
  NOR2_X1 U10486 ( .A1(n9197), .A2(n9196), .ZN(n9198) );
  AND3_X1 U10487 ( .A1(n9199), .A2(n9198), .A3(n9594), .ZN(n9200) );
  NAND2_X1 U10488 ( .A1(n9201), .A2(n9200), .ZN(n9302) );
  OR2_X1 U10489 ( .A1(n9203), .A2(n4895), .ZN(n9204) );
  NAND2_X1 U10490 ( .A1(n9204), .A2(n9206), .ZN(n9298) );
  NAND3_X1 U10491 ( .A1(n7054), .A2(n9293), .A3(n9298), .ZN(n9213) );
  AND2_X1 U10492 ( .A1(n9206), .A2(n9205), .ZN(n9296) );
  NAND2_X1 U10493 ( .A1(n9291), .A2(n9295), .ZN(n9208) );
  NAND2_X1 U10494 ( .A1(n9296), .A2(n9209), .ZN(n9210) );
  NAND2_X1 U10495 ( .A1(n9210), .A2(n4894), .ZN(n9212) );
  INV_X1 U10496 ( .A(n9299), .ZN(n9211) );
  AOI21_X1 U10497 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(n9214) );
  NOR2_X1 U10498 ( .A1(n9302), .A2(n9214), .ZN(n9215) );
  NOR2_X1 U10499 ( .A1(n9304), .A2(n9215), .ZN(n9219) );
  AND2_X1 U10500 ( .A1(n9217), .A2(n9216), .ZN(n9282) );
  OAI211_X1 U10501 ( .C1(n9219), .C2(n9306), .A(n9218), .B(n9282), .ZN(n9220)
         );
  NAND2_X1 U10502 ( .A1(n9221), .A2(n9220), .ZN(n9222) );
  NAND4_X1 U10503 ( .A1(n9457), .A2(n9223), .A3(n9222), .A4(n9315), .ZN(n9233)
         );
  NAND2_X1 U10504 ( .A1(n9457), .A2(n9242), .ZN(n9224) );
  NAND3_X1 U10505 ( .A1(n9226), .A2(n9225), .A3(n9224), .ZN(n9230) );
  AND2_X1 U10506 ( .A1(n9228), .A2(n9227), .ZN(n9229) );
  OAI211_X1 U10507 ( .C1(n9320), .C2(n9233), .A(n9318), .B(n9232), .ZN(n9234)
         );
  NAND2_X1 U10508 ( .A1(n9235), .A2(n9234), .ZN(n9238) );
  AND2_X1 U10509 ( .A1(n9236), .A2(n9284), .ZN(n9237) );
  NAND2_X1 U10510 ( .A1(n9238), .A2(n9237), .ZN(n9277) );
  NAND2_X1 U10511 ( .A1(n9277), .A2(n9440), .ZN(n9274) );
  NAND2_X1 U10512 ( .A1(n9725), .A2(n9241), .ZN(n9317) );
  INV_X1 U10513 ( .A(n9242), .ZN(n9243) );
  NOR2_X1 U10514 ( .A1(n9283), .A2(n9249), .ZN(n9250) );
  NAND4_X1 U10515 ( .A1(n9252), .A2(n4897), .A3(n9251), .A4(n9250), .ZN(n9254)
         );
  NOR2_X1 U10516 ( .A1(n9254), .A2(n9253), .ZN(n9258) );
  NAND4_X1 U10517 ( .A1(n9258), .A2(n9257), .A3(n9256), .A4(n9255), .ZN(n9260)
         );
  NOR2_X1 U10518 ( .A1(n9260), .A2(n9259), .ZN(n9262) );
  AND4_X1 U10519 ( .A1(n6141), .A2(n9263), .A3(n9262), .A4(n9261), .ZN(n9264)
         );
  NAND4_X1 U10520 ( .A1(n9684), .A2(n4911), .A3(n9265), .A4(n9264), .ZN(n9266)
         );
  NOR2_X1 U10521 ( .A1(n9650), .A2(n9266), .ZN(n9267) );
  NAND4_X1 U10522 ( .A1(n9607), .A2(n9637), .A3(n9618), .A4(n9267), .ZN(n9268)
         );
  NOR2_X1 U10523 ( .A1(n9576), .A2(n9268), .ZN(n9269) );
  NAND4_X1 U10524 ( .A1(n9530), .A2(n9544), .A3(n9566), .A4(n9269), .ZN(n9270)
         );
  NOR2_X1 U10525 ( .A1(n9485), .A2(n9271), .ZN(n9272) );
  NAND3_X1 U10526 ( .A1(n9277), .A2(n9284), .A3(n9440), .ZN(n9278) );
  INV_X1 U10527 ( .A(n9281), .ZN(n9313) );
  INV_X1 U10528 ( .A(n9282), .ZN(n9308) );
  INV_X1 U10529 ( .A(n9283), .ZN(n9285) );
  AND2_X1 U10530 ( .A1(n9285), .A2(n9284), .ZN(n9289) );
  OAI211_X1 U10531 ( .C1(n9289), .C2(n9288), .A(n9287), .B(n9286), .ZN(n9292)
         );
  NAND3_X1 U10532 ( .A1(n9292), .A2(n9291), .A3(n9290), .ZN(n9294) );
  NAND2_X1 U10533 ( .A1(n9294), .A2(n9293), .ZN(n9297) );
  NAND3_X1 U10534 ( .A1(n9297), .A2(n9296), .A3(n9295), .ZN(n9300) );
  AND3_X1 U10535 ( .A1(n9300), .A2(n9299), .A3(n9298), .ZN(n9301) );
  NOR2_X1 U10536 ( .A1(n9302), .A2(n9301), .ZN(n9303) );
  NOR2_X1 U10537 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  NOR2_X1 U10538 ( .A1(n9306), .A2(n9305), .ZN(n9307) );
  NOR2_X1 U10539 ( .A1(n9308), .A2(n9307), .ZN(n9309) );
  NOR2_X1 U10540 ( .A1(n9310), .A2(n9309), .ZN(n9312) );
  OAI21_X1 U10541 ( .B1(n9313), .B2(n9312), .A(n9311), .ZN(n9314) );
  NAND3_X1 U10542 ( .A1(n9316), .A2(n9315), .A3(n9314), .ZN(n9319) );
  OAI211_X1 U10543 ( .C1(n9320), .C2(n9319), .A(n9318), .B(n9317), .ZN(n9322)
         );
  AOI21_X1 U10544 ( .B1(n4281), .B2(n9322), .A(n9321), .ZN(n9328) );
  INV_X1 U10545 ( .A(n9323), .ZN(n9327) );
  NAND2_X1 U10546 ( .A1(n9328), .A2(n9324), .ZN(n9326) );
  OAI211_X1 U10547 ( .C1(n9328), .C2(n9327), .A(n9326), .B(n9325), .ZN(n9335)
         );
  NOR3_X1 U10548 ( .A1(n9331), .A2(n9330), .A3(n9329), .ZN(n9334) );
  OAI21_X1 U10549 ( .B1(n6379), .B2(n9332), .A(P1_B_REG_SCAN_IN), .ZN(n9333)
         );
  MUX2_X1 U10550 ( .A(n9337), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9336), .Z(
        P1_U3586) );
  MUX2_X1 U10551 ( .A(n9338), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9336), .Z(
        P1_U3585) );
  MUX2_X1 U10552 ( .A(n9462), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9336), .Z(
        P1_U3584) );
  MUX2_X1 U10553 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8051), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10554 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9463), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10555 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9339), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10556 ( .A(n9340), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9336), .Z(
        P1_U3580) );
  MUX2_X1 U10557 ( .A(n9341), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9336), .Z(
        P1_U3579) );
  MUX2_X1 U10558 ( .A(n9342), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9336), .Z(
        P1_U3578) );
  MUX2_X1 U10559 ( .A(n9560), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9336), .Z(
        P1_U3577) );
  MUX2_X1 U10560 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9343), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10561 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9598), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10562 ( .A(n9344), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9336), .Z(
        P1_U3574) );
  MUX2_X1 U10563 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9597), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10564 ( .A(n9345), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9336), .Z(
        P1_U3572) );
  MUX2_X1 U10565 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9686), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10566 ( .A(n9704), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9336), .Z(
        P1_U3570) );
  MUX2_X1 U10567 ( .A(n9685), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9336), .Z(
        P1_U3569) );
  MUX2_X1 U10568 ( .A(n9706), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9336), .Z(
        P1_U3568) );
  MUX2_X1 U10569 ( .A(n9346), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9336), .Z(
        P1_U3567) );
  MUX2_X1 U10570 ( .A(n9347), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9336), .Z(
        P1_U3566) );
  MUX2_X1 U10571 ( .A(n9348), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9336), .Z(
        P1_U3565) );
  MUX2_X1 U10572 ( .A(n9349), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9336), .Z(
        P1_U3564) );
  MUX2_X1 U10573 ( .A(n9350), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9336), .Z(
        P1_U3563) );
  MUX2_X1 U10574 ( .A(n9351), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9336), .Z(
        P1_U3562) );
  MUX2_X1 U10575 ( .A(n9352), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9336), .Z(
        P1_U3561) );
  MUX2_X1 U10576 ( .A(n9353), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9336), .Z(
        P1_U3560) );
  MUX2_X1 U10577 ( .A(n9354), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9336), .Z(
        P1_U3559) );
  MUX2_X1 U10578 ( .A(n9355), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9336), .Z(
        P1_U3558) );
  MUX2_X1 U10579 ( .A(n9356), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9336), .Z(
        P1_U3557) );
  MUX2_X1 U10580 ( .A(n9357), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9336), .Z(
        P1_U3556) );
  MUX2_X1 U10581 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6334), .S(P1_U4006), .Z(
        P1_U3555) );
  INV_X1 U10582 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9358) );
  XNOR2_X1 U10583 ( .A(n9378), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9373) );
  XNOR2_X1 U10584 ( .A(n9374), .B(n9373), .ZN(n9371) );
  NAND2_X1 U10585 ( .A1(n9927), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n9363) );
  OAI211_X1 U10586 ( .C1(n9366), .C2(n9918), .A(n9363), .B(n9362), .ZN(n9370)
         );
  XNOR2_X1 U10587 ( .A(n9376), .B(n9366), .ZN(n9368) );
  INV_X1 U10588 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9367) );
  NOR2_X1 U10589 ( .A1(n9368), .A2(n9367), .ZN(n9377) );
  AOI211_X1 U10590 ( .C1(n9368), .C2(n9367), .A(n9438), .B(n9377), .ZN(n9369)
         );
  AOI211_X1 U10591 ( .C1(n9410), .C2(n9371), .A(n9370), .B(n9369), .ZN(n9372)
         );
  INV_X1 U10592 ( .A(n9372), .ZN(P1_U3255) );
  OAI22_X1 U10593 ( .A1(n9374), .A2(n9373), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9378), .ZN(n9387) );
  XNOR2_X1 U10594 ( .A(n9387), .B(n9389), .ZN(n9375) );
  OAI21_X1 U10595 ( .B1(n9375), .B2(P1_REG1_REG_15__SCAN_IN), .A(n9410), .ZN(
        n9386) );
  INV_X1 U10596 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9379) );
  AOI211_X1 U10597 ( .C1(n9380), .C2(n9379), .A(n9395), .B(n9438), .ZN(n9381)
         );
  INV_X1 U10598 ( .A(n9381), .ZN(n9385) );
  NOR2_X1 U10599 ( .A1(n9918), .A2(n9393), .ZN(n9382) );
  AOI211_X1 U10600 ( .C1(n9927), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n9383), .B(
        n9382), .ZN(n9384) );
  OAI211_X1 U10601 ( .C1(n9388), .C2(n9386), .A(n9385), .B(n9384), .ZN(
        P1_U3256) );
  INV_X1 U10602 ( .A(n9387), .ZN(n9390) );
  XNOR2_X1 U10603 ( .A(n9400), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9391) );
  NOR2_X1 U10604 ( .A1(n9392), .A2(n9391), .ZN(n9407) );
  AOI211_X1 U10605 ( .C1(n9392), .C2(n9391), .A(n9407), .B(n9923), .ZN(n9405)
         );
  NAND2_X1 U10606 ( .A1(n9400), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9397) );
  OAI21_X1 U10607 ( .B1(n9400), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9397), .ZN(
        n9398) );
  AOI211_X1 U10608 ( .C1(n4313), .C2(n9398), .A(n9413), .B(n9438), .ZN(n9404)
         );
  INV_X1 U10609 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9402) );
  AOI21_X1 U10610 ( .B1(n9418), .B2(n9400), .A(n9399), .ZN(n9401) );
  OAI21_X1 U10611 ( .B1(n9442), .B2(n9402), .A(n9401), .ZN(n9403) );
  OR3_X1 U10612 ( .A1(n9405), .A2(n9404), .A3(n9403), .ZN(P1_U3257) );
  INV_X1 U10613 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9424) );
  XNOR2_X1 U10614 ( .A(n9429), .B(n9406), .ZN(n9412) );
  INV_X1 U10615 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9409) );
  INV_X1 U10616 ( .A(n9407), .ZN(n9408) );
  OAI21_X1 U10617 ( .B1(n9415), .B2(n9409), .A(n9408), .ZN(n9411) );
  NAND2_X1 U10618 ( .A1(n9412), .A2(n9411), .ZN(n9426) );
  OAI211_X1 U10619 ( .C1(n9412), .C2(n9411), .A(n9410), .B(n9426), .ZN(n9422)
         );
  INV_X1 U10620 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10117) );
  XNOR2_X1 U10621 ( .A(n9429), .B(n10117), .ZN(n9417) );
  INV_X1 U10622 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9669) );
  INV_X1 U10623 ( .A(n9413), .ZN(n9414) );
  OAI21_X1 U10624 ( .B1(n9415), .B2(n9669), .A(n9414), .ZN(n9416) );
  NAND2_X1 U10625 ( .A1(n9417), .A2(n9416), .ZN(n9431) );
  OAI211_X1 U10626 ( .C1(n9417), .C2(n9416), .A(n9913), .B(n9431), .ZN(n9421)
         );
  NAND2_X1 U10627 ( .A1(n9418), .A2(n9429), .ZN(n9419) );
  OAI21_X1 U10628 ( .B1(n9442), .B2(n9424), .A(n9423), .ZN(P1_U3258) );
  NAND2_X1 U10629 ( .A1(n9429), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U10630 ( .A1(n9426), .A2(n9425), .ZN(n9922) );
  XNOR2_X1 U10631 ( .A(n9911), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9921) );
  OR2_X1 U10632 ( .A1(n9911), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U10633 ( .A1(n9429), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U10634 ( .A1(n9431), .A2(n9430), .ZN(n9914) );
  NAND2_X1 U10635 ( .A1(n9911), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9433) );
  OR2_X1 U10636 ( .A1(n9911), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9432) );
  AND2_X1 U10637 ( .A1(n9433), .A2(n9432), .ZN(n9915) );
  NAND2_X1 U10638 ( .A1(n9914), .A2(n9915), .ZN(n9912) );
  INV_X1 U10639 ( .A(n9436), .ZN(n9437) );
  INV_X1 U10640 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9446) );
  NOR2_X1 U10641 ( .A1(n9445), .A2(n9444), .ZN(n9724) );
  NAND2_X1 U10642 ( .A1(n9724), .A2(n9670), .ZN(n9450) );
  OAI21_X1 U10643 ( .B1(n9670), .B2(n9446), .A(n9450), .ZN(n9447) );
  AOI21_X1 U10644 ( .B1(n9721), .B2(n9672), .A(n9447), .ZN(n9448) );
  OAI21_X1 U10645 ( .B1(n9723), .B2(n9645), .A(n9448), .ZN(P1_U3261) );
  XNOR2_X1 U10646 ( .A(n9449), .B(n9725), .ZN(n9727) );
  INV_X1 U10647 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9451) );
  OAI21_X1 U10648 ( .B1(n9670), .B2(n9451), .A(n9450), .ZN(n9452) );
  AOI21_X1 U10649 ( .B1(n9725), .B2(n9672), .A(n9452), .ZN(n9453) );
  OAI21_X1 U10650 ( .B1(n9727), .B2(n9645), .A(n9453), .ZN(P1_U3262) );
  AOI21_X1 U10651 ( .B1(n9459), .B2(n9455), .A(n9454), .ZN(n9456) );
  INV_X1 U10652 ( .A(n9456), .ZN(n9739) );
  AOI22_X1 U10653 ( .A1(n9463), .A2(n9705), .B1(n9703), .B2(n9462), .ZN(n9464)
         );
  INV_X1 U10654 ( .A(n9738), .ZN(n9473) );
  NAND2_X1 U10655 ( .A1(n9465), .A2(n9736), .ZN(n9466) );
  NAND2_X1 U10656 ( .A1(n9466), .A2(n10008), .ZN(n9467) );
  NOR2_X1 U10657 ( .A1(n9468), .A2(n9467), .ZN(n9735) );
  NAND2_X1 U10658 ( .A1(n9735), .A2(n9719), .ZN(n9471) );
  AOI22_X1 U10659 ( .A1(n9712), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9469), .B2(
        n9710), .ZN(n9470) );
  OAI211_X1 U10660 ( .C1(n4473), .C2(n9714), .A(n9471), .B(n9470), .ZN(n9472)
         );
  NAND2_X1 U10661 ( .A1(n9474), .A2(n9672), .ZN(n9476) );
  NAND2_X1 U10662 ( .A1(n9694), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9475) );
  OAI211_X1 U10663 ( .C1(n9667), .C2(n9477), .A(n9476), .B(n9475), .ZN(n9478)
         );
  AOI21_X1 U10664 ( .B1(n9479), .B2(n9719), .A(n9478), .ZN(n9482) );
  NAND2_X1 U10665 ( .A1(n9480), .A2(n9670), .ZN(n9481) );
  OAI211_X1 U10666 ( .C1(n9483), .C2(n9716), .A(n9482), .B(n9481), .ZN(
        P1_U3264) );
  XNOR2_X1 U10667 ( .A(n9484), .B(n9485), .ZN(n9746) );
  XNOR2_X1 U10668 ( .A(n9486), .B(n9485), .ZN(n9487) );
  OAI222_X1 U10669 ( .A1(n9654), .A2(n9516), .B1(n9656), .B2(n9488), .C1(n9557), .C2(n9487), .ZN(n9741) );
  AOI21_X1 U10670 ( .B1(n9503), .B2(n9742), .A(n10000), .ZN(n9490) );
  AND2_X1 U10671 ( .A1(n9490), .A2(n9489), .ZN(n9744) );
  NAND2_X1 U10672 ( .A1(n9744), .A2(n9719), .ZN(n9493) );
  AOI22_X1 U10673 ( .A1(n9712), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9491), .B2(
        n9710), .ZN(n9492) );
  OAI211_X1 U10674 ( .C1(n9494), .C2(n9714), .A(n9493), .B(n9492), .ZN(n9495)
         );
  AOI21_X1 U10675 ( .B1(n9741), .B2(n9670), .A(n9495), .ZN(n9496) );
  OAI21_X1 U10676 ( .B1(n9746), .B2(n9716), .A(n9496), .ZN(P1_U3265) );
  XOR2_X1 U10677 ( .A(n9497), .B(n9499), .Z(n9754) );
  OR2_X1 U10678 ( .A1(n9518), .A2(n9501), .ZN(n9502) );
  NAND2_X1 U10679 ( .A1(n9751), .A2(n9719), .ZN(n9508) );
  INV_X1 U10680 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9504) );
  OAI22_X1 U10681 ( .A1(n9505), .A2(n9667), .B1(n9504), .B2(n9670), .ZN(n9506)
         );
  AOI21_X1 U10682 ( .B1(n9752), .B2(n9672), .A(n9506), .ZN(n9507) );
  NAND2_X1 U10683 ( .A1(n9508), .A2(n9507), .ZN(n9509) );
  AOI21_X1 U10684 ( .B1(n9750), .B2(n9670), .A(n9509), .ZN(n9510) );
  OAI21_X1 U10685 ( .B1(n9754), .B2(n9716), .A(n9510), .ZN(P1_U3266) );
  XNOR2_X1 U10686 ( .A(n9512), .B(n9511), .ZN(n9760) );
  XNOR2_X1 U10687 ( .A(n9514), .B(n9513), .ZN(n9515) );
  OAI222_X1 U10688 ( .A1(n9656), .A2(n9516), .B1(n9654), .B2(n9548), .C1(n9557), .C2(n9515), .ZN(n9756) );
  OAI21_X1 U10689 ( .B1(n9526), .B2(n9517), .A(n10008), .ZN(n9519) );
  OR2_X1 U10690 ( .A1(n9519), .A2(n9518), .ZN(n9755) );
  AOI22_X1 U10691 ( .A1(n9520), .A2(n9710), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9694), .ZN(n9522) );
  NAND2_X1 U10692 ( .A1(n9758), .A2(n9672), .ZN(n9521) );
  OAI211_X1 U10693 ( .C1(n9755), .C2(n9675), .A(n9522), .B(n9521), .ZN(n9523)
         );
  AOI21_X1 U10694 ( .B1(n9756), .B2(n9670), .A(n9523), .ZN(n9524) );
  OAI21_X1 U10695 ( .B1(n9716), .B2(n9760), .A(n9524), .ZN(P1_U3267) );
  XNOR2_X1 U10696 ( .A(n9525), .B(n9530), .ZN(n9765) );
  AOI21_X1 U10697 ( .B1(n9761), .B2(n4380), .A(n9526), .ZN(n9762) );
  AOI22_X1 U10698 ( .A1(n9527), .A2(n9710), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9712), .ZN(n9528) );
  OAI21_X1 U10699 ( .B1(n4421), .B2(n9714), .A(n9528), .ZN(n9539) );
  NAND2_X1 U10700 ( .A1(n9529), .A2(n9566), .ZN(n9565) );
  NAND3_X1 U10701 ( .A1(n9565), .A2(n9544), .A3(n9545), .ZN(n9543) );
  AOI21_X1 U10702 ( .B1(n9543), .B2(n9531), .A(n9530), .ZN(n9533) );
  NOR3_X1 U10703 ( .A1(n9533), .A2(n9557), .A3(n9532), .ZN(n9537) );
  OAI22_X1 U10704 ( .A1(n9535), .A2(n9656), .B1(n9534), .B2(n9654), .ZN(n9536)
         );
  NOR2_X1 U10705 ( .A1(n9537), .A2(n9536), .ZN(n9764) );
  NOR2_X1 U10706 ( .A1(n9764), .A2(n9694), .ZN(n9538) );
  AOI211_X1 U10707 ( .C1(n9762), .C2(n9700), .A(n9539), .B(n9538), .ZN(n9540)
         );
  OAI21_X1 U10708 ( .B1(n9716), .B2(n9765), .A(n9540), .ZN(P1_U3268) );
  XNOR2_X1 U10709 ( .A(n9542), .B(n9541), .ZN(n9770) );
  INV_X1 U10710 ( .A(n9543), .ZN(n9547) );
  AOI21_X1 U10711 ( .B1(n9565), .B2(n9545), .A(n9544), .ZN(n9546) );
  AOI21_X1 U10712 ( .B1(n4311), .B2(n9768), .A(n10000), .ZN(n9549) );
  AND2_X1 U10713 ( .A1(n9549), .A2(n4380), .ZN(n9767) );
  NAND2_X1 U10714 ( .A1(n9767), .A2(n9719), .ZN(n9553) );
  INV_X1 U10715 ( .A(n9550), .ZN(n9551) );
  AOI22_X1 U10716 ( .A1(n9551), .A2(n9710), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9694), .ZN(n9552) );
  OAI211_X1 U10717 ( .C1(n9554), .C2(n9714), .A(n9553), .B(n9552), .ZN(n9555)
         );
  AOI21_X1 U10718 ( .B1(n9766), .B2(n9670), .A(n9555), .ZN(n9556) );
  OAI21_X1 U10719 ( .B1(n9716), .B2(n9770), .A(n9556), .ZN(P1_U3269) );
  INV_X1 U10720 ( .A(n9566), .ZN(n9558) );
  AOI21_X1 U10721 ( .B1(n9559), .B2(n9558), .A(n9557), .ZN(n9564) );
  NAND2_X1 U10722 ( .A1(n9560), .A2(n9703), .ZN(n9561) );
  OAI21_X1 U10723 ( .B1(n9562), .B2(n9654), .A(n9561), .ZN(n9563) );
  AOI21_X1 U10724 ( .B1(n9565), .B2(n9564), .A(n9563), .ZN(n9776) );
  NAND2_X1 U10725 ( .A1(n9567), .A2(n9566), .ZN(n9568) );
  AND2_X1 U10726 ( .A1(n9569), .A2(n9568), .ZN(n9774) );
  OAI211_X1 U10727 ( .C1(n9585), .C2(n9772), .A(n10008), .B(n4311), .ZN(n9771)
         );
  AOI22_X1 U10728 ( .A1(n9570), .A2(n9710), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9694), .ZN(n9573) );
  NAND2_X1 U10729 ( .A1(n9571), .A2(n9672), .ZN(n9572) );
  OAI211_X1 U10730 ( .C1(n9771), .C2(n9675), .A(n9573), .B(n9572), .ZN(n9574)
         );
  AOI21_X1 U10731 ( .B1(n9774), .B2(n9677), .A(n9574), .ZN(n9575) );
  OAI21_X1 U10732 ( .B1(n9776), .B2(n9694), .A(n9575), .ZN(P1_U3270) );
  XNOR2_X1 U10733 ( .A(n9577), .B(n9582), .ZN(n9580) );
  OAI22_X1 U10734 ( .A1(n9578), .A2(n9656), .B1(n9615), .B2(n9654), .ZN(n9579)
         );
  AOI21_X1 U10735 ( .B1(n9580), .B2(n9708), .A(n9579), .ZN(n9784) );
  XNOR2_X1 U10736 ( .A(n9583), .B(n9582), .ZN(n9782) );
  NOR2_X1 U10737 ( .A1(n9600), .A2(n9779), .ZN(n9584) );
  OR2_X1 U10738 ( .A1(n9585), .A2(n9584), .ZN(n9780) );
  AOI22_X1 U10739 ( .A1(n9712), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9586), .B2(
        n9710), .ZN(n9589) );
  NAND2_X1 U10740 ( .A1(n9587), .A2(n9672), .ZN(n9588) );
  OAI211_X1 U10741 ( .C1(n9780), .C2(n9645), .A(n9589), .B(n9588), .ZN(n9590)
         );
  AOI21_X1 U10742 ( .B1(n9782), .B2(n9677), .A(n9590), .ZN(n9591) );
  OAI21_X1 U10743 ( .B1(n9784), .B2(n9694), .A(n9591), .ZN(P1_U3271) );
  INV_X1 U10744 ( .A(n9607), .ZN(n9593) );
  NAND3_X1 U10745 ( .A1(n9595), .A2(n9594), .A3(n9593), .ZN(n9596) );
  NAND2_X1 U10746 ( .A1(n9592), .A2(n9596), .ZN(n9599) );
  AOI222_X1 U10747 ( .A1(n9708), .A2(n9599), .B1(n9598), .B2(n9703), .C1(n9597), .C2(n9705), .ZN(n9788) );
  AOI21_X1 U10748 ( .B1(n9785), .B2(n5044), .A(n9600), .ZN(n9786) );
  INV_X1 U10749 ( .A(n9785), .ZN(n9604) );
  INV_X1 U10750 ( .A(n9601), .ZN(n9602) );
  AOI22_X1 U10751 ( .A1(n9712), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9602), .B2(
        n9710), .ZN(n9603) );
  OAI21_X1 U10752 ( .B1(n9604), .B2(n9714), .A(n9603), .ZN(n9609) );
  XOR2_X1 U10753 ( .A(n9606), .B(n9607), .Z(n9789) );
  NOR2_X1 U10754 ( .A1(n9789), .A2(n9716), .ZN(n9608) );
  AOI211_X1 U10755 ( .C1(n9786), .C2(n9700), .A(n9609), .B(n9608), .ZN(n9610)
         );
  OAI21_X1 U10756 ( .B1(n9788), .B2(n9694), .A(n9610), .ZN(P1_U3272) );
  NAND2_X1 U10757 ( .A1(n9612), .A2(n9611), .ZN(n9614) );
  INV_X1 U10758 ( .A(n9618), .ZN(n9613) );
  XNOR2_X1 U10759 ( .A(n9614), .B(n9613), .ZN(n9617) );
  OAI22_X1 U10760 ( .A1(n9615), .A2(n9656), .B1(n9657), .B2(n9654), .ZN(n9616)
         );
  AOI21_X1 U10761 ( .B1(n9617), .B2(n9708), .A(n9616), .ZN(n9795) );
  NAND2_X1 U10762 ( .A1(n9619), .A2(n9618), .ZN(n9620) );
  AND2_X1 U10763 ( .A1(n9621), .A2(n9620), .ZN(n9793) );
  AOI21_X1 U10764 ( .B1(n9640), .B2(n9624), .A(n10000), .ZN(n9622) );
  NAND2_X1 U10765 ( .A1(n9622), .A2(n5044), .ZN(n9790) );
  AOI22_X1 U10766 ( .A1(n9694), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9623), .B2(
        n9710), .ZN(n9626) );
  NAND2_X1 U10767 ( .A1(n9624), .A2(n9672), .ZN(n9625) );
  OAI211_X1 U10768 ( .C1(n9790), .C2(n9675), .A(n9626), .B(n9625), .ZN(n9627)
         );
  AOI21_X1 U10769 ( .B1(n9793), .B2(n9677), .A(n9627), .ZN(n9628) );
  OAI21_X1 U10770 ( .B1(n9795), .B2(n9694), .A(n9628), .ZN(P1_U3273) );
  XNOR2_X1 U10771 ( .A(n9629), .B(n9637), .ZN(n9630) );
  NAND2_X1 U10772 ( .A1(n9630), .A2(n9708), .ZN(n9635) );
  OAI22_X1 U10773 ( .A1(n9632), .A2(n9656), .B1(n9631), .B2(n9654), .ZN(n9633)
         );
  INV_X1 U10774 ( .A(n9633), .ZN(n9634) );
  NAND2_X1 U10775 ( .A1(n9635), .A2(n9634), .ZN(n9801) );
  INV_X1 U10776 ( .A(n9801), .ZN(n9648) );
  XNOR2_X1 U10777 ( .A(n9638), .B(n9637), .ZN(n9796) );
  OR2_X1 U10778 ( .A1(n9665), .A2(n9797), .ZN(n9639) );
  NAND2_X1 U10779 ( .A1(n9640), .A2(n9639), .ZN(n9798) );
  AOI22_X1 U10780 ( .A1(n9694), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9641), .B2(
        n9710), .ZN(n9644) );
  NAND2_X1 U10781 ( .A1(n9642), .A2(n9672), .ZN(n9643) );
  OAI211_X1 U10782 ( .C1(n9798), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9646)
         );
  AOI21_X1 U10783 ( .B1(n9796), .B2(n9677), .A(n9646), .ZN(n9647) );
  OAI21_X1 U10784 ( .B1(n9648), .B2(n9694), .A(n9647), .ZN(P1_U3274) );
  NAND2_X1 U10785 ( .A1(n9651), .A2(n9650), .ZN(n9652) );
  NAND2_X1 U10786 ( .A1(n9649), .A2(n9652), .ZN(n9653) );
  NAND2_X1 U10787 ( .A1(n9653), .A2(n9708), .ZN(n9660) );
  OAI22_X1 U10788 ( .A1(n9657), .A2(n9656), .B1(n9655), .B2(n9654), .ZN(n9658)
         );
  INV_X1 U10789 ( .A(n9658), .ZN(n9659) );
  NAND2_X1 U10790 ( .A1(n9660), .A2(n9659), .ZN(n9806) );
  INV_X1 U10791 ( .A(n9806), .ZN(n9679) );
  XNOR2_X1 U10792 ( .A(n9662), .B(n9663), .ZN(n9802) );
  NAND2_X1 U10793 ( .A1(n9691), .A2(n9673), .ZN(n9664) );
  NAND2_X1 U10794 ( .A1(n9664), .A2(n10008), .ZN(n9666) );
  OR2_X1 U10795 ( .A1(n9666), .A2(n9665), .ZN(n9803) );
  OAI22_X1 U10796 ( .A1(n9670), .A2(n9669), .B1(n9668), .B2(n9667), .ZN(n9671)
         );
  AOI21_X1 U10797 ( .B1(n9673), .B2(n9672), .A(n9671), .ZN(n9674) );
  OAI21_X1 U10798 ( .B1(n9803), .B2(n9675), .A(n9674), .ZN(n9676) );
  AOI21_X1 U10799 ( .B1(n9802), .B2(n9677), .A(n9676), .ZN(n9678) );
  OAI21_X1 U10800 ( .B1(n9679), .B2(n9694), .A(n9678), .ZN(P1_U3275) );
  INV_X1 U10801 ( .A(n9684), .ZN(n9680) );
  XNOR2_X1 U10802 ( .A(n9681), .B(n9680), .ZN(n9812) );
  OAI211_X1 U10803 ( .C1(n9684), .C2(n9683), .A(n9682), .B(n9708), .ZN(n9688)
         );
  AOI22_X1 U10804 ( .A1(n9686), .A2(n9703), .B1(n9705), .B2(n9685), .ZN(n9687)
         );
  OAI211_X1 U10805 ( .C1(n9812), .C2(n9689), .A(n9688), .B(n9687), .ZN(n9690)
         );
  INV_X1 U10806 ( .A(n9690), .ZN(n9810) );
  AOI21_X1 U10807 ( .B1(n9807), .B2(n9709), .A(n4443), .ZN(n9808) );
  INV_X1 U10808 ( .A(n9692), .ZN(n9693) );
  AOI22_X1 U10809 ( .A1(n9694), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9693), .B2(
        n9710), .ZN(n9695) );
  OAI21_X1 U10810 ( .B1(n9696), .B2(n9714), .A(n9695), .ZN(n9699) );
  NOR2_X1 U10811 ( .A1(n9812), .A2(n9697), .ZN(n9698) );
  AOI211_X1 U10812 ( .C1(n9808), .C2(n9700), .A(n9699), .B(n9698), .ZN(n9701)
         );
  OAI21_X1 U10813 ( .B1(n9810), .B2(n9712), .A(n9701), .ZN(P1_U3276) );
  XNOR2_X1 U10814 ( .A(n9702), .B(n4911), .ZN(n9707) );
  AOI222_X1 U10815 ( .A1(n9708), .A2(n9707), .B1(n9706), .B2(n9705), .C1(n9704), .C2(n9703), .ZN(n9816) );
  AOI211_X1 U10816 ( .C1(n4411), .C2(n4369), .A(n10000), .B(n4868), .ZN(n9813)
         );
  AOI22_X1 U10817 ( .A1(n9712), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9711), .B2(
        n9710), .ZN(n9713) );
  OAI21_X1 U10818 ( .B1(n4873), .B2(n9714), .A(n9713), .ZN(n9718) );
  XNOR2_X1 U10819 ( .A(n9715), .B(n4911), .ZN(n9817) );
  NOR2_X1 U10820 ( .A1(n9817), .A2(n9716), .ZN(n9717) );
  AOI211_X1 U10821 ( .C1(n9719), .C2(n9813), .A(n9718), .B(n9717), .ZN(n9720)
         );
  OAI21_X1 U10822 ( .B1(n9816), .B2(n9694), .A(n9720), .ZN(P1_U3277) );
  AOI21_X1 U10823 ( .B1(n9721), .B2(n9957), .A(n9724), .ZN(n9722) );
  OAI21_X1 U10824 ( .B1(n9723), .B2(n10000), .A(n9722), .ZN(n9828) );
  MUX2_X1 U10825 ( .A(n9828), .B(P1_REG1_REG_31__SCAN_IN), .S(n10026), .Z(
        P1_U3554) );
  AOI21_X1 U10826 ( .B1(n9725), .B2(n9957), .A(n9724), .ZN(n9726) );
  OAI21_X1 U10827 ( .B1(n9727), .B2(n10000), .A(n9726), .ZN(n9829) );
  MUX2_X1 U10828 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9829), .S(n10029), .Z(
        P1_U3553) );
  INV_X1 U10829 ( .A(n9728), .ZN(n9733) );
  OAI22_X1 U10830 ( .A1(n9730), .A2(n10000), .B1(n9729), .B2(n9998), .ZN(n9731) );
  OAI211_X1 U10831 ( .C1(n9734), .C2(n9961), .A(n9733), .B(n9732), .ZN(n9830)
         );
  MUX2_X1 U10832 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9830), .S(n10029), .Z(
        P1_U3552) );
  AOI21_X1 U10833 ( .B1(n9957), .B2(n9736), .A(n9735), .ZN(n9737) );
  MUX2_X1 U10834 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9831), .S(n10029), .Z(
        P1_U3551) );
  MUX2_X1 U10835 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9740), .S(n10029), .Z(
        P1_U3550) );
  MUX2_X1 U10836 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9832), .S(n10029), .Z(
        P1_U3549) );
  AOI211_X1 U10837 ( .C1(n9957), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9753)
         );
  OAI21_X1 U10838 ( .B1(n9961), .B2(n9754), .A(n9753), .ZN(n9833) );
  MUX2_X1 U10839 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9833), .S(n10029), .Z(
        P1_U3548) );
  INV_X1 U10840 ( .A(n9755), .ZN(n9757) );
  AOI211_X1 U10841 ( .C1(n9957), .C2(n9758), .A(n9757), .B(n9756), .ZN(n9759)
         );
  OAI21_X1 U10842 ( .B1(n9961), .B2(n9760), .A(n9759), .ZN(n9834) );
  MUX2_X1 U10843 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9834), .S(n10029), .Z(
        P1_U3547) );
  AOI22_X1 U10844 ( .A1(n9762), .A2(n10008), .B1(n9957), .B2(n9761), .ZN(n9763) );
  OAI211_X1 U10845 ( .C1(n9961), .C2(n9765), .A(n9764), .B(n9763), .ZN(n9835)
         );
  MUX2_X1 U10846 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9835), .S(n10029), .Z(
        P1_U3546) );
  OAI21_X1 U10847 ( .B1(n9961), .B2(n9770), .A(n9769), .ZN(n9836) );
  MUX2_X1 U10848 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9836), .S(n10029), .Z(
        P1_U3545) );
  OAI21_X1 U10849 ( .B1(n9772), .B2(n9998), .A(n9771), .ZN(n9773) );
  AOI21_X1 U10850 ( .B1(n9774), .B2(n10010), .A(n9773), .ZN(n9775) );
  AND2_X1 U10851 ( .A1(n9776), .A2(n9775), .ZN(n9837) );
  MUX2_X1 U10852 ( .A(n9777), .B(n9837), .S(n10029), .Z(n9778) );
  INV_X1 U10853 ( .A(n9778), .ZN(P1_U3544) );
  OAI22_X1 U10854 ( .A1(n9780), .A2(n10000), .B1(n9779), .B2(n9998), .ZN(n9781) );
  AOI21_X1 U10855 ( .B1(n9782), .B2(n10010), .A(n9781), .ZN(n9783) );
  NAND2_X1 U10856 ( .A1(n9784), .A2(n9783), .ZN(n9839) );
  MUX2_X1 U10857 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9839), .S(n10029), .Z(
        P1_U3543) );
  AOI22_X1 U10858 ( .A1(n9786), .A2(n10008), .B1(n9957), .B2(n9785), .ZN(n9787) );
  OAI211_X1 U10859 ( .C1(n9961), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9840)
         );
  MUX2_X1 U10860 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9840), .S(n10029), .Z(
        P1_U3542) );
  OAI21_X1 U10861 ( .B1(n9791), .B2(n9998), .A(n9790), .ZN(n9792) );
  AOI21_X1 U10862 ( .B1(n9793), .B2(n10010), .A(n9792), .ZN(n9794) );
  NAND2_X1 U10863 ( .A1(n9795), .A2(n9794), .ZN(n9841) );
  MUX2_X1 U10864 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9841), .S(n10029), .Z(
        P1_U3541) );
  AND2_X1 U10865 ( .A1(n9796), .A2(n10010), .ZN(n9800) );
  OAI22_X1 U10866 ( .A1(n9798), .A2(n10000), .B1(n9797), .B2(n9998), .ZN(n9799) );
  MUX2_X1 U10867 ( .A(n9842), .B(P1_REG1_REG_17__SCAN_IN), .S(n10026), .Z(
        P1_U3540) );
  NAND2_X1 U10868 ( .A1(n9802), .A2(n10010), .ZN(n9804) );
  OAI211_X1 U10869 ( .C1(n4442), .C2(n9998), .A(n9804), .B(n9803), .ZN(n9805)
         );
  MUX2_X1 U10870 ( .A(n9843), .B(P1_REG1_REG_16__SCAN_IN), .S(n10026), .Z(
        P1_U3539) );
  AOI22_X1 U10871 ( .A1(n9808), .A2(n10008), .B1(n9957), .B2(n9807), .ZN(n9809) );
  OAI211_X1 U10872 ( .C1(n9812), .C2(n9811), .A(n9810), .B(n9809), .ZN(n9844)
         );
  MUX2_X1 U10873 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9844), .S(n10029), .Z(
        P1_U3538) );
  AOI21_X1 U10874 ( .B1(n9957), .B2(n4411), .A(n9813), .ZN(n9815) );
  OAI211_X1 U10875 ( .C1(n9961), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9845)
         );
  MUX2_X1 U10876 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9845), .S(n10029), .Z(
        P1_U3537) );
  AOI22_X1 U10877 ( .A1(n9819), .A2(n10008), .B1(n9957), .B2(n9818), .ZN(n9820) );
  OAI211_X1 U10878 ( .C1(n9961), .C2(n9822), .A(n9821), .B(n9820), .ZN(n9846)
         );
  MUX2_X1 U10879 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9846), .S(n10029), .Z(
        P1_U3536) );
  AOI21_X1 U10880 ( .B1(n9957), .B2(n9824), .A(n9823), .ZN(n9825) );
  OAI211_X1 U10881 ( .C1(n9961), .C2(n9827), .A(n9826), .B(n9825), .ZN(n9847)
         );
  MUX2_X1 U10882 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9847), .S(n10029), .Z(
        P1_U3535) );
  MUX2_X1 U10883 ( .A(n9828), .B(P1_REG0_REG_31__SCAN_IN), .S(n10015), .Z(
        P1_U3522) );
  MUX2_X1 U10884 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9829), .S(n10017), .Z(
        P1_U3521) );
  MUX2_X1 U10885 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9830), .S(n10017), .Z(
        P1_U3520) );
  MUX2_X1 U10886 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9831), .S(n10017), .Z(
        P1_U3519) );
  MUX2_X1 U10887 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9832), .S(n10017), .Z(
        P1_U3517) );
  MUX2_X1 U10888 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9833), .S(n10017), .Z(
        P1_U3516) );
  MUX2_X1 U10889 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9834), .S(n10017), .Z(
        P1_U3515) );
  MUX2_X1 U10890 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9835), .S(n10017), .Z(
        P1_U3514) );
  MUX2_X1 U10891 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9836), .S(n10017), .Z(
        P1_U3513) );
  INV_X1 U10892 ( .A(n9837), .ZN(n9838) );
  MUX2_X1 U10893 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9838), .S(n10017), .Z(
        P1_U3512) );
  MUX2_X1 U10894 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9839), .S(n10017), .Z(
        P1_U3511) );
  MUX2_X1 U10895 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9840), .S(n10017), .Z(
        P1_U3510) );
  MUX2_X1 U10896 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9841), .S(n10017), .Z(
        P1_U3508) );
  MUX2_X1 U10897 ( .A(n9842), .B(P1_REG0_REG_17__SCAN_IN), .S(n10015), .Z(
        P1_U3505) );
  MUX2_X1 U10898 ( .A(n9843), .B(P1_REG0_REG_16__SCAN_IN), .S(n10015), .Z(
        P1_U3502) );
  MUX2_X1 U10899 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9844), .S(n10017), .Z(
        P1_U3499) );
  MUX2_X1 U10900 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9845), .S(n10017), .Z(
        P1_U3496) );
  MUX2_X1 U10901 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9846), .S(n10017), .Z(
        P1_U3493) );
  MUX2_X1 U10902 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9847), .S(n10017), .Z(
        P1_U3490) );
  NOR2_X1 U10903 ( .A1(n9849), .A2(n9848), .ZN(n9941) );
  MUX2_X1 U10904 ( .A(P1_D_REG_0__SCAN_IN), .B(n9850), .S(n9954), .Z(P1_U3440)
         );
  NOR4_X1 U10905 ( .A1(n5984), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5993), .ZN(n9851) );
  AOI21_X1 U10906 ( .B1(n9864), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9851), .ZN(
        n9852) );
  OAI21_X1 U10907 ( .B1(n9853), .B2(n9866), .A(n9852), .ZN(P1_U3322) );
  AOI22_X1 U10908 ( .A1(n9854), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9864), .ZN(n9855) );
  OAI21_X1 U10909 ( .B1(n9856), .B2(n9866), .A(n9855), .ZN(P1_U3323) );
  AOI22_X1 U10910 ( .A1(n4670), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9864), .ZN(n9857) );
  OAI21_X1 U10911 ( .B1(n9858), .B2(n9866), .A(n9857), .ZN(P1_U3324) );
  INV_X1 U10912 ( .A(n9859), .ZN(n9862) );
  AOI21_X1 U10913 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(n9864), .A(n9860), .ZN(
        n9861) );
  OAI21_X1 U10914 ( .B1(n9862), .B2(n9866), .A(n9861), .ZN(P1_U3325) );
  AOI21_X1 U10915 ( .B1(n9864), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9863), .ZN(
        n9865) );
  OAI21_X1 U10916 ( .B1(n9867), .B2(n9866), .A(n9865), .ZN(P1_U3326) );
  MUX2_X1 U10917 ( .A(n9868), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10918 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10276) );
  NOR2_X1 U10919 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9869) );
  AOI21_X1 U10920 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9869), .ZN(n10091) );
  NOR2_X1 U10921 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9870) );
  AOI21_X1 U10922 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9870), .ZN(n10094) );
  NOR2_X1 U10923 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9871) );
  AOI21_X1 U10924 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9871), .ZN(n10097) );
  NOR2_X1 U10925 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9872) );
  AOI21_X1 U10926 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9872), .ZN(n10100) );
  NOR2_X1 U10927 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9873) );
  AOI21_X1 U10928 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9873), .ZN(n10103) );
  NOR2_X1 U10929 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9880) );
  XOR2_X1 U10930 ( .A(n9874), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10289) );
  NAND2_X1 U10931 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9878) );
  XOR2_X1 U10932 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10287) );
  NAND2_X1 U10933 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9876) );
  XNOR2_X1 U10934 ( .A(n10195), .B(P1_ADDR_REG_2__SCAN_IN), .ZN(n10285) );
  AOI21_X1 U10935 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10085) );
  NAND3_X1 U10936 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10087) );
  OAI21_X1 U10937 ( .B1(n10085), .B2(n10219), .A(n10087), .ZN(n10284) );
  NAND2_X1 U10938 ( .A1(n10285), .A2(n10284), .ZN(n9875) );
  NAND2_X1 U10939 ( .A1(n9876), .A2(n9875), .ZN(n10286) );
  NAND2_X1 U10940 ( .A1(n10287), .A2(n10286), .ZN(n9877) );
  NAND2_X1 U10941 ( .A1(n9878), .A2(n9877), .ZN(n10288) );
  NOR2_X1 U10942 ( .A1(n10289), .A2(n10288), .ZN(n9879) );
  NOR2_X1 U10943 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9881), .ZN(n10271) );
  NAND2_X1 U10944 ( .A1(n9883), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U10945 ( .A1(n10269), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9884) );
  NAND2_X1 U10946 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9886), .ZN(n9889) );
  INV_X1 U10947 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U10948 ( .A1(n10273), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9888) );
  AND2_X1 U10949 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9890), .ZN(n9891) );
  INV_X1 U10950 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10279) );
  INV_X1 U10951 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10192) );
  NOR2_X1 U10952 ( .A1(n9892), .A2(n10192), .ZN(n9893) );
  INV_X1 U10953 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10283) );
  XOR2_X1 U10954 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9892), .Z(n10282) );
  NAND2_X1 U10955 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9894) );
  OAI21_X1 U10956 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9894), .ZN(n10111) );
  NAND2_X1 U10957 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9895) );
  OAI21_X1 U10958 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9895), .ZN(n10108) );
  NOR2_X1 U10959 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9896) );
  AOI21_X1 U10960 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9896), .ZN(n10105) );
  NAND2_X1 U10961 ( .A1(n10100), .A2(n10099), .ZN(n10098) );
  NAND2_X1 U10962 ( .A1(n10094), .A2(n10093), .ZN(n10092) );
  OAI21_X1 U10963 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10092), .ZN(n10090) );
  NAND2_X1 U10964 ( .A1(n10091), .A2(n10090), .ZN(n10089) );
  OAI21_X2 U10965 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10089), .ZN(n10275) );
  NOR2_X1 U10966 ( .A1(n10276), .A2(n10275), .ZN(n9897) );
  NAND2_X1 U10967 ( .A1(n10276), .A2(n10275), .ZN(n10274) );
  XNOR2_X1 U10968 ( .A(n9898), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n9899) );
  XNOR2_X1 U10969 ( .A(n9900), .B(n9899), .ZN(ADD_1071_U4) );
  INV_X1 U10970 ( .A(n9901), .ZN(n9903) );
  OAI22_X1 U10971 ( .A1(n9903), .A2(n10000), .B1(n9902), .B2(n9998), .ZN(n9906) );
  INV_X1 U10972 ( .A(n9904), .ZN(n9905) );
  AOI211_X1 U10973 ( .C1(n9907), .C2(n10010), .A(n9906), .B(n9905), .ZN(n9910)
         );
  AOI22_X1 U10974 ( .A1(n10029), .A2(n9910), .B1(n9908), .B2(n10026), .ZN(
        P1_U3534) );
  INV_X1 U10975 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U10976 ( .A1(n10017), .A2(n9910), .B1(n9909), .B2(n10015), .ZN(
        P1_U3487) );
  INV_X1 U10977 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10237) );
  XOR2_X1 U10978 ( .A(n10237), .B(P2_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U10979 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10980 ( .A(n9911), .ZN(n9919) );
  OAI211_X1 U10981 ( .C1(n9915), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9917)
         );
  OAI211_X1 U10982 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9920)
         );
  INV_X1 U10983 ( .A(n9920), .ZN(n9929) );
  NAND2_X1 U10984 ( .A1(n9922), .A2(n9921), .ZN(n9924) );
  AOI21_X1 U10985 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9926) );
  AOI21_X1 U10986 ( .B1(n9927), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9926), .ZN(
        n9928) );
  NAND2_X1 U10987 ( .A1(n9929), .A2(n9928), .ZN(P1_U3259) );
  INV_X1 U10988 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9930) );
  NOR2_X1 U10989 ( .A1(n9941), .A2(n9930), .ZN(P1_U3292) );
  INV_X1 U10990 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10173) );
  NOR2_X1 U10991 ( .A1(n9941), .A2(n10173), .ZN(P1_U3293) );
  INV_X1 U10992 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9931) );
  NOR2_X1 U10993 ( .A1(n9954), .A2(n9931), .ZN(P1_U3294) );
  INV_X1 U10994 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U10995 ( .A1(n9954), .A2(n9932), .ZN(P1_U3295) );
  INV_X1 U10996 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9933) );
  NOR2_X1 U10997 ( .A1(n9954), .A2(n9933), .ZN(P1_U3296) );
  INV_X1 U10998 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9934) );
  NOR2_X1 U10999 ( .A1(n9954), .A2(n9934), .ZN(P1_U3297) );
  INV_X1 U11000 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9935) );
  NOR2_X1 U11001 ( .A1(n9954), .A2(n9935), .ZN(P1_U3298) );
  INV_X1 U11002 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U11003 ( .A1(n9954), .A2(n10222), .ZN(P1_U3299) );
  INV_X1 U11004 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U11005 ( .A1(n9954), .A2(n10208), .ZN(P1_U3300) );
  INV_X1 U11006 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9936) );
  NOR2_X1 U11007 ( .A1(n9941), .A2(n9936), .ZN(P1_U3301) );
  INV_X1 U11008 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9937) );
  NOR2_X1 U11009 ( .A1(n9941), .A2(n9937), .ZN(P1_U3302) );
  INV_X1 U11010 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10253) );
  NOR2_X1 U11011 ( .A1(n9941), .A2(n10253), .ZN(P1_U3303) );
  INV_X1 U11012 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10228) );
  NOR2_X1 U11013 ( .A1(n9941), .A2(n10228), .ZN(P1_U3304) );
  INV_X1 U11014 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9938) );
  NOR2_X1 U11015 ( .A1(n9941), .A2(n9938), .ZN(P1_U3305) );
  INV_X1 U11016 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9939) );
  NOR2_X1 U11017 ( .A1(n9941), .A2(n9939), .ZN(P1_U3306) );
  INV_X1 U11018 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10162) );
  NOR2_X1 U11019 ( .A1(n9941), .A2(n10162), .ZN(P1_U3307) );
  INV_X1 U11020 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9940) );
  NOR2_X1 U11021 ( .A1(n9941), .A2(n9940), .ZN(P1_U3308) );
  INV_X1 U11022 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9942) );
  NOR2_X1 U11023 ( .A1(n9954), .A2(n9942), .ZN(P1_U3309) );
  INV_X1 U11024 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9943) );
  NOR2_X1 U11025 ( .A1(n9954), .A2(n9943), .ZN(P1_U3310) );
  INV_X1 U11026 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9944) );
  NOR2_X1 U11027 ( .A1(n9954), .A2(n9944), .ZN(P1_U3311) );
  INV_X1 U11028 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9945) );
  NOR2_X1 U11029 ( .A1(n9954), .A2(n9945), .ZN(P1_U3312) );
  INV_X1 U11030 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10255) );
  NOR2_X1 U11031 ( .A1(n9954), .A2(n10255), .ZN(P1_U3313) );
  INV_X1 U11032 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9946) );
  NOR2_X1 U11033 ( .A1(n9954), .A2(n9946), .ZN(P1_U3314) );
  INV_X1 U11034 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9947) );
  NOR2_X1 U11035 ( .A1(n9954), .A2(n9947), .ZN(P1_U3315) );
  INV_X1 U11036 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9948) );
  NOR2_X1 U11037 ( .A1(n9954), .A2(n9948), .ZN(P1_U3316) );
  INV_X1 U11038 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9949) );
  NOR2_X1 U11039 ( .A1(n9954), .A2(n9949), .ZN(P1_U3317) );
  INV_X1 U11040 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9950) );
  NOR2_X1 U11041 ( .A1(n9954), .A2(n9950), .ZN(P1_U3318) );
  INV_X1 U11042 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9951) );
  NOR2_X1 U11043 ( .A1(n9954), .A2(n9951), .ZN(P1_U3319) );
  INV_X1 U11044 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9952) );
  NOR2_X1 U11045 ( .A1(n9954), .A2(n9952), .ZN(P1_U3320) );
  INV_X1 U11046 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9953) );
  NOR2_X1 U11047 ( .A1(n9954), .A2(n9953), .ZN(P1_U3321) );
  AOI21_X1 U11048 ( .B1(n9957), .B2(n9956), .A(n9955), .ZN(n9958) );
  OAI211_X1 U11049 ( .C1(n9961), .C2(n9960), .A(n9959), .B(n9958), .ZN(n9962)
         );
  INV_X1 U11050 ( .A(n9962), .ZN(n10018) );
  INV_X1 U11051 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U11052 ( .A1(n10017), .A2(n10018), .B1(n10224), .B2(n10015), .ZN(
        P1_U3457) );
  INV_X1 U11053 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U11054 ( .A1(n10017), .A2(n9964), .B1(n9963), .B2(n10015), .ZN(
        P1_U3460) );
  INV_X1 U11055 ( .A(n9965), .ZN(n9969) );
  OAI22_X1 U11056 ( .A1(n9966), .A2(n10000), .B1(n4860), .B2(n9998), .ZN(n9968) );
  AOI211_X1 U11057 ( .C1(n10005), .C2(n9969), .A(n9968), .B(n9967), .ZN(n10019) );
  INV_X1 U11058 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11059 ( .A1(n10017), .A2(n10019), .B1(n9970), .B2(n10015), .ZN(
        P1_U3463) );
  INV_X1 U11060 ( .A(n9971), .ZN(n9976) );
  OAI22_X1 U11061 ( .A1(n9973), .A2(n10000), .B1(n9972), .B2(n9998), .ZN(n9975) );
  AOI211_X1 U11062 ( .C1(n10005), .C2(n9976), .A(n9975), .B(n9974), .ZN(n10020) );
  INV_X1 U11063 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U11064 ( .A1(n10017), .A2(n10020), .B1(n9977), .B2(n10015), .ZN(
        P1_U3466) );
  NAND3_X1 U11065 ( .A1(n9979), .A2(n10010), .A3(n9978), .ZN(n9981) );
  OAI211_X1 U11066 ( .C1(n9982), .C2(n9998), .A(n9981), .B(n9980), .ZN(n9983)
         );
  NOR2_X1 U11067 ( .A1(n9984), .A2(n9983), .ZN(n10021) );
  INV_X1 U11068 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U11069 ( .A1(n10017), .A2(n10021), .B1(n9985), .B2(n10015), .ZN(
        P1_U3469) );
  INV_X1 U11070 ( .A(n9986), .ZN(n9990) );
  OAI22_X1 U11071 ( .A1(n9987), .A2(n10000), .B1(n4520), .B2(n9998), .ZN(n9989) );
  AOI211_X1 U11072 ( .C1(n10005), .C2(n9990), .A(n9989), .B(n9988), .ZN(n10022) );
  INV_X1 U11073 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U11074 ( .A1(n10017), .A2(n10022), .B1(n9991), .B2(n10015), .ZN(
        P1_U3472) );
  OAI211_X1 U11075 ( .C1(n9994), .C2(n9998), .A(n9993), .B(n9992), .ZN(n9995)
         );
  AOI21_X1 U11076 ( .B1(n10010), .B2(n9996), .A(n9995), .ZN(n10024) );
  INV_X1 U11077 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9997) );
  AOI22_X1 U11078 ( .A1(n10017), .A2(n10024), .B1(n9997), .B2(n10015), .ZN(
        P1_U3475) );
  OAI22_X1 U11079 ( .A1(n10001), .A2(n10000), .B1(n9999), .B2(n9998), .ZN(
        n10003) );
  AOI211_X1 U11080 ( .C1(n10005), .C2(n10004), .A(n10003), .B(n10002), .ZN(
        n10025) );
  INV_X1 U11081 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10006) );
  AOI22_X1 U11082 ( .A1(n10017), .A2(n10025), .B1(n10006), .B2(n10015), .ZN(
        P1_U3478) );
  AOI21_X1 U11083 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(n10013) );
  NAND2_X1 U11084 ( .A1(n10011), .A2(n10010), .ZN(n10012) );
  AND3_X1 U11085 ( .A1(n10014), .A2(n10013), .A3(n10012), .ZN(n10028) );
  INV_X1 U11086 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10016) );
  AOI22_X1 U11087 ( .A1(n10017), .A2(n10028), .B1(n10016), .B2(n10015), .ZN(
        P1_U3481) );
  AOI22_X1 U11088 ( .A1(n10029), .A2(n10018), .B1(n6511), .B2(n10026), .ZN(
        P1_U3524) );
  AOI22_X1 U11089 ( .A1(n10029), .A2(n10019), .B1(n6514), .B2(n10026), .ZN(
        P1_U3526) );
  AOI22_X1 U11090 ( .A1(n10029), .A2(n10020), .B1(n6515), .B2(n10026), .ZN(
        P1_U3527) );
  AOI22_X1 U11091 ( .A1(n10029), .A2(n10021), .B1(n6516), .B2(n10026), .ZN(
        P1_U3528) );
  AOI22_X1 U11092 ( .A1(n10029), .A2(n10022), .B1(n10116), .B2(n10026), .ZN(
        P1_U3529) );
  INV_X1 U11093 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10023) );
  AOI22_X1 U11094 ( .A1(n10029), .A2(n10024), .B1(n10023), .B2(n10026), .ZN(
        P1_U3530) );
  AOI22_X1 U11095 ( .A1(n10029), .A2(n10025), .B1(n6542), .B2(n10026), .ZN(
        P1_U3531) );
  INV_X1 U11096 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10027) );
  AOI22_X1 U11097 ( .A1(n10029), .A2(n10028), .B1(n10027), .B2(n10026), .ZN(
        P1_U3532) );
  AND2_X1 U11098 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n4271), .ZN(P2_U3297) );
  AND2_X1 U11099 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n4271), .ZN(P2_U3298) );
  AND2_X1 U11100 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n4271), .ZN(P2_U3299) );
  AND2_X1 U11101 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n4271), .ZN(P2_U3300) );
  AND2_X1 U11102 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n4271), .ZN(P2_U3301) );
  AND2_X1 U11103 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n4271), .ZN(P2_U3302) );
  AND2_X1 U11104 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n4271), .ZN(P2_U3303) );
  AND2_X1 U11105 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n4271), .ZN(P2_U3304) );
  AND2_X1 U11106 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n4271), .ZN(P2_U3305) );
  AND2_X1 U11107 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n4271), .ZN(P2_U3306) );
  AND2_X1 U11108 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n4271), .ZN(P2_U3307) );
  AND2_X1 U11109 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n4271), .ZN(P2_U3308) );
  AND2_X1 U11110 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n4271), .ZN(P2_U3309) );
  AND2_X1 U11111 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n4271), .ZN(P2_U3311) );
  AND2_X1 U11112 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n4271), .ZN(P2_U3312) );
  AND2_X1 U11113 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n4271), .ZN(P2_U3313) );
  AND2_X1 U11114 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n4271), .ZN(P2_U3314) );
  AND2_X1 U11115 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n4271), .ZN(P2_U3315) );
  AND2_X1 U11116 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n4271), .ZN(P2_U3316) );
  AND2_X1 U11117 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n4271), .ZN(P2_U3317) );
  AND2_X1 U11118 ( .A1(n4271), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3318) );
  AND2_X1 U11119 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n4271), .ZN(P2_U3319) );
  AND2_X1 U11120 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n4271), .ZN(P2_U3320) );
  AND2_X1 U11121 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n4271), .ZN(P2_U3321) );
  AND2_X1 U11122 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n4271), .ZN(P2_U3322) );
  AND2_X1 U11123 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n4271), .ZN(P2_U3323) );
  AND2_X1 U11124 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n4271), .ZN(P2_U3324) );
  AND2_X1 U11125 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n4271), .ZN(P2_U3325) );
  AND2_X1 U11126 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n4271), .ZN(P2_U3326) );
  INV_X1 U11127 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10034) );
  AOI22_X1 U11128 ( .A1(n10034), .A2(n4271), .B1(n10037), .B2(n10033), .ZN(
        P2_U3437) );
  AOI22_X1 U11129 ( .A1(n10037), .A2(n10036), .B1(n10035), .B2(n4271), .ZN(
        P2_U3438) );
  INV_X1 U11130 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U11131 ( .A1(n10076), .A2(n10039), .B1(n10038), .B2(n10074), .ZN(
        P2_U3451) );
  INV_X1 U11132 ( .A(n10040), .ZN(n10042) );
  INV_X1 U11133 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U11134 ( .A1(n10076), .A2(n10042), .B1(n10041), .B2(n10074), .ZN(
        P2_U3457) );
  OAI22_X1 U11135 ( .A1(n10044), .A2(n10052), .B1(n10043), .B2(n10070), .ZN(
        n10045) );
  INV_X1 U11136 ( .A(n10045), .ZN(n10048) );
  NAND2_X1 U11137 ( .A1(n10046), .A2(n10066), .ZN(n10047) );
  AND3_X1 U11138 ( .A1(n10049), .A2(n10048), .A3(n10047), .ZN(n10077) );
  INV_X1 U11139 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U11140 ( .A1(n10076), .A2(n10077), .B1(n10146), .B2(n10074), .ZN(
        P2_U3463) );
  INV_X1 U11141 ( .A(n10050), .ZN(n10057) );
  OAI22_X1 U11142 ( .A1(n10053), .A2(n10052), .B1(n10051), .B2(n10070), .ZN(
        n10056) );
  INV_X1 U11143 ( .A(n10054), .ZN(n10055) );
  AOI211_X1 U11144 ( .C1(n10066), .C2(n10057), .A(n10056), .B(n10055), .ZN(
        n10079) );
  INV_X1 U11145 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10058) );
  AOI22_X1 U11146 ( .A1(n10076), .A2(n10079), .B1(n10058), .B2(n10074), .ZN(
        P2_U3469) );
  INV_X1 U11147 ( .A(n10059), .ZN(n10065) );
  OAI21_X1 U11148 ( .B1(n10061), .B2(n10070), .A(n10060), .ZN(n10064) );
  INV_X1 U11149 ( .A(n10062), .ZN(n10063) );
  AOI211_X1 U11150 ( .C1(n10066), .C2(n10065), .A(n10064), .B(n10063), .ZN(
        n10080) );
  INV_X1 U11151 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U11152 ( .A1(n10076), .A2(n10080), .B1(n10254), .B2(n10074), .ZN(
        P2_U3472) );
  NAND3_X1 U11153 ( .A1(n7655), .A2(n10067), .A3(n10066), .ZN(n10069) );
  OAI211_X1 U11154 ( .C1(n10071), .C2(n10070), .A(n10069), .B(n10068), .ZN(
        n10072) );
  NOR2_X1 U11155 ( .A1(n10073), .A2(n10072), .ZN(n10083) );
  INV_X1 U11156 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10075) );
  AOI22_X1 U11157 ( .A1(n10076), .A2(n10083), .B1(n10075), .B2(n10074), .ZN(
        P2_U3475) );
  AOI22_X1 U11158 ( .A1(n10084), .A2(n10077), .B1(n6827), .B2(n10081), .ZN(
        P2_U3524) );
  INV_X1 U11159 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10078) );
  AOI22_X1 U11160 ( .A1(n10084), .A2(n10079), .B1(n10078), .B2(n10081), .ZN(
        P2_U3526) );
  AOI22_X1 U11161 ( .A1(n10084), .A2(n10080), .B1(n6846), .B2(n10081), .ZN(
        P2_U3527) );
  INV_X1 U11162 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U11163 ( .A1(n10084), .A2(n10083), .B1(n10082), .B2(n10081), .ZN(
        P2_U3528) );
  INV_X1 U11164 ( .A(n10085), .ZN(n10086) );
  NAND2_X1 U11165 ( .A1(n10087), .A2(n10086), .ZN(n10088) );
  XOR2_X1 U11166 ( .A(n10219), .B(n10088), .Z(ADD_1071_U5) );
  XOR2_X1 U11167 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11168 ( .B1(n10091), .B2(n10090), .A(n10089), .ZN(ADD_1071_U56) );
  OAI21_X1 U11169 ( .B1(n10094), .B2(n10093), .A(n10092), .ZN(ADD_1071_U57) );
  OAI21_X1 U11170 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(ADD_1071_U58) );
  OAI21_X1 U11171 ( .B1(n10100), .B2(n10099), .A(n10098), .ZN(ADD_1071_U59) );
  OAI21_X1 U11172 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(ADD_1071_U60) );
  OAI21_X1 U11173 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(ADD_1071_U61) );
  AOI21_X1 U11174 ( .B1(n10109), .B2(n10108), .A(n10107), .ZN(ADD_1071_U62) );
  AOI21_X1 U11175 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(ADD_1071_U63) );
  NAND2_X1 U11176 ( .A1(n4271), .A2(P2_D_REG_18__SCAN_IN), .ZN(n10268) );
  NOR4_X1 U11177 ( .A1(SI_17_), .A2(P1_REG2_REG_24__SCAN_IN), .A3(
        P1_REG0_REG_20__SCAN_IN), .A4(n10194), .ZN(n10115) );
  NOR3_X1 U11178 ( .A1(SI_11_), .A2(P2_REG0_REG_28__SCAN_IN), .A3(n10197), 
        .ZN(n10114) );
  NOR4_X1 U11179 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_REG0_REG_1__SCAN_IN), 
        .A3(P2_REG2_REG_1__SCAN_IN), .A4(n7372), .ZN(n10113) );
  NAND4_X1 U11180 ( .A1(SI_14_), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(
        n10128) );
  NAND4_X1 U11181 ( .A1(n10236), .A2(SI_5_), .A3(SI_27_), .A4(
        P1_REG3_REG_15__SCAN_IN), .ZN(n10127) );
  NAND4_X1 U11182 ( .A1(n10117), .A2(n10116), .A3(n10254), .A4(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10126) );
  NAND4_X1 U11183 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_DATAO_REG_19__SCAN_IN), 
        .A3(P2_D_REG_10__SCAN_IN), .A4(P2_REG1_REG_14__SCAN_IN), .ZN(n10124)
         );
  INV_X1 U11184 ( .A(n10238), .ZN(n10122) );
  INV_X1 U11185 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10121) );
  INV_X1 U11186 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10118) );
  NOR3_X1 U11187 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(n10118), .A3(n6876), .ZN(
        n10119) );
  NAND4_X1 U11188 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10123) );
  OR4_X1 U11189 ( .A1(n10124), .A2(n10123), .A3(P1_D_REG_23__SCAN_IN), .A4(
        n10237), .ZN(n10125) );
  NOR4_X1 U11190 ( .A1(n10128), .A2(n10127), .A3(n10126), .A4(n10125), .ZN(
        n10266) );
  NAND4_X1 U11191 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .A3(n10192), .A4(n10219), .ZN(n10142) );
  NAND4_X1 U11192 ( .A1(n10157), .A2(n10130), .A3(P2_IR_REG_4__SCAN_IN), .A4(
        P2_IR_REG_20__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U11193 ( .A1(n10174), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n10131) );
  INV_X1 U11194 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10163) );
  NOR4_X1 U11195 ( .A1(n10132), .A2(n10131), .A3(P2_IR_REG_19__SCAN_IN), .A4(
        n10163), .ZN(n10133) );
  NAND2_X1 U11196 ( .A1(n10134), .A2(n10133), .ZN(n10141) );
  NAND4_X1 U11197 ( .A1(P2_REG0_REG_4__SCAN_IN), .A2(P2_REG2_REG_24__SCAN_IN), 
        .A3(n10149), .A4(n10148), .ZN(n10140) );
  NOR3_X1 U11198 ( .A1(SI_6_), .A2(P1_REG2_REG_23__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n10136) );
  INV_X1 U11199 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10172) );
  INV_X1 U11200 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10171) );
  NOR4_X1 U11201 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .A3(n10172), .A4(n10171), .ZN(n10135) );
  AND4_X1 U11202 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(
        P2_REG2_REG_6__SCAN_IN), .ZN(n10138) );
  NAND4_X1 U11203 ( .A1(n10138), .A2(P2_DATAO_REG_5__SCAN_IN), .A3(
        P1_REG2_REG_5__SCAN_IN), .A4(n10144), .ZN(n10139) );
  NOR4_X1 U11204 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n10265) );
  AOI22_X1 U11205 ( .A1(n5606), .A2(keyinput61), .B1(n10144), .B2(keyinput62), 
        .ZN(n10143) );
  OAI221_X1 U11206 ( .B1(n5606), .B2(keyinput61), .C1(n10144), .C2(keyinput62), 
        .A(n10143), .ZN(n10155) );
  AOI22_X1 U11207 ( .A1(n7290), .A2(keyinput32), .B1(keyinput8), .B2(n10146), 
        .ZN(n10145) );
  OAI221_X1 U11208 ( .B1(n7290), .B2(keyinput32), .C1(n10146), .C2(keyinput8), 
        .A(n10145), .ZN(n10154) );
  AOI22_X1 U11209 ( .A1(n10149), .A2(keyinput18), .B1(keyinput37), .B2(n10148), 
        .ZN(n10147) );
  OAI221_X1 U11210 ( .B1(n10149), .B2(keyinput18), .C1(n10148), .C2(keyinput37), .A(n10147), .ZN(n10153) );
  XOR2_X1 U11211 ( .A(n6261), .B(keyinput27), .Z(n10151) );
  XNOR2_X1 U11212 ( .A(SI_6_), .B(keyinput53), .ZN(n10150) );
  NAND2_X1 U11213 ( .A1(n10151), .A2(n10150), .ZN(n10152) );
  NOR4_X1 U11214 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10206) );
  INV_X1 U11215 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U11216 ( .A1(n10158), .A2(keyinput51), .B1(keyinput56), .B2(n10157), 
        .ZN(n10156) );
  OAI221_X1 U11217 ( .B1(n10158), .B2(keyinput51), .C1(n10157), .C2(keyinput56), .A(n10156), .ZN(n10161) );
  XOR2_X1 U11218 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput55), .Z(n10160) );
  XNOR2_X1 U11219 ( .A(keyinput35), .B(n7441), .ZN(n10159) );
  OR3_X1 U11220 ( .A1(n10161), .A2(n10160), .A3(n10159), .ZN(n10169) );
  XNOR2_X1 U11221 ( .A(n10162), .B(keyinput38), .ZN(n10168) );
  XNOR2_X1 U11222 ( .A(keyinput2), .B(n10163), .ZN(n10167) );
  XNOR2_X1 U11223 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput7), .ZN(n10165) );
  XNOR2_X1 U11224 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput28), .ZN(n10164) );
  NAND2_X1 U11225 ( .A1(n10165), .A2(n10164), .ZN(n10166) );
  NOR4_X1 U11226 ( .A1(n10169), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n10205) );
  AOI22_X1 U11227 ( .A1(n10172), .A2(keyinput21), .B1(keyinput12), .B2(n10171), 
        .ZN(n10170) );
  OAI221_X1 U11228 ( .B1(n10172), .B2(keyinput21), .C1(n10171), .C2(keyinput12), .A(n10170), .ZN(n10177) );
  XNOR2_X1 U11229 ( .A(n10173), .B(keyinput26), .ZN(n10176) );
  XNOR2_X1 U11230 ( .A(n10174), .B(keyinput31), .ZN(n10175) );
  OR3_X1 U11231 ( .A1(n10177), .A2(n10176), .A3(n10175), .ZN(n10186) );
  INV_X1 U11232 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U11233 ( .A1(n10180), .A2(keyinput63), .B1(keyinput57), .B2(n10179), 
        .ZN(n10178) );
  OAI221_X1 U11234 ( .B1(n10180), .B2(keyinput63), .C1(n10179), .C2(keyinput57), .A(n10178), .ZN(n10185) );
  AOI22_X1 U11235 ( .A1(n10183), .A2(keyinput48), .B1(keyinput14), .B2(n10182), 
        .ZN(n10181) );
  OAI221_X1 U11236 ( .B1(n10183), .B2(keyinput48), .C1(n10182), .C2(keyinput14), .A(n10181), .ZN(n10184) );
  NOR3_X1 U11237 ( .A1(n10186), .A2(n10185), .A3(n10184), .ZN(n10204) );
  AOI22_X1 U11238 ( .A1(n10189), .A2(keyinput29), .B1(n10188), .B2(keyinput16), 
        .ZN(n10187) );
  OAI221_X1 U11239 ( .B1(n10189), .B2(keyinput29), .C1(n10188), .C2(keyinput16), .A(n10187), .ZN(n10202) );
  AOI22_X1 U11240 ( .A1(n10192), .A2(keyinput0), .B1(n10191), .B2(keyinput59), 
        .ZN(n10190) );
  OAI221_X1 U11241 ( .B1(n10192), .B2(keyinput0), .C1(n10191), .C2(keyinput59), 
        .A(n10190), .ZN(n10201) );
  AOI22_X1 U11242 ( .A1(n10195), .A2(keyinput22), .B1(n10194), .B2(keyinput1), 
        .ZN(n10193) );
  OAI221_X1 U11243 ( .B1(n10195), .B2(keyinput22), .C1(n10194), .C2(keyinput1), 
        .A(n10193), .ZN(n10200) );
  INV_X1 U11244 ( .A(SI_14_), .ZN(n10198) );
  AOI22_X1 U11245 ( .A1(n10198), .A2(keyinput4), .B1(n10197), .B2(keyinput6), 
        .ZN(n10196) );
  OAI221_X1 U11246 ( .B1(n10198), .B2(keyinput4), .C1(n10197), .C2(keyinput6), 
        .A(n10196), .ZN(n10199) );
  NOR4_X1 U11247 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10203) );
  NAND4_X1 U11248 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10264) );
  AOI22_X1 U11249 ( .A1(n10116), .A2(keyinput10), .B1(n10208), .B2(keyinput45), 
        .ZN(n10207) );
  OAI221_X1 U11250 ( .B1(n10116), .B2(keyinput10), .C1(n10208), .C2(keyinput45), .A(n10207), .ZN(n10217) );
  AOI22_X1 U11251 ( .A1(n10283), .A2(keyinput23), .B1(n6876), .B2(keyinput24), 
        .ZN(n10209) );
  OAI221_X1 U11252 ( .B1(n10283), .B2(keyinput23), .C1(n6876), .C2(keyinput24), 
        .A(n10209), .ZN(n10216) );
  AOI22_X1 U11253 ( .A1(n7372), .A2(keyinput44), .B1(n10211), .B2(keyinput3), 
        .ZN(n10210) );
  OAI221_X1 U11254 ( .B1(n7372), .B2(keyinput44), .C1(n10211), .C2(keyinput3), 
        .A(n10210), .ZN(n10215) );
  XNOR2_X1 U11255 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput47), .ZN(n10213) );
  XNOR2_X1 U11256 ( .A(P1_REG0_REG_24__SCAN_IN), .B(keyinput17), .ZN(n10212)
         );
  NAND2_X1 U11257 ( .A1(n10213), .A2(n10212), .ZN(n10214) );
  NOR4_X1 U11258 ( .A1(n10217), .A2(n10216), .A3(n10215), .A4(n10214), .ZN(
        n10262) );
  INV_X1 U11259 ( .A(SI_11_), .ZN(n10220) );
  AOI22_X1 U11260 ( .A1(n10220), .A2(keyinput33), .B1(keyinput46), .B2(n10219), 
        .ZN(n10218) );
  OAI221_X1 U11261 ( .B1(n10220), .B2(keyinput33), .C1(n10219), .C2(keyinput46), .A(n10218), .ZN(n10232) );
  AOI22_X1 U11262 ( .A1(n10223), .A2(keyinput25), .B1(n10222), .B2(keyinput5), 
        .ZN(n10221) );
  OAI221_X1 U11263 ( .B1(n10223), .B2(keyinput25), .C1(n10222), .C2(keyinput5), 
        .A(n10221), .ZN(n10231) );
  XOR2_X1 U11264 ( .A(n10224), .B(keyinput60), .Z(n10227) );
  XNOR2_X1 U11265 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput42), .ZN(n10226) );
  XNOR2_X1 U11266 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput41), .ZN(n10225) );
  NAND3_X1 U11267 ( .A1(n10227), .A2(n10226), .A3(n10225), .ZN(n10230) );
  XNOR2_X1 U11268 ( .A(n10228), .B(keyinput40), .ZN(n10229) );
  NOR4_X1 U11269 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        n10261) );
  AOI22_X1 U11270 ( .A1(n10117), .A2(keyinput9), .B1(n10234), .B2(keyinput50), 
        .ZN(n10233) );
  OAI221_X1 U11271 ( .B1(n10117), .B2(keyinput9), .C1(n10234), .C2(keyinput50), 
        .A(n10233), .ZN(n10245) );
  AOI22_X1 U11272 ( .A1(P2_U3152), .A2(keyinput13), .B1(n10236), .B2(
        keyinput11), .ZN(n10235) );
  OAI221_X1 U11273 ( .B1(P2_U3152), .B2(keyinput13), .C1(n10236), .C2(
        keyinput11), .A(n10235), .ZN(n10244) );
  XOR2_X1 U11274 ( .A(n10237), .B(keyinput43), .Z(n10242) );
  XNOR2_X1 U11275 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput30), .ZN(n10241) );
  XNOR2_X1 U11276 ( .A(n10238), .B(keyinput20), .ZN(n10240) );
  XNOR2_X1 U11277 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput58), .ZN(n10239) );
  NAND4_X1 U11278 ( .A1(n10242), .A2(n10241), .A3(n10240), .A4(n10239), .ZN(
        n10243) );
  NOR3_X1 U11279 ( .A1(n10245), .A2(n10244), .A3(n10243), .ZN(n10260) );
  XOR2_X1 U11280 ( .A(SI_5_), .B(keyinput15), .Z(n10248) );
  XOR2_X1 U11281 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput52), .Z(n10247) );
  XNOR2_X1 U11282 ( .A(n5272), .B(keyinput19), .ZN(n10246) );
  NOR3_X1 U11283 ( .A1(n10248), .A2(n10247), .A3(n10246), .ZN(n10251) );
  XNOR2_X1 U11284 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput54), .ZN(n10250) );
  XNOR2_X1 U11285 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput36), .ZN(n10249)
         );
  NAND3_X1 U11286 ( .A1(n10251), .A2(n10250), .A3(n10249), .ZN(n10258) );
  AOI22_X1 U11287 ( .A1(n10254), .A2(keyinput34), .B1(n10253), .B2(keyinput49), 
        .ZN(n10252) );
  OAI221_X1 U11288 ( .B1(n10254), .B2(keyinput34), .C1(n10253), .C2(keyinput49), .A(n10252), .ZN(n10257) );
  XNOR2_X1 U11289 ( .A(n10255), .B(keyinput39), .ZN(n10256) );
  NOR3_X1 U11290 ( .A1(n10258), .A2(n10257), .A3(n10256), .ZN(n10259) );
  NAND4_X1 U11291 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10263) );
  AOI211_X1 U11292 ( .C1(n10266), .C2(n10265), .A(n10264), .B(n10263), .ZN(
        n10267) );
  XNOR2_X1 U11293 ( .A(n10268), .B(n10267), .ZN(P2_U3310) );
  XOR2_X1 U11294 ( .A(n10269), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11295 ( .A1(n10271), .A2(n10270), .ZN(n10272) );
  XOR2_X1 U11296 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10272), .Z(ADD_1071_U51) );
  XOR2_X1 U11297 ( .A(n10273), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11298 ( .B1(n10276), .B2(n10275), .A(n10274), .ZN(n10277) );
  XNOR2_X1 U11299 ( .A(n10277), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11300 ( .B1(n10280), .B2(n10279), .A(n10278), .ZN(ADD_1071_U48) );
  AOI21_X1 U11301 ( .B1(n10283), .B2(n10282), .A(n10281), .ZN(ADD_1071_U47) );
  XOR2_X1 U11302 ( .A(n10285), .B(n10284), .Z(ADD_1071_U54) );
  XOR2_X1 U11303 ( .A(n10286), .B(n10287), .Z(ADD_1071_U53) );
  XNOR2_X1 U11304 ( .A(n10289), .B(n10288), .ZN(ADD_1071_U52) );
  CLKBUF_X3 U5003 ( .A(n5294), .Z(n4277) );
  INV_X1 U4775 ( .A(n8620), .ZN(n8637) );
  NOR2_X1 U4789 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5180) );
  CLKBUF_X1 U4796 ( .A(n5214), .Z(n5321) );
  CLKBUF_X1 U4808 ( .A(n5449), .Z(n10130) );
  CLKBUF_X1 U4852 ( .A(n8588), .Z(n4425) );
  AND4_X1 U5026 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n7768)
         );
  CLKBUF_X2 U5278 ( .A(n6044), .Z(n6424) );
  CLKBUF_X1 U5943 ( .A(n9941), .Z(n9954) );
  AND2_X1 U6913 ( .A1(n10031), .A2(n10030), .ZN(n10293) );
endmodule

