

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419;

  INV_X1 U2513 ( .A(n2478), .ZN(n2480) );
  INV_X1 U2514 ( .A(n2611), .ZN(n4103) );
  INV_X1 U2515 ( .A(n3090), .ZN(n4273) );
  INV_X2 U2516 ( .A(n3093), .ZN(n3296) );
  INV_X1 U2517 ( .A(n2478), .ZN(n2479) );
  NAND2_X1 U2518 ( .A1(n3340), .A2(n4729), .ZN(n4672) );
  NAND2_X1 U2519 ( .A1(n4661), .A2(n4658), .ZN(n3269) );
  INV_X1 U2520 ( .A(n2934), .ZN(n5151) );
  NAND2_X1 U2521 ( .A1(n3342), .A2(n4672), .ZN(n4610) );
  NAND2_X1 U2522 ( .A1(n2756), .A2(n5098), .ZN(n2478) );
  XNOR2_X2 U2523 ( .A(n3231), .B(n5109), .ZN(n3233) );
  OR2_X4 U2524 ( .A1(n2487), .A2(n3037), .ZN(n3231) );
  NAND2_X2 U2525 ( .A1(n2532), .A2(n2514), .ZN(n4313) );
  OR2_X2 U2526 ( .A1(n2855), .A2(n2856), .ZN(n2820) );
  XNOR2_X2 U2527 ( .A(n2815), .B(n5112), .ZN(n2855) );
  OAI21_X1 U2528 ( .B1(n4553), .B2(n2488), .A(n2662), .ZN(n4453) );
  AND2_X1 U2529 ( .A1(n2518), .A2(n2517), .ZN(n4758) );
  OR2_X1 U2530 ( .A1(n4240), .A2(n2661), .ZN(n2634) );
  NAND2_X1 U2531 ( .A1(n2653), .A2(n2509), .ZN(n4537) );
  AND2_X1 U2532 ( .A1(n2525), .A2(n4139), .ZN(n4154) );
  NOR2_X1 U2533 ( .A1(n4149), .A2(n4148), .ZN(n4167) );
  NAND2_X1 U2534 ( .A1(n3429), .A2(REG2_REG_10__SCAN_IN), .ZN(n3487) );
  NOR2_X2 U2535 ( .A1(n2486), .A2(n4796), .ZN(n4799) );
  XNOR2_X1 U2536 ( .A(n4128), .B(n3535), .ZN(n4127) );
  NAND2_X1 U2537 ( .A1(n3534), .A2(n3533), .ZN(n4128) );
  AND2_X1 U2538 ( .A1(n3277), .A2(n2663), .ZN(n3116) );
  NAND2_X1 U2539 ( .A1(n3041), .A2(n3040), .ZN(n3042) );
  NAND2_X1 U2540 ( .A1(n2522), .A2(n2521), .ZN(n3041) );
  NOR2_X2 U2541 ( .A1(n2834), .A2(n2833), .ZN(n5143) );
  NOR2_X1 U2542 ( .A1(n3008), .A2(n3375), .ZN(n3007) );
  NAND4_X1 U2543 ( .A1(n3089), .A2(n3088), .A3(n3087), .A4(n3086), .ZN(n4729)
         );
  NOR2_X1 U2544 ( .A1(n2818), .A2(n5111), .ZN(n2819) );
  AND2_X1 U2545 ( .A1(n5111), .A2(n2818), .ZN(n2816) );
  NAND2_X1 U2546 ( .A1(n2739), .A2(IR_REG_31__SCAN_IN), .ZN(n2740) );
  AND2_X2 U2547 ( .A1(n5097), .A2(n5098), .ZN(n4287) );
  BUF_X4 U2548 ( .A(n2738), .Z(n2481) );
  AOI21_X1 U2549 ( .B1(n2851), .B2(REG1_REG_3__SCAN_IN), .A(n2844), .ZN(n2845)
         );
  XOR2_X1 U2550 ( .A(n5112), .B(n2843), .Z(n2851) );
  NAND2_X1 U2551 ( .A1(n2531), .A2(n2530), .ZN(n2881) );
  NAND2_X1 U2552 ( .A1(n2529), .A2(n2497), .ZN(n2531) );
  NAND2_X1 U2553 ( .A1(n2679), .A2(IR_REG_31__SCAN_IN), .ZN(n2680) );
  AND4_X1 U2554 ( .A1(n2541), .A2(n2540), .A3(n2698), .A4(n3915), .ZN(n2674)
         );
  INV_X1 U2555 ( .A(IR_REG_7__SCAN_IN), .ZN(n2698) );
  INV_X1 U2556 ( .A(IR_REG_1__SCAN_IN), .ZN(n2536) );
  INV_X2 U2557 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U2558 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2541)
         );
  NOR2_X1 U2559 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2540)
         );
  NOR2_X2 U2560 ( .A1(n4161), .A2(n3529), .ZN(n4178) );
  OAI22_X2 U2561 ( .A1(n3235), .A2(n3234), .B1(n3233), .B2(n3232), .ZN(n3238)
         );
  INV_X1 U2562 ( .A(IR_REG_22__SCAN_IN), .ZN(n2744) );
  AND2_X1 U2563 ( .A1(n2741), .A2(n2656), .ZN(n2745) );
  AND4_X1 U2564 ( .A1(n2674), .A2(n2673), .A3(n2492), .A4(n2657), .ZN(n2656)
         );
  INV_X1 U2565 ( .A(IR_REG_21__SCAN_IN), .ZN(n2657) );
  AOI21_X1 U2566 ( .B1(n2622), .B2(n2620), .A(n2507), .ZN(n2619) );
  INV_X1 U2567 ( .A(n2662), .ZN(n2620) );
  OAI22_X1 U2568 ( .A1(n2617), .A2(n2616), .B1(n4292), .B2(n2619), .ZN(n2615)
         );
  NOR2_X1 U2569 ( .A1(n2622), .A2(n4292), .ZN(n2616) );
  NAND2_X1 U2570 ( .A1(n2628), .A2(n2626), .ZN(n4503) );
  AND2_X1 U2571 ( .A1(n4504), .A2(n2627), .ZN(n2626) );
  NAND2_X1 U2572 ( .A1(n4240), .A2(n2629), .ZN(n2628) );
  AOI22_X1 U2573 ( .A1(n2661), .A2(n2633), .B1(n2632), .B2(n2631), .ZN(n2627)
         );
  AOI22_X1 U2574 ( .A1(n2838), .A2(REG2_REG_2__SCAN_IN), .B1(n2839), .B2(n2812), .ZN(n2883) );
  INV_X1 U2575 ( .A(n5098), .ZN(n2757) );
  NAND2_X1 U2576 ( .A1(n3442), .A2(n4643), .ZN(n2560) );
  AND2_X1 U2577 ( .A1(n3764), .A2(n2770), .ZN(n2669) );
  NOR2_X1 U2578 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2771)
         );
  AND2_X1 U2579 ( .A1(n2745), .A2(n2744), .ZN(n2773) );
  AND2_X1 U2580 ( .A1(n2660), .A2(n2666), .ZN(n2741) );
  AND3_X1 U2581 ( .A1(n2727), .A2(n2715), .A3(n2668), .ZN(n2666) );
  NAND2_X1 U2582 ( .A1(n4537), .A2(n4209), .ZN(n4473) );
  INV_X1 U2583 ( .A(n3106), .ZN(n4285) );
  INV_X1 U2584 ( .A(n4287), .ZN(n4267) );
  INV_X1 U2585 ( .A(n2883), .ZN(n2530) );
  INV_X1 U2586 ( .A(n3024), .ZN(n3022) );
  NAND2_X1 U2587 ( .A1(n3487), .A2(n2665), .ZN(n3492) );
  NOR2_X2 U2588 ( .A1(n4135), .A2(n4133), .ZN(n4149) );
  INV_X1 U2589 ( .A(n4132), .ZN(n4133) );
  AOI21_X1 U2590 ( .B1(n4152), .B2(REG1_REG_13__SCAN_IN), .A(n4131), .ZN(n4132) );
  NOR2_X1 U2591 ( .A1(n4749), .A2(n4750), .ZN(n4748) );
  NAND2_X1 U2592 ( .A1(n3248), .A2(REG3_REG_21__SCAN_IN), .ZN(n4196) );
  INV_X1 U2593 ( .A(n4115), .ZN(n3248) );
  NAND2_X1 U2594 ( .A1(n2511), .A2(n2591), .ZN(n2588) );
  NOR2_X1 U2595 ( .A1(n2752), .A2(IR_REG_29__SCAN_IN), .ZN(n2754) );
  XNOR2_X1 U2596 ( .A(n2606), .B(n3774), .ZN(n2756) );
  OR2_X1 U2597 ( .A1(n2754), .A2(n5094), .ZN(n2606) );
  NAND2_X1 U2598 ( .A1(n4553), .A2(n2613), .ZN(n2612) );
  AND2_X1 U2599 ( .A1(n2615), .A2(n2494), .ZN(n2613) );
  INV_X1 U2600 ( .A(keyinput_56), .ZN(n2533) );
  INV_X1 U2601 ( .A(keyinput_184), .ZN(n2534) );
  INV_X1 U2602 ( .A(n2896), .ZN(n2898) );
  OR2_X1 U2603 ( .A1(n3343), .A2(n4610), .ZN(n3347) );
  INV_X1 U2604 ( .A(n4051), .ZN(n2652) );
  NOR2_X1 U2605 ( .A1(n2652), .A2(n2649), .ZN(n2648) );
  INV_X1 U2606 ( .A(n3636), .ZN(n2649) );
  INV_X1 U2607 ( .A(n4242), .ZN(n2632) );
  OR2_X1 U2608 ( .A1(n4804), .A2(n4803), .ZN(n4806) );
  NAND2_X1 U2609 ( .A1(n2489), .A2(n4647), .ZN(n3515) );
  INV_X1 U2610 ( .A(n4677), .ZN(n2559) );
  OR2_X1 U2611 ( .A1(n5252), .A2(n3395), .ZN(n3442) );
  NAND2_X1 U2612 ( .A1(n2496), .A2(n3336), .ZN(n2594) );
  NAND2_X1 U2613 ( .A1(n4379), .A2(n4868), .ZN(n2591) );
  OR2_X1 U2614 ( .A1(n3415), .A2(n3414), .ZN(n3416) );
  AND2_X1 U2615 ( .A1(n3413), .A2(n3412), .ZN(n3414) );
  NOR2_X1 U2616 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2715)
         );
  INV_X1 U2617 ( .A(IR_REG_2__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U2618 ( .A1(n2635), .A2(n2638), .ZN(n4460) );
  INV_X1 U2619 ( .A(n2639), .ZN(n2638) );
  OAI21_X1 U2620 ( .B1(n5311), .B2(n2640), .A(n4462), .ZN(n2639) );
  OAI21_X1 U2621 ( .B1(n3131), .B2(n2645), .A(n3203), .ZN(n2644) );
  NAND2_X1 U2622 ( .A1(n2986), .A2(n4735), .ZN(n2609) );
  INV_X1 U2623 ( .A(n4540), .ZN(n2655) );
  INV_X1 U2624 ( .A(n2956), .ZN(n2529) );
  NAND2_X1 U2625 ( .A1(n2523), .A2(n2495), .ZN(n2522) );
  INV_X1 U2626 ( .A(n3028), .ZN(n2523) );
  INV_X1 U2627 ( .A(n3031), .ZN(n2521) );
  AND2_X1 U2628 ( .A1(n5110), .A2(REG1_REG_7__SCAN_IN), .ZN(n3037) );
  NOR2_X1 U2629 ( .A1(n3044), .A2(n3045), .ZN(n3228) );
  NAND2_X1 U2630 ( .A1(n3539), .A2(n2527), .ZN(n3541) );
  NOR2_X1 U2631 ( .A1(n5107), .A2(n2528), .ZN(n2527) );
  INV_X1 U2632 ( .A(n3538), .ZN(n2528) );
  AND2_X1 U2633 ( .A1(n4152), .A2(REG1_REG_13__SCAN_IN), .ZN(n4148) );
  INV_X1 U2634 ( .A(n4320), .ZN(n2517) );
  AND2_X1 U2635 ( .A1(n4799), .A2(n4781), .ZN(n4787) );
  NAND2_X1 U2636 ( .A1(n2574), .A2(n2573), .ZN(n2572) );
  INV_X1 U2637 ( .A(n2575), .ZN(n2574) );
  NOR2_X1 U2638 ( .A1(n4874), .A2(n4830), .ZN(n2573) );
  INV_X1 U2639 ( .A(n4083), .ZN(n3247) );
  OR2_X1 U2640 ( .A1(n4971), .A2(n4962), .ZN(n4963) );
  AND2_X1 U2641 ( .A1(n4565), .A2(n4036), .ZN(n4031) );
  NAND2_X1 U2642 ( .A1(n3503), .A2(n2493), .ZN(n2581) );
  OR2_X1 U2643 ( .A1(n2503), .A2(n2580), .ZN(n2579) );
  INV_X1 U2644 ( .A(n2583), .ZN(n2580) );
  NAND2_X1 U2645 ( .A1(n3450), .A2(n3449), .ZN(n2600) );
  OAI21_X1 U2646 ( .B1(n3357), .B2(n4611), .A(n4671), .ZN(n4340) );
  INV_X1 U2647 ( .A(n4732), .ZN(n3368) );
  NAND2_X1 U2648 ( .A1(n2595), .A2(n4608), .ZN(n3337) );
  NAND2_X1 U2649 ( .A1(n2590), .A2(n4360), .ZN(n4421) );
  OAI21_X1 U2650 ( .B1(n4881), .B2(n2587), .A(n2585), .ZN(n2590) );
  AND2_X1 U2651 ( .A1(n2586), .A2(n4359), .ZN(n2585) );
  INV_X1 U2652 ( .A(n2603), .ZN(n4911) );
  OAI21_X1 U2653 ( .B1(n4921), .B2(n2510), .A(n2604), .ZN(n2603) );
  NAND2_X1 U2654 ( .A1(n4372), .A2(n4945), .ZN(n2604) );
  NAND4_X1 U2655 ( .A1(n2742), .A2(n2741), .A3(n2500), .A4(n2671), .ZN(n2752)
         );
  AND2_X1 U2656 ( .A1(n2771), .A2(n2770), .ZN(n2772) );
  INV_X1 U2657 ( .A(IR_REG_23__SCAN_IN), .ZN(n3952) );
  INV_X1 U2658 ( .A(IR_REG_3__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U2659 ( .A1(n2537), .A2(n2536), .ZN(n2679) );
  NAND2_X1 U2660 ( .A1(n2615), .A2(n2498), .ZN(n2614) );
  INV_X1 U2661 ( .A(n4292), .ZN(n2618) );
  NAND2_X1 U2662 ( .A1(n3637), .A2(n3638), .ZN(n4052) );
  OR2_X1 U2663 ( .A1(n4250), .A2(n4249), .ZN(n4251) );
  OR2_X1 U2664 ( .A1(n4801), .A2(n4267), .ZN(n4272) );
  NAND2_X1 U2665 ( .A1(n4216), .A2(n4215), .ZN(n4896) );
  NAND2_X1 U2666 ( .A1(n4202), .A2(n4201), .ZN(n4903) );
  OR2_X1 U2667 ( .A1(n4886), .A2(n4267), .ZN(n4202) );
  NAND4_X1 U2668 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n4726)
         );
  NOR2_X1 U2669 ( .A1(n4301), .A2(n4736), .ZN(n4746) );
  AOI21_X1 U2670 ( .B1(n4321), .B2(n4320), .A(n4773), .ZN(n4326) );
  NAND2_X1 U2671 ( .A1(n4323), .A2(n2658), .ZN(n4324) );
  NAND2_X1 U2672 ( .A1(n2739), .A2(n2737), .ZN(n4767) );
  OR2_X1 U2673 ( .A1(n5146), .A2(n2999), .ZN(n4768) );
  NAND2_X1 U2674 ( .A1(n2566), .A2(IR_REG_31__SCAN_IN), .ZN(n2565) );
  XNOR2_X1 U2675 ( .A(n2533), .B(IR_REG_1__SCAN_IN), .ZN(n3729) );
  XNOR2_X1 U2676 ( .A(n2534), .B(IR_REG_1__SCAN_IN), .ZN(n3911) );
  NOR2_X1 U2677 ( .A1(n4701), .A2(n2555), .ZN(n2554) );
  INV_X1 U2678 ( .A(n4640), .ZN(n2555) );
  NOR2_X1 U2679 ( .A1(n3405), .A2(n5243), .ZN(n3415) );
  INV_X1 U2680 ( .A(IR_REG_26__SCAN_IN), .ZN(n3764) );
  INV_X1 U2681 ( .A(IR_REG_13__SCAN_IN), .ZN(n3934) );
  INV_X1 U2682 ( .A(n2682), .ZN(n2673) );
  OR2_X1 U2683 ( .A1(n3100), .A2(n3169), .ZN(n3122) );
  AND2_X1 U2684 ( .A1(n3147), .A2(n3122), .ZN(n3277) );
  INV_X1 U2685 ( .A(n3607), .ZN(n2640) );
  NOR2_X1 U2686 ( .A1(n2640), .A2(n2637), .ZN(n2636) );
  INV_X1 U2687 ( .A(n5313), .ZN(n2637) );
  NAND2_X1 U2688 ( .A1(n4241), .A2(n4528), .ZN(n2629) );
  NAND2_X1 U2689 ( .A1(n2761), .A2(n5137), .ZN(n2738) );
  OAI21_X1 U2690 ( .B1(n5178), .B2(n2838), .A(n2842), .ZN(n2843) );
  NAND2_X1 U2691 ( .A1(n2970), .A2(n2659), .ZN(n3019) );
  INV_X1 U2692 ( .A(IR_REG_18__SCAN_IN), .ZN(n3755) );
  INV_X1 U2693 ( .A(n4638), .ZN(n2546) );
  NAND2_X1 U2694 ( .A1(n2557), .A2(n2553), .ZN(n4804) );
  NOR2_X1 U2695 ( .A1(n2556), .A2(n2554), .ZN(n2553) );
  NAND2_X1 U2696 ( .A1(n4428), .A2(n4581), .ZN(n2557) );
  INV_X1 U2697 ( .A(n4600), .ZN(n2556) );
  NAND2_X1 U2698 ( .A1(n4851), .A2(n4362), .ZN(n2575) );
  OAI21_X1 U2699 ( .B1(n4902), .B2(n4561), .A(n4378), .ZN(n4845) );
  OR2_X1 U2700 ( .A1(n4889), .A2(n4888), .ZN(n4891) );
  AND2_X1 U2701 ( .A1(n4368), .A2(n4602), .ZN(n4690) );
  NAND2_X1 U2702 ( .A1(n4723), .A2(n5320), .ZN(n2583) );
  INV_X1 U2703 ( .A(n2551), .ZN(n2550) );
  OAI21_X1 U2704 ( .B1(n4653), .B2(n2552), .A(n4651), .ZN(n2551) );
  AND2_X1 U2705 ( .A1(n4719), .A2(n4789), .ZN(n4589) );
  OR2_X1 U2706 ( .A1(n2504), .A2(n2587), .ZN(n2586) );
  INV_X1 U2707 ( .A(n2588), .ZN(n2587) );
  AND2_X1 U2708 ( .A1(n5242), .A2(n4627), .ZN(n5243) );
  AND2_X1 U2709 ( .A1(n3348), .A2(n3349), .ZN(n3413) );
  INV_X1 U2710 ( .A(IR_REG_25__SCAN_IN), .ZN(n2770) );
  NOR2_X1 U2711 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2727)
         );
  INV_X1 U2712 ( .A(n2619), .ZN(n2617) );
  INV_X1 U2713 ( .A(n4454), .ZN(n2623) );
  AND2_X1 U2714 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n3073) );
  XNOR2_X1 U2715 ( .A(n3119), .B(n3117), .ZN(n3147) );
  NOR2_X1 U2716 ( .A1(n3549), .A2(n4519), .ZN(n3568) );
  OR2_X1 U2717 ( .A1(n4240), .A2(n2632), .ZN(n2625) );
  NAND2_X1 U2718 ( .A1(n3130), .A2(n3131), .ZN(n3185) );
  NAND2_X1 U2719 ( .A1(n4187), .A2(n2508), .ZN(n2653) );
  INV_X1 U2720 ( .A(n4186), .ZN(n2654) );
  XNOR2_X1 U2721 ( .A(n2911), .B(n3093), .ZN(n2914) );
  NAND2_X1 U2722 ( .A1(n2647), .A2(n2650), .ZN(n4079) );
  INV_X1 U2723 ( .A(n2651), .ZN(n2650) );
  OAI21_X1 U2724 ( .B1(n3638), .B2(n2652), .A(n4063), .ZN(n2651) );
  NAND2_X1 U2725 ( .A1(n3568), .A2(REG3_REG_17__SCAN_IN), .ZN(n3639) );
  NOR2_X1 U2726 ( .A1(n3505), .A2(n4150), .ZN(n3518) );
  NAND2_X1 U2727 ( .A1(n3518), .A2(REG3_REG_15__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U2728 ( .A1(n2839), .A2(REG1_REG_2__SCAN_IN), .B1(n5178), .B2(n2838), .ZN(n2880) );
  NAND2_X1 U2729 ( .A1(n2881), .A2(n2813), .ZN(n2815) );
  OR2_X1 U2730 ( .A1(n5214), .A2(n3011), .ZN(n3009) );
  INV_X1 U2731 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3083) );
  INV_X1 U2732 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3239) );
  NOR2_X1 U2733 ( .A1(n3427), .A2(n2512), .ZN(n3486) );
  XNOR2_X1 U2734 ( .A(n3479), .B(n3428), .ZN(n3436) );
  INV_X1 U2735 ( .A(n3494), .ZN(n3491) );
  NAND2_X1 U2736 ( .A1(n3435), .A2(n3434), .ZN(n3479) );
  AND2_X1 U2737 ( .A1(n4159), .A2(n4158), .ZN(n4160) );
  OR2_X1 U2738 ( .A1(n4181), .A2(n4180), .ZN(n2532) );
  OAI22_X1 U2739 ( .A1(n4169), .A2(n4168), .B1(n4167), .B2(n4166), .ZN(n4172)
         );
  NAND2_X1 U2740 ( .A1(n4172), .A2(n4171), .ZN(n4299) );
  XNOR2_X1 U2741 ( .A(n4313), .B(n5379), .ZN(n4739) );
  NAND2_X1 U2742 ( .A1(n4299), .A2(n4298), .ZN(n4300) );
  OR2_X1 U2743 ( .A1(n4748), .A2(n4317), .ZN(n2518) );
  INV_X1 U2744 ( .A(IR_REG_19__SCAN_IN), .ZN(n3754) );
  INV_X1 U2745 ( .A(n2544), .ZN(n2543) );
  OAI22_X1 U2746 ( .A1(n4779), .A2(n2545), .B1(n4431), .B2(n2546), .ZN(n2544)
         );
  NAND2_X1 U2747 ( .A1(n4431), .A2(n2546), .ZN(n2545) );
  NAND2_X1 U2748 ( .A1(n4778), .A2(n4779), .ZN(n4777) );
  OR2_X1 U2749 ( .A1(n4428), .A2(n4640), .ZN(n4817) );
  NOR3_X1 U2750 ( .A1(n4883), .A2(n4874), .A3(n4532), .ZN(n4839) );
  NOR2_X1 U2751 ( .A1(n4883), .A2(n4874), .ZN(n4873) );
  OR2_X1 U2752 ( .A1(n4210), .A2(n4476), .ZN(n4228) );
  NAND2_X1 U2753 ( .A1(n4925), .A2(n4914), .ZN(n4913) );
  OR2_X1 U2754 ( .A1(n4913), .A2(n4882), .ZN(n4883) );
  NAND2_X1 U2755 ( .A1(n2563), .A2(n4562), .ZN(n4902) );
  NAND2_X1 U2756 ( .A1(n4930), .A2(n4690), .ZN(n2563) );
  NOR2_X1 U2757 ( .A1(n4963), .A2(n4922), .ZN(n4925) );
  NAND2_X1 U2758 ( .A1(n3246), .A2(REG3_REG_19__SCAN_IN), .ZN(n4083) );
  INV_X1 U2759 ( .A(n4069), .ZN(n3246) );
  NAND2_X1 U2760 ( .A1(n4992), .A2(n2513), .ZN(n4971) );
  NAND2_X1 U2761 ( .A1(n4992), .A2(n5001), .ZN(n4994) );
  OR2_X1 U2762 ( .A1(n4998), .A2(n4518), .ZN(n4347) );
  AND2_X1 U2763 ( .A1(n4042), .A2(n4349), .ZN(n4992) );
  AND2_X1 U2764 ( .A1(n2577), .A2(n3558), .ZN(n2576) );
  NAND2_X1 U2765 ( .A1(n3510), .A2(n3526), .ZN(n3558) );
  OR2_X1 U2766 ( .A1(n2579), .A2(n2578), .ZN(n2577) );
  NOR2_X1 U2767 ( .A1(n3560), .A2(n5365), .ZN(n4042) );
  NAND2_X1 U2768 ( .A1(n5324), .A2(n5331), .ZN(n5323) );
  OR2_X1 U2769 ( .A1(n5323), .A2(n4464), .ZN(n3560) );
  NAND2_X1 U2770 ( .A1(n2549), .A2(n2548), .ZN(n4035) );
  AOI21_X1 U2771 ( .B1(n2550), .B2(n2552), .A(n4609), .ZN(n2548) );
  NAND2_X1 U2772 ( .A1(n3515), .A2(n2550), .ZN(n2549) );
  OAI21_X1 U2773 ( .B1(n3515), .B2(n2552), .A(n2550), .ZN(n4564) );
  NAND2_X1 U2774 ( .A1(n3459), .A2(REG3_REG_13__SCAN_IN), .ZN(n3505) );
  NAND2_X1 U2775 ( .A1(n3515), .A2(n4653), .ZN(n5326) );
  AND2_X1 U2776 ( .A1(n3307), .A2(REG3_REG_12__SCAN_IN), .ZN(n3459) );
  AND2_X1 U2777 ( .A1(n3213), .A2(REG3_REG_11__SCAN_IN), .ZN(n3307) );
  NOR2_X1 U2778 ( .A1(n3473), .A2(n4495), .ZN(n5324) );
  NAND2_X1 U2779 ( .A1(n5247), .A2(n2567), .ZN(n3473) );
  AND2_X1 U2780 ( .A1(n2569), .A2(n2568), .ZN(n2567) );
  NOR2_X1 U2781 ( .A1(n4400), .A2(n3469), .ZN(n2568) );
  NAND2_X1 U2782 ( .A1(n2560), .A2(n2558), .ZN(n2561) );
  NOR2_X1 U2783 ( .A1(n3444), .A2(n2559), .ZN(n2558) );
  OAI21_X1 U2784 ( .B1(n3450), .B2(n2599), .A(n2596), .ZN(n2601) );
  AOI21_X1 U2785 ( .B1(n2598), .B2(n2597), .A(n2602), .ZN(n2596) );
  AND2_X1 U2786 ( .A1(n4725), .A2(n4400), .ZN(n2602) );
  AND2_X1 U2787 ( .A1(n3186), .A2(REG3_REG_10__SCAN_IN), .ZN(n3213) );
  NOR2_X1 U2788 ( .A1(n3133), .A2(n3239), .ZN(n3186) );
  NAND2_X1 U2789 ( .A1(n2560), .A2(n4677), .ZN(n4405) );
  AND2_X1 U2790 ( .A1(n3400), .A2(n5256), .ZN(n2569) );
  NAND2_X1 U2791 ( .A1(n3103), .A2(REG3_REG_7__SCAN_IN), .ZN(n3105) );
  OR2_X1 U2792 ( .A1(n3105), .A2(n3141), .ZN(n3133) );
  AND2_X1 U2793 ( .A1(n5247), .A2(n5256), .ZN(n5248) );
  OAI21_X1 U2794 ( .B1(n4340), .B2(n3326), .A(n3342), .ZN(n3327) );
  AND2_X1 U2795 ( .A1(n4674), .A2(n4642), .ZN(n4628) );
  INV_X1 U2796 ( .A(n5184), .ZN(n5302) );
  NOR2_X1 U2797 ( .A1(n4334), .A2(n3404), .ZN(n5247) );
  OR2_X1 U2798 ( .A1(n4336), .A2(n4342), .ZN(n4334) );
  NAND2_X1 U2799 ( .A1(n3325), .A2(n4668), .ZN(n3357) );
  NAND2_X1 U2800 ( .A1(n2482), .A2(n3361), .ZN(n4336) );
  OAI211_X1 U2801 ( .C1(n2595), .C2(n2594), .A(n2499), .B(n2593), .ZN(n3372)
         );
  NAND2_X1 U2802 ( .A1(n2592), .A2(n3321), .ZN(n2593) );
  INV_X1 U2803 ( .A(n2594), .ZN(n2592) );
  NAND2_X1 U2804 ( .A1(n2610), .A2(n2945), .ZN(n3266) );
  INV_X1 U2805 ( .A(n2940), .ZN(n2610) );
  NAND2_X1 U2806 ( .A1(n2483), .A2(n2681), .ZN(n5194) );
  NAND2_X1 U2807 ( .A1(n2562), .A2(n4662), .ZN(n5183) );
  NAND2_X1 U2808 ( .A1(n3322), .A2(n3321), .ZN(n2562) );
  NAND2_X1 U2809 ( .A1(n3385), .A2(n3270), .ZN(n3272) );
  NAND2_X1 U2810 ( .A1(n2681), .A2(n3335), .ZN(n5196) );
  OAI21_X1 U2811 ( .B1(n3269), .B2(n4657), .A(n4661), .ZN(n3322) );
  INV_X1 U2812 ( .A(n5330), .ZN(n5396) );
  OR2_X1 U2813 ( .A1(n2864), .A2(n5149), .ZN(n5330) );
  AOI211_X1 U2814 ( .C1(n4789), .C2(n4788), .A(n5390), .B(n4787), .ZN(n5012)
         );
  OR2_X1 U2815 ( .A1(n4584), .A2(n4589), .ZN(n4775) );
  AOI21_X1 U2816 ( .B1(n4827), .B2(n4423), .A(n4422), .ZN(n4795) );
  NAND2_X1 U2817 ( .A1(n2605), .A2(n4356), .ZN(n4921) );
  NAND2_X1 U2818 ( .A1(n4959), .A2(n4355), .ZN(n2605) );
  NAND2_X1 U2819 ( .A1(n4371), .A2(n4956), .ZN(n4355) );
  AOI22_X1 U2820 ( .A1(n4970), .A2(n4978), .B1(n4354), .B2(n4353), .ZN(n4959)
         );
  INV_X1 U2821 ( .A(n5406), .ZN(n5390) );
  NAND2_X1 U2822 ( .A1(n2774), .A2(n2775), .ZN(n2781) );
  MUX2_X1 U2823 ( .A(IR_REG_31__SCAN_IN), .B(n2769), .S(IR_REG_25__SCAN_IN), 
        .Z(n2774) );
  NAND2_X1 U2824 ( .A1(n2746), .A2(n2607), .ZN(n4361) );
  INV_X1 U2825 ( .A(n2773), .ZN(n2607) );
  INV_X1 U2826 ( .A(IR_REG_20__SCAN_IN), .ZN(n3947) );
  AND2_X1 U2827 ( .A1(n2724), .A2(n2725), .ZN(n4310) );
  INV_X1 U2828 ( .A(IR_REG_5__SCAN_IN), .ZN(n2691) );
  XNOR2_X1 U2829 ( .A(n2689), .B(IR_REG_5__SCAN_IN), .ZN(n2836) );
  NAND2_X1 U2830 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2677)
         );
  INV_X1 U2831 ( .A(n4727), .ZN(n3403) );
  NAND2_X1 U2832 ( .A1(n5317), .A2(n3607), .ZN(n4461) );
  OAI22_X1 U2833 ( .A1(n3130), .A2(n2642), .B1(n2643), .B2(n3202), .ZN(n3211)
         );
  NAND2_X1 U2834 ( .A1(n2646), .A2(n3184), .ZN(n2642) );
  INV_X1 U2835 ( .A(n2644), .ZN(n2643) );
  NAND2_X1 U2836 ( .A1(n3211), .A2(n3210), .ZN(n3584) );
  INV_X1 U2837 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3141) );
  INV_X1 U2838 ( .A(n3387), .ZN(n4420) );
  XNOR2_X1 U2839 ( .A(n2914), .B(n2915), .ZN(n4415) );
  NAND2_X1 U2840 ( .A1(n4187), .A2(n4186), .ZN(n4486) );
  OR2_X1 U2841 ( .A1(n4833), .A2(n4267), .ZN(n4260) );
  INV_X1 U2842 ( .A(n3448), .ZN(n3400) );
  NAND2_X1 U2843 ( .A1(n3185), .A2(n3184), .ZN(n3204) );
  NAND2_X1 U2844 ( .A1(n2641), .A2(n5311), .ZN(n5317) );
  NAND2_X1 U2845 ( .A1(n5314), .A2(n5313), .ZN(n2641) );
  NAND2_X1 U2846 ( .A1(n2653), .A2(n4483), .ZN(n4539) );
  NAND2_X1 U2847 ( .A1(n4052), .A2(n4051), .ZN(n4062) );
  AND2_X1 U2848 ( .A1(n2939), .A2(n2938), .ZN(n5359) );
  INV_X1 U2849 ( .A(n4809), .ZN(n4720) );
  INV_X1 U2850 ( .A(n4821), .ZN(n4853) );
  NAND2_X1 U2851 ( .A1(n4234), .A2(n4233), .ZN(n4870) );
  OR2_X1 U2852 ( .A1(n4842), .A2(n4267), .ZN(n4234) );
  NAND2_X1 U2853 ( .A1(n4121), .A2(n4120), .ZN(n4947) );
  NAND2_X1 U2854 ( .A1(n4089), .A2(n4088), .ZN(n4905) );
  OR2_X1 U2855 ( .A1(n4926), .A2(n4267), .ZN(n4089) );
  NAND4_X1 U2856 ( .A1(n2933), .A2(n2932), .A3(n2931), .A4(n2930), .ZN(n4732)
         );
  NAND4_X1 U2857 ( .A1(n2893), .A2(n2892), .A3(n2891), .A4(n2890), .ZN(n4733)
         );
  NAND4_X1 U2858 ( .A1(n2863), .A2(n2862), .A3(n2861), .A4(n2860), .ZN(n4735)
         );
  INV_X1 U2859 ( .A(n2531), .ZN(n2884) );
  XNOR2_X1 U2860 ( .A(n2845), .B(n3014), .ZN(n3011) );
  NOR2_X1 U2861 ( .A1(n3007), .A2(n2823), .ZN(n2968) );
  NOR2_X1 U2862 ( .A1(n2968), .A2(n2967), .ZN(n2966) );
  NOR2_X1 U2863 ( .A1(n3030), .A2(n2519), .ZN(n3033) );
  OAI21_X1 U2864 ( .B1(n2522), .B2(n2521), .A(n2520), .ZN(n2519) );
  INV_X1 U2865 ( .A(n4773), .ZN(n2520) );
  NOR2_X1 U2866 ( .A1(n3228), .A2(n3227), .ZN(n3229) );
  NOR2_X1 U2867 ( .A1(n3229), .A2(n3230), .ZN(n3427) );
  AND2_X1 U2868 ( .A1(n2525), .A2(n2524), .ZN(n3544) );
  AND2_X1 U2869 ( .A1(n4130), .A2(n4129), .ZN(n4135) );
  XNOR2_X1 U2870 ( .A(n4167), .B(n4166), .ZN(n4169) );
  INV_X1 U2871 ( .A(n2532), .ZN(n4311) );
  XNOR2_X1 U2872 ( .A(n4300), .B(n4312), .ZN(n4737) );
  NOR2_X1 U2873 ( .A1(n4758), .A2(n2515), .ZN(n4761) );
  NOR2_X1 U2874 ( .A1(n2516), .A2(n4319), .ZN(n2515) );
  AOI21_X1 U2875 ( .B1(REG1_REG_18__SCAN_IN), .B2(n5104), .A(n4762), .ZN(n4764) );
  XNOR2_X1 U2876 ( .A(n2571), .B(n4577), .ZN(n5416) );
  AND2_X1 U2877 ( .A1(n2485), .A2(n5400), .ZN(n2570) );
  AND2_X1 U2878 ( .A1(n4282), .A2(n4281), .ZN(n4790) );
  NAND2_X1 U2879 ( .A1(n3511), .A2(n4609), .ZN(n3559) );
  NAND2_X1 U2880 ( .A1(n2581), .A2(n2579), .ZN(n3511) );
  AND2_X1 U2881 ( .A1(n2582), .A2(n2491), .ZN(n5322) );
  NAND2_X1 U2882 ( .A1(n3503), .A2(n4620), .ZN(n2582) );
  AND2_X1 U2883 ( .A1(n2600), .A2(n2598), .ZN(n4399) );
  AND2_X1 U2884 ( .A1(n2600), .A2(n2490), .ZN(n4397) );
  NAND2_X1 U2885 ( .A1(n5247), .A2(n2569), .ZN(n5272) );
  NAND2_X1 U2886 ( .A1(n3337), .A2(n3336), .ZN(n5181) );
  NAND2_X1 U2887 ( .A1(n2584), .A2(n2588), .ZN(n4838) );
  NAND2_X1 U2888 ( .A1(n4881), .A2(n2504), .ZN(n2584) );
  AND2_X1 U2889 ( .A1(n2589), .A2(n2506), .ZN(n4858) );
  NAND2_X1 U2890 ( .A1(n4881), .A2(n4888), .ZN(n2589) );
  INV_X1 U2891 ( .A(n2756), .ZN(n5097) );
  AND2_X1 U2892 ( .A1(n2755), .A2(n5095), .ZN(n5098) );
  MUX2_X1 U2893 ( .A(IR_REG_31__SCAN_IN), .B(n2753), .S(IR_REG_29__SCAN_IN), 
        .Z(n2755) );
  XNOR2_X1 U2894 ( .A(n2776), .B(IR_REG_26__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U2895 ( .A1(n2775), .A2(IR_REG_31__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U2896 ( .A1(n2766), .A2(IR_REG_31__SCAN_IN), .ZN(n2767) );
  AND2_X1 U2897 ( .A1(n2994), .A2(STATE_REG_SCAN_IN), .ZN(n2810) );
  INV_X1 U2898 ( .A(n4361), .ZN(n5102) );
  INV_X1 U2899 ( .A(n4592), .ZN(n5103) );
  NOR2_X1 U2900 ( .A1(n2717), .A2(n2716), .ZN(n4152) );
  AND2_X1 U2901 ( .A1(n2701), .A2(n2700), .ZN(n5110) );
  AND2_X1 U2902 ( .A1(n2686), .A2(n2685), .ZN(n5112) );
  OAI211_X1 U2903 ( .C1(n4553), .C2(n2614), .A(n2612), .B(n5366), .ZN(n2624)
         );
  AOI21_X1 U2904 ( .B1(n4326), .B2(n4325), .A(n4324), .ZN(n4327) );
  OR2_X1 U2905 ( .A1(n4452), .A2(n5051), .ZN(n2539) );
  OR2_X1 U2906 ( .A1(n4452), .A2(n5092), .ZN(n2538) );
  AND3_X1 U2907 ( .A1(n2681), .A2(n2483), .A3(n3324), .ZN(n2482) );
  AND2_X1 U2908 ( .A1(n2608), .A2(n3266), .ZN(n2986) );
  AND2_X1 U2909 ( .A1(n3338), .A2(n3335), .ZN(n2483) );
  AND2_X1 U2910 ( .A1(n2634), .A2(n2633), .ZN(n2484) );
  AND2_X2 U2911 ( .A1(n2896), .A2(n2865), .ZN(n3090) );
  INV_X1 U2912 ( .A(n3449), .ZN(n2597) );
  OAI21_X1 U2913 ( .B1(n2733), .B2(IR_REG_17__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2734) );
  AND2_X1 U2914 ( .A1(n4439), .A2(n4781), .ZN(n2485) );
  OR2_X1 U2915 ( .A1(n4883), .A2(n2572), .ZN(n2486) );
  NAND3_X1 U2916 ( .A1(n2778), .A2(n5101), .A3(n5100), .ZN(n2865) );
  INV_X1 U2917 ( .A(n2839), .ZN(n2838) );
  AND2_X1 U2918 ( .A1(n3023), .A2(n3022), .ZN(n2487) );
  NOR2_X1 U2919 ( .A1(n4262), .A2(n4263), .ZN(n2488) );
  NAND4_X1 U2920 ( .A1(n2908), .A2(n2907), .A3(n2906), .A4(n2905), .ZN(n2934)
         );
  AND2_X1 U2921 ( .A1(n2561), .A2(n4646), .ZN(n2489) );
  OR2_X1 U2922 ( .A1(n4726), .A2(n3448), .ZN(n2490) );
  NAND2_X1 U2923 ( .A1(n3502), .A2(n3501), .ZN(n2491) );
  NOR2_X1 U2924 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2492)
         );
  AND2_X1 U2925 ( .A1(n4620), .A2(n2583), .ZN(n2493) );
  OR2_X1 U2926 ( .A1(n2617), .A2(n4292), .ZN(n2494) );
  OR2_X1 U2927 ( .A1(n3027), .A2(n2826), .ZN(n2495) );
  INV_X1 U2928 ( .A(n2622), .ZN(n2621) );
  AOI21_X1 U2929 ( .B1(n2488), .B2(n2662), .A(n2623), .ZN(n2622) );
  INV_X1 U2930 ( .A(n2518), .ZN(n4321) );
  INV_X1 U2931 ( .A(n2630), .ZN(n4526) );
  OR2_X1 U2932 ( .A1(n4732), .A2(n5197), .ZN(n2496) );
  INV_X1 U2933 ( .A(n3184), .ZN(n2645) );
  AND2_X1 U2934 ( .A1(n4361), .A2(n4592), .ZN(n2945) );
  NAND2_X1 U2935 ( .A1(n2841), .A2(REG2_REG_1__SCAN_IN), .ZN(n2497) );
  OR2_X1 U2936 ( .A1(n2621), .A2(n2618), .ZN(n2498) );
  OR2_X1 U2937 ( .A1(n3368), .A2(n3338), .ZN(n2499) );
  AND2_X1 U2938 ( .A1(n2675), .A2(n3959), .ZN(n2500) );
  INV_X1 U2939 ( .A(n2599), .ZN(n2598) );
  NAND2_X1 U2940 ( .A1(n4404), .A2(n2490), .ZN(n2599) );
  AND2_X1 U2941 ( .A1(n2625), .A2(n2631), .ZN(n2501) );
  INV_X1 U2942 ( .A(IR_REG_31__SCAN_IN), .ZN(n5094) );
  AND2_X1 U2943 ( .A1(n4779), .A2(n4638), .ZN(n2502) );
  AND2_X1 U2944 ( .A1(n3504), .A2(n2491), .ZN(n2503) );
  INV_X1 U2945 ( .A(IR_REG_4__SCAN_IN), .ZN(n3915) );
  INV_X1 U2946 ( .A(n4609), .ZN(n2578) );
  AND3_X1 U2947 ( .A1(n2674), .A2(n2492), .A3(n2673), .ZN(n2742) );
  OAI211_X1 U2948 ( .C1(n4285), .C2(n5086), .A(n4072), .B(n4071), .ZN(n4943)
         );
  NAND2_X1 U2949 ( .A1(n2674), .A2(n2673), .ZN(n2703) );
  AND2_X1 U2950 ( .A1(n2591), .A2(n4888), .ZN(n2504) );
  OR2_X1 U2951 ( .A1(n2773), .A2(n5094), .ZN(n2777) );
  OR3_X1 U2952 ( .A1(n4883), .A2(n2575), .A3(n4874), .ZN(n2505) );
  NAND2_X1 U2953 ( .A1(n4903), .A2(n4882), .ZN(n2506) );
  AND2_X1 U2954 ( .A1(n4278), .A2(n4277), .ZN(n2507) );
  NAND2_X1 U2955 ( .A1(n4513), .A2(n3636), .ZN(n3637) );
  NOR2_X1 U2956 ( .A1(n4482), .A2(n2654), .ZN(n2508) );
  AND2_X1 U2957 ( .A1(n2655), .A2(n4483), .ZN(n2509) );
  AND2_X1 U2958 ( .A1(n4905), .A2(n4922), .ZN(n2510) );
  INV_X1 U2959 ( .A(n4241), .ZN(n2631) );
  NAND2_X1 U2960 ( .A1(n3492), .A2(n3491), .ZN(n3539) );
  INV_X1 U2961 ( .A(n3202), .ZN(n2646) );
  NAND2_X1 U2962 ( .A1(n4358), .A2(n2506), .ZN(n2511) );
  NAND2_X1 U2963 ( .A1(n2898), .A2(n2865), .ZN(n2611) );
  XNOR2_X1 U2964 ( .A(n2767), .B(IR_REG_24__SCAN_IN), .ZN(n2778) );
  BUF_X1 U2965 ( .A(n2986), .Z(n4239) );
  OAI21_X1 U2966 ( .B1(n2581), .B2(n2578), .A(n2576), .ZN(n4033) );
  AND2_X1 U2967 ( .A1(n3426), .A2(REG2_REG_9__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U2968 ( .A1(n2535), .A2(n3226), .ZN(n3044) );
  INV_X1 U2969 ( .A(n2601), .ZN(n3451) );
  AND2_X1 U2970 ( .A1(n5001), .A2(n4353), .ZN(n2513) );
  INV_X1 U2971 ( .A(n4650), .ZN(n2552) );
  INV_X1 U2972 ( .A(IR_REG_16__SCAN_IN), .ZN(n3935) );
  NAND2_X1 U2973 ( .A1(n2866), .A2(n2609), .ZN(n2872) );
  AND2_X1 U2974 ( .A1(n4662), .A2(n4665), .ZN(n3321) );
  NAND2_X1 U2975 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4310), .ZN(n2514) );
  INV_X1 U2976 ( .A(n4627), .ZN(n5251) );
  INV_X1 U2977 ( .A(n5104), .ZN(n2516) );
  AOI21_X1 U2978 ( .B1(n3542), .B2(n3543), .A(n4773), .ZN(n2524) );
  NAND2_X1 U2979 ( .A1(n2526), .A2(REG2_REG_12__SCAN_IN), .ZN(n2525) );
  INV_X1 U2980 ( .A(n3542), .ZN(n2526) );
  NAND2_X1 U2981 ( .A1(n3539), .A2(n3538), .ZN(n3540) );
  NOR2_X1 U2982 ( .A1(n4178), .A2(n4177), .ZN(n4181) );
  XNOR2_X2 U2983 ( .A(n2677), .B(IR_REG_1__SCAN_IN), .ZN(n2841) );
  NAND2_X1 U2984 ( .A1(n3042), .A2(n5109), .ZN(n3226) );
  NAND2_X1 U2985 ( .A1(n3043), .A2(n3234), .ZN(n2535) );
  INV_X1 U2986 ( .A(n2820), .ZN(n2854) );
  NAND3_X1 U2987 ( .A1(n2537), .A2(n2536), .A3(n2672), .ZN(n2682) );
  INV_X1 U2988 ( .A(IR_REG_0__SCAN_IN), .ZN(n2537) );
  OAI21_X1 U2989 ( .B1(n5106), .B2(n4176), .A(n4160), .ZN(n4161) );
  NAND2_X1 U2990 ( .A1(n4127), .A2(REG1_REG_12__SCAN_IN), .ZN(n4130) );
  NAND2_X1 U2991 ( .A1(n4739), .A2(n4044), .ZN(n4738) );
  NAND2_X1 U2992 ( .A1(n4451), .A2(n2538), .ZN(U3515) );
  NAND2_X1 U2993 ( .A1(n4441), .A2(n2539), .ZN(U3547) );
  OAI211_X1 U2994 ( .C1(n4778), .C2(n2545), .A(n2543), .B(n2542), .ZN(n2547)
         );
  NAND2_X1 U2995 ( .A1(n4778), .A2(n2502), .ZN(n2542) );
  AOI21_X1 U2996 ( .B1(n2547), .B2(n5333), .A(n4438), .ZN(n4442) );
  NAND2_X1 U2997 ( .A1(n2566), .A2(n2564), .ZN(n5137) );
  OR2_X1 U2998 ( .A1(n2676), .A2(n3959), .ZN(n2564) );
  XNOR2_X1 U2999 ( .A(n2565), .B(n2675), .ZN(n2761) );
  NAND2_X1 U3000 ( .A1(n2676), .A2(n3959), .ZN(n2566) );
  NAND2_X1 U3001 ( .A1(n4799), .A2(n2485), .ZN(n5401) );
  NAND2_X1 U3002 ( .A1(n4799), .A2(n2570), .ZN(n2571) );
  INV_X1 U3003 ( .A(n3272), .ZN(n2595) );
  NAND2_X1 U3004 ( .A1(n3451), .A2(n4617), .ZN(n3472) );
  NAND3_X1 U3005 ( .A1(n2742), .A2(n2741), .A3(n2671), .ZN(n2751) );
  AND2_X2 U3006 ( .A1(n2757), .A2(n2756), .ZN(n3106) );
  INV_X1 U3007 ( .A(n2611), .ZN(n2608) );
  NAND2_X1 U3008 ( .A1(n2624), .A2(n4297), .ZN(U3217) );
  OR2_X1 U3009 ( .A1(n2484), .A2(n2501), .ZN(n2630) );
  INV_X1 U3010 ( .A(n4240), .ZN(n4474) );
  INV_X1 U3011 ( .A(n2634), .ZN(n4530) );
  INV_X1 U3012 ( .A(n4528), .ZN(n2633) );
  NAND2_X1 U3013 ( .A1(n5314), .A2(n2636), .ZN(n2635) );
  NAND2_X1 U3014 ( .A1(n4513), .A2(n2648), .ZN(n2647) );
  NAND2_X1 U3015 ( .A1(n2742), .A2(n2741), .ZN(n2747) );
  INV_X1 U3016 ( .A(n5165), .ZN(n2681) );
  NAND2_X1 U3017 ( .A1(n2678), .A2(n4420), .ZN(n5165) );
  NOR2_X1 U3018 ( .A1(n2966), .A2(n2825), .ZN(n3027) );
  AOI21_X1 U3019 ( .B1(n4790), .B2(n4287), .A(n4286), .ZN(n4719) );
  AOI22_X2 U3020 ( .A1(n4421), .A2(n4640), .B1(n4506), .B2(n4853), .ZN(n4827)
         );
  OR2_X1 U3021 ( .A1(STATE_REG_SCAN_IN), .A2(n4322), .ZN(n2658) );
  INV_X1 U3022 ( .A(n3480), .ZN(n3428) );
  OR2_X1 U3023 ( .A1(n5218), .A2(n2837), .ZN(n2659) );
  AND4_X1 U3024 ( .A1(n3755), .A2(n3942), .A3(n3934), .A4(n3935), .ZN(n2660)
         );
  INV_X1 U3025 ( .A(n5107), .ZN(n3535) );
  INV_X1 U3026 ( .A(n5225), .ZN(n2826) );
  NAND2_X1 U3027 ( .A1(n4241), .A2(n4242), .ZN(n2661) );
  OR2_X1 U3028 ( .A1(n4551), .A2(n4550), .ZN(n2662) );
  AND2_X1 U3029 ( .A1(n3146), .A2(n3126), .ZN(n2663) );
  OR2_X1 U3030 ( .A1(n2903), .A2(n3296), .ZN(n2664) );
  INV_X1 U3031 ( .A(n4604), .ZN(n2678) );
  OR2_X1 U3032 ( .A1(n3486), .A2(n3428), .ZN(n2665) );
  OR2_X1 U3033 ( .A1(n4154), .A2(n4155), .ZN(n4153) );
  NOR2_X1 U3034 ( .A1(n4155), .A2(n4166), .ZN(n2667) );
  INV_X1 U3035 ( .A(n3469), .ZN(n3470) );
  NOR2_X1 U3036 ( .A1(n2670), .A2(IR_REG_21__SCAN_IN), .ZN(n2671) );
  NOR2_X1 U3037 ( .A1(n3158), .A2(n3071), .ZN(n3072) );
  AND2_X2 U3038 ( .A1(n2864), .A2(n5103), .ZN(n2896) );
  INV_X1 U3039 ( .A(n4228), .ZN(n3249) );
  INV_X1 U3040 ( .A(n3639), .ZN(n3245) );
  AND2_X1 U3041 ( .A1(n2843), .A2(n5112), .ZN(n2844) );
  AND2_X1 U3042 ( .A1(n2836), .A2(REG2_REG_5__SCAN_IN), .ZN(n2825) );
  OR3_X1 U3043 ( .A1(n4254), .A2(n4253), .A3(n4252), .ZN(n4265) );
  OR2_X1 U3044 ( .A1(n4196), .A2(n4541), .ZN(n4210) );
  NAND2_X1 U3045 ( .A1(n3247), .A2(REG3_REG_20__SCAN_IN), .ZN(n4115) );
  OR2_X1 U3046 ( .A1(n4350), .A2(n4349), .ZN(n4351) );
  INV_X1 U3047 ( .A(IR_REG_27__SCAN_IN), .ZN(n3959) );
  INV_X1 U3048 ( .A(n4723), .ZN(n4465) );
  NAND2_X1 U3049 ( .A1(n3249), .A2(REG3_REG_24__SCAN_IN), .ZN(n4254) );
  NAND2_X1 U3050 ( .A1(n3635), .A2(n3634), .ZN(n5361) );
  NAND2_X1 U3051 ( .A1(n3245), .A2(REG3_REG_18__SCAN_IN), .ZN(n4069) );
  NOR2_X1 U3052 ( .A1(n3084), .A2(n3083), .ZN(n3103) );
  INV_X1 U3053 ( .A(n5186), .ZN(n5304) );
  OR2_X1 U3054 ( .A1(n4280), .A2(n4279), .ZN(n4282) );
  AOI22_X1 U3055 ( .A1(n2840), .A2(REG2_REG_1__SCAN_IN), .B1(n3389), .B2(n2841), .ZN(n2955) );
  XNOR2_X1 U3056 ( .A(n3019), .B(n2826), .ZN(n2846) );
  INV_X1 U3057 ( .A(n4369), .ZN(n5001) );
  INV_X1 U3058 ( .A(n5320), .ZN(n5331) );
  INV_X1 U3059 ( .A(n3339), .ZN(n3361) );
  OR2_X1 U3060 ( .A1(n4903), .A2(n4894), .ZN(n4863) );
  NAND2_X1 U3061 ( .A1(n4943), .A2(n4962), .ZN(n4356) );
  INV_X1 U3062 ( .A(n4518), .ZN(n4349) );
  INV_X1 U3063 ( .A(n5250), .ZN(n5256) );
  INV_X1 U3064 ( .A(n2945), .ZN(n5149) );
  MUX2_X1 U3065 ( .A(n5107), .B(DATAI_12_), .S(n2481), .Z(n4495) );
  NAND2_X1 U3066 ( .A1(n3073), .A2(REG3_REG_5__SCAN_IN), .ZN(n3084) );
  AND2_X1 U3067 ( .A1(n5359), .A2(n2999), .ZN(n4558) );
  INV_X1 U3068 ( .A(n5315), .ZN(n5366) );
  OR2_X1 U3069 ( .A1(n4916), .A2(n4267), .ZN(n4121) );
  NOR2_X1 U3070 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4737), .ZN(n4736) );
  AND2_X1 U3071 ( .A1(n2864), .A2(n5265), .ZN(n5154) );
  INV_X1 U3072 ( .A(n4877), .ZN(n4976) );
  INV_X1 U3073 ( .A(n4991), .ZN(n5345) );
  OR2_X1 U3074 ( .A1(n4587), .A2(n4429), .ZN(n4803) );
  AND2_X1 U3075 ( .A1(n2864), .A2(n2945), .ZN(n5406) );
  AND2_X1 U3076 ( .A1(n2796), .A2(n2795), .ZN(n2800) );
  AND2_X1 U3077 ( .A1(n2865), .A2(n2810), .ZN(n2946) );
  AND2_X1 U3078 ( .A1(n2696), .A2(n2697), .ZN(n5225) );
  INV_X1 U3079 ( .A(n4870), .ZN(n4508) );
  AND2_X1 U3080 ( .A1(n4260), .A2(n4259), .ZN(n4809) );
  AND2_X1 U3081 ( .A1(n4247), .A2(n4246), .ZN(n4821) );
  NAND2_X1 U3082 ( .A1(n4272), .A2(n4271), .ZN(n4820) );
  NAND4_X1 U3083 ( .A1(n3465), .A2(n3464), .A3(n3463), .A4(n3462), .ZN(n4723)
         );
  OR2_X1 U3084 ( .A1(n5146), .A2(n2829), .ZN(n4773) );
  NAND2_X1 U3085 ( .A1(n2947), .A2(n5154), .ZN(n5339) );
  NAND2_X1 U3086 ( .A1(n3257), .A2(n5339), .ZN(n5341) );
  INV_X1 U3087 ( .A(n5410), .ZN(n5408) );
  INV_X1 U3088 ( .A(n5414), .ZN(n5411) );
  INV_X1 U3089 ( .A(n5130), .ZN(n5136) );
  AND2_X1 U3090 ( .A1(n2708), .A2(n2711), .ZN(n5108) );
  INV_X1 U3091 ( .A(n2836), .ZN(n5218) );
  INV_X1 U3092 ( .A(IR_REG_17__SCAN_IN), .ZN(n3942) );
  NOR2_X1 U3093 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2668)
         );
  NAND3_X1 U3094 ( .A1(n2669), .A2(n2744), .A3(n2771), .ZN(n2670) );
  NAND2_X1 U3095 ( .A1(n2751), .A2(IR_REG_31__SCAN_IN), .ZN(n2676) );
  INV_X1 U3096 ( .A(IR_REG_28__SCAN_IN), .ZN(n2675) );
  MUX2_X1 U3097 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2481), .Z(n4604) );
  MUX2_X1 U3098 ( .A(n2841), .B(DATAI_1_), .S(n2481), .Z(n3387) );
  XNOR2_X2 U3099 ( .A(n2680), .B(IR_REG_2__SCAN_IN), .ZN(n2839) );
  MUX2_X1 U3100 ( .A(n2839), .B(DATAI_2_), .S(n2481), .Z(n3264) );
  NAND2_X1 U3101 ( .A1(n2682), .A2(IR_REG_31__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3102 ( .A1(n2684), .A2(n2683), .ZN(n2686) );
  OR2_X1 U3103 ( .A1(n2684), .A2(n2683), .ZN(n2685) );
  MUX2_X1 U3104 ( .A(n5112), .B(DATAI_3_), .S(n2481), .Z(n5197) );
  NAND2_X1 U3105 ( .A1(n2686), .A2(IR_REG_31__SCAN_IN), .ZN(n2687) );
  XNOR2_X1 U3106 ( .A(n2687), .B(IR_REG_4__SCAN_IN), .ZN(n5111) );
  MUX2_X1 U3107 ( .A(n5111), .B(DATAI_4_), .S(n2481), .Z(n3373) );
  NAND2_X1 U3108 ( .A1(n3915), .A2(n2683), .ZN(n2688) );
  OR2_X1 U3109 ( .A1(n2682), .A2(n2688), .ZN(n2690) );
  NAND2_X1 U3110 ( .A1(n2690), .A2(IR_REG_31__SCAN_IN), .ZN(n2689) );
  MUX2_X1 U3111 ( .A(n2836), .B(DATAI_5_), .S(n2481), .Z(n3339) );
  INV_X1 U3112 ( .A(n2690), .ZN(n2692) );
  NAND2_X1 U3113 ( .A1(n2692), .A2(n2691), .ZN(n2694) );
  NAND2_X1 U3114 ( .A1(n2694), .A2(IR_REG_31__SCAN_IN), .ZN(n2693) );
  MUX2_X1 U3115 ( .A(IR_REG_31__SCAN_IN), .B(n2693), .S(IR_REG_6__SCAN_IN), 
        .Z(n2696) );
  INV_X1 U3116 ( .A(n2694), .ZN(n2695) );
  INV_X1 U3117 ( .A(IR_REG_6__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U3118 ( .A1(n2695), .A2(n3922), .ZN(n2697) );
  MUX2_X1 U3119 ( .A(n5225), .B(DATAI_6_), .S(n2481), .Z(n4342) );
  NAND2_X1 U3120 ( .A1(n2697), .A2(IR_REG_31__SCAN_IN), .ZN(n2699) );
  NAND2_X1 U3121 ( .A1(n2699), .A2(n2698), .ZN(n2701) );
  OR2_X1 U3122 ( .A1(n2699), .A2(n2698), .ZN(n2700) );
  MUX2_X1 U3123 ( .A(n5110), .B(DATAI_7_), .S(n2481), .Z(n3404) );
  NAND2_X1 U3124 ( .A1(n2701), .A2(IR_REG_31__SCAN_IN), .ZN(n2702) );
  XNOR2_X1 U3125 ( .A(n2702), .B(IR_REG_8__SCAN_IN), .ZN(n5109) );
  MUX2_X1 U3126 ( .A(n5109), .B(DATAI_8_), .S(n2481), .Z(n5250) );
  NAND2_X1 U3127 ( .A1(n2703), .A2(IR_REG_31__SCAN_IN), .ZN(n2704) );
  XNOR2_X1 U3128 ( .A(n2704), .B(IR_REG_9__SCAN_IN), .ZN(n3426) );
  MUX2_X1 U3129 ( .A(n3426), .B(DATAI_9_), .S(n2481), .Z(n3448) );
  NOR2_X1 U3130 ( .A1(n2742), .A2(n5094), .ZN(n2705) );
  NAND2_X1 U3131 ( .A1(n2705), .A2(IR_REG_11__SCAN_IN), .ZN(n2708) );
  INV_X1 U3132 ( .A(n2705), .ZN(n2707) );
  INV_X1 U3133 ( .A(IR_REG_11__SCAN_IN), .ZN(n2706) );
  NAND2_X1 U3134 ( .A1(n2707), .A2(n2706), .ZN(n2711) );
  MUX2_X1 U3135 ( .A(n5108), .B(DATAI_11_), .S(n2481), .Z(n3469) );
  NOR2_X1 U3136 ( .A1(n2703), .A2(IR_REG_9__SCAN_IN), .ZN(n2709) );
  OR2_X1 U3137 ( .A1(n2709), .A2(n5094), .ZN(n2710) );
  XNOR2_X1 U3138 ( .A(n2710), .B(IR_REG_10__SCAN_IN), .ZN(n3480) );
  MUX2_X1 U3139 ( .A(n3480), .B(DATAI_10_), .S(n2481), .Z(n4400) );
  NAND2_X1 U3140 ( .A1(n2711), .A2(IR_REG_31__SCAN_IN), .ZN(n2712) );
  XNOR2_X1 U3141 ( .A(n2712), .B(IR_REG_12__SCAN_IN), .ZN(n5107) );
  AND2_X1 U3142 ( .A1(n2742), .A2(n2715), .ZN(n2713) );
  NOR2_X1 U3143 ( .A1(n2713), .A2(n5094), .ZN(n2714) );
  MUX2_X1 U3144 ( .A(n5094), .B(n2714), .S(IR_REG_13__SCAN_IN), .Z(n2717) );
  AND2_X1 U3145 ( .A1(n2715), .A2(n3934), .ZN(n2728) );
  NAND2_X1 U3146 ( .A1(n2742), .A2(n2728), .ZN(n2719) );
  INV_X1 U3147 ( .A(n2719), .ZN(n2716) );
  MUX2_X1 U31480 ( .A(n4152), .B(DATAI_13_), .S(n2481), .Z(n5320) );
  NAND2_X1 U31490 ( .A1(n2719), .A2(IR_REG_31__SCAN_IN), .ZN(n2718) );
  XNOR2_X1 U3150 ( .A(n2718), .B(IR_REG_14__SCAN_IN), .ZN(n5106) );
  MUX2_X1 U3151 ( .A(n5106), .B(DATAI_14_), .S(n2481), .Z(n4464) );
  OR2_X1 U3152 ( .A1(n2719), .A2(IR_REG_14__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U3153 ( .A1(n2720), .A2(IR_REG_31__SCAN_IN), .ZN(n2723) );
  INV_X1 U3154 ( .A(n2723), .ZN(n2721) );
  NAND2_X1 U3155 ( .A1(n2721), .A2(IR_REG_15__SCAN_IN), .ZN(n2724) );
  INV_X1 U3156 ( .A(IR_REG_15__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U3157 ( .A1(n2723), .A2(n2722), .ZN(n2725) );
  MUX2_X1 U3158 ( .A(n4310), .B(DATAI_15_), .S(n2481), .Z(n5365) );
  NAND2_X1 U3159 ( .A1(n2725), .A2(IR_REG_31__SCAN_IN), .ZN(n2726) );
  XNOR2_X1 U3160 ( .A(n2726), .B(IR_REG_16__SCAN_IN), .ZN(n4312) );
  MUX2_X1 U3161 ( .A(n4312), .B(DATAI_16_), .S(n2481), .Z(n4518) );
  NAND2_X1 U3162 ( .A1(n2727), .A2(n3935), .ZN(n2730) );
  INV_X1 U3163 ( .A(n2728), .ZN(n2729) );
  NOR2_X1 U3164 ( .A1(n2730), .A2(n2729), .ZN(n2731) );
  NAND2_X1 U3165 ( .A1(n2731), .A2(n2742), .ZN(n2733) );
  NAND2_X1 U3166 ( .A1(n2733), .A2(IR_REG_31__SCAN_IN), .ZN(n2732) );
  XNOR2_X1 U3167 ( .A(n2732), .B(IR_REG_17__SCAN_IN), .ZN(n5105) );
  MUX2_X1 U3168 ( .A(n5105), .B(DATAI_17_), .S(n2481), .Z(n4369) );
  XNOR2_X1 U3169 ( .A(n2734), .B(IR_REG_18__SCAN_IN), .ZN(n5104) );
  MUX2_X1 U3170 ( .A(n5104), .B(DATAI_18_), .S(n2481), .Z(n4984) );
  NAND2_X1 U3171 ( .A1(n2734), .A2(n3755), .ZN(n2735) );
  NAND2_X1 U3172 ( .A1(n2735), .A2(IR_REG_31__SCAN_IN), .ZN(n2736) );
  NAND2_X1 U3173 ( .A1(n2736), .A2(n3754), .ZN(n2739) );
  OR2_X1 U3174 ( .A1(n2736), .A2(n3754), .ZN(n2737) );
  INV_X1 U3175 ( .A(n4767), .ZN(n5265) );
  MUX2_X1 U3176 ( .A(n5265), .B(DATAI_19_), .S(n2481), .Z(n4962) );
  NAND2_X1 U3177 ( .A1(n2481), .A2(DATAI_20_), .ZN(n4945) );
  INV_X1 U3178 ( .A(n4945), .ZN(n4922) );
  NAND2_X1 U3179 ( .A1(n2481), .A2(DATAI_21_), .ZN(n4914) );
  NAND2_X1 U3180 ( .A1(n2481), .A2(DATAI_22_), .ZN(n4894) );
  INV_X1 U3181 ( .A(n4894), .ZN(n4882) );
  NAND2_X1 U3182 ( .A1(n2481), .A2(DATAI_23_), .ZN(n4868) );
  INV_X1 U3183 ( .A(n4868), .ZN(n4874) );
  NAND2_X1 U3184 ( .A1(n2481), .A2(DATAI_24_), .ZN(n4851) );
  NAND2_X1 U3185 ( .A1(n2481), .A2(DATAI_25_), .ZN(n4362) );
  NAND2_X1 U3186 ( .A1(n2481), .A2(DATAI_26_), .ZN(n4824) );
  INV_X1 U3187 ( .A(n4824), .ZN(n4830) );
  NAND2_X1 U3188 ( .A1(n2481), .A2(DATAI_27_), .ZN(n4808) );
  INV_X1 U3189 ( .A(n4808), .ZN(n4796) );
  NAND2_X1 U3190 ( .A1(n2481), .A2(DATAI_28_), .ZN(n4781) );
  AND2_X1 U3191 ( .A1(n2481), .A2(DATAI_29_), .ZN(n4435) );
  INV_X1 U3192 ( .A(n4435), .ZN(n4439) );
  AND2_X1 U3193 ( .A1(n2481), .A2(DATAI_30_), .ZN(n5397) );
  AND2_X1 U3194 ( .A1(n2481), .A2(DATAI_31_), .ZN(n4597) );
  XNOR2_X2 U3195 ( .A(n2740), .B(n3947), .ZN(n2864) );
  INV_X1 U3196 ( .A(n2745), .ZN(n2749) );
  NAND2_X1 U3197 ( .A1(n2749), .A2(IR_REG_31__SCAN_IN), .ZN(n2743) );
  MUX2_X1 U3198 ( .A(IR_REG_31__SCAN_IN), .B(n2743), .S(IR_REG_22__SCAN_IN), 
        .Z(n2746) );
  NAND2_X1 U3199 ( .A1(n2747), .A2(IR_REG_31__SCAN_IN), .ZN(n2748) );
  MUX2_X1 U3200 ( .A(IR_REG_31__SCAN_IN), .B(n2748), .S(IR_REG_21__SCAN_IN), 
        .Z(n2750) );
  NAND2_X1 U3201 ( .A1(n2750), .A2(n2749), .ZN(n4592) );
  INV_X1 U3202 ( .A(IR_REG_30__SCAN_IN), .ZN(n3774) );
  NAND2_X1 U3203 ( .A1(n2752), .A2(IR_REG_31__SCAN_IN), .ZN(n2753) );
  INV_X1 U3204 ( .A(n2754), .ZN(n5095) );
  NAND2_X1 U3205 ( .A1(n2479), .A2(REG1_REG_31__SCAN_IN), .ZN(n2760) );
  AND2_X2 U3206 ( .A1(n5097), .A2(n2757), .ZN(n3212) );
  NAND2_X1 U3207 ( .A1(n3212), .A2(REG2_REG_31__SCAN_IN), .ZN(n2759) );
  NAND2_X1 U3208 ( .A1(n3106), .A2(REG0_REG_31__SCAN_IN), .ZN(n2758) );
  AND3_X1 U3209 ( .A1(n2760), .A2(n2759), .A3(n2758), .ZN(n4594) );
  INV_X1 U32100 ( .A(n4594), .ZN(n4717) );
  AND2_X1 U32110 ( .A1(n5102), .A2(n5103), .ZN(n2935) );
  NAND2_X1 U32120 ( .A1(n2761), .A2(n2935), .ZN(n5184) );
  INV_X1 U32130 ( .A(B_REG_SCAN_IN), .ZN(n2762) );
  NOR2_X1 U32140 ( .A1(n5137), .A2(n2762), .ZN(n2763) );
  NOR2_X1 U32150 ( .A1(n5184), .A2(n2763), .ZN(n4436) );
  NAND2_X1 U32160 ( .A1(n4717), .A2(n4436), .ZN(n5399) );
  NAND2_X1 U32170 ( .A1(n4597), .A2(n5396), .ZN(n2764) );
  AND2_X1 U32180 ( .A1(n5399), .A2(n2764), .ZN(n5418) );
  INV_X1 U32190 ( .A(n5418), .ZN(n2765) );
  AOI21_X1 U32200 ( .B1(n5416), .B2(n5406), .A(n2765), .ZN(n2802) );
  NAND2_X1 U32210 ( .A1(n2864), .A2(n4767), .ZN(n2940) );
  NAND2_X1 U32220 ( .A1(n2940), .A2(n2935), .ZN(n2995) );
  NAND2_X1 U32230 ( .A1(n2777), .A2(n3952), .ZN(n2766) );
  NAND2_X1 U32240 ( .A1(n2773), .A2(n2771), .ZN(n2768) );
  NAND2_X1 U32250 ( .A1(n2768), .A2(IR_REG_31__SCAN_IN), .ZN(n2769) );
  NAND2_X1 U32260 ( .A1(n2773), .A2(n2772), .ZN(n2775) );
  INV_X1 U32270 ( .A(n2781), .ZN(n5101) );
  XNOR2_X1 U32280 ( .A(n2777), .B(n3952), .ZN(n2994) );
  NAND2_X1 U32290 ( .A1(n2995), .A2(n2946), .ZN(n2943) );
  NAND2_X1 U32300 ( .A1(n2781), .A2(B_REG_SCAN_IN), .ZN(n2779) );
  MUX2_X1 U32310 ( .A(n2779), .B(B_REG_SCAN_IN), .S(n2778), .Z(n2780) );
  NAND2_X1 U32320 ( .A1(n2780), .A2(n5100), .ZN(n2927) );
  INV_X1 U32330 ( .A(n5100), .ZN(n2798) );
  NAND2_X1 U32340 ( .A1(n2798), .A2(n2781), .ZN(n2925) );
  OAI21_X1 U32350 ( .B1(n2927), .B2(D_REG_1__SCAN_IN), .A(n2925), .ZN(n2782)
         );
  INV_X1 U32360 ( .A(n2782), .ZN(n2783) );
  NOR2_X1 U32370 ( .A1(n2943), .A2(n2783), .ZN(n2796) );
  INV_X1 U32380 ( .A(n2927), .ZN(n2794) );
  NOR4_X1 U32390 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2787) );
  NOR4_X1 U32400 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2786) );
  NOR4_X1 U32410 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2785) );
  NOR4_X1 U32420 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2784) );
  AND4_X1 U32430 ( .A1(n2787), .A2(n2786), .A3(n2785), .A4(n2784), .ZN(n2793)
         );
  NOR2_X1 U32440 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_12__SCAN_IN), .ZN(n2791)
         );
  NOR4_X1 U32450 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2790) );
  NOR4_X1 U32460 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2789) );
  NOR4_X1 U32470 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2788) );
  AND4_X1 U32480 ( .A1(n2791), .A2(n2790), .A3(n2789), .A4(n2788), .ZN(n2792)
         );
  NAND2_X1 U32490 ( .A1(n2793), .A2(n2792), .ZN(n2924) );
  AOI22_X1 U32500 ( .A1(n2945), .A2(n5154), .B1(n2794), .B2(n2924), .ZN(n2795)
         );
  INV_X1 U32510 ( .A(n2778), .ZN(n2797) );
  NAND2_X1 U32520 ( .A1(n2798), .A2(n2797), .ZN(n2807) );
  OAI21_X1 U32530 ( .B1(n2927), .B2(D_REG_0__SCAN_IN), .A(n2807), .ZN(n3255)
         );
  INV_X1 U32540 ( .A(n3255), .ZN(n2928) );
  AND2_X2 U32550 ( .A1(n2800), .A2(n2928), .ZN(n5410) );
  NOR2_X1 U32560 ( .A1(n5410), .A2(REG1_REG_31__SCAN_IN), .ZN(n2799) );
  AOI21_X1 U32570 ( .B1(n2802), .B2(n5410), .A(n2799), .ZN(U3549) );
  AND2_X2 U32580 ( .A1(n2800), .A2(n3255), .ZN(n5414) );
  NOR2_X1 U32590 ( .A1(n5414), .A2(REG0_REG_31__SCAN_IN), .ZN(n2801) );
  AOI21_X1 U32600 ( .B1(n2802), .B2(n5414), .A(n2801), .ZN(U3517) );
  INV_X1 U32610 ( .A(n2810), .ZN(n2803) );
  NOR2_X1 U32620 ( .A1(n2865), .A2(n2803), .ZN(U4043) );
  INV_X1 U32630 ( .A(DATAI_28_), .ZN(n2804) );
  MUX2_X1 U32640 ( .A(n2804), .B(n2761), .S(STATE_REG_SCAN_IN), .Z(n2805) );
  INV_X1 U32650 ( .A(n2805), .ZN(U3324) );
  INV_X1 U32660 ( .A(DATAI_23_), .ZN(n2806) );
  AOI21_X1 U32670 ( .B1(n2806), .B2(U3149), .A(n2810), .ZN(U3329) );
  NAND2_X1 U32680 ( .A1(n2946), .A2(n2927), .ZN(n5130) );
  INV_X1 U32690 ( .A(D_REG_0__SCAN_IN), .ZN(n2809) );
  INV_X1 U32700 ( .A(n2807), .ZN(n2808) );
  AOI22_X1 U32710 ( .A1(n5130), .A2(n2809), .B1(n2808), .B2(n2810), .ZN(U3458)
         );
  INV_X1 U32720 ( .A(D_REG_1__SCAN_IN), .ZN(n2923) );
  INV_X1 U32730 ( .A(n2925), .ZN(n2811) );
  AOI22_X1 U32740 ( .A1(n5130), .A2(n2923), .B1(n2811), .B2(n2810), .ZN(U3459)
         );
  INV_X1 U32750 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2831) );
  NAND2_X1 U32760 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(
        n2957) );
  INV_X1 U32770 ( .A(n2841), .ZN(n2840) );
  INV_X1 U32780 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3389) );
  NOR2_X1 U32790 ( .A1(n2957), .A2(n2955), .ZN(n2956) );
  INV_X1 U32800 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2812) );
  NAND2_X1 U32810 ( .A1(n2839), .A2(REG2_REG_2__SCAN_IN), .ZN(n2813) );
  INV_X1 U32820 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2856) );
  OR2_X1 U32830 ( .A1(n2856), .A2(n3014), .ZN(n2814) );
  NOR2_X1 U32840 ( .A1(n2855), .A2(n2814), .ZN(n2817) );
  AND2_X1 U32850 ( .A1(n2815), .A2(n5112), .ZN(n2818) );
  NOR2_X1 U32860 ( .A1(n2817), .A2(n2816), .ZN(n2822) );
  NAND2_X1 U32870 ( .A1(n2820), .A2(n2819), .ZN(n2821) );
  NAND2_X1 U32880 ( .A1(n2822), .A2(n2821), .ZN(n3008) );
  INV_X1 U32890 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3375) );
  INV_X1 U32900 ( .A(n2822), .ZN(n2823) );
  INV_X1 U32910 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2824) );
  AOI22_X1 U32920 ( .A1(n2836), .A2(n2824), .B1(REG2_REG_5__SCAN_IN), .B2(
        n5218), .ZN(n2967) );
  XNOR2_X1 U32930 ( .A(n3027), .B(n2826), .ZN(n2830) );
  NOR2_X2 U32940 ( .A1(n2830), .A2(n2831), .ZN(n3028) );
  NAND2_X1 U32950 ( .A1(n2935), .A2(n2994), .ZN(n2827) );
  NAND2_X1 U32960 ( .A1(n2481), .A2(n2827), .ZN(n2832) );
  OR2_X1 U32970 ( .A1(n2994), .A2(U3149), .ZN(n4715) );
  INV_X1 U32980 ( .A(n4715), .ZN(n2828) );
  NOR2_X1 U32990 ( .A1(n2946), .A2(n2828), .ZN(n2833) );
  OR2_X1 U33000 ( .A1(n2832), .A2(n2833), .ZN(n5146) );
  OR2_X1 U33010 ( .A1(n2761), .A2(n5137), .ZN(n2829) );
  AOI211_X1 U33020 ( .C1(n2831), .C2(n2830), .A(n3028), .B(n4773), .ZN(n2850)
         );
  INV_X1 U33030 ( .A(n2761), .ZN(n2999) );
  INV_X1 U33040 ( .A(n2832), .ZN(n2834) );
  NOR2_X1 U33050 ( .A1(STATE_REG_SCAN_IN), .A2(n3083), .ZN(n2835) );
  AOI21_X1 U33060 ( .B1(n5143), .B2(ADDR_REG_6__SCAN_IN), .A(n2835), .ZN(n2848) );
  INV_X1 U33070 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2837) );
  MUX2_X1 U33080 ( .A(REG1_REG_5__SCAN_IN), .B(n2837), .S(n2836), .Z(n2971) );
  INV_X1 U33090 ( .A(REG1_REG_2__SCAN_IN), .ZN(n5178) );
  INV_X1 U33100 ( .A(REG1_REG_1__SCAN_IN), .ZN(n5170) );
  MUX2_X1 U33110 ( .A(REG1_REG_1__SCAN_IN), .B(n5170), .S(n2841), .Z(n2960) );
  NAND3_X1 U33120 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .A3(
        n2960), .ZN(n2959) );
  OAI21_X1 U33130 ( .B1(n5170), .B2(n2840), .A(n2959), .ZN(n2879) );
  NAND2_X1 U33140 ( .A1(n2880), .A2(n2879), .ZN(n2842) );
  INV_X1 U33150 ( .A(n5111), .ZN(n3014) );
  INV_X1 U33160 ( .A(REG1_REG_4__SCAN_IN), .ZN(n5214) );
  OAI21_X1 U33170 ( .B1(n2845), .B2(n3014), .A(n3009), .ZN(n2972) );
  NAND2_X1 U33180 ( .A1(n2971), .A2(n2972), .ZN(n2970) );
  INV_X1 U33190 ( .A(n5137), .ZN(n5099) );
  OR2_X1 U33200 ( .A1(n5146), .A2(n5099), .ZN(n4756) );
  INV_X1 U33210 ( .A(n4756), .ZN(n4770) );
  NAND2_X1 U33220 ( .A1(REG1_REG_6__SCAN_IN), .A2(n2846), .ZN(n3021) );
  OAI211_X1 U33230 ( .C1(REG1_REG_6__SCAN_IN), .C2(n2846), .A(n4770), .B(n3021), .ZN(n2847) );
  OAI211_X1 U33240 ( .C1(n4768), .C2(n2826), .A(n2848), .B(n2847), .ZN(n2849)
         );
  OR2_X1 U33250 ( .A1(n2850), .A2(n2849), .ZN(U3246) );
  INV_X1 U33260 ( .A(n4768), .ZN(n4753) );
  XNOR2_X1 U33270 ( .A(n2851), .B(REG1_REG_3__SCAN_IN), .ZN(n2853) );
  INV_X1 U33280 ( .A(REG3_REG_3__SCAN_IN), .ZN(n5203) );
  NOR2_X1 U33290 ( .A1(n5203), .A2(STATE_REG_SCAN_IN), .ZN(n3000) );
  AOI21_X1 U33300 ( .B1(n5143), .B2(ADDR_REG_3__SCAN_IN), .A(n3000), .ZN(n2852) );
  OAI21_X1 U33310 ( .B1(n2853), .B2(n4756), .A(n2852), .ZN(n2858) );
  AOI211_X1 U33320 ( .C1(n2856), .C2(n2855), .A(n2854), .B(n4773), .ZN(n2857)
         );
  AOI211_X1 U33330 ( .C1(n4753), .C2(n5112), .A(n2858), .B(n2857), .ZN(n2859)
         );
  INV_X1 U33340 ( .A(n2859), .ZN(U3243) );
  NOR2_X1 U33350 ( .A1(n5143), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U33360 ( .A1(n4287), .A2(REG3_REG_0__SCAN_IN), .ZN(n2863) );
  NAND2_X1 U33370 ( .A1(n3106), .A2(REG0_REG_0__SCAN_IN), .ZN(n2862) );
  NAND2_X1 U33380 ( .A1(n2480), .A2(REG1_REG_0__SCAN_IN), .ZN(n2861) );
  NAND2_X1 U33390 ( .A1(n3212), .A2(REG2_REG_0__SCAN_IN), .ZN(n2860) );
  NAND2_X1 U33400 ( .A1(n4604), .A2(n3090), .ZN(n2866) );
  NAND2_X1 U33410 ( .A1(n4735), .A2(n3090), .ZN(n2868) );
  NAND2_X1 U33420 ( .A1(n4604), .A2(n4103), .ZN(n2867) );
  NAND2_X1 U33430 ( .A1(n2868), .A2(n2867), .ZN(n2903) );
  NAND2_X1 U33440 ( .A1(n2872), .A2(n2903), .ZN(n2871) );
  INV_X1 U33450 ( .A(n2865), .ZN(n2869) );
  NAND3_X1 U33460 ( .A1(n2869), .A2(IR_REG_0__SCAN_IN), .A3(
        REG1_REG_0__SCAN_IN), .ZN(n2870) );
  NAND2_X1 U33470 ( .A1(n2871), .A2(n2870), .ZN(n2902) );
  INV_X1 U33480 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2873) );
  AOI21_X1 U33490 ( .B1(n5148), .B2(n2873), .A(n2865), .ZN(n2874) );
  NOR3_X1 U33500 ( .A1(n2903), .A2(n2872), .A3(n2874), .ZN(n2875) );
  OR2_X1 U33510 ( .A1(n2902), .A2(n2875), .ZN(n2954) );
  INV_X1 U33520 ( .A(n2957), .ZN(n2876) );
  MUX2_X1 U3353 ( .A(n2954), .B(n2876), .S(n5099), .Z(n2878) );
  INV_X1 U33540 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2877) );
  AOI21_X1 U3355 ( .B1(n5099), .B2(n2877), .A(n2761), .ZN(n5139) );
  INV_X1 U3356 ( .A(IR_REG_0__SCAN_IN), .ZN(n5148) );
  NOR2_X1 U3357 ( .A1(n5139), .A2(IR_REG_0__SCAN_IN), .ZN(n5138) );
  INV_X2 U3358 ( .A(U4043), .ZN(n4734) );
  AOI211_X1 U3359 ( .C1(n2878), .C2(n2999), .A(n5138), .B(n4734), .ZN(n3018)
         );
  XOR2_X1 U3360 ( .A(n2880), .B(n2879), .Z(n2886) );
  INV_X1 U3361 ( .A(n2881), .ZN(n2882) );
  AOI211_X1 U3362 ( .C1(n2884), .C2(n2883), .A(n2882), .B(n4773), .ZN(n2885)
         );
  AOI21_X1 U3363 ( .B1(n2886), .B2(n4770), .A(n2885), .ZN(n2888) );
  AOI22_X1 U3364 ( .A1(n5143), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2887) );
  OAI211_X1 U3365 ( .C1(n2838), .C2(n4768), .A(n2888), .B(n2887), .ZN(n2889)
         );
  OR2_X1 U3366 ( .A1(n3018), .A2(n2889), .ZN(U3242) );
  NAND2_X1 U3367 ( .A1(n2480), .A2(REG1_REG_2__SCAN_IN), .ZN(n2893) );
  NAND2_X1 U3368 ( .A1(n3212), .A2(REG2_REG_2__SCAN_IN), .ZN(n2892) );
  NAND2_X1 U3369 ( .A1(n4287), .A2(REG3_REG_2__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U3370 ( .A1(n3106), .A2(REG0_REG_2__SCAN_IN), .ZN(n2890) );
  NAND2_X1 U3371 ( .A1(n4733), .A2(n3090), .ZN(n2895) );
  NAND2_X1 U3372 ( .A1(n3264), .A2(n4103), .ZN(n2894) );
  NAND2_X1 U3373 ( .A1(n2895), .A2(n2894), .ZN(n2899) );
  XNOR2_X1 U3374 ( .A(n2896), .B(n4361), .ZN(n2897) );
  NAND2_X1 U3375 ( .A1(n2897), .A2(n4767), .ZN(n3273) );
  AND2_X4 U3376 ( .A1(n2898), .A2(n3273), .ZN(n3093) );
  XNOR2_X1 U3377 ( .A(n2899), .B(n3296), .ZN(n2977) );
  NAND2_X1 U3378 ( .A1(n4733), .A2(n2986), .ZN(n2901) );
  INV_X4 U3379 ( .A(n4273), .ZN(n4235) );
  NAND2_X1 U3380 ( .A1(n3264), .A2(n4235), .ZN(n2900) );
  NAND2_X1 U3381 ( .A1(n2901), .A2(n2900), .ZN(n2978) );
  XNOR2_X1 U3382 ( .A(n2977), .B(n2978), .ZN(n2922) );
  INV_X1 U3383 ( .A(n2902), .ZN(n2904) );
  NAND2_X1 U3384 ( .A1(n2904), .A2(n2664), .ZN(n4413) );
  NAND2_X1 U3385 ( .A1(n4287), .A2(REG3_REG_1__SCAN_IN), .ZN(n2908) );
  NAND2_X1 U3386 ( .A1(n3212), .A2(REG2_REG_1__SCAN_IN), .ZN(n2907) );
  NAND2_X1 U3387 ( .A1(n2480), .A2(REG1_REG_1__SCAN_IN), .ZN(n2906) );
  NAND2_X1 U3388 ( .A1(n3106), .A2(REG0_REG_1__SCAN_IN), .ZN(n2905) );
  NAND2_X1 U3389 ( .A1(n2934), .A2(n3090), .ZN(n2910) );
  NAND2_X1 U3390 ( .A1(n3387), .A2(n2608), .ZN(n2909) );
  NAND2_X1 U3391 ( .A1(n2910), .A2(n2909), .ZN(n2911) );
  NAND2_X1 U3392 ( .A1(n2934), .A2(n2986), .ZN(n2913) );
  NAND2_X1 U3393 ( .A1(n3387), .A2(n3090), .ZN(n2912) );
  NAND2_X1 U3394 ( .A1(n2913), .A2(n2912), .ZN(n2915) );
  NAND2_X1 U3395 ( .A1(n4413), .A2(n4415), .ZN(n4414) );
  INV_X1 U3396 ( .A(n2914), .ZN(n2916) );
  NAND2_X1 U3397 ( .A1(n2916), .A2(n2915), .ZN(n2917) );
  NAND2_X1 U3398 ( .A1(n4414), .A2(n2917), .ZN(n2921) );
  INV_X1 U3399 ( .A(n2922), .ZN(n2919) );
  INV_X1 U3400 ( .A(n2921), .ZN(n2918) );
  NAND2_X1 U3401 ( .A1(n2919), .A2(n2918), .ZN(n2982) );
  INV_X1 U3402 ( .A(n2982), .ZN(n2920) );
  AOI21_X1 U3403 ( .B1(n2922), .B2(n2921), .A(n2920), .ZN(n2951) );
  NOR2_X1 U3404 ( .A1(n2924), .A2(n2923), .ZN(n2926) );
  OAI21_X1 U3405 ( .B1(n2927), .B2(n2926), .A(n2925), .ZN(n2936) );
  INV_X1 U3406 ( .A(n2936), .ZN(n3256) );
  AND3_X1 U3407 ( .A1(n2928), .A2(n3256), .A3(n2946), .ZN(n2944) );
  AOI21_X1 U3408 ( .B1(n2940), .B2(n2945), .A(n2935), .ZN(n2929) );
  NAND2_X1 U3409 ( .A1(n2944), .A2(n2929), .ZN(n5315) );
  NAND2_X1 U3410 ( .A1(n2480), .A2(REG1_REG_3__SCAN_IN), .ZN(n2933) );
  NAND2_X1 U3411 ( .A1(n3212), .A2(REG2_REG_3__SCAN_IN), .ZN(n2932) );
  NAND2_X1 U3412 ( .A1(n4287), .A2(n5203), .ZN(n2931) );
  NAND2_X1 U3413 ( .A1(n3106), .A2(REG0_REG_3__SCAN_IN), .ZN(n2930) );
  INV_X1 U3414 ( .A(n2935), .ZN(n2937) );
  OR2_X1 U3415 ( .A1(n2761), .A2(n2937), .ZN(n5186) );
  OAI22_X1 U3416 ( .A1(n3368), .A2(n5184), .B1(n5151), .B2(n5186), .ZN(n3261)
         );
  OR2_X1 U3417 ( .A1(n3255), .A2(n2936), .ZN(n2942) );
  INV_X1 U3418 ( .A(n2942), .ZN(n2939) );
  NOR2_X1 U3419 ( .A1(n2943), .A2(n2937), .ZN(n2938) );
  NAND2_X1 U3420 ( .A1(n5406), .A2(n2940), .ZN(n2941) );
  NAND2_X1 U3421 ( .A1(n2942), .A2(n2941), .ZN(n2997) );
  INV_X1 U3422 ( .A(n2943), .ZN(n4712) );
  NAND2_X1 U3423 ( .A1(n2997), .A2(n4712), .ZN(n4416) );
  AOI22_X1 U3424 ( .A1(n3261), .A2(n5359), .B1(REG3_REG_2__SCAN_IN), .B2(n4416), .ZN(n2950) );
  NAND2_X1 U3425 ( .A1(n2944), .A2(n5396), .ZN(n2948) );
  AND2_X1 U3426 ( .A1(n2946), .A2(n2945), .ZN(n2947) );
  NAND2_X1 U3427 ( .A1(n2948), .A2(n5339), .ZN(n5364) );
  NAND2_X1 U3428 ( .A1(n5364), .A2(n3264), .ZN(n2949) );
  OAI211_X1 U3429 ( .C1(n2951), .C2(n5315), .A(n2950), .B(n2949), .ZN(U3234)
         );
  NAND2_X1 U3430 ( .A1(n5359), .A2(n2761), .ZN(n4555) );
  INV_X1 U3431 ( .A(n4555), .ZN(n4547) );
  AOI22_X1 U3432 ( .A1(n4547), .A2(n2934), .B1(REG3_REG_0__SCAN_IN), .B2(n4416), .ZN(n2953) );
  NAND2_X1 U3433 ( .A1(n5364), .A2(n4604), .ZN(n2952) );
  OAI211_X1 U3434 ( .C1(n2954), .C2(n5315), .A(n2953), .B(n2952), .ZN(U3229)
         );
  AOI211_X1 U3435 ( .C1(n2957), .C2(n2955), .A(n2956), .B(n4773), .ZN(n2965)
         );
  INV_X1 U3436 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3388) );
  NOR2_X1 U3437 ( .A1(STATE_REG_SCAN_IN), .A2(n3388), .ZN(n2958) );
  AOI21_X1 U3438 ( .B1(n5143), .B2(ADDR_REG_1__SCAN_IN), .A(n2958), .ZN(n2963)
         );
  NOR2_X1 U3439 ( .A1(n5148), .A2(n2873), .ZN(n2961) );
  OAI211_X1 U3440 ( .C1(n2961), .C2(n2960), .A(n4770), .B(n2959), .ZN(n2962)
         );
  OAI211_X1 U3441 ( .C1(n4768), .C2(n2840), .A(n2963), .B(n2962), .ZN(n2964)
         );
  OR2_X1 U3442 ( .A1(n2965), .A2(n2964), .ZN(U3241) );
  AOI211_X1 U3443 ( .C1(n2968), .C2(n2967), .A(n2966), .B(n4773), .ZN(n2976)
         );
  INV_X1 U3444 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3149) );
  NOR2_X1 U3445 ( .A1(STATE_REG_SCAN_IN), .A2(n3149), .ZN(n2969) );
  AOI21_X1 U3446 ( .B1(n5143), .B2(ADDR_REG_5__SCAN_IN), .A(n2969), .ZN(n2974)
         );
  OAI211_X1 U3447 ( .C1(n2972), .C2(n2971), .A(n4770), .B(n2970), .ZN(n2973)
         );
  OAI211_X1 U3448 ( .C1(n4768), .C2(n5218), .A(n2974), .B(n2973), .ZN(n2975)
         );
  OR2_X1 U3449 ( .A1(n2976), .A2(n2975), .ZN(U3245) );
  INV_X1 U3450 ( .A(n2977), .ZN(n2980) );
  INV_X1 U3451 ( .A(n2978), .ZN(n2979) );
  NAND2_X1 U3452 ( .A1(n2980), .A2(n2979), .ZN(n2981) );
  NAND2_X1 U3453 ( .A1(n2982), .A2(n2981), .ZN(n3062) );
  NAND2_X1 U3454 ( .A1(n4732), .A2(n4235), .ZN(n2984) );
  NAND2_X1 U3455 ( .A1(n5197), .A2(n4103), .ZN(n2983) );
  NAND2_X1 U3456 ( .A1(n2984), .A2(n2983), .ZN(n2985) );
  XNOR2_X1 U3457 ( .A(n2985), .B(n3093), .ZN(n3070) );
  NAND2_X1 U34580 ( .A1(n4732), .A2(n4239), .ZN(n2988) );
  NAND2_X1 U34590 ( .A1(n5197), .A2(n3090), .ZN(n2987) );
  NAND2_X1 U3460 ( .A1(n2988), .A2(n2987), .ZN(n3068) );
  XNOR2_X1 U3461 ( .A(n3070), .B(n3068), .ZN(n3061) );
  XNOR2_X1 U3462 ( .A(n3062), .B(n3061), .ZN(n3005) );
  INV_X1 U3463 ( .A(n5364), .ZN(n4542) );
  INV_X1 U3464 ( .A(n5197), .ZN(n3338) );
  NAND2_X1 U3465 ( .A1(n3212), .A2(REG2_REG_4__SCAN_IN), .ZN(n2993) );
  NOR2_X1 U3466 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2989) );
  NOR2_X1 U34670 ( .A1(n3073), .A2(n2989), .ZN(n3159) );
  NAND2_X1 U3468 ( .A1(n4287), .A2(n3159), .ZN(n2992) );
  NAND2_X1 U34690 ( .A1(n2480), .A2(REG1_REG_4__SCAN_IN), .ZN(n2991) );
  NAND2_X1 U3470 ( .A1(n3106), .A2(REG0_REG_4__SCAN_IN), .ZN(n2990) );
  NAND4_X1 U34710 ( .A1(n2993), .A2(n2992), .A3(n2991), .A4(n2990), .ZN(n4731)
         );
  INV_X1 U3472 ( .A(n4731), .ZN(n5185) );
  OAI22_X1 U34730 ( .A1(n4542), .A2(n3338), .B1(n4555), .B2(n5185), .ZN(n3004)
         );
  AND3_X1 U3474 ( .A1(n2995), .A2(n2865), .A3(n2994), .ZN(n2996) );
  NAND2_X1 U34750 ( .A1(n2997), .A2(n2996), .ZN(n2998) );
  NAND2_X1 U3476 ( .A1(n2998), .A2(STATE_REG_SCAN_IN), .ZN(n5370) );
  NAND2_X1 U34770 ( .A1(n4558), .A2(n4733), .ZN(n3002) );
  INV_X1 U3478 ( .A(n3000), .ZN(n3001) );
  OAI211_X1 U34790 ( .C1(REG3_REG_3__SCAN_IN), .C2(n5370), .A(n3002), .B(n3001), .ZN(n3003) );
  AOI211_X1 U3480 ( .C1(n3005), .C2(n5366), .A(n3004), .B(n3003), .ZN(n3006)
         );
  INV_X1 U34810 ( .A(n3006), .ZN(U3215) );
  AOI211_X1 U3482 ( .C1(n3375), .C2(n3008), .A(n3007), .B(n4773), .ZN(n3017)
         );
  INV_X1 U34830 ( .A(n3009), .ZN(n3010) );
  AOI211_X1 U3484 ( .C1(n5214), .C2(n3011), .A(n3010), .B(n4756), .ZN(n3016)
         );
  INV_X1 U34850 ( .A(REG3_REG_4__SCAN_IN), .ZN(n3012) );
  NOR2_X1 U3486 ( .A1(n3012), .A2(STATE_REG_SCAN_IN), .ZN(n3160) );
  AOI21_X1 U34870 ( .B1(n5143), .B2(ADDR_REG_4__SCAN_IN), .A(n3160), .ZN(n3013) );
  OAI21_X1 U3488 ( .B1(n3014), .B2(n4768), .A(n3013), .ZN(n3015) );
  OR4_X1 U34890 ( .A1(n3018), .A2(n3017), .A3(n3016), .A4(n3015), .ZN(U3244)
         );
  INV_X1 U3490 ( .A(n5110), .ZN(n3036) );
  NAND2_X1 U34910 ( .A1(n5225), .A2(n3019), .ZN(n3020) );
  NAND2_X1 U3492 ( .A1(n3021), .A2(n3020), .ZN(n3023) );
  INV_X1 U34930 ( .A(n3023), .ZN(n3025) );
  INV_X1 U3494 ( .A(REG1_REG_7__SCAN_IN), .ZN(n5239) );
  MUX2_X1 U34950 ( .A(n5239), .B(REG1_REG_7__SCAN_IN), .S(n5110), .Z(n3024) );
  AOI211_X1 U3496 ( .C1(n3025), .C2(n3024), .A(n4756), .B(n2487), .ZN(n3026)
         );
  INV_X1 U34970 ( .A(n3026), .ZN(n3035) );
  INV_X1 U3498 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3029) );
  MUX2_X1 U34990 ( .A(n3029), .B(REG2_REG_7__SCAN_IN), .S(n5110), .Z(n3031) );
  INV_X1 U3500 ( .A(n3041), .ZN(n3030) );
  NAND2_X1 U35010 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n3286) );
  INV_X1 U3502 ( .A(n3286), .ZN(n3032) );
  AOI211_X1 U35030 ( .C1(n5143), .C2(ADDR_REG_7__SCAN_IN), .A(n3033), .B(n3032), .ZN(n3034) );
  OAI211_X1 U3504 ( .C1(n4768), .C2(n3036), .A(n3035), .B(n3034), .ZN(U3247)
         );
  XNOR2_X1 U35050 ( .A(n3233), .B(REG1_REG_8__SCAN_IN), .ZN(n3048) );
  INV_X1 U35060 ( .A(n5109), .ZN(n3234) );
  NOR2_X1 U35070 ( .A1(STATE_REG_SCAN_IN), .A2(n3141), .ZN(n3038) );
  AOI21_X1 U35080 ( .B1(n5143), .B2(ADDR_REG_8__SCAN_IN), .A(n3038), .ZN(n3039) );
  OAI21_X1 U35090 ( .B1(n3234), .B2(n4768), .A(n3039), .ZN(n3047) );
  INV_X1 U35100 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3045) );
  NAND2_X1 U35110 ( .A1(n5110), .A2(REG2_REG_7__SCAN_IN), .ZN(n3040) );
  INV_X1 U35120 ( .A(n3042), .ZN(n3043) );
  AOI211_X1 U35130 ( .C1(n3045), .C2(n3044), .A(n3228), .B(n4773), .ZN(n3046)
         );
  AOI211_X1 U35140 ( .C1(n4770), .C2(n3048), .A(n3047), .B(n3046), .ZN(n3049)
         );
  INV_X1 U35150 ( .A(n3049), .ZN(U3248) );
  NAND2_X1 U35160 ( .A1(n3105), .A2(n3141), .ZN(n3050) );
  NAND2_X1 U35170 ( .A1(n3133), .A2(n3050), .ZN(n5269) );
  NAND2_X1 U35180 ( .A1(n2479), .A2(REG1_REG_8__SCAN_IN), .ZN(n3055) );
  NAND2_X1 U35190 ( .A1(n3212), .A2(REG2_REG_8__SCAN_IN), .ZN(n3054) );
  INV_X1 U35200 ( .A(n5269), .ZN(n3051) );
  NAND2_X1 U35210 ( .A1(n4287), .A2(n3051), .ZN(n3053) );
  NAND2_X1 U35220 ( .A1(n3106), .A2(REG0_REG_8__SCAN_IN), .ZN(n3052) );
  NAND4_X1 U35230 ( .A1(n3055), .A2(n3054), .A3(n3053), .A4(n3052), .ZN(n4727)
         );
  NAND2_X1 U35240 ( .A1(n4727), .A2(n3090), .ZN(n3057) );
  NAND2_X1 U35250 ( .A1(n5250), .A2(n4103), .ZN(n3056) );
  NAND2_X1 U35260 ( .A1(n3057), .A2(n3056), .ZN(n3058) );
  XNOR2_X1 U35270 ( .A(n3058), .B(n3093), .ZN(n3183) );
  NAND2_X1 U35280 ( .A1(n4727), .A2(n4239), .ZN(n3060) );
  NAND2_X1 U35290 ( .A1(n5250), .A2(n3090), .ZN(n3059) );
  NAND2_X1 U35300 ( .A1(n3060), .A2(n3059), .ZN(n3181) );
  XNOR2_X1 U35310 ( .A(n3183), .B(n3181), .ZN(n3131) );
  NAND2_X1 U35320 ( .A1(n3062), .A2(n3061), .ZN(n3155) );
  NAND2_X1 U35330 ( .A1(n4731), .A2(n4235), .ZN(n3064) );
  NAND2_X1 U35340 ( .A1(n3373), .A2(n4103), .ZN(n3063) );
  NAND2_X1 U35350 ( .A1(n3064), .A2(n3063), .ZN(n3065) );
  XNOR2_X1 U35360 ( .A(n3065), .B(n3296), .ZN(n3102) );
  NAND2_X1 U35370 ( .A1(n4731), .A2(n4239), .ZN(n3067) );
  NAND2_X1 U35380 ( .A1(n3373), .A2(n3090), .ZN(n3066) );
  NAND2_X1 U35390 ( .A1(n3067), .A2(n3066), .ZN(n3101) );
  XNOR2_X1 U35400 ( .A(n3102), .B(n3101), .ZN(n3158) );
  INV_X1 U35410 ( .A(n3068), .ZN(n3069) );
  NAND2_X1 U35420 ( .A1(n3070), .A2(n3069), .ZN(n3154) );
  INV_X1 U35430 ( .A(n3154), .ZN(n3071) );
  NAND2_X1 U35440 ( .A1(n3155), .A2(n3072), .ZN(n3145) );
  NAND2_X1 U35450 ( .A1(n2479), .A2(REG1_REG_5__SCAN_IN), .ZN(n3077) );
  NAND2_X1 U35460 ( .A1(n3212), .A2(REG2_REG_5__SCAN_IN), .ZN(n3076) );
  OAI21_X1 U35470 ( .B1(n3073), .B2(REG3_REG_5__SCAN_IN), .A(n3084), .ZN(n3153) );
  INV_X1 U35480 ( .A(n3153), .ZN(n3362) );
  NAND2_X1 U35490 ( .A1(n4287), .A2(n3362), .ZN(n3075) );
  NAND2_X1 U35500 ( .A1(n3106), .A2(REG0_REG_5__SCAN_IN), .ZN(n3074) );
  NAND4_X1 U35510 ( .A1(n3077), .A2(n3076), .A3(n3075), .A4(n3074), .ZN(n4730)
         );
  NAND2_X1 U35520 ( .A1(n4730), .A2(n4235), .ZN(n3079) );
  NAND2_X1 U35530 ( .A1(n3339), .A2(n4103), .ZN(n3078) );
  NAND2_X1 U35540 ( .A1(n3079), .A2(n3078), .ZN(n3080) );
  XNOR2_X1 U35550 ( .A(n3080), .B(n3093), .ZN(n3119) );
  NAND2_X1 U35560 ( .A1(n4730), .A2(n4239), .ZN(n3082) );
  NAND2_X1 U35570 ( .A1(n3339), .A2(n3090), .ZN(n3081) );
  NAND2_X1 U35580 ( .A1(n3082), .A2(n3081), .ZN(n3117) );
  AND2_X1 U35590 ( .A1(n3084), .A2(n3083), .ZN(n3085) );
  NOR2_X1 U35600 ( .A1(n3103), .A2(n3085), .ZN(n4337) );
  NAND2_X1 U35610 ( .A1(n4287), .A2(n4337), .ZN(n3089) );
  NAND2_X1 U35620 ( .A1(n3212), .A2(REG2_REG_6__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U35630 ( .A1(n2479), .A2(REG1_REG_6__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U35640 ( .A1(n3106), .A2(REG0_REG_6__SCAN_IN), .ZN(n3086) );
  NAND2_X1 U35650 ( .A1(n4729), .A2(n3090), .ZN(n3092) );
  NAND2_X1 U35660 ( .A1(n4342), .A2(n4103), .ZN(n3091) );
  NAND2_X1 U35670 ( .A1(n3092), .A2(n3091), .ZN(n3094) );
  XNOR2_X1 U35680 ( .A(n3094), .B(n3093), .ZN(n3099) );
  NAND2_X1 U35690 ( .A1(n4729), .A2(n2986), .ZN(n3096) );
  NAND2_X1 U35700 ( .A1(n4342), .A2(n3090), .ZN(n3095) );
  NAND2_X1 U35710 ( .A1(n3096), .A2(n3095), .ZN(n3098) );
  INV_X1 U35720 ( .A(n3098), .ZN(n3097) );
  NAND2_X1 U35730 ( .A1(n3099), .A2(n3097), .ZN(n3120) );
  INV_X1 U35740 ( .A(n3120), .ZN(n3100) );
  XNOR2_X1 U35750 ( .A(n3099), .B(n3098), .ZN(n3169) );
  NAND2_X1 U35760 ( .A1(n3102), .A2(n3101), .ZN(n3146) );
  NAND2_X1 U35770 ( .A1(n2480), .A2(REG1_REG_7__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U35780 ( .A1(n3212), .A2(REG2_REG_7__SCAN_IN), .ZN(n3109) );
  OR2_X1 U35790 ( .A1(n3103), .A2(REG3_REG_7__SCAN_IN), .ZN(n3104) );
  AND2_X1 U35800 ( .A1(n3105), .A2(n3104), .ZN(n3285) );
  NAND2_X1 U35810 ( .A1(n4287), .A2(n3285), .ZN(n3108) );
  NAND2_X1 U3582 ( .A1(n3106), .A2(REG0_REG_7__SCAN_IN), .ZN(n3107) );
  NAND4_X1 U3583 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .ZN(n4728)
         );
  NAND2_X1 U3584 ( .A1(n4728), .A2(n3090), .ZN(n3112) );
  NAND2_X1 U3585 ( .A1(n3404), .A2(n4103), .ZN(n3111) );
  NAND2_X1 U3586 ( .A1(n3112), .A2(n3111), .ZN(n3113) );
  XNOR2_X1 U3587 ( .A(n3113), .B(n3296), .ZN(n3124) );
  NAND2_X1 U3588 ( .A1(n4728), .A2(n4239), .ZN(n3115) );
  NAND2_X1 U3589 ( .A1(n3404), .A2(n3090), .ZN(n3114) );
  NAND2_X1 U3590 ( .A1(n3115), .A2(n3114), .ZN(n3123) );
  NAND2_X1 U3591 ( .A1(n3124), .A2(n3123), .ZN(n3126) );
  NAND2_X1 U3592 ( .A1(n3145), .A2(n3116), .ZN(n3129) );
  INV_X1 U3593 ( .A(n3117), .ZN(n3118) );
  NAND2_X1 U3594 ( .A1(n3119), .A2(n3118), .ZN(n3166) );
  NAND2_X1 U3595 ( .A1(n3166), .A2(n3120), .ZN(n3121) );
  NAND2_X1 U3596 ( .A1(n3122), .A2(n3121), .ZN(n3279) );
  XNOR2_X1 U3597 ( .A(n3124), .B(n3123), .ZN(n3284) );
  INV_X1 U3598 ( .A(n3284), .ZN(n3125) );
  AND2_X1 U3599 ( .A1(n3279), .A2(n3125), .ZN(n3281) );
  INV_X1 U3600 ( .A(n3281), .ZN(n3127) );
  NAND2_X1 U3601 ( .A1(n3127), .A2(n3126), .ZN(n3128) );
  NAND2_X1 U3602 ( .A1(n3129), .A2(n3128), .ZN(n3130) );
  OAI21_X1 U3603 ( .B1(n3131), .B2(n3130), .A(n3185), .ZN(n3132) );
  NAND2_X1 U3604 ( .A1(n3132), .A2(n5366), .ZN(n3144) );
  NAND2_X1 U3605 ( .A1(n2480), .A2(REG1_REG_9__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U3606 ( .A1(n3212), .A2(REG2_REG_9__SCAN_IN), .ZN(n3137) );
  AND2_X1 U3607 ( .A1(n3133), .A2(n3239), .ZN(n3134) );
  NOR2_X1 U3608 ( .A1(n3186), .A2(n3134), .ZN(n3419) );
  NAND2_X1 U3609 ( .A1(n4287), .A2(n3419), .ZN(n3136) );
  NAND2_X1 U3610 ( .A1(n3106), .A2(REG0_REG_9__SCAN_IN), .ZN(n3135) );
  NAND2_X1 U3611 ( .A1(n4726), .A2(n5302), .ZN(n3140) );
  NAND2_X1 U3612 ( .A1(n4728), .A2(n5304), .ZN(n3139) );
  AND2_X1 U3613 ( .A1(n3140), .A2(n3139), .ZN(n5254) );
  INV_X1 U3614 ( .A(n5359), .ZN(n5310) );
  OAI22_X1 U3615 ( .A1(n5254), .A2(n5310), .B1(STATE_REG_SCAN_IN), .B2(n3141), 
        .ZN(n3142) );
  AOI21_X1 U3616 ( .B1(n5250), .B2(n5364), .A(n3142), .ZN(n3143) );
  OAI211_X1 U3617 ( .C1(n5370), .C2(n5269), .A(n3144), .B(n3143), .ZN(U3218)
         );
  AND2_X1 U3618 ( .A1(n3145), .A2(n3146), .ZN(n3278) );
  NAND2_X1 U3619 ( .A1(n3278), .A2(n3147), .ZN(n3167) );
  OAI21_X1 U3620 ( .B1(n3147), .B2(n3278), .A(n3167), .ZN(n3148) );
  NAND2_X1 U3621 ( .A1(n3148), .A2(n5366), .ZN(n3152) );
  AOI22_X1 U3622 ( .A1(n5302), .A2(n4729), .B1(n4731), .B2(n5304), .ZN(n3358)
         );
  OAI22_X1 U3623 ( .A1(n3358), .A2(n5310), .B1(STATE_REG_SCAN_IN), .B2(n3149), 
        .ZN(n3150) );
  AOI21_X1 U3624 ( .B1(n3339), .B2(n5364), .A(n3150), .ZN(n3151) );
  OAI211_X1 U3625 ( .C1(n5370), .C2(n3153), .A(n3152), .B(n3151), .ZN(U3224)
         );
  NAND2_X1 U3626 ( .A1(n3155), .A2(n3154), .ZN(n3157) );
  INV_X1 U3627 ( .A(n3145), .ZN(n3156) );
  AOI211_X1 U3628 ( .C1(n3158), .C2(n3157), .A(n5315), .B(n3156), .ZN(n3165)
         );
  INV_X1 U3629 ( .A(n3373), .ZN(n3324) );
  INV_X1 U3630 ( .A(n4730), .ZN(n3367) );
  OAI22_X1 U3631 ( .A1(n4542), .A2(n3324), .B1(n4555), .B2(n3367), .ZN(n3164)
         );
  INV_X1 U3632 ( .A(n3159), .ZN(n3374) );
  NAND2_X1 U3633 ( .A1(n4558), .A2(n4732), .ZN(n3162) );
  INV_X1 U3634 ( .A(n3160), .ZN(n3161) );
  OAI211_X1 U3635 ( .C1(n5370), .C2(n3374), .A(n3162), .B(n3161), .ZN(n3163)
         );
  OR3_X1 U3636 ( .A1(n3165), .A2(n3164), .A3(n3163), .ZN(U3227) );
  NAND2_X1 U3637 ( .A1(n3167), .A2(n3166), .ZN(n3168) );
  XOR2_X1 U3638 ( .A(n3169), .B(n3168), .Z(n3175) );
  INV_X1 U3639 ( .A(n5370), .ZN(n4522) );
  INV_X1 U3640 ( .A(n4342), .ZN(n3340) );
  NAND2_X1 U3641 ( .A1(n4728), .A2(n5302), .ZN(n3171) );
  NAND2_X1 U3642 ( .A1(n4730), .A2(n5304), .ZN(n3170) );
  NAND2_X1 U3643 ( .A1(n3171), .A2(n3170), .ZN(n4341) );
  AOI22_X1 U3644 ( .A1(n4341), .A2(n5359), .B1(REG3_REG_6__SCAN_IN), .B2(U3149), .ZN(n3172) );
  OAI21_X1 U3645 ( .B1(n4542), .B2(n3340), .A(n3172), .ZN(n3173) );
  AOI21_X1 U3646 ( .B1(n4337), .B2(n4522), .A(n3173), .ZN(n3174) );
  OAI21_X1 U3647 ( .B1(n3175), .B2(n5315), .A(n3174), .ZN(U3236) );
  NAND2_X1 U3648 ( .A1(n4726), .A2(n3090), .ZN(n3177) );
  NAND2_X1 U3649 ( .A1(n3448), .A2(n4103), .ZN(n3176) );
  NAND2_X1 U3650 ( .A1(n3177), .A2(n3176), .ZN(n3178) );
  XNOR2_X1 U3651 ( .A(n3178), .B(n3093), .ZN(n3201) );
  NAND2_X1 U3652 ( .A1(n3448), .A2(n3090), .ZN(n3180) );
  NAND2_X1 U3653 ( .A1(n4726), .A2(n4239), .ZN(n3179) );
  NAND2_X1 U3654 ( .A1(n3180), .A2(n3179), .ZN(n3199) );
  XNOR2_X1 U3655 ( .A(n3201), .B(n3199), .ZN(n3203) );
  INV_X1 U3656 ( .A(n3181), .ZN(n3182) );
  NAND2_X1 U3657 ( .A1(n3183), .A2(n3182), .ZN(n3184) );
  XOR2_X1 U3658 ( .A(n3203), .B(n3204), .Z(n3198) );
  NAND2_X1 U3659 ( .A1(n2479), .A2(REG1_REG_10__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U3660 ( .A1(n3212), .A2(REG2_REG_10__SCAN_IN), .ZN(n3191) );
  NOR2_X1 U3661 ( .A1(n3186), .A2(REG3_REG_10__SCAN_IN), .ZN(n3187) );
  OR2_X1 U3662 ( .A1(n3213), .A2(n3187), .ZN(n4401) );
  INV_X1 U3663 ( .A(n4401), .ZN(n3188) );
  NAND2_X1 U3664 ( .A1(n4287), .A2(n3188), .ZN(n3190) );
  NAND2_X1 U3665 ( .A1(n3106), .A2(REG0_REG_10__SCAN_IN), .ZN(n3189) );
  NAND4_X1 U3666 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n4725)
         );
  NAND2_X1 U3667 ( .A1(n4725), .A2(n5302), .ZN(n3194) );
  NAND2_X1 U3668 ( .A1(n4727), .A2(n5304), .ZN(n3193) );
  NAND2_X1 U3669 ( .A1(n3194), .A2(n3193), .ZN(n3398) );
  AOI22_X1 U3670 ( .A1(n3398), .A2(n5359), .B1(REG3_REG_9__SCAN_IN), .B2(U3149), .ZN(n3195) );
  OAI21_X1 U3671 ( .B1(n4542), .B2(n3400), .A(n3195), .ZN(n3196) );
  AOI21_X1 U3672 ( .B1(n3419), .B2(n4522), .A(n3196), .ZN(n3197) );
  OAI21_X1 U3673 ( .B1(n3198), .B2(n5315), .A(n3197), .ZN(U3228) );
  INV_X1 U3674 ( .A(n3199), .ZN(n3200) );
  AND2_X1 U3675 ( .A1(n3201), .A2(n3200), .ZN(n3202) );
  NAND2_X1 U3676 ( .A1(n4725), .A2(n3090), .ZN(n3206) );
  NAND2_X1 U3677 ( .A1(n4400), .A2(n4103), .ZN(n3205) );
  NAND2_X1 U3678 ( .A1(n3206), .A2(n3205), .ZN(n3207) );
  XNOR2_X1 U3679 ( .A(n3207), .B(n3093), .ZN(n3291) );
  NAND2_X1 U3680 ( .A1(n4725), .A2(n4239), .ZN(n3209) );
  NAND2_X1 U3681 ( .A1(n4400), .A2(n3090), .ZN(n3208) );
  NAND2_X1 U3682 ( .A1(n3209), .A2(n3208), .ZN(n3292) );
  XNOR2_X1 U3683 ( .A(n3291), .B(n3292), .ZN(n3210) );
  OAI211_X1 U3684 ( .C1(n3211), .C2(n3210), .A(n3584), .B(n5366), .ZN(n3225)
         );
  INV_X1 U3685 ( .A(n4400), .ZN(n4409) );
  NAND2_X1 U3686 ( .A1(n2480), .A2(REG1_REG_11__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U3687 ( .A1(n3212), .A2(REG2_REG_11__SCAN_IN), .ZN(n3217) );
  NOR2_X1 U3688 ( .A1(n3213), .A2(REG3_REG_11__SCAN_IN), .ZN(n3214) );
  OR2_X1 U3689 ( .A1(n3307), .A2(n3214), .ZN(n3453) );
  INV_X1 U3690 ( .A(n3453), .ZN(n3317) );
  NAND2_X1 U3691 ( .A1(n4287), .A2(n3317), .ZN(n3216) );
  NAND2_X1 U3692 ( .A1(n3106), .A2(REG0_REG_11__SCAN_IN), .ZN(n3215) );
  NAND4_X1 U3693 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n4724)
         );
  INV_X1 U3694 ( .A(n4724), .ZN(n4496) );
  OAI22_X1 U3695 ( .A1(n4542), .A2(n4409), .B1(n4555), .B2(n4496), .ZN(n3223)
         );
  NAND2_X1 U3696 ( .A1(n4558), .A2(n4726), .ZN(n3221) );
  INV_X1 U3697 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3219) );
  NOR2_X1 U3698 ( .A1(n3219), .A2(STATE_REG_SCAN_IN), .ZN(n3433) );
  INV_X1 U3699 ( .A(n3433), .ZN(n3220) );
  OAI211_X1 U3700 ( .C1(n5370), .C2(n4401), .A(n3221), .B(n3220), .ZN(n3222)
         );
  NOR2_X1 U3701 ( .A1(n3223), .A2(n3222), .ZN(n3224) );
  NAND2_X1 U3702 ( .A1(n3225), .A2(n3224), .ZN(U3214) );
  INV_X1 U3703 ( .A(n3226), .ZN(n3227) );
  INV_X1 U3704 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3421) );
  INV_X1 U3705 ( .A(n3426), .ZN(n5271) );
  AOI22_X1 U3706 ( .A1(n3426), .A2(n3421), .B1(REG2_REG_9__SCAN_IN), .B2(n5271), .ZN(n3230) );
  AOI211_X1 U3707 ( .C1(n3229), .C2(n3230), .A(n3427), .B(n4773), .ZN(n3244)
         );
  INV_X1 U3708 ( .A(n3231), .ZN(n3235) );
  INV_X1 U3709 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3232) );
  OR2_X1 U3710 ( .A1(n3426), .A2(REG1_REG_9__SCAN_IN), .ZN(n3236) );
  NAND2_X1 U3711 ( .A1(n3426), .A2(REG1_REG_9__SCAN_IN), .ZN(n3434) );
  AND2_X1 U3712 ( .A1(n3236), .A2(n3434), .ZN(n3237) );
  NAND2_X1 U3713 ( .A1(n3237), .A2(n3238), .ZN(n3435) );
  OAI211_X1 U3714 ( .C1(n3238), .C2(n3237), .A(n4770), .B(n3435), .ZN(n3242)
         );
  NOR2_X1 U3715 ( .A1(STATE_REG_SCAN_IN), .A2(n3239), .ZN(n3240) );
  AOI21_X1 U3716 ( .B1(n5143), .B2(ADDR_REG_9__SCAN_IN), .A(n3240), .ZN(n3241)
         );
  OAI211_X1 U3717 ( .C1(n4768), .C2(n5271), .A(n3242), .B(n3241), .ZN(n3243)
         );
  OR2_X1 U3718 ( .A1(n3244), .A2(n3243), .ZN(U3249) );
  INV_X1 U3719 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4150) );
  INV_X1 U3720 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4519) );
  INV_X1 U3721 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4541) );
  INV_X1 U3722 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4476) );
  INV_X1 U3723 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4253) );
  INV_X1 U3724 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4252) );
  INV_X1 U3725 ( .A(n4265), .ZN(n3250) );
  NAND2_X1 U3726 ( .A1(n3250), .A2(REG3_REG_27__SCAN_IN), .ZN(n4280) );
  INV_X1 U3727 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4279) );
  INV_X1 U3728 ( .A(n4282), .ZN(n4443) );
  INV_X1 U3729 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U3730 ( .A1(n3212), .A2(REG2_REG_29__SCAN_IN), .ZN(n3252) );
  NAND2_X1 U3731 ( .A1(n2479), .A2(REG1_REG_29__SCAN_IN), .ZN(n3251) );
  OAI211_X1 U3732 ( .C1(n4450), .C2(n4285), .A(n3252), .B(n3251), .ZN(n3253)
         );
  AOI21_X1 U3733 ( .B1(n4443), .B2(n4287), .A(n3253), .ZN(n4782) );
  NAND2_X1 U3734 ( .A1(n4734), .A2(DATAO_REG_29__SCAN_IN), .ZN(n3254) );
  OAI21_X1 U3735 ( .B1(n4782), .B2(n4734), .A(n3254), .ZN(U3579) );
  NAND3_X1 U3736 ( .A1(n4712), .A2(n3256), .A3(n3255), .ZN(n3257) );
  NAND2_X1 U3737 ( .A1(n5151), .A2(n3387), .ZN(n4661) );
  NAND2_X1 U3738 ( .A1(n4420), .A2(n2934), .ZN(n4658) );
  INV_X1 U3739 ( .A(n4735), .ZN(n3258) );
  NAND2_X1 U3740 ( .A1(n3258), .A2(n4604), .ZN(n4657) );
  INV_X1 U3741 ( .A(n4733), .ZN(n5187) );
  NAND2_X1 U3742 ( .A1(n5187), .A2(n3264), .ZN(n4662) );
  INV_X1 U3743 ( .A(n3264), .ZN(n3335) );
  NAND2_X1 U3744 ( .A1(n3335), .A2(n4733), .ZN(n4665) );
  INV_X1 U3745 ( .A(n3321), .ZN(n4608) );
  XNOR2_X1 U3746 ( .A(n3322), .B(n4608), .ZN(n3263) );
  OR2_X1 U3747 ( .A1(n2864), .A2(n4592), .ZN(n3260) );
  OR2_X1 U3748 ( .A1(n4767), .A2(n4361), .ZN(n3259) );
  NAND2_X1 U3749 ( .A1(n3260), .A2(n3259), .ZN(n5333) );
  INV_X1 U3750 ( .A(n5333), .ZN(n5190) );
  AOI21_X1 U3751 ( .B1(n3264), .B2(n5396), .A(n3261), .ZN(n3262) );
  OAI21_X1 U3752 ( .B1(n3263), .B2(n5190), .A(n3262), .ZN(n5176) );
  NAND2_X1 U3753 ( .A1(n5165), .A2(n3264), .ZN(n3265) );
  NAND2_X1 U3754 ( .A1(n5196), .A2(n3265), .ZN(n5174) );
  INV_X1 U3755 ( .A(n3266), .ZN(n3267) );
  AND2_X1 U3756 ( .A1(n5341), .A2(n3267), .ZN(n5415) );
  INV_X1 U3757 ( .A(n5415), .ZN(n5010) );
  INV_X1 U3758 ( .A(n5339), .ZN(n5204) );
  AOI22_X1 U3759 ( .A1(n5402), .A2(REG2_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(n5204), .ZN(n3268) );
  OAI21_X1 U3760 ( .B1(n5174), .B2(n5010), .A(n3268), .ZN(n3275) );
  AND2_X1 U3761 ( .A1(n4735), .A2(n4604), .ZN(n3386) );
  NAND2_X1 U3762 ( .A1(n3269), .A2(n3386), .ZN(n3385) );
  NAND2_X1 U3763 ( .A1(n2934), .A2(n3387), .ZN(n3270) );
  INV_X1 U3764 ( .A(n3337), .ZN(n3271) );
  AOI21_X1 U3765 ( .B1(n3321), .B2(n3272), .A(n3271), .ZN(n5175) );
  INV_X2 U3766 ( .A(n5402), .ZN(n5262) );
  NAND2_X1 U3767 ( .A1(n5154), .A2(n5103), .ZN(n5158) );
  NAND2_X1 U3768 ( .A1(n3273), .A2(n5158), .ZN(n5260) );
  NAND2_X1 U3769 ( .A1(n5262), .A2(n5260), .ZN(n4991) );
  NOR2_X1 U3770 ( .A1(n5175), .A2(n4991), .ZN(n3274) );
  AOI211_X1 U3771 ( .C1(n5341), .C2(n5176), .A(n3275), .B(n3274), .ZN(n3276)
         );
  INV_X1 U3772 ( .A(n3276), .ZN(U3288) );
  NAND2_X1 U3773 ( .A1(n3278), .A2(n3277), .ZN(n3280) );
  NAND2_X1 U3774 ( .A1(n3280), .A2(n3279), .ZN(n3283) );
  AND2_X1 U3775 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  AOI211_X1 U3776 ( .C1(n3284), .C2(n3283), .A(n5315), .B(n3282), .ZN(n3290)
         );
  INV_X1 U3777 ( .A(n3404), .ZN(n3331) );
  OAI22_X1 U3778 ( .A1(n4542), .A2(n3331), .B1(n4555), .B2(n3403), .ZN(n3289)
         );
  INV_X1 U3779 ( .A(n3285), .ZN(n3334) );
  NAND2_X1 U3780 ( .A1(n4558), .A2(n4729), .ZN(n3287) );
  OAI211_X1 U3781 ( .C1(n5370), .C2(n3334), .A(n3287), .B(n3286), .ZN(n3288)
         );
  OR3_X1 U3782 ( .A1(n3290), .A2(n3289), .A3(n3288), .ZN(U3210) );
  INV_X1 U3783 ( .A(n3291), .ZN(n3293) );
  NAND2_X1 U3784 ( .A1(n3293), .A2(n3292), .ZN(n3581) );
  NAND2_X1 U3785 ( .A1(n3584), .A2(n3581), .ZN(n3306) );
  NAND2_X1 U3786 ( .A1(n4724), .A2(n4235), .ZN(n3295) );
  NAND2_X1 U3787 ( .A1(n3469), .A2(n4103), .ZN(n3294) );
  NAND2_X1 U3788 ( .A1(n3295), .A2(n3294), .ZN(n3297) );
  XNOR2_X1 U3789 ( .A(n3297), .B(n3296), .ZN(n3303) );
  INV_X1 U3790 ( .A(n3303), .ZN(n3301) );
  NAND2_X1 U3791 ( .A1(n4724), .A2(n4239), .ZN(n3299) );
  NAND2_X1 U3792 ( .A1(n3469), .A2(n3090), .ZN(n3298) );
  NAND2_X1 U3793 ( .A1(n3299), .A2(n3298), .ZN(n3302) );
  INV_X1 U3794 ( .A(n3302), .ZN(n3300) );
  NAND2_X1 U3795 ( .A1(n3301), .A2(n3300), .ZN(n3585) );
  INV_X1 U3796 ( .A(n3585), .ZN(n3304) );
  AND2_X1 U3797 ( .A1(n3303), .A2(n3302), .ZN(n3580) );
  NOR2_X1 U3798 ( .A1(n3304), .A2(n3580), .ZN(n3305) );
  XNOR2_X1 U3799 ( .A(n3306), .B(n3305), .ZN(n3319) );
  NAND2_X1 U3800 ( .A1(n2479), .A2(REG1_REG_12__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U3801 ( .A1(n3212), .A2(REG2_REG_12__SCAN_IN), .ZN(n3311) );
  NOR2_X1 U3802 ( .A1(n3307), .A2(REG3_REG_12__SCAN_IN), .ZN(n3308) );
  NOR2_X1 U3803 ( .A1(n3459), .A2(n3308), .ZN(n4499) );
  NAND2_X1 U3804 ( .A1(n4287), .A2(n4499), .ZN(n3310) );
  NAND2_X1 U3805 ( .A1(n3106), .A2(REG0_REG_12__SCAN_IN), .ZN(n3309) );
  NAND4_X1 U3806 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n5305)
         );
  NAND2_X1 U3807 ( .A1(n5305), .A2(n5302), .ZN(n3314) );
  NAND2_X1 U3808 ( .A1(n4725), .A2(n5304), .ZN(n3313) );
  NAND2_X1 U3809 ( .A1(n3314), .A2(n3313), .ZN(n3445) );
  AOI22_X1 U3810 ( .A1(n3445), .A2(n5359), .B1(REG3_REG_11__SCAN_IN), .B2(
        U3149), .ZN(n3315) );
  OAI21_X1 U3811 ( .B1(n4542), .B2(n3470), .A(n3315), .ZN(n3316) );
  AOI21_X1 U3812 ( .B1(n3317), .B2(n4522), .A(n3316), .ZN(n3318) );
  OAI21_X1 U3813 ( .B1(n3319), .B2(n5315), .A(n3318), .ZN(U3233) );
  INV_X1 U3814 ( .A(n4728), .ZN(n3320) );
  NAND2_X1 U3815 ( .A1(n3320), .A2(n3404), .ZN(n4674) );
  NAND2_X1 U3816 ( .A1(n3331), .A2(n4728), .ZN(n4642) );
  NAND2_X1 U3817 ( .A1(n3368), .A2(n5197), .ZN(n4667) );
  NAND2_X1 U3818 ( .A1(n3338), .A2(n4732), .ZN(n4664) );
  AND2_X1 U3819 ( .A1(n4667), .A2(n4664), .ZN(n4606) );
  NAND2_X1 U3820 ( .A1(n5183), .A2(n4606), .ZN(n3323) );
  NAND2_X1 U3821 ( .A1(n3323), .A2(n4667), .ZN(n3366) );
  NAND2_X1 U3822 ( .A1(n3324), .A2(n4731), .ZN(n4670) );
  NAND2_X1 U3823 ( .A1(n3366), .A2(n4670), .ZN(n3325) );
  NAND2_X1 U3824 ( .A1(n5185), .A2(n3373), .ZN(n4668) );
  NAND2_X1 U3825 ( .A1(n3361), .A2(n4730), .ZN(n4671) );
  NAND2_X1 U3826 ( .A1(n3367), .A2(n3339), .ZN(n4644) );
  NAND2_X1 U3827 ( .A1(n4671), .A2(n4644), .ZN(n4611) );
  INV_X1 U3828 ( .A(n4672), .ZN(n3326) );
  INV_X1 U3829 ( .A(n4729), .ZN(n3341) );
  NAND2_X1 U3830 ( .A1(n3341), .A2(n4342), .ZN(n3342) );
  NAND2_X1 U3831 ( .A1(n3327), .A2(n4628), .ZN(n3394) );
  OAI21_X1 U3832 ( .B1(n4628), .B2(n3327), .A(n3394), .ZN(n3328) );
  NAND2_X1 U3833 ( .A1(n3328), .A2(n5333), .ZN(n3330) );
  AOI22_X1 U3834 ( .A1(n5304), .A2(n4729), .B1(n4727), .B2(n5302), .ZN(n3329)
         );
  OAI211_X1 U3835 ( .C1(n5330), .C2(n3331), .A(n3330), .B(n3329), .ZN(n5236)
         );
  INV_X1 U3836 ( .A(n5236), .ZN(n3356) );
  NAND2_X1 U3837 ( .A1(n5262), .A2(n4767), .ZN(n4877) );
  NAND2_X1 U3838 ( .A1(n4334), .A2(n3404), .ZN(n3332) );
  NAND2_X1 U3839 ( .A1(n3332), .A2(n5406), .ZN(n3333) );
  NOR2_X1 U3840 ( .A1(n5247), .A2(n3333), .ZN(n5237) );
  OAI22_X1 U3841 ( .A1(n5341), .A2(n3029), .B1(n3334), .B2(n5339), .ZN(n3354)
         );
  NAND2_X1 U3842 ( .A1(n5187), .A2(n3335), .ZN(n3336) );
  NAND2_X1 U3843 ( .A1(n4668), .A2(n4670), .ZN(n4607) );
  NAND2_X1 U3844 ( .A1(n3372), .A2(n4607), .ZN(n3410) );
  NAND2_X1 U3845 ( .A1(n4731), .A2(n3373), .ZN(n3407) );
  NAND2_X1 U3846 ( .A1(n3410), .A2(n3407), .ZN(n4330) );
  AND2_X1 U3847 ( .A1(n4730), .A2(n3339), .ZN(n4329) );
  NAND2_X1 U3848 ( .A1(n3341), .A2(n3340), .ZN(n3345) );
  INV_X1 U3849 ( .A(n3345), .ZN(n3343) );
  INV_X1 U3850 ( .A(n3347), .ZN(n3344) );
  OR2_X1 U3851 ( .A1(n4329), .A2(n3344), .ZN(n3406) );
  OR2_X1 U3852 ( .A1(n4330), .A2(n3406), .ZN(n3350) );
  INV_X1 U3853 ( .A(n4628), .ZN(n3348) );
  NAND2_X1 U3854 ( .A1(n3367), .A2(n3361), .ZN(n4331) );
  NAND2_X1 U3855 ( .A1(n4331), .A2(n3345), .ZN(n3346) );
  NAND2_X1 U3856 ( .A1(n3347), .A2(n3346), .ZN(n3349) );
  NAND2_X1 U3857 ( .A1(n3350), .A2(n3413), .ZN(n5244) );
  INV_X1 U3858 ( .A(n5244), .ZN(n3352) );
  NAND2_X1 U3859 ( .A1(n3350), .A2(n3349), .ZN(n3351) );
  AND2_X1 U3860 ( .A1(n3351), .A2(n4628), .ZN(n5235) );
  NOR3_X1 U3861 ( .A1(n3352), .A2(n5235), .A3(n4991), .ZN(n3353) );
  AOI211_X1 U3862 ( .C1(n4976), .C2(n5237), .A(n3354), .B(n3353), .ZN(n3355)
         );
  OAI21_X1 U3863 ( .B1(n5419), .B2(n3356), .A(n3355), .ZN(U3283) );
  XOR2_X1 U3864 ( .A(n4611), .B(n3357), .Z(n3360) );
  OAI21_X1 U3865 ( .B1(n3361), .B2(n5330), .A(n3358), .ZN(n3359) );
  AOI21_X1 U3866 ( .B1(n3360), .B2(n5333), .A(n3359), .ZN(n5219) );
  XOR2_X1 U3867 ( .A(n4611), .B(n4330), .Z(n5222) );
  OAI21_X1 U3868 ( .B1(n2482), .B2(n3361), .A(n4336), .ZN(n5220) );
  AOI22_X1 U3869 ( .A1(n5419), .A2(REG2_REG_5__SCAN_IN), .B1(n3362), .B2(n5204), .ZN(n3363) );
  OAI21_X1 U3870 ( .B1(n5220), .B2(n5010), .A(n3363), .ZN(n3364) );
  AOI21_X1 U3871 ( .B1(n5222), .B2(n5345), .A(n3364), .ZN(n3365) );
  OAI21_X1 U3872 ( .B1(n5419), .B2(n5219), .A(n3365), .ZN(U3285) );
  XNOR2_X1 U3873 ( .A(n3366), .B(n4607), .ZN(n3371) );
  OAI22_X1 U3874 ( .A1(n3368), .A2(n5186), .B1(n3367), .B2(n5184), .ZN(n3369)
         );
  AOI21_X1 U3875 ( .B1(n3373), .B2(n5396), .A(n3369), .ZN(n3370) );
  OAI21_X1 U3876 ( .B1(n3371), .B2(n5190), .A(n3370), .ZN(n5211) );
  INV_X1 U3877 ( .A(n5211), .ZN(n3379) );
  XOR2_X1 U3878 ( .A(n3372), .B(n4607), .Z(n5213) );
  NAND2_X1 U3879 ( .A1(n5213), .A2(n5345), .ZN(n3378) );
  AOI211_X1 U3880 ( .C1(n3373), .C2(n5194), .A(n5390), .B(n2482), .ZN(n5212)
         );
  OAI22_X1 U3881 ( .A1(n5341), .A2(n3375), .B1(n3374), .B2(n5339), .ZN(n3376)
         );
  AOI21_X1 U3882 ( .B1(n5212), .B2(n4976), .A(n3376), .ZN(n3377) );
  OAI211_X1 U3883 ( .C1(n5419), .C2(n3379), .A(n3378), .B(n3377), .ZN(U3286)
         );
  XNOR2_X1 U3884 ( .A(n3269), .B(n4657), .ZN(n3384) );
  NAND2_X1 U3885 ( .A1(n4735), .A2(n5304), .ZN(n3381) );
  NAND2_X1 U3886 ( .A1(n4733), .A2(n5302), .ZN(n3380) );
  NAND2_X1 U3887 ( .A1(n3381), .A2(n3380), .ZN(n4417) );
  INV_X1 U3888 ( .A(n4417), .ZN(n3382) );
  OAI21_X1 U3889 ( .B1(n4420), .B2(n5330), .A(n3382), .ZN(n3383) );
  AOI21_X1 U3890 ( .B1(n3384), .B2(n5333), .A(n3383), .ZN(n5167) );
  OAI21_X1 U3891 ( .B1(n3269), .B2(n3386), .A(n3385), .ZN(n5168) );
  INV_X1 U3892 ( .A(n5168), .ZN(n3392) );
  NAND2_X1 U3893 ( .A1(n3387), .A2(n4604), .ZN(n5164) );
  AND3_X1 U3894 ( .A1(n5415), .A2(n5165), .A3(n5164), .ZN(n3391) );
  OAI22_X1 U3895 ( .A1(n5341), .A2(n3389), .B1(n3388), .B2(n5339), .ZN(n3390)
         );
  AOI211_X1 U3896 ( .C1(n3392), .C2(n5345), .A(n3391), .B(n3390), .ZN(n3393)
         );
  OAI21_X1 U3897 ( .B1(n5419), .B2(n5167), .A(n3393), .ZN(U3289) );
  NAND2_X1 U3898 ( .A1(n3394), .A2(n4674), .ZN(n5252) );
  NAND2_X1 U3899 ( .A1(n3403), .A2(n5250), .ZN(n4676) );
  INV_X1 U3900 ( .A(n4676), .ZN(n3395) );
  NAND2_X1 U3901 ( .A1(n5256), .A2(n4727), .ZN(n3441) );
  NAND2_X1 U3902 ( .A1(n3442), .A2(n3441), .ZN(n3397) );
  INV_X1 U3903 ( .A(n4726), .ZN(n3396) );
  NAND2_X1 U3904 ( .A1(n3396), .A2(n3448), .ZN(n4677) );
  NAND2_X1 U3905 ( .A1(n3400), .A2(n4726), .ZN(n4679) );
  NAND2_X1 U3906 ( .A1(n4677), .A2(n4679), .ZN(n3449) );
  XNOR2_X1 U3907 ( .A(n3397), .B(n3449), .ZN(n3402) );
  INV_X1 U3908 ( .A(n3398), .ZN(n3399) );
  OAI21_X1 U3909 ( .B1(n3400), .B2(n5330), .A(n3399), .ZN(n3401) );
  AOI21_X1 U3910 ( .B1(n3402), .B2(n5333), .A(n3401), .ZN(n5275) );
  NAND2_X1 U3911 ( .A1(n3403), .A2(n5256), .ZN(n3412) );
  INV_X1 U3912 ( .A(n3412), .ZN(n3405) );
  NAND2_X1 U3913 ( .A1(n4728), .A2(n3404), .ZN(n5242) );
  NAND2_X1 U3914 ( .A1(n4676), .A2(n3441), .ZN(n4627) );
  OR2_X1 U3915 ( .A1(n3406), .A2(n3415), .ZN(n3409) );
  INV_X1 U3916 ( .A(n3407), .ZN(n3408) );
  NOR2_X1 U3917 ( .A1(n3409), .A2(n3408), .ZN(n3411) );
  NAND2_X1 U3918 ( .A1(n3411), .A2(n3410), .ZN(n3417) );
  NAND2_X1 U3919 ( .A1(n3417), .A2(n3416), .ZN(n3450) );
  XNOR2_X1 U3920 ( .A(n3450), .B(n2597), .ZN(n5276) );
  INV_X1 U3921 ( .A(n5276), .ZN(n3424) );
  INV_X1 U3922 ( .A(n5248), .ZN(n3418) );
  NAND2_X1 U3923 ( .A1(n3418), .A2(n3448), .ZN(n5273) );
  AND3_X1 U3924 ( .A1(n5273), .A2(n5415), .A3(n5272), .ZN(n3423) );
  INV_X1 U3925 ( .A(n3419), .ZN(n3420) );
  OAI22_X1 U3926 ( .A1(n5341), .A2(n3421), .B1(n3420), .B2(n5339), .ZN(n3422)
         );
  AOI211_X1 U3927 ( .C1(n3424), .C2(n5345), .A(n3423), .B(n3422), .ZN(n3425)
         );
  OAI21_X1 U3928 ( .B1(n5419), .B2(n5275), .A(n3425), .ZN(U3281) );
  INV_X1 U3929 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3432) );
  XNOR2_X1 U3930 ( .A(n3486), .B(n3428), .ZN(n3431) );
  INV_X1 U3931 ( .A(n3431), .ZN(n3429) );
  INV_X1 U3932 ( .A(n3487), .ZN(n3430) );
  AOI211_X1 U3933 ( .C1(n3432), .C2(n3431), .A(n3430), .B(n4773), .ZN(n3440)
         );
  AOI21_X1 U3934 ( .B1(n5143), .B2(ADDR_REG_10__SCAN_IN), .A(n3433), .ZN(n3438) );
  NAND2_X1 U3935 ( .A1(REG1_REG_10__SCAN_IN), .A2(n3436), .ZN(n3481) );
  OAI211_X1 U3936 ( .C1(REG1_REG_10__SCAN_IN), .C2(n3436), .A(n4770), .B(n3481), .ZN(n3437) );
  OAI211_X1 U3937 ( .C1(n4768), .C2(n3428), .A(n3438), .B(n3437), .ZN(n3439)
         );
  OR2_X1 U3938 ( .A1(n3440), .A2(n3439), .ZN(U3250) );
  AND2_X1 U3939 ( .A1(n4679), .A2(n3441), .ZN(n4643) );
  INV_X1 U3940 ( .A(n4725), .ZN(n3443) );
  NAND2_X1 U3941 ( .A1(n3443), .A2(n4400), .ZN(n4648) );
  INV_X1 U3942 ( .A(n4648), .ZN(n3444) );
  NAND2_X1 U3943 ( .A1(n4409), .A2(n4725), .ZN(n4646) );
  NAND2_X1 U3944 ( .A1(n4496), .A2(n3469), .ZN(n3514) );
  NAND2_X1 U3945 ( .A1(n3470), .A2(n4724), .ZN(n4647) );
  NAND2_X1 U3946 ( .A1(n3514), .A2(n4647), .ZN(n4617) );
  XNOR2_X1 U3947 ( .A(n2489), .B(n4617), .ZN(n3447) );
  AOI21_X1 U3948 ( .B1(n3469), .B2(n5396), .A(n3445), .ZN(n3446) );
  OAI21_X1 U3949 ( .B1(n3447), .B2(n5190), .A(n3446), .ZN(n5290) );
  INV_X1 U3950 ( .A(n5290), .ZN(n3457) );
  NAND2_X1 U3951 ( .A1(n4648), .A2(n4646), .ZN(n4404) );
  OAI21_X1 U3952 ( .B1(n3451), .B2(n4617), .A(n3472), .ZN(n5292) );
  OAI21_X1 U3953 ( .B1(n5272), .B2(n4400), .A(n3469), .ZN(n3452) );
  NAND2_X1 U3954 ( .A1(n3452), .A2(n3473), .ZN(n5289) );
  NOR2_X1 U3955 ( .A1(n5289), .A2(n5010), .ZN(n3455) );
  INV_X1 U3956 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3488) );
  OAI22_X1 U3957 ( .A1(n5262), .A2(n3488), .B1(n3453), .B2(n5339), .ZN(n3454)
         );
  AOI211_X1 U3958 ( .C1(n5292), .C2(n5345), .A(n3455), .B(n3454), .ZN(n3456)
         );
  OAI21_X1 U3959 ( .B1(n5419), .B2(n3457), .A(n3456), .ZN(U3279) );
  NAND2_X1 U3960 ( .A1(n3515), .A2(n3514), .ZN(n3458) );
  INV_X1 U3961 ( .A(n5305), .ZN(n3502) );
  NAND2_X1 U3962 ( .A1(n3502), .A2(n4495), .ZN(n3513) );
  INV_X1 U3963 ( .A(n4495), .ZN(n3501) );
  NAND2_X1 U3964 ( .A1(n3501), .A2(n5305), .ZN(n5325) );
  NAND2_X1 U3965 ( .A1(n3513), .A2(n5325), .ZN(n4620) );
  XNOR2_X1 U3966 ( .A(n3458), .B(n4620), .ZN(n3468) );
  NAND2_X1 U3967 ( .A1(n2480), .A2(REG1_REG_13__SCAN_IN), .ZN(n3465) );
  NAND2_X1 U3968 ( .A1(n3212), .A2(REG2_REG_13__SCAN_IN), .ZN(n3464) );
  OR2_X1 U3969 ( .A1(n3459), .A2(REG3_REG_13__SCAN_IN), .ZN(n3460) );
  NAND2_X1 U3970 ( .A1(n3460), .A2(n3505), .ZN(n5340) );
  INV_X1 U3971 ( .A(n5340), .ZN(n3461) );
  NAND2_X1 U3972 ( .A1(n4287), .A2(n3461), .ZN(n3463) );
  NAND2_X1 U3973 ( .A1(n3106), .A2(REG0_REG_13__SCAN_IN), .ZN(n3462) );
  OAI22_X1 U3974 ( .A1(n4496), .A2(n5186), .B1(n4465), .B2(n5184), .ZN(n3466)
         );
  AOI21_X1 U3975 ( .B1(n4495), .B2(n5396), .A(n3466), .ZN(n3467) );
  OAI21_X1 U3976 ( .B1(n3468), .B2(n5190), .A(n3467), .ZN(n5296) );
  AOI21_X1 U3977 ( .B1(n4499), .B2(n5204), .A(n5296), .ZN(n3478) );
  NAND2_X1 U3978 ( .A1(n4496), .A2(n3470), .ZN(n3471) );
  NAND2_X1 U3979 ( .A1(n3472), .A2(n3471), .ZN(n3503) );
  XNOR2_X1 U3980 ( .A(n3503), .B(n4620), .ZN(n5298) );
  NAND2_X1 U3981 ( .A1(n5298), .A2(n5345), .ZN(n3477) );
  NAND2_X1 U3982 ( .A1(n3473), .A2(n4495), .ZN(n3474) );
  NAND2_X1 U3983 ( .A1(n3474), .A2(n5406), .ZN(n3475) );
  NOR2_X1 U3984 ( .A1(n5324), .A2(n3475), .ZN(n5297) );
  INV_X1 U3985 ( .A(n5341), .ZN(n5402) );
  AOI22_X1 U3986 ( .A1(n5297), .A2(n4976), .B1(REG2_REG_12__SCAN_IN), .B2(
        n5402), .ZN(n3476) );
  OAI211_X1 U3987 ( .C1(n5419), .C2(n3478), .A(n3477), .B(n3476), .ZN(U3278)
         );
  INV_X1 U3988 ( .A(n5108), .ZN(n3500) );
  NAND2_X1 U3989 ( .A1(n3480), .A2(n3479), .ZN(n3482) );
  NAND2_X1 U3990 ( .A1(n3482), .A2(n3481), .ZN(n3485) );
  NAND2_X1 U3991 ( .A1(n3500), .A2(REG1_REG_11__SCAN_IN), .ZN(n3483) );
  OAI21_X1 U3992 ( .B1(n3500), .B2(REG1_REG_11__SCAN_IN), .A(n3483), .ZN(n3484) );
  NAND2_X1 U3993 ( .A1(n5108), .A2(REG1_REG_11__SCAN_IN), .ZN(n3533) );
  OAI211_X1 U3994 ( .C1(n5108), .C2(REG1_REG_11__SCAN_IN), .A(n3485), .B(n3533), .ZN(n3534) );
  OAI211_X1 U3995 ( .C1(n3485), .C2(n3484), .A(n3534), .B(n4770), .ZN(n3499)
         );
  INV_X1 U3996 ( .A(n3492), .ZN(n3495) );
  NAND2_X1 U3997 ( .A1(n3500), .A2(REG2_REG_11__SCAN_IN), .ZN(n3490) );
  NAND2_X1 U3998 ( .A1(n5108), .A2(n3488), .ZN(n3489) );
  AND2_X1 U3999 ( .A1(n3490), .A2(n3489), .ZN(n3494) );
  INV_X1 U4000 ( .A(n3539), .ZN(n3493) );
  AOI211_X1 U4001 ( .C1(n3495), .C2(n3494), .A(n3493), .B(n4773), .ZN(n3497)
         );
  AND2_X1 U4002 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3496) );
  AOI211_X1 U4003 ( .C1(n5143), .C2(ADDR_REG_11__SCAN_IN), .A(n3497), .B(n3496), .ZN(n3498) );
  OAI211_X1 U4004 ( .C1(n4768), .C2(n3500), .A(n3499), .B(n3498), .ZN(U3251)
         );
  NAND2_X1 U4005 ( .A1(n4465), .A2(n5331), .ZN(n3504) );
  NAND2_X1 U4006 ( .A1(n2480), .A2(REG1_REG_14__SCAN_IN), .ZN(n3509) );
  NAND2_X1 U4007 ( .A1(n3212), .A2(REG2_REG_14__SCAN_IN), .ZN(n3508) );
  AOI21_X1 U4008 ( .B1(n3505), .B2(n4150), .A(n3518), .ZN(n4468) );
  NAND2_X1 U4009 ( .A1(n4287), .A2(n4468), .ZN(n3507) );
  NAND2_X1 U4010 ( .A1(n3106), .A2(REG0_REG_14__SCAN_IN), .ZN(n3506) );
  NAND4_X1 U4011 ( .A1(n3509), .A2(n3508), .A3(n3507), .A4(n3506), .ZN(n5303)
         );
  INV_X1 U4012 ( .A(n5303), .ZN(n3510) );
  NAND2_X1 U4013 ( .A1(n3510), .A2(n4464), .ZN(n4566) );
  INV_X1 U4014 ( .A(n4464), .ZN(n3526) );
  NAND2_X1 U4015 ( .A1(n3526), .A2(n5303), .ZN(n4569) );
  NAND2_X1 U4016 ( .A1(n4566), .A2(n4569), .ZN(n4609) );
  OAI21_X1 U4017 ( .B1(n3511), .B2(n4609), .A(n3559), .ZN(n3512) );
  INV_X1 U4018 ( .A(n3512), .ZN(n5351) );
  AND2_X1 U4019 ( .A1(n3514), .A2(n3513), .ZN(n4653) );
  NAND2_X1 U4020 ( .A1(n5331), .A2(n4723), .ZN(n3516) );
  AND2_X1 U4021 ( .A1(n5325), .A2(n3516), .ZN(n4650) );
  NAND2_X1 U4022 ( .A1(n4465), .A2(n5320), .ZN(n4651) );
  OAI21_X1 U4023 ( .B1(n2578), .B2(n4564), .A(n4035), .ZN(n3517) );
  NAND2_X1 U4024 ( .A1(n3517), .A2(n5333), .ZN(n3525) );
  NAND2_X1 U4025 ( .A1(n3212), .A2(REG2_REG_15__SCAN_IN), .ZN(n3523) );
  NAND2_X1 U4026 ( .A1(n2479), .A2(REG1_REG_15__SCAN_IN), .ZN(n3522) );
  OAI21_X1 U4027 ( .B1(n3518), .B2(REG3_REG_15__SCAN_IN), .A(n3549), .ZN(n5371) );
  INV_X1 U4028 ( .A(n5371), .ZN(n3519) );
  NAND2_X1 U4029 ( .A1(n4287), .A2(n3519), .ZN(n3521) );
  NAND2_X1 U4030 ( .A1(n3106), .A2(REG0_REG_15__SCAN_IN), .ZN(n3520) );
  NAND4_X1 U4031 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n4722)
         );
  AOI22_X1 U4032 ( .A1(n5304), .A2(n4723), .B1(n4722), .B2(n5302), .ZN(n3524)
         );
  OAI211_X1 U4033 ( .C1(n5330), .C2(n3526), .A(n3525), .B(n3524), .ZN(n5353)
         );
  INV_X1 U4034 ( .A(n5323), .ZN(n3527) );
  OAI21_X1 U4035 ( .B1(n3527), .B2(n3526), .A(n3560), .ZN(n5350) );
  NOR2_X1 U4036 ( .A1(n5350), .A2(n5010), .ZN(n3531) );
  INV_X1 U4037 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3529) );
  INV_X1 U4038 ( .A(n4468), .ZN(n3528) );
  OAI22_X1 U4039 ( .A1(n5262), .A2(n3529), .B1(n3528), .B2(n5339), .ZN(n3530)
         );
  AOI211_X1 U4040 ( .C1(n5353), .C2(n5262), .A(n3531), .B(n3530), .ZN(n3532)
         );
  OAI21_X1 U4041 ( .B1(n5351), .B2(n4991), .A(n3532), .ZN(U3276) );
  XOR2_X1 U4042 ( .A(n4127), .B(REG1_REG_12__SCAN_IN), .Z(n3546) );
  INV_X1 U40430 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3536) );
  NOR2_X1 U4044 ( .A1(STATE_REG_SCAN_IN), .A2(n3536), .ZN(n4498) );
  AOI21_X1 U4045 ( .B1(n5143), .B2(ADDR_REG_12__SCAN_IN), .A(n4498), .ZN(n3537) );
  OAI21_X1 U4046 ( .B1(n3535), .B2(n4768), .A(n3537), .ZN(n3545) );
  INV_X1 U4047 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3543) );
  NAND2_X1 U4048 ( .A1(n5108), .A2(REG2_REG_11__SCAN_IN), .ZN(n3538) );
  NAND2_X1 U4049 ( .A1(n3540), .A2(n5107), .ZN(n4139) );
  NAND2_X1 U4050 ( .A1(n4139), .A2(n3541), .ZN(n3542) );
  AOI211_X1 U4051 ( .C1(n4770), .C2(n3546), .A(n3545), .B(n3544), .ZN(n3547)
         );
  INV_X1 U4052 ( .A(n3547), .ZN(U3252) );
  XNOR2_X1 U4053 ( .A(n5365), .B(n4722), .ZN(n4633) );
  NAND2_X1 U4054 ( .A1(n4035), .A2(n4566), .ZN(n3548) );
  XOR2_X1 U4055 ( .A(n4633), .B(n3548), .Z(n3557) );
  NAND2_X1 U4056 ( .A1(n3212), .A2(REG2_REG_16__SCAN_IN), .ZN(n3553) );
  AOI21_X1 U4057 ( .B1(n3549), .B2(n4519), .A(n3568), .ZN(n4521) );
  NAND2_X1 U4058 ( .A1(n4287), .A2(n4521), .ZN(n3552) );
  NAND2_X1 U4059 ( .A1(n2480), .A2(REG1_REG_16__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U4060 ( .A1(n3106), .A2(REG0_REG_16__SCAN_IN), .ZN(n3550) );
  NAND4_X1 U4061 ( .A1(n3553), .A2(n3552), .A3(n3551), .A4(n3550), .ZN(n4998)
         );
  NAND2_X1 U4062 ( .A1(n4998), .A2(n5302), .ZN(n3555) );
  NAND2_X1 U4063 ( .A1(n5303), .A2(n5304), .ZN(n3554) );
  NAND2_X1 U4064 ( .A1(n3555), .A2(n3554), .ZN(n5358) );
  AOI21_X1 U4065 ( .B1(n5365), .B2(n5396), .A(n5358), .ZN(n3556) );
  OAI21_X1 U4066 ( .B1(n3557), .B2(n5190), .A(n3556), .ZN(n5372) );
  INV_X1 U4067 ( .A(n5372), .ZN(n3567) );
  XOR2_X1 U4068 ( .A(n4633), .B(n4033), .Z(n5374) );
  NAND2_X1 U4069 ( .A1(n5374), .A2(n5345), .ZN(n3566) );
  NAND2_X1 U4070 ( .A1(n3560), .A2(n5365), .ZN(n3561) );
  NAND2_X1 U4071 ( .A1(n3561), .A2(n5406), .ZN(n3562) );
  NOR2_X1 U4072 ( .A1(n4042), .A2(n3562), .ZN(n5373) );
  INV_X1 U4073 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3563) );
  OAI22_X1 U4074 ( .A1(n5262), .A2(n3563), .B1(n5371), .B2(n5339), .ZN(n3564)
         );
  AOI21_X1 U4075 ( .B1(n5373), .B2(n4976), .A(n3564), .ZN(n3565) );
  OAI211_X1 U4076 ( .C1(n5419), .C2(n3567), .A(n3566), .B(n3565), .ZN(U3275)
         );
  NAND2_X1 U4077 ( .A1(n2479), .A2(REG1_REG_17__SCAN_IN), .ZN(n3574) );
  NAND2_X1 U4078 ( .A1(n3212), .A2(REG2_REG_17__SCAN_IN), .ZN(n3573) );
  OR2_X1 U4079 ( .A1(n3568), .A2(REG3_REG_17__SCAN_IN), .ZN(n3569) );
  NAND2_X1 U4080 ( .A1(n3639), .A2(n3569), .ZN(n5004) );
  INV_X1 U4081 ( .A(n5004), .ZN(n3570) );
  NAND2_X1 U4082 ( .A1(n4287), .A2(n3570), .ZN(n3572) );
  NAND2_X1 U4083 ( .A1(n3106), .A2(REG0_REG_17__SCAN_IN), .ZN(n3571) );
  NAND4_X1 U4084 ( .A1(n3574), .A2(n3573), .A3(n3572), .A4(n3571), .ZN(n4721)
         );
  NAND2_X1 U4085 ( .A1(n4721), .A2(n4235), .ZN(n3576) );
  NAND2_X1 U4086 ( .A1(n4369), .A2(n4103), .ZN(n3575) );
  NAND2_X1 U4087 ( .A1(n3576), .A2(n3575), .ZN(n3577) );
  XNOR2_X1 U4088 ( .A(n3577), .B(n3093), .ZN(n4050) );
  NAND2_X1 U4089 ( .A1(n4721), .A2(n4239), .ZN(n3579) );
  NAND2_X1 U4090 ( .A1(n4369), .A2(n4235), .ZN(n3578) );
  NAND2_X1 U4091 ( .A1(n3579), .A2(n3578), .ZN(n4048) );
  XNOR2_X1 U4092 ( .A(n4050), .B(n4048), .ZN(n3638) );
  INV_X1 U4093 ( .A(n3580), .ZN(n3582) );
  AND2_X1 U4094 ( .A1(n3582), .A2(n3581), .ZN(n3583) );
  NAND2_X1 U4095 ( .A1(n3584), .A2(n3583), .ZN(n3586) );
  NAND2_X1 U4096 ( .A1(n3586), .A2(n3585), .ZN(n4492) );
  NAND2_X1 U4097 ( .A1(n5305), .A2(n3090), .ZN(n3588) );
  NAND2_X1 U4098 ( .A1(n4495), .A2(n4103), .ZN(n3587) );
  NAND2_X1 U4099 ( .A1(n3588), .A2(n3587), .ZN(n3589) );
  XNOR2_X1 U4100 ( .A(n3589), .B(n3093), .ZN(n3592) );
  NAND2_X1 U4101 ( .A1(n5305), .A2(n4239), .ZN(n3591) );
  NAND2_X1 U4102 ( .A1(n4495), .A2(n3090), .ZN(n3590) );
  AND2_X1 U4103 ( .A1(n3591), .A2(n3590), .ZN(n3593) );
  NAND2_X1 U4104 ( .A1(n3592), .A2(n3593), .ZN(n5313) );
  INV_X1 U4105 ( .A(n3592), .ZN(n3595) );
  INV_X1 U4106 ( .A(n3593), .ZN(n3594) );
  NAND2_X1 U4107 ( .A1(n3595), .A2(n3594), .ZN(n3596) );
  AND2_X1 U4108 ( .A1(n5313), .A2(n3596), .ZN(n4493) );
  NAND2_X1 U4109 ( .A1(n4492), .A2(n4493), .ZN(n5314) );
  NAND2_X1 U4110 ( .A1(n4723), .A2(n3090), .ZN(n3598) );
  NAND2_X1 U4111 ( .A1(n5320), .A2(n4103), .ZN(n3597) );
  NAND2_X1 U4112 ( .A1(n3598), .A2(n3597), .ZN(n3599) );
  XNOR2_X1 U4113 ( .A(n3599), .B(n3093), .ZN(n3602) );
  NAND2_X1 U4114 ( .A1(n4723), .A2(n4239), .ZN(n3601) );
  NAND2_X1 U4115 ( .A1(n5320), .A2(n3090), .ZN(n3600) );
  AND2_X1 U4116 ( .A1(n3601), .A2(n3600), .ZN(n3603) );
  NAND2_X1 U4117 ( .A1(n3602), .A2(n3603), .ZN(n3607) );
  INV_X1 U4118 ( .A(n3602), .ZN(n3605) );
  INV_X1 U4119 ( .A(n3603), .ZN(n3604) );
  NAND2_X1 U4120 ( .A1(n3605), .A2(n3604), .ZN(n3606) );
  AND2_X1 U4121 ( .A1(n3607), .A2(n3606), .ZN(n5311) );
  NAND2_X1 U4122 ( .A1(n5303), .A2(n4235), .ZN(n3609) );
  NAND2_X1 U4123 ( .A1(n4464), .A2(n4103), .ZN(n3608) );
  NAND2_X1 U4124 ( .A1(n3609), .A2(n3608), .ZN(n3610) );
  XNOR2_X1 U4125 ( .A(n3610), .B(n3093), .ZN(n3615) );
  NAND2_X1 U4126 ( .A1(n5303), .A2(n2986), .ZN(n3612) );
  NAND2_X1 U4127 ( .A1(n4464), .A2(n4235), .ZN(n3611) );
  NAND2_X1 U4128 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  XNOR2_X1 U4129 ( .A(n3615), .B(n3613), .ZN(n4462) );
  INV_X1 U4130 ( .A(n3613), .ZN(n3614) );
  NAND2_X1 U4131 ( .A1(n3615), .A2(n3614), .ZN(n3616) );
  NAND2_X1 U4132 ( .A1(n4460), .A2(n3616), .ZN(n3632) );
  NAND2_X1 U4133 ( .A1(n4722), .A2(n4235), .ZN(n3618) );
  NAND2_X1 U4134 ( .A1(n5365), .A2(n4103), .ZN(n3617) );
  NAND2_X1 U4135 ( .A1(n3618), .A2(n3617), .ZN(n3619) );
  XNOR2_X1 U4136 ( .A(n3619), .B(n3093), .ZN(n3633) );
  NAND2_X1 U4137 ( .A1(n3632), .A2(n3633), .ZN(n5360) );
  NAND2_X1 U4138 ( .A1(n4722), .A2(n4239), .ZN(n3621) );
  NAND2_X1 U4139 ( .A1(n5365), .A2(n4235), .ZN(n3620) );
  NAND2_X1 U4140 ( .A1(n3621), .A2(n3620), .ZN(n5362) );
  NAND2_X1 U4141 ( .A1(n5360), .A2(n5362), .ZN(n4515) );
  NAND2_X1 U4142 ( .A1(n4998), .A2(n4235), .ZN(n3623) );
  NAND2_X1 U4143 ( .A1(n4518), .A2(n4103), .ZN(n3622) );
  NAND2_X1 U4144 ( .A1(n3623), .A2(n3622), .ZN(n3624) );
  XNOR2_X1 U4145 ( .A(n3624), .B(n3093), .ZN(n3627) );
  NAND2_X1 U4146 ( .A1(n4998), .A2(n4239), .ZN(n3626) );
  NAND2_X1 U4147 ( .A1(n4518), .A2(n4235), .ZN(n3625) );
  AND2_X1 U4148 ( .A1(n3626), .A2(n3625), .ZN(n3628) );
  NAND2_X1 U4149 ( .A1(n3627), .A2(n3628), .ZN(n3636) );
  INV_X1 U4150 ( .A(n3627), .ZN(n3630) );
  INV_X1 U4151 ( .A(n3628), .ZN(n3629) );
  NAND2_X1 U4152 ( .A1(n3630), .A2(n3629), .ZN(n3631) );
  AND2_X1 U4153 ( .A1(n3636), .A2(n3631), .ZN(n4514) );
  INV_X1 U4154 ( .A(n3632), .ZN(n3635) );
  INV_X1 U4155 ( .A(n3633), .ZN(n3634) );
  NAND3_X1 U4156 ( .A1(n4515), .A2(n4514), .A3(n5361), .ZN(n4513) );
  OAI21_X1 U4157 ( .B1(n3638), .B2(n3637), .A(n4052), .ZN(n3649) );
  INV_X1 U4158 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4322) );
  NAND2_X1 U4159 ( .A1(n3639), .A2(n4322), .ZN(n3640) );
  AND2_X1 U4160 ( .A1(n4069), .A2(n3640), .ZN(n4973) );
  NAND2_X1 U4161 ( .A1(n4973), .A2(n4287), .ZN(n3644) );
  NAND2_X1 U4162 ( .A1(n3106), .A2(REG0_REG_18__SCAN_IN), .ZN(n3643) );
  NAND2_X1 U4163 ( .A1(n2480), .A2(REG1_REG_18__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U4164 ( .A1(n3212), .A2(REG2_REG_18__SCAN_IN), .ZN(n3641) );
  NAND4_X1 U4165 ( .A1(n3644), .A2(n3643), .A3(n3642), .A4(n3641), .ZN(n4999)
         );
  AOI22_X1 U4166 ( .A1(n4547), .A2(n4999), .B1(n4369), .B2(n5364), .ZN(n3647)
         );
  INV_X1 U4167 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3645) );
  NOR2_X1 U4168 ( .A1(STATE_REG_SCAN_IN), .A2(n3645), .ZN(n4752) );
  AOI21_X1 U4169 ( .B1(n4558), .B2(n4998), .A(n4752), .ZN(n3646) );
  OAI211_X1 U4170 ( .C1(n5004), .C2(n5370), .A(n3647), .B(n3646), .ZN(n3648)
         );
  AOI21_X1 U4171 ( .B1(n3649), .B2(n5366), .A(n3648), .ZN(n3650) );
  INV_X1 U4172 ( .A(n3650), .ZN(U3225) );
  XNOR2_X1 U4173 ( .A(DATAI_31_), .B(keyinput_0), .ZN(n3653) );
  XNOR2_X1 U4174 ( .A(DATAI_30_), .B(keyinput_1), .ZN(n3652) );
  XNOR2_X1 U4175 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n3651) );
  OAI21_X1 U4176 ( .B1(n3653), .B2(n3652), .A(n3651), .ZN(n3659) );
  XNOR2_X1 U4177 ( .A(DATAI_28_), .B(keyinput_3), .ZN(n3658) );
  XOR2_X1 U4178 ( .A(DATAI_26_), .B(keyinput_5), .Z(n3656) );
  XOR2_X1 U4179 ( .A(DATAI_25_), .B(keyinput_6), .Z(n3655) );
  XNOR2_X1 U4180 ( .A(DATAI_27_), .B(keyinput_4), .ZN(n3654) );
  NAND3_X1 U4181 ( .A1(n3656), .A2(n3655), .A3(n3654), .ZN(n3657) );
  AOI21_X1 U4182 ( .B1(n3659), .B2(n3658), .A(n3657), .ZN(n3662) );
  XOR2_X1 U4183 ( .A(DATAI_23_), .B(keyinput_8), .Z(n3661) );
  XNOR2_X1 U4184 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n3660) );
  NOR3_X1 U4185 ( .A1(n3662), .A2(n3661), .A3(n3660), .ZN(n3665) );
  XOR2_X1 U4186 ( .A(DATAI_22_), .B(keyinput_9), .Z(n3664) );
  XNOR2_X1 U4187 ( .A(DATAI_21_), .B(keyinput_10), .ZN(n3663) );
  NOR3_X1 U4188 ( .A1(n3665), .A2(n3664), .A3(n3663), .ZN(n3668) );
  XOR2_X1 U4189 ( .A(DATAI_19_), .B(keyinput_12), .Z(n3667) );
  XNOR2_X1 U4190 ( .A(DATAI_20_), .B(keyinput_11), .ZN(n3666) );
  NOR3_X1 U4191 ( .A1(n3668), .A2(n3667), .A3(n3666), .ZN(n3671) );
  XNOR2_X1 U4192 ( .A(DATAI_17_), .B(keyinput_14), .ZN(n3670) );
  XNOR2_X1 U4193 ( .A(DATAI_18_), .B(keyinput_13), .ZN(n3669) );
  NOR3_X1 U4194 ( .A1(n3671), .A2(n3670), .A3(n3669), .ZN(n3674) );
  INV_X1 U4195 ( .A(DATAI_16_), .ZN(n5378) );
  XNOR2_X1 U4196 ( .A(n5378), .B(keyinput_15), .ZN(n3673) );
  XNOR2_X1 U4197 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n3672) );
  OAI21_X1 U4198 ( .B1(n3674), .B2(n3673), .A(n3672), .ZN(n3677) );
  XOR2_X1 U4199 ( .A(DATAI_14_), .B(keyinput_17), .Z(n3676) );
  XNOR2_X1 U4200 ( .A(DATAI_13_), .B(keyinput_18), .ZN(n3675) );
  NAND3_X1 U4201 ( .A1(n3677), .A2(n3676), .A3(n3675), .ZN(n3680) );
  XOR2_X1 U4202 ( .A(DATAI_12_), .B(keyinput_19), .Z(n3679) );
  XNOR2_X1 U4203 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n3678) );
  AOI21_X1 U4204 ( .B1(n3680), .B2(n3679), .A(n3678), .ZN(n3683) );
  INV_X1 U4205 ( .A(DATAI_9_), .ZN(n5270) );
  XNOR2_X1 U4206 ( .A(n5270), .B(keyinput_22), .ZN(n3682) );
  XNOR2_X1 U4207 ( .A(DATAI_10_), .B(keyinput_21), .ZN(n3681) );
  NOR3_X1 U4208 ( .A1(n3683), .A2(n3682), .A3(n3681), .ZN(n3686) );
  XNOR2_X1 U4209 ( .A(DATAI_8_), .B(keyinput_23), .ZN(n3685) );
  XNOR2_X1 U4210 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n3684) );
  NOR3_X1 U4211 ( .A1(n3686), .A2(n3685), .A3(n3684), .ZN(n3690) );
  XOR2_X1 U4212 ( .A(DATAI_4_), .B(keyinput_27), .Z(n3689) );
  XNOR2_X1 U4213 ( .A(DATAI_5_), .B(keyinput_26), .ZN(n3688) );
  XNOR2_X1 U4214 ( .A(DATAI_6_), .B(keyinput_25), .ZN(n3687) );
  NOR4_X1 U4215 ( .A1(n3690), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3693)
         );
  XOR2_X1 U4216 ( .A(DATAI_3_), .B(keyinput_28), .Z(n3692) );
  XNOR2_X1 U4217 ( .A(DATAI_2_), .B(keyinput_29), .ZN(n3691) );
  OAI21_X1 U4218 ( .B1(n3693), .B2(n3692), .A(n3691), .ZN(n3696) );
  XNOR2_X1 U4219 ( .A(DATAI_1_), .B(keyinput_30), .ZN(n3695) );
  XNOR2_X1 U4220 ( .A(DATAI_0_), .B(keyinput_31), .ZN(n3694) );
  AOI21_X1 U4221 ( .B1(n3696), .B2(n3695), .A(n3694), .ZN(n3699) );
  XNOR2_X1 U4222 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_33), .ZN(n3698) );
  XNOR2_X1 U4223 ( .A(STATE_REG_SCAN_IN), .B(keyinput_32), .ZN(n3697) );
  NOR3_X1 U4224 ( .A1(n3699), .A2(n3698), .A3(n3697), .ZN(n3702) );
  XOR2_X1 U4225 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_35), .Z(n3701) );
  XNOR2_X1 U4226 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_34), .ZN(n3700) );
  NOR3_X1 U4227 ( .A1(n3702), .A2(n3701), .A3(n3700), .ZN(n3706) );
  XNOR2_X1 U4228 ( .A(n4476), .B(keyinput_36), .ZN(n3705) );
  XOR2_X1 U4229 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_37), .Z(n3704) );
  XNOR2_X1 U4230 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_38), .ZN(n3703) );
  OAI211_X1 U4231 ( .C1(n3706), .C2(n3705), .A(n3704), .B(n3703), .ZN(n3709)
         );
  INV_X1 U4232 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4068) );
  XNOR2_X1 U4233 ( .A(n4068), .B(keyinput_39), .ZN(n3708) );
  XNOR2_X1 U4234 ( .A(n4279), .B(keyinput_40), .ZN(n3707) );
  AOI21_X1 U4235 ( .B1(n3709), .B2(n3708), .A(n3707), .ZN(n3713) );
  XNOR2_X1 U4236 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_41), .ZN(n3712) );
  XOR2_X1 U4237 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .Z(n3711) );
  XNOR2_X1 U4238 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_43), .ZN(n3710) );
  OAI211_X1 U4239 ( .C1(n3713), .C2(n3712), .A(n3711), .B(n3710), .ZN(n3716)
         );
  XOR2_X1 U4240 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_44), .Z(n3715) );
  XOR2_X1 U4241 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_45), .Z(n3714) );
  NAND3_X1 U4242 ( .A1(n3716), .A2(n3715), .A3(n3714), .ZN(n3720) );
  XNOR2_X1 U4243 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_46), .ZN(n3719) );
  XOR2_X1 U4244 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_48), .Z(n3718) );
  XOR2_X1 U4245 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_47), .Z(n3717) );
  AOI211_X1 U4246 ( .C1(n3720), .C2(n3719), .A(n3718), .B(n3717), .ZN(n3723)
         );
  XOR2_X1 U4247 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_50), .Z(n3722) );
  INV_X1 U4248 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4227) );
  XNOR2_X1 U4249 ( .A(n4227), .B(keyinput_49), .ZN(n3721) );
  NOR3_X1 U4250 ( .A1(n3723), .A2(n3722), .A3(n3721), .ZN(n3732) );
  INV_X1 U4251 ( .A(keyinput_52), .ZN(n3724) );
  XNOR2_X1 U4252 ( .A(n3724), .B(REG3_REG_0__SCAN_IN), .ZN(n3728) );
  XNOR2_X1 U4253 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_54), .ZN(n3727) );
  XNOR2_X1 U4254 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_53), .ZN(n3726) );
  XNOR2_X1 U4255 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput_51), .ZN(n3725) );
  NAND4_X1 U4256 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3731)
         );
  XOR2_X1 U4257 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_55), .Z(n3730) );
  OAI211_X1 U4258 ( .C1(n3732), .C2(n3731), .A(n3730), .B(n3729), .ZN(n3747)
         );
  XNOR2_X1 U4259 ( .A(n2683), .B(keyinput_58), .ZN(n3736) );
  XNOR2_X1 U4260 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n3735) );
  XNOR2_X1 U4261 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_57), .ZN(n3734) );
  XNOR2_X1 U4262 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_59), .ZN(n3733) );
  NOR4_X1 U4263 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3746)
         );
  XOR2_X1 U4264 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_64), .Z(n3739) );
  XNOR2_X1 U4265 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_67), .ZN(n3738) );
  XNOR2_X1 U4266 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .ZN(n3737) );
  NAND3_X1 U4267 ( .A1(n3739), .A2(n3738), .A3(n3737), .ZN(n3745) );
  XNOR2_X1 U4268 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_65), .ZN(n3743) );
  XNOR2_X1 U4269 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_66), .ZN(n3742) );
  XNOR2_X1 U4270 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n3741) );
  XNOR2_X1 U4271 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_62), .ZN(n3740) );
  NAND4_X1 U4272 ( .A1(n3743), .A2(n3742), .A3(n3741), .A4(n3740), .ZN(n3744)
         );
  AOI211_X1 U4273 ( .C1(n3747), .C2(n3746), .A(n3745), .B(n3744), .ZN(n3753)
         );
  XNOR2_X1 U4274 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_71), .ZN(n3749) );
  XNOR2_X1 U4275 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_68), .ZN(n3748) );
  NAND2_X1 U4276 ( .A1(n3749), .A2(n3748), .ZN(n3752) );
  XNOR2_X1 U4277 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_69), .ZN(n3751) );
  XNOR2_X1 U4278 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_70), .ZN(n3750) );
  NOR4_X1 U4279 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3759)
         );
  XNOR2_X1 U4280 ( .A(n3754), .B(keyinput_74), .ZN(n3758) );
  XNOR2_X1 U4281 ( .A(n3755), .B(keyinput_73), .ZN(n3757) );
  XNOR2_X1 U4282 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_72), .ZN(n3756) );
  NOR4_X1 U4283 ( .A1(n3759), .A2(n3758), .A3(n3757), .A4(n3756), .ZN(n3763)
         );
  XNOR2_X1 U4284 ( .A(n3947), .B(keyinput_75), .ZN(n3762) );
  XOR2_X1 U4285 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_76), .Z(n3761) );
  XNOR2_X1 U4286 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_77), .ZN(n3760) );
  OAI211_X1 U4287 ( .C1(n3763), .C2(n3762), .A(n3761), .B(n3760), .ZN(n3770)
         );
  XNOR2_X1 U4288 ( .A(n3952), .B(keyinput_78), .ZN(n3769) );
  XNOR2_X1 U4289 ( .A(n3764), .B(keyinput_81), .ZN(n3767) );
  XNOR2_X1 U4290 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_79), .ZN(n3766) );
  XNOR2_X1 U4291 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_80), .ZN(n3765) );
  NAND3_X1 U4292 ( .A1(n3767), .A2(n3766), .A3(n3765), .ZN(n3768) );
  AOI21_X1 U4293 ( .B1(n3770), .B2(n3769), .A(n3768), .ZN(n3773) );
  XNOR2_X1 U4294 ( .A(n3959), .B(keyinput_82), .ZN(n3772) );
  XNOR2_X1 U4295 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_83), .ZN(n3771) );
  OAI21_X1 U4296 ( .B1(n3773), .B2(n3772), .A(n3771), .ZN(n3778) );
  XOR2_X1 U4297 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_84), .Z(n3777) );
  XNOR2_X1 U4298 ( .A(n3774), .B(keyinput_85), .ZN(n3776) );
  XNOR2_X1 U4299 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_86), .ZN(n3775) );
  AOI211_X1 U4300 ( .C1(n3778), .C2(n3777), .A(n3776), .B(n3775), .ZN(n3782)
         );
  XNOR2_X1 U4301 ( .A(D_REG_0__SCAN_IN), .B(keyinput_87), .ZN(n3781) );
  INV_X1 U4302 ( .A(D_REG_2__SCAN_IN), .ZN(n5113) );
  XNOR2_X1 U4303 ( .A(n5113), .B(keyinput_89), .ZN(n3780) );
  XNOR2_X1 U4304 ( .A(D_REG_1__SCAN_IN), .B(keyinput_88), .ZN(n3779) );
  OAI211_X1 U4305 ( .C1(n3782), .C2(n3781), .A(n3780), .B(n3779), .ZN(n3785)
         );
  XOR2_X1 U4306 ( .A(D_REG_3__SCAN_IN), .B(keyinput_90), .Z(n3784) );
  XNOR2_X1 U4307 ( .A(D_REG_4__SCAN_IN), .B(keyinput_91), .ZN(n3783) );
  NAND3_X1 U4308 ( .A1(n3785), .A2(n3784), .A3(n3783), .ZN(n3792) );
  XOR2_X1 U4309 ( .A(D_REG_5__SCAN_IN), .B(keyinput_92), .Z(n3791) );
  XOR2_X1 U4310 ( .A(D_REG_6__SCAN_IN), .B(keyinput_93), .Z(n3789) );
  XNOR2_X1 U4311 ( .A(D_REG_9__SCAN_IN), .B(keyinput_96), .ZN(n3788) );
  XNOR2_X1 U4312 ( .A(D_REG_8__SCAN_IN), .B(keyinput_95), .ZN(n3787) );
  XNOR2_X1 U4313 ( .A(D_REG_7__SCAN_IN), .B(keyinput_94), .ZN(n3786) );
  NAND4_X1 U4314 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3790)
         );
  AOI21_X1 U4315 ( .B1(n3792), .B2(n3791), .A(n3790), .ZN(n3795) );
  INV_X1 U4316 ( .A(D_REG_10__SCAN_IN), .ZN(n5118) );
  XNOR2_X1 U4317 ( .A(n5118), .B(keyinput_97), .ZN(n3794) );
  XNOR2_X1 U4318 ( .A(D_REG_11__SCAN_IN), .B(keyinput_98), .ZN(n3793) );
  NOR3_X1 U4319 ( .A1(n3795), .A2(n3794), .A3(n3793), .ZN(n3798) );
  INV_X1 U4320 ( .A(D_REG_12__SCAN_IN), .ZN(n5119) );
  XNOR2_X1 U4321 ( .A(n5119), .B(keyinput_99), .ZN(n3797) );
  XNOR2_X1 U4322 ( .A(D_REG_13__SCAN_IN), .B(keyinput_100), .ZN(n3796) );
  OAI21_X1 U4323 ( .B1(n3798), .B2(n3797), .A(n3796), .ZN(n3802) );
  XNOR2_X1 U4324 ( .A(D_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n3801) );
  XNOR2_X1 U4325 ( .A(D_REG_15__SCAN_IN), .B(keyinput_102), .ZN(n3800) );
  XNOR2_X1 U4326 ( .A(D_REG_16__SCAN_IN), .B(keyinput_103), .ZN(n3799) );
  NAND4_X1 U4327 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n3806)
         );
  XOR2_X1 U4328 ( .A(D_REG_17__SCAN_IN), .B(keyinput_104), .Z(n3805) );
  INV_X1 U4329 ( .A(D_REG_19__SCAN_IN), .ZN(n5125) );
  XNOR2_X1 U4330 ( .A(n5125), .B(keyinput_106), .ZN(n3804) );
  INV_X1 U4331 ( .A(D_REG_18__SCAN_IN), .ZN(n5124) );
  XNOR2_X1 U4332 ( .A(n5124), .B(keyinput_105), .ZN(n3803) );
  AOI211_X1 U4333 ( .C1(n3806), .C2(n3805), .A(n3804), .B(n3803), .ZN(n3809)
         );
  INV_X1 U4334 ( .A(D_REG_20__SCAN_IN), .ZN(n5126) );
  XNOR2_X1 U4335 ( .A(n5126), .B(keyinput_107), .ZN(n3808) );
  INV_X1 U4336 ( .A(D_REG_21__SCAN_IN), .ZN(n5127) );
  XNOR2_X1 U4337 ( .A(n5127), .B(keyinput_108), .ZN(n3807) );
  NOR3_X1 U4338 ( .A1(n3809), .A2(n3808), .A3(n3807), .ZN(n3817) );
  XOR2_X1 U4339 ( .A(D_REG_24__SCAN_IN), .B(keyinput_111), .Z(n3813) );
  XOR2_X1 U4340 ( .A(D_REG_25__SCAN_IN), .B(keyinput_112), .Z(n3812) );
  XNOR2_X1 U4341 ( .A(D_REG_23__SCAN_IN), .B(keyinput_110), .ZN(n3811) );
  XNOR2_X1 U4342 ( .A(D_REG_22__SCAN_IN), .B(keyinput_109), .ZN(n3810) );
  NAND4_X1 U4343 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3816)
         );
  INV_X1 U4344 ( .A(D_REG_27__SCAN_IN), .ZN(n5131) );
  XNOR2_X1 U4345 ( .A(n5131), .B(keyinput_114), .ZN(n3815) );
  XOR2_X1 U4346 ( .A(D_REG_26__SCAN_IN), .B(keyinput_113), .Z(n3814) );
  OAI211_X1 U4347 ( .C1(n3817), .C2(n3816), .A(n3815), .B(n3814), .ZN(n3821)
         );
  INV_X1 U4348 ( .A(D_REG_28__SCAN_IN), .ZN(n5132) );
  XNOR2_X1 U4349 ( .A(n5132), .B(keyinput_115), .ZN(n3820) );
  XNOR2_X1 U4350 ( .A(D_REG_29__SCAN_IN), .B(keyinput_116), .ZN(n3819) );
  XNOR2_X1 U4351 ( .A(D_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n3818) );
  NAND4_X1 U4352 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3824)
         );
  XOR2_X1 U4353 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_119), .Z(n3823) );
  XNOR2_X1 U4354 ( .A(D_REG_31__SCAN_IN), .B(keyinput_118), .ZN(n3822) );
  NAND3_X1 U4355 ( .A1(n3824), .A2(n3823), .A3(n3822), .ZN(n3827) );
  XNOR2_X1 U4356 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_120), .ZN(n3826) );
  XOR2_X1 U4357 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_121), .Z(n3825) );
  AOI21_X1 U4358 ( .B1(n3827), .B2(n3826), .A(n3825), .ZN(n3830) );
  XOR2_X1 U4359 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_122), .Z(n3829) );
  XNOR2_X1 U4360 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_123), .ZN(n3828) );
  NOR3_X1 U4361 ( .A1(n3830), .A2(n3829), .A3(n3828), .ZN(n4028) );
  XOR2_X1 U4362 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_124), .Z(n4027) );
  XNOR2_X1 U4363 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_125), .ZN(n3833) );
  XNOR2_X1 U4364 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_127), .ZN(n3832) );
  XNOR2_X1 U4365 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_126), .ZN(n3831) );
  NOR3_X1 U4366 ( .A1(n3833), .A2(n3832), .A3(n3831), .ZN(n4026) );
  XNOR2_X1 U4367 ( .A(DATAI_30_), .B(keyinput_129), .ZN(n3836) );
  XNOR2_X1 U4368 ( .A(DATAI_31_), .B(keyinput_128), .ZN(n3835) );
  XOR2_X1 U4369 ( .A(DATAI_29_), .B(keyinput_130), .Z(n3834) );
  OAI21_X1 U4370 ( .B1(n3836), .B2(n3835), .A(n3834), .ZN(n3842) );
  XNOR2_X1 U4371 ( .A(DATAI_28_), .B(keyinput_131), .ZN(n3841) );
  XOR2_X1 U4372 ( .A(DATAI_25_), .B(keyinput_134), .Z(n3839) );
  XNOR2_X1 U4373 ( .A(DATAI_27_), .B(keyinput_132), .ZN(n3838) );
  XNOR2_X1 U4374 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n3837) );
  NAND3_X1 U4375 ( .A1(n3839), .A2(n3838), .A3(n3837), .ZN(n3840) );
  AOI21_X1 U4376 ( .B1(n3842), .B2(n3841), .A(n3840), .ZN(n3845) );
  XNOR2_X1 U4377 ( .A(DATAI_23_), .B(keyinput_136), .ZN(n3844) );
  XNOR2_X1 U4378 ( .A(DATAI_24_), .B(keyinput_135), .ZN(n3843) );
  NOR3_X1 U4379 ( .A1(n3845), .A2(n3844), .A3(n3843), .ZN(n3848) );
  XOR2_X1 U4380 ( .A(DATAI_22_), .B(keyinput_137), .Z(n3847) );
  XOR2_X1 U4381 ( .A(DATAI_21_), .B(keyinput_138), .Z(n3846) );
  NOR3_X1 U4382 ( .A1(n3848), .A2(n3847), .A3(n3846), .ZN(n3851) );
  XOR2_X1 U4383 ( .A(DATAI_20_), .B(keyinput_139), .Z(n3850) );
  XOR2_X1 U4384 ( .A(DATAI_19_), .B(keyinput_140), .Z(n3849) );
  NOR3_X1 U4385 ( .A1(n3851), .A2(n3850), .A3(n3849), .ZN(n3854) );
  XOR2_X1 U4386 ( .A(DATAI_18_), .B(keyinput_141), .Z(n3853) );
  XNOR2_X1 U4387 ( .A(DATAI_17_), .B(keyinput_142), .ZN(n3852) );
  NOR3_X1 U4388 ( .A1(n3854), .A2(n3853), .A3(n3852), .ZN(n3857) );
  XNOR2_X1 U4389 ( .A(n5378), .B(keyinput_143), .ZN(n3856) );
  INV_X1 U4390 ( .A(DATAI_15_), .ZN(n5356) );
  XNOR2_X1 U4391 ( .A(n5356), .B(keyinput_144), .ZN(n3855) );
  OAI21_X1 U4392 ( .B1(n3857), .B2(n3856), .A(n3855), .ZN(n3860) );
  XNOR2_X1 U4393 ( .A(DATAI_14_), .B(keyinput_145), .ZN(n3859) );
  XNOR2_X1 U4394 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n3858) );
  NAND3_X1 U4395 ( .A1(n3860), .A2(n3859), .A3(n3858), .ZN(n3863) );
  XOR2_X1 U4396 ( .A(DATAI_12_), .B(keyinput_147), .Z(n3862) );
  XNOR2_X1 U4397 ( .A(DATAI_11_), .B(keyinput_148), .ZN(n3861) );
  AOI21_X1 U4398 ( .B1(n3863), .B2(n3862), .A(n3861), .ZN(n3866) );
  XNOR2_X1 U4399 ( .A(n5270), .B(keyinput_150), .ZN(n3865) );
  INV_X1 U4400 ( .A(DATAI_10_), .ZN(n5281) );
  XNOR2_X1 U4401 ( .A(n5281), .B(keyinput_149), .ZN(n3864) );
  NOR3_X1 U4402 ( .A1(n3866), .A2(n3865), .A3(n3864), .ZN(n3869) );
  XOR2_X1 U4403 ( .A(DATAI_8_), .B(keyinput_151), .Z(n3868) );
  XNOR2_X1 U4404 ( .A(DATAI_7_), .B(keyinput_152), .ZN(n3867) );
  NOR3_X1 U4405 ( .A1(n3869), .A2(n3868), .A3(n3867), .ZN(n3873) );
  XOR2_X1 U4406 ( .A(DATAI_4_), .B(keyinput_155), .Z(n3872) );
  INV_X1 U4407 ( .A(DATAI_5_), .ZN(n5217) );
  XNOR2_X1 U4408 ( .A(n5217), .B(keyinput_154), .ZN(n3871) );
  XNOR2_X1 U4409 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n3870) );
  NOR4_X1 U4410 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3876)
         );
  XOR2_X1 U4411 ( .A(DATAI_3_), .B(keyinput_156), .Z(n3875) );
  XNOR2_X1 U4412 ( .A(DATAI_2_), .B(keyinput_157), .ZN(n3874) );
  OAI21_X1 U4413 ( .B1(n3876), .B2(n3875), .A(n3874), .ZN(n3879) );
  INV_X1 U4414 ( .A(DATAI_1_), .ZN(n5163) );
  XNOR2_X1 U4415 ( .A(n5163), .B(keyinput_158), .ZN(n3878) );
  XNOR2_X1 U4416 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n3877) );
  AOI21_X1 U4417 ( .B1(n3879), .B2(n3878), .A(n3877), .ZN(n3882) );
  XNOR2_X1 U4418 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_161), .ZN(n3881) );
  XNOR2_X1 U4419 ( .A(STATE_REG_SCAN_IN), .B(keyinput_160), .ZN(n3880) );
  NOR3_X1 U4420 ( .A1(n3882), .A2(n3881), .A3(n3880), .ZN(n3885) );
  INV_X1 U4421 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4264) );
  XNOR2_X1 U4422 ( .A(n4264), .B(keyinput_162), .ZN(n3884) );
  XOR2_X1 U4423 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_163), .Z(n3883) );
  NOR3_X1 U4424 ( .A1(n3885), .A2(n3884), .A3(n3883), .ZN(n3889) );
  XNOR2_X1 U4425 ( .A(n4476), .B(keyinput_164), .ZN(n3888) );
  XNOR2_X1 U4426 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_166), .ZN(n3887) );
  XNOR2_X1 U4427 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_165), .ZN(n3886) );
  OAI211_X1 U4428 ( .C1(n3889), .C2(n3888), .A(n3887), .B(n3886), .ZN(n3892)
         );
  XNOR2_X1 U4429 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_167), .ZN(n3891) );
  XNOR2_X1 U4430 ( .A(n4279), .B(keyinput_168), .ZN(n3890) );
  AOI21_X1 U4431 ( .B1(n3892), .B2(n3891), .A(n3890), .ZN(n3896) );
  XNOR2_X1 U4432 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_169), .ZN(n3895) );
  XNOR2_X1 U4433 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_170), .ZN(n3894) );
  XNOR2_X1 U4434 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_171), .ZN(n3893) );
  OAI211_X1 U4435 ( .C1(n3896), .C2(n3895), .A(n3894), .B(n3893), .ZN(n3899)
         );
  XOR2_X1 U4436 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_172), .Z(n3898) );
  XOR2_X1 U4437 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_173), .Z(n3897) );
  NAND3_X1 U4438 ( .A1(n3899), .A2(n3898), .A3(n3897), .ZN(n3903) );
  XNOR2_X1 U4439 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_174), .ZN(n3902) );
  XOR2_X1 U4440 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_176), .Z(n3901) );
  XOR2_X1 U4441 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_175), .Z(n3900) );
  AOI211_X1 U4442 ( .C1(n3903), .C2(n3902), .A(n3901), .B(n3900), .ZN(n3906)
         );
  XNOR2_X1 U4443 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_178), .ZN(n3905) );
  XNOR2_X1 U4444 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_177), .ZN(n3904) );
  NOR3_X1 U4445 ( .A1(n3906), .A2(n3905), .A3(n3904), .ZN(n3914) );
  XOR2_X1 U4446 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .Z(n3910) );
  INV_X1 U4447 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4138) );
  XNOR2_X1 U4448 ( .A(n4138), .B(keyinput_182), .ZN(n3909) );
  XNOR2_X1 U4449 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_181), .ZN(n3908) );
  XNOR2_X1 U4450 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput_179), .ZN(n3907) );
  NAND4_X1 U4451 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3913)
         );
  XOR2_X1 U4452 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_183), .Z(n3912) );
  OAI211_X1 U4453 ( .C1(n3914), .C2(n3913), .A(n3912), .B(n3911), .ZN(n3933)
         );
  XNOR2_X1 U4454 ( .A(n3915), .B(keyinput_187), .ZN(n3919) );
  XNOR2_X1 U4455 ( .A(n2683), .B(keyinput_186), .ZN(n3918) );
  XNOR2_X1 U4456 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_185), .ZN(n3917) );
  XNOR2_X1 U4457 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_188), .ZN(n3916) );
  NOR4_X1 U4458 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3932)
         );
  INV_X1 U4459 ( .A(IR_REG_10__SCAN_IN), .ZN(n3926) );
  INV_X1 U4460 ( .A(keyinput_193), .ZN(n3925) );
  AOI22_X1 U4461 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput_194), .B1(
        IR_REG_10__SCAN_IN), .B2(keyinput_193), .ZN(n3921) );
  AOI22_X1 U4462 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput_192), .B1(n3922), .B2(
        keyinput_189), .ZN(n3920) );
  OAI211_X1 U4463 ( .C1(IR_REG_9__SCAN_IN), .C2(keyinput_192), .A(n3921), .B(
        n3920), .ZN(n3924) );
  OAI22_X1 U4464 ( .A1(n3922), .A2(keyinput_189), .B1(IR_REG_11__SCAN_IN), 
        .B2(keyinput_194), .ZN(n3923) );
  AOI211_X1 U4465 ( .C1(n3926), .C2(n3925), .A(n3924), .B(n3923), .ZN(n3930)
         );
  XNOR2_X1 U4466 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_191), .ZN(n3929) );
  XNOR2_X1 U4467 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_195), .ZN(n3928) );
  XNOR2_X1 U4468 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_190), .ZN(n3927) );
  NAND4_X1 U4469 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3931)
         );
  AOI21_X1 U4470 ( .B1(n3933), .B2(n3932), .A(n3931), .ZN(n3941) );
  XNOR2_X1 U4471 ( .A(n3934), .B(keyinput_196), .ZN(n3939) );
  XNOR2_X1 U4472 ( .A(n3935), .B(keyinput_199), .ZN(n3938) );
  XNOR2_X1 U4473 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_198), .ZN(n3937) );
  XNOR2_X1 U4474 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_197), .ZN(n3936) );
  NAND4_X1 U4475 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3940)
         );
  NOR2_X1 U4476 ( .A1(n3941), .A2(n3940), .ZN(n3946) );
  XNOR2_X1 U4477 ( .A(n3942), .B(keyinput_200), .ZN(n3945) );
  XNOR2_X1 U4478 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_202), .ZN(n3944) );
  XNOR2_X1 U4479 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_201), .ZN(n3943) );
  NOR4_X1 U4480 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3951)
         );
  XNOR2_X1 U4481 ( .A(n3947), .B(keyinput_203), .ZN(n3950) );
  XOR2_X1 U4482 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_204), .Z(n3949) );
  XNOR2_X1 U4483 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_205), .ZN(n3948) );
  OAI211_X1 U4484 ( .C1(n3951), .C2(n3950), .A(n3949), .B(n3948), .ZN(n3958)
         );
  XNOR2_X1 U4485 ( .A(n3952), .B(keyinput_206), .ZN(n3957) );
  XOR2_X1 U4486 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_207), .Z(n3955) );
  XOR2_X1 U4487 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_208), .Z(n3954) );
  XNOR2_X1 U4488 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_209), .ZN(n3953) );
  NAND3_X1 U4489 ( .A1(n3955), .A2(n3954), .A3(n3953), .ZN(n3956) );
  AOI21_X1 U4490 ( .B1(n3958), .B2(n3957), .A(n3956), .ZN(n3962) );
  XNOR2_X1 U4491 ( .A(n3959), .B(keyinput_210), .ZN(n3961) );
  XNOR2_X1 U4492 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_211), .ZN(n3960) );
  OAI21_X1 U4493 ( .B1(n3962), .B2(n3961), .A(n3960), .ZN(n3966) );
  XNOR2_X1 U4494 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_212), .ZN(n3965) );
  XOR2_X1 U4495 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_214), .Z(n3964) );
  XNOR2_X1 U4496 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_213), .ZN(n3963) );
  AOI211_X1 U4497 ( .C1(n3966), .C2(n3965), .A(n3964), .B(n3963), .ZN(n3970)
         );
  XNOR2_X1 U4498 ( .A(D_REG_0__SCAN_IN), .B(keyinput_215), .ZN(n3969) );
  XNOR2_X1 U4499 ( .A(D_REG_1__SCAN_IN), .B(keyinput_216), .ZN(n3968) );
  XNOR2_X1 U4500 ( .A(D_REG_2__SCAN_IN), .B(keyinput_217), .ZN(n3967) );
  OAI211_X1 U4501 ( .C1(n3970), .C2(n3969), .A(n3968), .B(n3967), .ZN(n3973)
         );
  XOR2_X1 U4502 ( .A(D_REG_3__SCAN_IN), .B(keyinput_218), .Z(n3972) );
  INV_X1 U4503 ( .A(D_REG_4__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U4504 ( .A(n5114), .B(keyinput_219), .ZN(n3971) );
  NAND3_X1 U4505 ( .A1(n3973), .A2(n3972), .A3(n3971), .ZN(n3980) );
  XNOR2_X1 U4506 ( .A(D_REG_5__SCAN_IN), .B(keyinput_220), .ZN(n3979) );
  XOR2_X1 U4507 ( .A(D_REG_6__SCAN_IN), .B(keyinput_221), .Z(n3977) );
  XNOR2_X1 U4508 ( .A(D_REG_8__SCAN_IN), .B(keyinput_223), .ZN(n3976) );
  XNOR2_X1 U4509 ( .A(D_REG_9__SCAN_IN), .B(keyinput_224), .ZN(n3975) );
  XNOR2_X1 U4510 ( .A(D_REG_7__SCAN_IN), .B(keyinput_222), .ZN(n3974) );
  NAND4_X1 U4511 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3978)
         );
  AOI21_X1 U4512 ( .B1(n3980), .B2(n3979), .A(n3978), .ZN(n3983) );
  XNOR2_X1 U4513 ( .A(n5118), .B(keyinput_225), .ZN(n3982) );
  XNOR2_X1 U4514 ( .A(D_REG_11__SCAN_IN), .B(keyinput_226), .ZN(n3981) );
  NOR3_X1 U4515 ( .A1(n3983), .A2(n3982), .A3(n3981), .ZN(n3986) );
  XNOR2_X1 U4516 ( .A(n5119), .B(keyinput_227), .ZN(n3985) );
  XNOR2_X1 U4517 ( .A(D_REG_13__SCAN_IN), .B(keyinput_228), .ZN(n3984) );
  OAI21_X1 U4518 ( .B1(n3986), .B2(n3985), .A(n3984), .ZN(n3990) );
  INV_X1 U4519 ( .A(D_REG_14__SCAN_IN), .ZN(n5121) );
  XNOR2_X1 U4520 ( .A(n5121), .B(keyinput_229), .ZN(n3989) );
  INV_X1 U4521 ( .A(D_REG_15__SCAN_IN), .ZN(n5122) );
  XNOR2_X1 U4522 ( .A(n5122), .B(keyinput_230), .ZN(n3988) );
  XNOR2_X1 U4523 ( .A(D_REG_16__SCAN_IN), .B(keyinput_231), .ZN(n3987) );
  NAND4_X1 U4524 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n3994)
         );
  XOR2_X1 U4525 ( .A(D_REG_17__SCAN_IN), .B(keyinput_232), .Z(n3993) );
  XNOR2_X1 U4526 ( .A(n5124), .B(keyinput_233), .ZN(n3992) );
  XNOR2_X1 U4527 ( .A(D_REG_19__SCAN_IN), .B(keyinput_234), .ZN(n3991) );
  AOI211_X1 U4528 ( .C1(n3994), .C2(n3993), .A(n3992), .B(n3991), .ZN(n3997)
         );
  XNOR2_X1 U4529 ( .A(n5126), .B(keyinput_235), .ZN(n3996) );
  XNOR2_X1 U4530 ( .A(n5127), .B(keyinput_236), .ZN(n3995) );
  NOR3_X1 U4531 ( .A1(n3997), .A2(n3996), .A3(n3995), .ZN(n4005) );
  XOR2_X1 U4532 ( .A(D_REG_25__SCAN_IN), .B(keyinput_240), .Z(n4001) );
  XOR2_X1 U4533 ( .A(D_REG_24__SCAN_IN), .B(keyinput_239), .Z(n4000) );
  INV_X1 U4534 ( .A(D_REG_23__SCAN_IN), .ZN(n5129) );
  XNOR2_X1 U4535 ( .A(n5129), .B(keyinput_238), .ZN(n3999) );
  XNOR2_X1 U4536 ( .A(D_REG_22__SCAN_IN), .B(keyinput_237), .ZN(n3998) );
  NAND4_X1 U4537 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4004)
         );
  XOR2_X1 U4538 ( .A(D_REG_26__SCAN_IN), .B(keyinput_241), .Z(n4003) );
  XNOR2_X1 U4539 ( .A(D_REG_27__SCAN_IN), .B(keyinput_242), .ZN(n4002) );
  OAI211_X1 U4540 ( .C1(n4005), .C2(n4004), .A(n4003), .B(n4002), .ZN(n4009)
         );
  XNOR2_X1 U4541 ( .A(D_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n4008) );
  XNOR2_X1 U4542 ( .A(D_REG_28__SCAN_IN), .B(keyinput_243), .ZN(n4007) );
  XNOR2_X1 U4543 ( .A(D_REG_29__SCAN_IN), .B(keyinput_244), .ZN(n4006) );
  NAND4_X1 U4544 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4012)
         );
  XOR2_X1 U4545 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_247), .Z(n4011) );
  XNOR2_X1 U4546 ( .A(D_REG_31__SCAN_IN), .B(keyinput_246), .ZN(n4010) );
  NAND3_X1 U4547 ( .A1(n4012), .A2(n4011), .A3(n4010), .ZN(n4015) );
  XNOR2_X1 U4548 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_248), .ZN(n4014) );
  XOR2_X1 U4549 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_249), .Z(n4013) );
  AOI21_X1 U4550 ( .B1(n4015), .B2(n4014), .A(n4013), .ZN(n4018) );
  XOR2_X1 U4551 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_250), .Z(n4017) );
  XOR2_X1 U4552 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_251), .Z(n4016) );
  NOR3_X1 U4553 ( .A1(n4018), .A2(n4017), .A3(n4016), .ZN(n4024) );
  XOR2_X1 U4554 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_252), .Z(n4023) );
  XOR2_X1 U4555 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_254), .Z(n4021) );
  XNOR2_X1 U4556 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .ZN(n4020) );
  XNOR2_X1 U4557 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_255), .ZN(n4019) );
  NOR3_X1 U4558 ( .A1(n4021), .A2(n4020), .A3(n4019), .ZN(n4022) );
  OAI21_X1 U4559 ( .B1(n4024), .B2(n4023), .A(n4022), .ZN(n4025) );
  OAI211_X1 U4560 ( .C1(n4028), .C2(n4027), .A(n4026), .B(n4025), .ZN(n4030)
         );
  MUX2_X1 U4561 ( .A(n4152), .B(DATAI_13_), .S(U3149), .Z(n4029) );
  XNOR2_X1 U4562 ( .A(n4030), .B(n4029), .ZN(U3339) );
  NAND2_X1 U4563 ( .A1(n4722), .A2(n5365), .ZN(n4032) );
  INV_X1 U4564 ( .A(n4722), .ZN(n4565) );
  INV_X1 U4565 ( .A(n5365), .ZN(n4036) );
  AOI21_X1 U4566 ( .B1(n4033), .B2(n4032), .A(n4031), .ZN(n4348) );
  INV_X1 U4567 ( .A(n4998), .ZN(n4350) );
  AND2_X1 U4568 ( .A1(n4350), .A2(n4518), .ZN(n4691) );
  NAND2_X1 U4569 ( .A1(n4349), .A2(n4998), .ZN(n4929) );
  INV_X1 U4570 ( .A(n4929), .ZN(n4034) );
  NOR2_X1 U4571 ( .A1(n4691), .A2(n4034), .ZN(n4364) );
  INV_X1 U4572 ( .A(n4364), .ZN(n4605) );
  XNOR2_X1 U4573 ( .A(n4348), .B(n4605), .ZN(n5382) );
  NAND3_X1 U4574 ( .A1(n4035), .A2(n4633), .A3(n4566), .ZN(n4037) );
  NAND2_X1 U4575 ( .A1(n4036), .A2(n4722), .ZN(n4568) );
  NAND2_X1 U4576 ( .A1(n4037), .A2(n4568), .ZN(n4365) );
  XNOR2_X1 U4577 ( .A(n4365), .B(n4605), .ZN(n4038) );
  NAND2_X1 U4578 ( .A1(n4038), .A2(n5333), .ZN(n4040) );
  AOI22_X1 U4579 ( .A1(n5302), .A2(n4721), .B1(n4722), .B2(n5304), .ZN(n4039)
         );
  OAI211_X1 U4580 ( .C1(n5330), .C2(n4349), .A(n4040), .B(n4039), .ZN(n5384)
         );
  INV_X1 U4581 ( .A(n4992), .ZN(n4041) );
  OAI21_X1 U4582 ( .B1(n4042), .B2(n4349), .A(n4041), .ZN(n5380) );
  NOR2_X1 U4583 ( .A1(n5380), .A2(n5010), .ZN(n4046) );
  INV_X1 U4584 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4044) );
  INV_X1 U4585 ( .A(n4521), .ZN(n4043) );
  OAI22_X1 U4586 ( .A1(n5262), .A2(n4044), .B1(n4043), .B2(n5339), .ZN(n4045)
         );
  AOI211_X1 U4587 ( .C1(n5384), .C2(n5262), .A(n4046), .B(n4045), .ZN(n4047)
         );
  OAI21_X1 U4588 ( .B1(n5382), .B2(n4991), .A(n4047), .ZN(U3274) );
  INV_X1 U4589 ( .A(n4048), .ZN(n4049) );
  NAND2_X1 U4590 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  NAND2_X1 U4591 ( .A1(n4999), .A2(n4235), .ZN(n4054) );
  NAND2_X1 U4592 ( .A1(n4984), .A2(n4103), .ZN(n4053) );
  NAND2_X1 U4593 ( .A1(n4054), .A2(n4053), .ZN(n4055) );
  XNOR2_X1 U4594 ( .A(n4055), .B(n3296), .ZN(n4058) );
  NAND2_X1 U4595 ( .A1(n4999), .A2(n4239), .ZN(n4057) );
  NAND2_X1 U4596 ( .A1(n4984), .A2(n4235), .ZN(n4056) );
  NAND2_X1 U4597 ( .A1(n4057), .A2(n4056), .ZN(n4059) );
  NAND2_X1 U4598 ( .A1(n4058), .A2(n4059), .ZN(n4063) );
  INV_X1 U4599 ( .A(n4079), .ZN(n4065) );
  INV_X1 U4600 ( .A(n4058), .ZN(n4061) );
  INV_X1 U4601 ( .A(n4059), .ZN(n4060) );
  NAND2_X1 U4602 ( .A1(n4061), .A2(n4060), .ZN(n4078) );
  AOI21_X1 U4603 ( .B1(n4063), .B2(n4078), .A(n4062), .ZN(n4064) );
  AOI21_X1 U4604 ( .B1(n4065), .B2(n4078), .A(n4064), .ZN(n4077) );
  INV_X1 U4605 ( .A(REG0_REG_19__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U4606 ( .A1(n2480), .A2(REG1_REG_19__SCAN_IN), .ZN(n4067) );
  NAND2_X1 U4607 ( .A1(n3212), .A2(REG2_REG_19__SCAN_IN), .ZN(n4066) );
  AND2_X1 U4608 ( .A1(n4067), .A2(n4066), .ZN(n4072) );
  NAND2_X1 U4609 ( .A1(n4069), .A2(n4068), .ZN(n4070) );
  NAND2_X1 U4610 ( .A1(n4083), .A2(n4070), .ZN(n4965) );
  OR2_X1 U4611 ( .A1(n4965), .A2(n4267), .ZN(n4071) );
  NAND2_X1 U4612 ( .A1(n4943), .A2(n5302), .ZN(n4074) );
  NAND2_X1 U4613 ( .A1(n4721), .A2(n5304), .ZN(n4073) );
  NAND2_X1 U4614 ( .A1(n4074), .A2(n4073), .ZN(n4986) );
  AOI22_X1 U4615 ( .A1(n4986), .A2(n5359), .B1(REG3_REG_18__SCAN_IN), .B2(
        U3149), .ZN(n4076) );
  AOI22_X1 U4616 ( .A1(n4973), .A2(n4522), .B1(n5364), .B2(n4984), .ZN(n4075)
         );
  OAI211_X1 U4617 ( .C1(n4077), .C2(n5315), .A(n4076), .B(n4075), .ZN(U3235)
         );
  NAND2_X1 U4618 ( .A1(n4079), .A2(n4078), .ZN(n4097) );
  NAND2_X1 U4619 ( .A1(n4943), .A2(n4235), .ZN(n4081) );
  NAND2_X1 U4620 ( .A1(n4962), .A2(n4103), .ZN(n4080) );
  NAND2_X1 U4621 ( .A1(n4081), .A2(n4080), .ZN(n4082) );
  XNOR2_X1 U4622 ( .A(n4082), .B(n3296), .ZN(n4098) );
  AOI22_X1 U4623 ( .A1(n4943), .A2(n4239), .B1(n4962), .B2(n4235), .ZN(n4099)
         );
  XNOR2_X1 U4624 ( .A(n4098), .B(n4099), .ZN(n4096) );
  XOR2_X1 U4625 ( .A(n4097), .B(n4096), .Z(n4095) );
  INV_X1 U4626 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4122) );
  NAND2_X1 U4627 ( .A1(n4083), .A2(n4122), .ZN(n4084) );
  NAND2_X1 U4628 ( .A1(n4115), .A2(n4084), .ZN(n4926) );
  INV_X1 U4629 ( .A(REG0_REG_20__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U4630 ( .A1(n2480), .A2(REG1_REG_20__SCAN_IN), .ZN(n4086) );
  NAND2_X1 U4631 ( .A1(n3212), .A2(REG2_REG_20__SCAN_IN), .ZN(n4085) );
  OAI211_X1 U4632 ( .C1(n5082), .C2(n4285), .A(n4086), .B(n4085), .ZN(n4087)
         );
  INV_X1 U4633 ( .A(n4087), .ZN(n4088) );
  NAND2_X1 U4634 ( .A1(n4905), .A2(n5302), .ZN(n4091) );
  NAND2_X1 U4635 ( .A1(n4999), .A2(n5304), .ZN(n4090) );
  NAND2_X1 U4636 ( .A1(n4091), .A2(n4090), .ZN(n4954) );
  NAND2_X1 U4637 ( .A1(n5364), .A2(n4962), .ZN(n4092) );
  NAND2_X1 U4638 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4765) );
  OAI211_X1 U4639 ( .C1(n5370), .C2(n4965), .A(n4092), .B(n4765), .ZN(n4093)
         );
  AOI21_X1 U4640 ( .B1(n5359), .B2(n4954), .A(n4093), .ZN(n4094) );
  OAI21_X1 U4641 ( .B1(n4095), .B2(n5315), .A(n4094), .ZN(U3216) );
  NAND2_X1 U4642 ( .A1(n4097), .A2(n4096), .ZN(n4102) );
  INV_X1 U4643 ( .A(n4098), .ZN(n4100) );
  NAND2_X1 U4644 ( .A1(n4100), .A2(n4099), .ZN(n4101) );
  NAND2_X1 U4645 ( .A1(n4102), .A2(n4101), .ZN(n4185) );
  NAND2_X1 U4646 ( .A1(n4905), .A2(n4235), .ZN(n4105) );
  OR2_X1 U4647 ( .A1(n4945), .A2(n2611), .ZN(n4104) );
  NAND2_X1 U4648 ( .A1(n4105), .A2(n4104), .ZN(n4106) );
  XNOR2_X1 U4649 ( .A(n4106), .B(n3296), .ZN(n4112) );
  INV_X1 U4650 ( .A(n4112), .ZN(n4110) );
  NAND2_X1 U4651 ( .A1(n4905), .A2(n4239), .ZN(n4108) );
  OR2_X1 U4652 ( .A1(n4273), .A2(n4945), .ZN(n4107) );
  NAND2_X1 U4653 ( .A1(n4108), .A2(n4107), .ZN(n4111) );
  INV_X1 U4654 ( .A(n4111), .ZN(n4109) );
  NAND2_X1 U4655 ( .A1(n4110), .A2(n4109), .ZN(n4186) );
  NAND2_X1 U4656 ( .A1(n4112), .A2(n4111), .ZN(n4184) );
  NAND2_X1 U4657 ( .A1(n4186), .A2(n4184), .ZN(n4113) );
  XNOR2_X1 U4658 ( .A(n4185), .B(n4113), .ZN(n4126) );
  INV_X1 U4659 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4114) );
  NAND2_X1 U4660 ( .A1(n4115), .A2(n4114), .ZN(n4116) );
  NAND2_X1 U4661 ( .A1(n4196), .A2(n4116), .ZN(n4916) );
  INV_X1 U4662 ( .A(REG0_REG_21__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U4663 ( .A1(n3212), .A2(REG2_REG_21__SCAN_IN), .ZN(n4118) );
  NAND2_X1 U4664 ( .A1(n2479), .A2(REG1_REG_21__SCAN_IN), .ZN(n4117) );
  OAI211_X1 U4665 ( .C1(n4285), .C2(n5078), .A(n4118), .B(n4117), .ZN(n4119)
         );
  INV_X1 U4666 ( .A(n4119), .ZN(n4120) );
  OAI22_X1 U4667 ( .A1(n4542), .A2(n4945), .B1(n4926), .B2(n5370), .ZN(n4124)
         );
  INV_X1 U4668 ( .A(n4558), .ZN(n4543) );
  INV_X1 U4669 ( .A(n4943), .ZN(n4371) );
  OAI22_X1 U4670 ( .A1(n4543), .A2(n4371), .B1(STATE_REG_SCAN_IN), .B2(n4122), 
        .ZN(n4123) );
  AOI211_X1 U4671 ( .C1(n4547), .C2(n4947), .A(n4124), .B(n4123), .ZN(n4125)
         );
  OAI21_X1 U4672 ( .B1(n4126), .B2(n5315), .A(n4125), .ZN(U3230) );
  INV_X1 U4673 ( .A(n4152), .ZN(n4147) );
  NAND2_X1 U4674 ( .A1(n4128), .A2(n5107), .ZN(n4129) );
  NOR2_X1 U4675 ( .A1(n4152), .A2(REG1_REG_13__SCAN_IN), .ZN(n4131) );
  INV_X1 U4676 ( .A(n4149), .ZN(n4137) );
  NAND2_X1 U4677 ( .A1(n4147), .A2(REG1_REG_13__SCAN_IN), .ZN(n4134) );
  OAI211_X1 U4678 ( .C1(REG1_REG_13__SCAN_IN), .C2(n4147), .A(n4135), .B(n4134), .ZN(n4136) );
  NAND3_X1 U4679 ( .A1(n4137), .A2(n4770), .A3(n4136), .ZN(n4146) );
  NOR2_X1 U4680 ( .A1(STATE_REG_SCAN_IN), .A2(n4138), .ZN(n5308) );
  INV_X1 U4681 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4140) );
  OR2_X1 U4682 ( .A1(n4152), .A2(n4140), .ZN(n4142) );
  NAND2_X1 U4683 ( .A1(n4152), .A2(n4140), .ZN(n4141) );
  AND2_X1 U4684 ( .A1(n4142), .A2(n4141), .ZN(n4155) );
  INV_X1 U4685 ( .A(n4153), .ZN(n4143) );
  AOI211_X1 U4686 ( .C1(n4154), .C2(n4155), .A(n4143), .B(n4773), .ZN(n4144)
         );
  AOI211_X1 U4687 ( .C1(n5143), .C2(ADDR_REG_13__SCAN_IN), .A(n5308), .B(n4144), .ZN(n4145) );
  OAI211_X1 U4688 ( .C1(n4768), .C2(n4147), .A(n4146), .B(n4145), .ZN(U3253)
         );
  XNOR2_X1 U4689 ( .A(n4169), .B(REG1_REG_14__SCAN_IN), .ZN(n4164) );
  INV_X1 U4690 ( .A(n5106), .ZN(n4166) );
  NOR2_X1 U4691 ( .A1(STATE_REG_SCAN_IN), .A2(n4150), .ZN(n4467) );
  AOI21_X1 U4692 ( .B1(n5143), .B2(ADDR_REG_14__SCAN_IN), .A(n4467), .ZN(n4151) );
  OAI21_X1 U4693 ( .B1(n4166), .B2(n4768), .A(n4151), .ZN(n4163) );
  NAND2_X1 U4694 ( .A1(n4152), .A2(REG2_REG_13__SCAN_IN), .ZN(n4157) );
  NAND2_X1 U4695 ( .A1(n4153), .A2(n4157), .ZN(n4176) );
  INV_X1 U4696 ( .A(n4154), .ZN(n4156) );
  NAND2_X1 U4697 ( .A1(n4156), .A2(n2667), .ZN(n4159) );
  OR2_X1 U4698 ( .A1(n4166), .A2(n4157), .ZN(n4158) );
  AOI211_X1 U4699 ( .C1(n3529), .C2(n4161), .A(n4178), .B(n4773), .ZN(n4162)
         );
  AOI211_X1 U4700 ( .C1(n4770), .C2(n4164), .A(n4163), .B(n4162), .ZN(n4165)
         );
  INV_X1 U4701 ( .A(n4165), .ZN(U3254) );
  INV_X1 U4702 ( .A(n4310), .ZN(n5357) );
  INV_X1 U4703 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4168) );
  INV_X1 U4704 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U4705 ( .A1(n4310), .A2(REG1_REG_15__SCAN_IN), .ZN(n4298) );
  INV_X1 U4706 ( .A(n4298), .ZN(n4170) );
  AOI21_X1 U4707 ( .B1(n5375), .B2(n5357), .A(n4170), .ZN(n4171) );
  OAI211_X1 U4708 ( .C1(n4172), .C2(n4171), .A(n4770), .B(n4299), .ZN(n4175)
         );
  AND2_X1 U4709 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4173) );
  AOI21_X1 U4710 ( .B1(n5143), .B2(ADDR_REG_15__SCAN_IN), .A(n4173), .ZN(n4174) );
  OAI211_X1 U4711 ( .C1(n4768), .C2(n5357), .A(n4175), .B(n4174), .ZN(n4183)
         );
  AND2_X1 U4712 ( .A1(n4176), .A2(n5106), .ZN(n4177) );
  NAND2_X1 U4713 ( .A1(n4310), .A2(REG2_REG_15__SCAN_IN), .ZN(n4179) );
  OAI21_X1 U4714 ( .B1(n4310), .B2(REG2_REG_15__SCAN_IN), .A(n4179), .ZN(n4180) );
  AOI211_X1 U4715 ( .C1(n4181), .C2(n4180), .A(n4311), .B(n4773), .ZN(n4182)
         );
  OR2_X1 U4716 ( .A1(n4183), .A2(n4182), .ZN(U3255) );
  NAND2_X1 U4717 ( .A1(n4185), .A2(n4184), .ZN(n4187) );
  NAND2_X1 U4718 ( .A1(n4947), .A2(n4235), .ZN(n4189) );
  OR2_X1 U4719 ( .A1(n4914), .A2(n2611), .ZN(n4188) );
  NAND2_X1 U4720 ( .A1(n4189), .A2(n4188), .ZN(n4190) );
  XNOR2_X1 U4721 ( .A(n4190), .B(n3093), .ZN(n4192) );
  NOR2_X1 U4722 ( .A1(n4914), .A2(n4273), .ZN(n4191) );
  AOI21_X1 U4723 ( .B1(n4947), .B2(n4239), .A(n4191), .ZN(n4193) );
  AND2_X1 U4724 ( .A1(n4192), .A2(n4193), .ZN(n4482) );
  INV_X1 U4725 ( .A(n4192), .ZN(n4195) );
  INV_X1 U4726 ( .A(n4193), .ZN(n4194) );
  NAND2_X1 U4727 ( .A1(n4195), .A2(n4194), .ZN(n4483) );
  NAND2_X1 U4728 ( .A1(n4196), .A2(n4541), .ZN(n4197) );
  NAND2_X1 U4729 ( .A1(n4210), .A2(n4197), .ZN(n4886) );
  INV_X1 U4730 ( .A(REG0_REG_22__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U4731 ( .A1(n3212), .A2(REG2_REG_22__SCAN_IN), .ZN(n4199) );
  NAND2_X1 U4732 ( .A1(n2479), .A2(REG1_REG_22__SCAN_IN), .ZN(n4198) );
  OAI211_X1 U4733 ( .C1(n5074), .C2(n4285), .A(n4199), .B(n4198), .ZN(n4200)
         );
  INV_X1 U4734 ( .A(n4200), .ZN(n4201) );
  NAND2_X1 U4735 ( .A1(n4903), .A2(n4235), .ZN(n4204) );
  OR2_X1 U4736 ( .A1(n4894), .A2(n2611), .ZN(n4203) );
  NAND2_X1 U4737 ( .A1(n4204), .A2(n4203), .ZN(n4205) );
  XNOR2_X1 U4738 ( .A(n4205), .B(n3093), .ZN(n4208) );
  NOR2_X1 U4739 ( .A1(n4894), .A2(n4273), .ZN(n4206) );
  AOI21_X1 U4740 ( .B1(n4903), .B2(n2986), .A(n4206), .ZN(n4207) );
  XNOR2_X1 U4741 ( .A(n4208), .B(n4207), .ZN(n4540) );
  NAND2_X1 U4742 ( .A1(n4208), .A2(n4207), .ZN(n4209) );
  NAND2_X1 U4743 ( .A1(n4210), .A2(n4476), .ZN(n4211) );
  AND2_X1 U4744 ( .A1(n4228), .A2(n4211), .ZN(n4875) );
  NAND2_X1 U4745 ( .A1(n4875), .A2(n4287), .ZN(n4216) );
  INV_X1 U4746 ( .A(REG0_REG_23__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U4747 ( .A1(n3212), .A2(REG2_REG_23__SCAN_IN), .ZN(n4213) );
  NAND2_X1 U4748 ( .A1(n2480), .A2(REG1_REG_23__SCAN_IN), .ZN(n4212) );
  OAI211_X1 U4749 ( .C1(n4285), .C2(n5070), .A(n4213), .B(n4212), .ZN(n4214)
         );
  INV_X1 U4750 ( .A(n4214), .ZN(n4215) );
  NAND2_X1 U4751 ( .A1(n4896), .A2(n4235), .ZN(n4218) );
  OR2_X1 U4752 ( .A1(n4868), .A2(n2611), .ZN(n4217) );
  NAND2_X1 U4753 ( .A1(n4218), .A2(n4217), .ZN(n4219) );
  XNOR2_X1 U4754 ( .A(n4219), .B(n3296), .ZN(n4222) );
  NAND2_X1 U4755 ( .A1(n4896), .A2(n4239), .ZN(n4221) );
  OR2_X1 U4756 ( .A1(n4273), .A2(n4868), .ZN(n4220) );
  NAND2_X1 U4757 ( .A1(n4221), .A2(n4220), .ZN(n4223) );
  NAND2_X1 U4758 ( .A1(n4222), .A2(n4223), .ZN(n4242) );
  INV_X1 U4759 ( .A(n4222), .ZN(n4225) );
  INV_X1 U4760 ( .A(n4223), .ZN(n4224) );
  NAND2_X1 U4761 ( .A1(n4225), .A2(n4224), .ZN(n4226) );
  NAND2_X1 U4762 ( .A1(n4242), .A2(n4226), .ZN(n4472) );
  NOR2_X2 U4763 ( .A1(n4473), .A2(n4472), .ZN(n4240) );
  NAND2_X1 U4764 ( .A1(n4228), .A2(n4227), .ZN(n4229) );
  NAND2_X1 U4765 ( .A1(n4254), .A2(n4229), .ZN(n4842) );
  INV_X1 U4766 ( .A(REG0_REG_24__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U4767 ( .A1(n3212), .A2(REG2_REG_24__SCAN_IN), .ZN(n4231) );
  NAND2_X1 U4768 ( .A1(n2480), .A2(REG1_REG_24__SCAN_IN), .ZN(n4230) );
  OAI211_X1 U4769 ( .C1(n5066), .C2(n4285), .A(n4231), .B(n4230), .ZN(n4232)
         );
  INV_X1 U4770 ( .A(n4232), .ZN(n4233) );
  NAND2_X1 U4771 ( .A1(n4870), .A2(n4235), .ZN(n4237) );
  OR2_X1 U4772 ( .A1(n4851), .A2(n2611), .ZN(n4236) );
  NAND2_X1 U4773 ( .A1(n4237), .A2(n4236), .ZN(n4238) );
  XNOR2_X1 U4774 ( .A(n4238), .B(n3093), .ZN(n4241) );
  INV_X1 U4775 ( .A(n4851), .ZN(n4532) );
  AOI22_X1 U4776 ( .A1(n4870), .A2(n4239), .B1(n3090), .B2(n4532), .ZN(n4528)
         );
  XNOR2_X1 U4777 ( .A(n4254), .B(REG3_REG_25__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U4778 ( .A1(n4510), .A2(n4287), .ZN(n4247) );
  INV_X1 U4779 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4385) );
  NAND2_X1 U4780 ( .A1(n3212), .A2(REG2_REG_25__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U4781 ( .A1(n2479), .A2(REG1_REG_25__SCAN_IN), .ZN(n4243) );
  OAI211_X1 U4782 ( .C1(n4385), .C2(n4285), .A(n4244), .B(n4243), .ZN(n4245)
         );
  INV_X1 U4783 ( .A(n4245), .ZN(n4246) );
  INV_X1 U4784 ( .A(n4239), .ZN(n4289) );
  OAI22_X1 U4785 ( .A1(n4821), .A2(n4289), .B1(n4273), .B2(n4362), .ZN(n4249)
         );
  OAI22_X1 U4786 ( .A1(n4821), .A2(n4273), .B1(n2611), .B2(n4362), .ZN(n4248)
         );
  XNOR2_X1 U4787 ( .A(n4248), .B(n3296), .ZN(n4250) );
  XOR2_X1 U4788 ( .A(n4249), .B(n4250), .Z(n4504) );
  NAND2_X1 U4789 ( .A1(n4503), .A2(n4251), .ZN(n4553) );
  OAI21_X1 U4790 ( .B1(n4254), .B2(n4253), .A(n4252), .ZN(n4255) );
  NAND2_X1 U4791 ( .A1(n4255), .A2(n4265), .ZN(n4833) );
  INV_X1 U4792 ( .A(REG0_REG_26__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U4793 ( .A1(n2479), .A2(REG1_REG_26__SCAN_IN), .ZN(n4257) );
  NAND2_X1 U4794 ( .A1(n3212), .A2(REG2_REG_26__SCAN_IN), .ZN(n4256) );
  OAI211_X1 U4795 ( .C1(n5062), .C2(n4285), .A(n4257), .B(n4256), .ZN(n4258)
         );
  INV_X1 U4796 ( .A(n4258), .ZN(n4259) );
  OAI22_X1 U4797 ( .A1(n4809), .A2(n4273), .B1(n2611), .B2(n4824), .ZN(n4261)
         );
  XOR2_X1 U4798 ( .A(n3296), .B(n4261), .Z(n4551) );
  INV_X1 U4799 ( .A(n4551), .ZN(n4262) );
  OAI22_X1 U4800 ( .A1(n4809), .A2(n4289), .B1(n4824), .B2(n4273), .ZN(n4263)
         );
  INV_X1 U4801 ( .A(n4263), .ZN(n4550) );
  NAND2_X1 U4802 ( .A1(n4265), .A2(n4264), .ZN(n4266) );
  NAND2_X1 U4803 ( .A1(n4280), .A2(n4266), .ZN(n4801) );
  INV_X1 U4804 ( .A(REG0_REG_27__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U4805 ( .A1(n3212), .A2(REG2_REG_27__SCAN_IN), .ZN(n4269) );
  NAND2_X1 U4806 ( .A1(n2480), .A2(REG1_REG_27__SCAN_IN), .ZN(n4268) );
  OAI211_X1 U4807 ( .C1(n5057), .C2(n4285), .A(n4269), .B(n4268), .ZN(n4270)
         );
  INV_X1 U4808 ( .A(n4270), .ZN(n4271) );
  INV_X1 U4809 ( .A(n4820), .ZN(n4786) );
  OAI22_X1 U4810 ( .A1(n4786), .A2(n4289), .B1(n4273), .B2(n4808), .ZN(n4277)
         );
  NAND2_X1 U4811 ( .A1(n4820), .A2(n3090), .ZN(n4275) );
  OR2_X1 U4812 ( .A1(n4808), .A2(n2611), .ZN(n4274) );
  NAND2_X1 U4813 ( .A1(n4275), .A2(n4274), .ZN(n4276) );
  XNOR2_X1 U4814 ( .A(n4276), .B(n3296), .ZN(n4278) );
  XOR2_X1 U4815 ( .A(n4277), .B(n4278), .Z(n4454) );
  NAND2_X1 U4816 ( .A1(n4280), .A2(n4279), .ZN(n4281) );
  INV_X1 U4817 ( .A(REG0_REG_28__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U4818 ( .A1(n3212), .A2(REG2_REG_28__SCAN_IN), .ZN(n4284) );
  NAND2_X1 U4819 ( .A1(n2479), .A2(REG1_REG_28__SCAN_IN), .ZN(n4283) );
  OAI211_X1 U4820 ( .C1(n5053), .C2(n4285), .A(n4284), .B(n4283), .ZN(n4286)
         );
  OAI22_X1 U4821 ( .A1(n4719), .A2(n4273), .B1(n2611), .B2(n4781), .ZN(n4288)
         );
  XNOR2_X1 U4822 ( .A(n4288), .B(n3296), .ZN(n4291) );
  OAI22_X1 U4823 ( .A1(n4719), .A2(n4289), .B1(n4273), .B2(n4781), .ZN(n4290)
         );
  XNOR2_X1 U4824 ( .A(n4291), .B(n4290), .ZN(n4292) );
  INV_X1 U4825 ( .A(n4790), .ZN(n4294) );
  INV_X1 U4826 ( .A(n4781), .ZN(n4789) );
  AOI22_X1 U4827 ( .A1(n5364), .A2(n4789), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n4293) );
  OAI21_X1 U4828 ( .B1(n4294), .B2(n5370), .A(n4293), .ZN(n4296) );
  NOR2_X1 U4829 ( .A1(n4782), .A2(n4555), .ZN(n4295) );
  AOI211_X1 U4830 ( .C1(n4558), .C2(n4820), .A(n4296), .B(n4295), .ZN(n4297)
         );
  NOR2_X1 U4831 ( .A1(n4312), .A2(n4300), .ZN(n4301) );
  INV_X1 U4832 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4302) );
  OR2_X1 U4833 ( .A1(n5105), .A2(n4302), .ZN(n4304) );
  NAND2_X1 U4834 ( .A1(n5105), .A2(n4302), .ZN(n4303) );
  AND2_X1 U4835 ( .A1(n4304), .A2(n4303), .ZN(n4747) );
  NOR2_X2 U4836 ( .A1(n4746), .A2(n4747), .ZN(n4305) );
  NOR2_X1 U4837 ( .A1(n5105), .A2(REG1_REG_17__SCAN_IN), .ZN(n4307) );
  XNOR2_X1 U4838 ( .A(n5104), .B(REG1_REG_18__SCAN_IN), .ZN(n4306) );
  NOR3_X2 U4839 ( .A1(n4305), .A2(n4307), .A3(n4306), .ZN(n4762) );
  INV_X1 U4840 ( .A(n4762), .ZN(n4309) );
  OAI21_X1 U4841 ( .B1(n4305), .B2(n4307), .A(n4306), .ZN(n4308) );
  NAND3_X1 U4842 ( .A1(n4309), .A2(n4770), .A3(n4308), .ZN(n4328) );
  INV_X1 U4843 ( .A(n4312), .ZN(n5379) );
  INV_X1 U4844 ( .A(n4313), .ZN(n4314) );
  NAND2_X1 U4845 ( .A1(n4314), .A2(n5379), .ZN(n4315) );
  NAND2_X1 U4846 ( .A1(n4738), .A2(n4315), .ZN(n4749) );
  NAND2_X1 U4847 ( .A1(n5105), .A2(REG2_REG_17__SCAN_IN), .ZN(n4316) );
  OAI21_X1 U4848 ( .B1(n5105), .B2(REG2_REG_17__SCAN_IN), .A(n4316), .ZN(n4750) );
  INV_X1 U4849 ( .A(n4316), .ZN(n4317) );
  INV_X1 U4850 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4319) );
  NOR2_X1 U4851 ( .A1(n5104), .A2(n4319), .ZN(n4318) );
  AOI21_X1 U4852 ( .B1(n5104), .B2(n4319), .A(n4318), .ZN(n4320) );
  INV_X1 U4853 ( .A(n4758), .ZN(n4325) );
  NAND2_X1 U4854 ( .A1(n5143), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4323) );
  OAI211_X1 U4855 ( .C1(n4768), .C2(n2516), .A(n4328), .B(n4327), .ZN(U3258)
         );
  OR2_X1 U4856 ( .A1(n4330), .A2(n4329), .ZN(n4332) );
  NAND2_X1 U4857 ( .A1(n4332), .A2(n4331), .ZN(n4333) );
  XOR2_X1 U4858 ( .A(n4610), .B(n4333), .Z(n5227) );
  INV_X1 U4859 ( .A(n4334), .ZN(n4335) );
  AOI21_X1 U4860 ( .B1(n4342), .B2(n4336), .A(n4335), .ZN(n5231) );
  INV_X1 U4861 ( .A(n4337), .ZN(n4338) );
  OAI22_X1 U4862 ( .A1(n5341), .A2(n2831), .B1(n4338), .B2(n5339), .ZN(n4339)
         );
  AOI21_X1 U4863 ( .B1(n5231), .B2(n5415), .A(n4339), .ZN(n4346) );
  XOR2_X1 U4864 ( .A(n4610), .B(n4340), .Z(n4344) );
  AOI21_X1 U4865 ( .B1(n4342), .B2(n5396), .A(n4341), .ZN(n4343) );
  OAI21_X1 U4866 ( .B1(n4344), .B2(n5190), .A(n4343), .ZN(n5230) );
  NAND2_X1 U4867 ( .A1(n5230), .A2(n5262), .ZN(n4345) );
  OAI211_X1 U4868 ( .C1(n5227), .C2(n4991), .A(n4346), .B(n4345), .ZN(U3284)
         );
  INV_X1 U4869 ( .A(n4947), .ZN(n4544) );
  INV_X1 U4870 ( .A(n4914), .ZN(n4904) );
  INV_X1 U4871 ( .A(n4905), .ZN(n4372) );
  NAND2_X1 U4872 ( .A1(n4348), .A2(n4347), .ZN(n4352) );
  NAND2_X1 U4873 ( .A1(n4352), .A2(n4351), .ZN(n4995) );
  AND2_X1 U4874 ( .A1(n4721), .A2(n4369), .ZN(n4621) );
  INV_X1 U4875 ( .A(n4721), .ZN(n4370) );
  NAND2_X1 U4876 ( .A1(n4370), .A2(n5001), .ZN(n4622) );
  OAI21_X2 U4877 ( .B1(n4995), .B2(n4621), .A(n4622), .ZN(n4970) );
  INV_X1 U4878 ( .A(n4999), .ZN(n4354) );
  NAND2_X1 U4879 ( .A1(n4354), .A2(n4984), .ZN(n4934) );
  INV_X1 U4880 ( .A(n4984), .ZN(n4353) );
  NAND2_X1 U4881 ( .A1(n4353), .A2(n4999), .ZN(n4977) );
  NAND2_X1 U4882 ( .A1(n4934), .A2(n4977), .ZN(n4978) );
  INV_X1 U4883 ( .A(n4962), .ZN(n4956) );
  OAI21_X1 U4884 ( .B1(n4904), .B2(n4947), .A(n4911), .ZN(n4357) );
  OAI21_X1 U4885 ( .B1(n4544), .B2(n4914), .A(n4357), .ZN(n4881) );
  NAND2_X1 U4886 ( .A1(n4903), .A2(n4894), .ZN(n4375) );
  NAND2_X1 U4887 ( .A1(n4863), .A2(n4375), .ZN(n4888) );
  NAND2_X1 U4888 ( .A1(n4896), .A2(n4874), .ZN(n4358) );
  INV_X1 U4889 ( .A(n4896), .ZN(n4379) );
  NAND2_X1 U4890 ( .A1(n4508), .A2(n4851), .ZN(n4359) );
  NAND2_X1 U4891 ( .A1(n4870), .A2(n4532), .ZN(n4360) );
  INV_X1 U4892 ( .A(n4362), .ZN(n4506) );
  OR2_X1 U4893 ( .A1(n4821), .A2(n4506), .ZN(n4693) );
  NAND2_X1 U4894 ( .A1(n4821), .A2(n4506), .ZN(n4816) );
  NAND2_X1 U4895 ( .A1(n4693), .A2(n4816), .ZN(n4640) );
  XNOR2_X1 U4896 ( .A(n4421), .B(n4640), .ZN(n4396) );
  NAND2_X1 U4897 ( .A1(n5154), .A2(n4361), .ZN(n5228) );
  NAND2_X1 U4898 ( .A1(n3273), .A2(n5228), .ZN(n5392) );
  NAND2_X1 U4899 ( .A1(n5414), .A2(n5392), .ZN(n5092) );
  OR2_X1 U4900 ( .A1(n4839), .A2(n4362), .ZN(n4363) );
  NAND2_X1 U4901 ( .A1(n2505), .A2(n4363), .ZN(n4392) );
  NAND2_X1 U4902 ( .A1(n4365), .A2(n4364), .ZN(n4930) );
  NAND2_X1 U4903 ( .A1(n4956), .A2(n4943), .ZN(n4366) );
  NAND2_X1 U4904 ( .A1(n4977), .A2(n4366), .ZN(n4935) );
  NAND2_X1 U4905 ( .A1(n5001), .A2(n4721), .ZN(n4932) );
  NAND2_X1 U4906 ( .A1(n4929), .A2(n4932), .ZN(n4367) );
  NOR2_X1 U4907 ( .A1(n4935), .A2(n4367), .ZN(n4368) );
  NAND2_X1 U4908 ( .A1(n4905), .A2(n4945), .ZN(n4602) );
  NAND2_X1 U4909 ( .A1(n4370), .A2(n4369), .ZN(n4931) );
  AND2_X1 U4910 ( .A1(n4934), .A2(n4931), .ZN(n4373) );
  NAND2_X1 U4911 ( .A1(n4371), .A2(n4962), .ZN(n4937) );
  NAND2_X1 U4912 ( .A1(n4372), .A2(n4922), .ZN(n4603) );
  OAI211_X1 U4913 ( .C1(n4373), .C2(n4935), .A(n4937), .B(n4603), .ZN(n4374)
         );
  NAND2_X1 U4914 ( .A1(n4374), .A2(n4602), .ZN(n4562) );
  OR2_X1 U4915 ( .A1(n4947), .A2(n4914), .ZN(n4859) );
  NAND2_X1 U4916 ( .A1(n4863), .A2(n4859), .ZN(n4561) );
  NAND2_X1 U4917 ( .A1(n4896), .A2(n4868), .ZN(n4377) );
  AND2_X1 U4918 ( .A1(n4947), .A2(n4914), .ZN(n4616) );
  NAND2_X1 U4919 ( .A1(n4863), .A2(n4616), .ZN(n4376) );
  NAND3_X1 U4920 ( .A1(n4377), .A2(n4376), .A3(n4375), .ZN(n4695) );
  INV_X1 U4921 ( .A(n4695), .ZN(n4378) );
  NAND2_X1 U4922 ( .A1(n4508), .A2(n4532), .ZN(n4601) );
  NAND2_X1 U4923 ( .A1(n4379), .A2(n4874), .ZN(n4844) );
  NAND2_X1 U4924 ( .A1(n4601), .A2(n4844), .ZN(n4575) );
  INV_X1 U4925 ( .A(n4575), .ZN(n4696) );
  NAND2_X1 U4926 ( .A1(n4845), .A2(n4696), .ZN(n4380) );
  NAND2_X1 U4927 ( .A1(n4870), .A2(n4851), .ZN(n4692) );
  NAND2_X1 U4928 ( .A1(n4380), .A2(n4692), .ZN(n4428) );
  XNOR2_X1 U4929 ( .A(n4428), .B(n4640), .ZN(n4383) );
  AOI22_X1 U4930 ( .A1(n4870), .A2(n5304), .B1(n4506), .B2(n5396), .ZN(n4381)
         );
  OAI21_X1 U4931 ( .B1(n4809), .B2(n5184), .A(n4381), .ZN(n4382) );
  AOI21_X1 U4932 ( .B1(n4383), .B2(n5333), .A(n4382), .ZN(n4390) );
  OAI21_X1 U4933 ( .B1(n5390), .B2(n4392), .A(n4390), .ZN(n4387) );
  INV_X1 U4934 ( .A(n4387), .ZN(n4384) );
  MUX2_X1 U4935 ( .A(n4385), .B(n4384), .S(n5414), .Z(n4386) );
  OAI21_X1 U4936 ( .B1(n4396), .B2(n5092), .A(n4386), .ZN(U3511) );
  NAND2_X1 U4937 ( .A1(n5410), .A2(n5392), .ZN(n5051) );
  MUX2_X1 U4938 ( .A(REG1_REG_25__SCAN_IN), .B(n4387), .S(n5410), .Z(n4388) );
  INV_X1 U4939 ( .A(n4388), .ZN(n4389) );
  OAI21_X1 U4940 ( .B1(n4396), .B2(n5051), .A(n4389), .ZN(U3543) );
  INV_X1 U4941 ( .A(n4390), .ZN(n4394) );
  AOI22_X1 U4942 ( .A1(n4510), .A2(n5204), .B1(REG2_REG_25__SCAN_IN), .B2(
        n5419), .ZN(n4391) );
  OAI21_X1 U4943 ( .B1(n4392), .B2(n5010), .A(n4391), .ZN(n4393) );
  AOI21_X1 U4944 ( .B1(n4394), .B2(n5262), .A(n4393), .ZN(n4395) );
  OAI21_X1 U4945 ( .B1(n4396), .B2(n4991), .A(n4395), .ZN(U3265) );
  NOR2_X1 U4946 ( .A1(n4397), .A2(n4404), .ZN(n4398) );
  OR2_X1 U4947 ( .A1(n4399), .A2(n4398), .ZN(n5283) );
  XNOR2_X1 U4948 ( .A(n5272), .B(n4400), .ZN(n5282) );
  INV_X1 U4949 ( .A(n5282), .ZN(n4403) );
  OAI22_X1 U4950 ( .A1(n5341), .A2(n3432), .B1(n4401), .B2(n5339), .ZN(n4402)
         );
  AOI21_X1 U4951 ( .B1(n4403), .B2(n5415), .A(n4402), .ZN(n4411) );
  INV_X1 U4952 ( .A(n4404), .ZN(n4629) );
  XNOR2_X1 U4953 ( .A(n4405), .B(n4629), .ZN(n4406) );
  NAND2_X1 U4954 ( .A1(n4406), .A2(n5333), .ZN(n4408) );
  AOI22_X1 U4955 ( .A1(n5304), .A2(n4726), .B1(n4724), .B2(n5302), .ZN(n4407)
         );
  OAI211_X1 U4956 ( .C1(n5330), .C2(n4409), .A(n4408), .B(n4407), .ZN(n5284)
         );
  NAND2_X1 U4957 ( .A1(n5284), .A2(n5262), .ZN(n4410) );
  OAI211_X1 U4958 ( .C1(n5283), .C2(n4991), .A(n4411), .B(n4410), .ZN(U3280)
         );
  INV_X1 U4959 ( .A(DATAI_20_), .ZN(n4412) );
  OAI22_X1 U4960 ( .A1(n2864), .A2(U3149), .B1(STATE_REG_SCAN_IN), .B2(n4412), 
        .ZN(U3332) );
  OAI211_X1 U4961 ( .C1(n4415), .C2(n4413), .A(n4414), .B(n5366), .ZN(n4419)
         );
  AOI22_X1 U4962 ( .A1(n4417), .A2(n5359), .B1(REG3_REG_1__SCAN_IN), .B2(n4416), .ZN(n4418) );
  OAI211_X1 U4963 ( .C1(n4542), .C2(n4420), .A(n4419), .B(n4418), .ZN(U3219)
         );
  NAND2_X1 U4964 ( .A1(n4720), .A2(n4830), .ZN(n4423) );
  NOR2_X1 U4965 ( .A1(n4720), .A2(n4830), .ZN(n4422) );
  OAI21_X1 U4966 ( .B1(n4796), .B2(n4820), .A(n4795), .ZN(n4425) );
  NAND2_X1 U4967 ( .A1(n4820), .A2(n4796), .ZN(n4424) );
  NAND2_X1 U4968 ( .A1(n4425), .A2(n4424), .ZN(n4776) );
  NOR2_X1 U4969 ( .A1(n4719), .A2(n4789), .ZN(n4584) );
  NOR2_X1 U4970 ( .A1(n4719), .A2(n4781), .ZN(n4426) );
  AOI21_X1 U4971 ( .B1(n4776), .B2(n4775), .A(n4426), .ZN(n4427) );
  OR2_X1 U4972 ( .A1(n4782), .A2(n4435), .ZN(n4583) );
  NAND2_X1 U4973 ( .A1(n4782), .A2(n4435), .ZN(n4578) );
  AND2_X1 U4974 ( .A1(n4583), .A2(n4578), .ZN(n4638) );
  XNOR2_X1 U4975 ( .A(n4427), .B(n4638), .ZN(n4452) );
  INV_X1 U4976 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4440) );
  NAND2_X1 U4977 ( .A1(n4809), .A2(n4830), .ZN(n4599) );
  NAND2_X1 U4978 ( .A1(n4599), .A2(n4816), .ZN(n4701) );
  INV_X1 U4979 ( .A(n4701), .ZN(n4581) );
  NAND2_X1 U4980 ( .A1(n4720), .A2(n4824), .ZN(n4600) );
  NOR2_X1 U4981 ( .A1(n4820), .A2(n4808), .ZN(n4587) );
  NAND2_X1 U4982 ( .A1(n4820), .A2(n4808), .ZN(n4699) );
  INV_X1 U4983 ( .A(n4699), .ZN(n4429) );
  INV_X1 U4984 ( .A(n4587), .ZN(n4430) );
  NAND2_X1 U4985 ( .A1(n4806), .A2(n4430), .ZN(n4778) );
  INV_X1 U4986 ( .A(n4775), .ZN(n4779) );
  INV_X1 U4987 ( .A(n4589), .ZN(n4431) );
  NAND2_X1 U4988 ( .A1(n2480), .A2(REG1_REG_30__SCAN_IN), .ZN(n4434) );
  NAND2_X1 U4989 ( .A1(n3212), .A2(REG2_REG_30__SCAN_IN), .ZN(n4433) );
  NAND2_X1 U4990 ( .A1(n3106), .A2(REG0_REG_30__SCAN_IN), .ZN(n4432) );
  NAND3_X1 U4991 ( .A1(n4434), .A2(n4433), .A3(n4432), .ZN(n4718) );
  AOI22_X1 U4992 ( .A1(n4718), .A2(n4436), .B1(n5396), .B2(n4435), .ZN(n4437)
         );
  OAI21_X1 U4993 ( .B1(n4719), .B2(n5186), .A(n4437), .ZN(n4438) );
  OAI211_X1 U4994 ( .C1(n4787), .C2(n4439), .A(n5406), .B(n5401), .ZN(n4445)
         );
  AND2_X1 U4995 ( .A1(n4442), .A2(n4445), .ZN(n4449) );
  MUX2_X1 U4996 ( .A(n4440), .B(n4449), .S(n5410), .Z(n4441) );
  INV_X1 U4997 ( .A(n4442), .ZN(n4447) );
  AOI22_X1 U4998 ( .A1(n4443), .A2(n5204), .B1(REG2_REG_29__SCAN_IN), .B2(
        n5419), .ZN(n4444) );
  OAI21_X1 U4999 ( .B1(n4445), .B2(n4877), .A(n4444), .ZN(n4446) );
  AOI21_X1 U5000 ( .B1(n4447), .B2(n5262), .A(n4446), .ZN(n4448) );
  OAI21_X1 U5001 ( .B1(n4452), .B2(n4991), .A(n4448), .ZN(U3354) );
  MUX2_X1 U5002 ( .A(n4450), .B(n4449), .S(n5414), .Z(n4451) );
  XNOR2_X1 U5003 ( .A(n4453), .B(n4454), .ZN(n4459) );
  AOI22_X1 U5004 ( .A1(n5364), .A2(n4796), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n4455) );
  OAI21_X1 U5005 ( .B1(n4801), .B2(n5370), .A(n4455), .ZN(n4457) );
  NOR2_X1 U5006 ( .A1(n4719), .A2(n4555), .ZN(n4456) );
  AOI211_X1 U5007 ( .C1(n4558), .C2(n4720), .A(n4457), .B(n4456), .ZN(n4458)
         );
  OAI21_X1 U5008 ( .B1(n4459), .B2(n5315), .A(n4458), .ZN(U3211) );
  OAI21_X1 U5009 ( .B1(n4462), .B2(n4461), .A(n4460), .ZN(n4463) );
  NAND2_X1 U5010 ( .A1(n4463), .A2(n5366), .ZN(n4471) );
  AOI22_X1 U5011 ( .A1(n4547), .A2(n4722), .B1(n4464), .B2(n5364), .ZN(n4470)
         );
  NOR2_X1 U5012 ( .A1(n4543), .A2(n4465), .ZN(n4466) );
  AOI211_X1 U5013 ( .C1(n4522), .C2(n4468), .A(n4467), .B(n4466), .ZN(n4469)
         );
  NAND3_X1 U5014 ( .A1(n4471), .A2(n4470), .A3(n4469), .ZN(U3212) );
  AOI21_X1 U5015 ( .B1(n4473), .B2(n4472), .A(n5315), .ZN(n4475) );
  NAND2_X1 U5016 ( .A1(n4475), .A2(n4474), .ZN(n4481) );
  OAI22_X1 U5017 ( .A1(n4542), .A2(n4868), .B1(STATE_REG_SCAN_IN), .B2(n4476), 
        .ZN(n4479) );
  INV_X1 U5018 ( .A(n4903), .ZN(n4477) );
  NOR2_X1 U5019 ( .A1(n4477), .A2(n4543), .ZN(n4478) );
  AOI211_X1 U5020 ( .C1(n4522), .C2(n4875), .A(n4479), .B(n4478), .ZN(n4480)
         );
  OAI211_X1 U5021 ( .C1(n4508), .C2(n4555), .A(n4481), .B(n4480), .ZN(U3213)
         );
  INV_X1 U5022 ( .A(n4482), .ZN(n4484) );
  NAND2_X1 U5023 ( .A1(n4484), .A2(n4483), .ZN(n4485) );
  XNOR2_X1 U5024 ( .A(n4486), .B(n4485), .ZN(n4491) );
  AOI22_X1 U5025 ( .A1(n4558), .A2(n4905), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n4488) );
  NAND2_X1 U5026 ( .A1(n5364), .A2(n4904), .ZN(n4487) );
  OAI211_X1 U5027 ( .C1(n5370), .C2(n4916), .A(n4488), .B(n4487), .ZN(n4489)
         );
  AOI21_X1 U5028 ( .B1(n4547), .B2(n4903), .A(n4489), .ZN(n4490) );
  OAI21_X1 U5029 ( .B1(n4491), .B2(n5315), .A(n4490), .ZN(U3220) );
  OAI21_X1 U5030 ( .B1(n4493), .B2(n4492), .A(n5314), .ZN(n4494) );
  NAND2_X1 U5031 ( .A1(n4494), .A2(n5366), .ZN(n4502) );
  AOI22_X1 U5032 ( .A1(n4547), .A2(n4723), .B1(n4495), .B2(n5364), .ZN(n4501)
         );
  NOR2_X1 U5033 ( .A1(n4543), .A2(n4496), .ZN(n4497) );
  AOI211_X1 U5034 ( .C1(n4522), .C2(n4499), .A(n4498), .B(n4497), .ZN(n4500)
         );
  NAND3_X1 U5035 ( .A1(n4502), .A2(n4501), .A3(n4500), .ZN(U3221) );
  OAI21_X1 U5036 ( .B1(n4504), .B2(n4526), .A(n4503), .ZN(n4505) );
  NAND2_X1 U5037 ( .A1(n4505), .A2(n5366), .ZN(n4512) );
  AOI22_X1 U5038 ( .A1(n5364), .A2(n4506), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n4507) );
  OAI21_X1 U5039 ( .B1(n4508), .B2(n4543), .A(n4507), .ZN(n4509) );
  AOI21_X1 U5040 ( .B1(n4510), .B2(n4522), .A(n4509), .ZN(n4511) );
  OAI211_X1 U5041 ( .C1(n4809), .C2(n4555), .A(n4512), .B(n4511), .ZN(U3222)
         );
  INV_X1 U5042 ( .A(n4513), .ZN(n4517) );
  AOI21_X1 U5043 ( .B1(n4515), .B2(n5361), .A(n4514), .ZN(n4516) );
  OAI21_X1 U5044 ( .B1(n4517), .B2(n4516), .A(n5366), .ZN(n4525) );
  AOI22_X1 U5045 ( .A1(n4547), .A2(n4721), .B1(n4518), .B2(n5364), .ZN(n4524)
         );
  NOR2_X1 U5046 ( .A1(STATE_REG_SCAN_IN), .A2(n4519), .ZN(n4742) );
  NOR2_X1 U5047 ( .A1(n4543), .A2(n4565), .ZN(n4520) );
  AOI211_X1 U5048 ( .C1(n4522), .C2(n4521), .A(n4742), .B(n4520), .ZN(n4523)
         );
  NAND3_X1 U5049 ( .A1(n4525), .A2(n4524), .A3(n4523), .ZN(U3223) );
  INV_X1 U5050 ( .A(n2484), .ZN(n4527) );
  NOR2_X1 U5051 ( .A1(n4527), .A2(n2501), .ZN(n4529) );
  OAI22_X1 U5052 ( .A1(n2630), .A2(n4530), .B1(n4529), .B2(n4528), .ZN(n4531)
         );
  NAND2_X1 U5053 ( .A1(n4531), .A2(n5366), .ZN(n4536) );
  AOI22_X1 U5054 ( .A1(n5364), .A2(n4532), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n4533) );
  OAI21_X1 U5055 ( .B1(n4842), .B2(n5370), .A(n4533), .ZN(n4534) );
  AOI21_X1 U5056 ( .B1(n4558), .B2(n4896), .A(n4534), .ZN(n4535) );
  OAI211_X1 U5057 ( .C1(n4821), .C2(n4555), .A(n4536), .B(n4535), .ZN(U3226)
         );
  INV_X1 U5058 ( .A(n4537), .ZN(n4538) );
  AOI21_X1 U5059 ( .B1(n4540), .B2(n4539), .A(n4538), .ZN(n4549) );
  OAI22_X1 U5060 ( .A1(n4542), .A2(n4894), .B1(STATE_REG_SCAN_IN), .B2(n4541), 
        .ZN(n4546) );
  OAI22_X1 U5061 ( .A1(n4544), .A2(n4543), .B1(n4886), .B2(n5370), .ZN(n4545)
         );
  AOI211_X1 U5062 ( .C1(n4547), .C2(n4896), .A(n4546), .B(n4545), .ZN(n4548)
         );
  OAI21_X1 U5063 ( .B1(n4549), .B2(n5315), .A(n4548), .ZN(U3232) );
  XNOR2_X1 U5064 ( .A(n4551), .B(n4550), .ZN(n4552) );
  XNOR2_X1 U5065 ( .A(n4553), .B(n4552), .ZN(n4560) );
  AOI22_X1 U5066 ( .A1(n5364), .A2(n4830), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4554) );
  OAI21_X1 U5067 ( .B1(n4833), .B2(n5370), .A(n4554), .ZN(n4557) );
  NOR2_X1 U5068 ( .A1(n4786), .A2(n4555), .ZN(n4556) );
  AOI211_X1 U5069 ( .C1(n4558), .C2(n4853), .A(n4557), .B(n4556), .ZN(n4559)
         );
  OAI21_X1 U5070 ( .B1(n4560), .B2(n5315), .A(n4559), .ZN(U3237) );
  INV_X1 U5071 ( .A(n4561), .ZN(n4563) );
  NAND2_X1 U5072 ( .A1(n4563), .A2(n4562), .ZN(n4688) );
  INV_X1 U5073 ( .A(n4688), .ZN(n4574) );
  INV_X1 U5074 ( .A(n4564), .ZN(n4571) );
  AND2_X1 U5075 ( .A1(n4565), .A2(n5365), .ZN(n4570) );
  INV_X1 U5076 ( .A(n4570), .ZN(n4567) );
  AND2_X1 U5077 ( .A1(n4567), .A2(n4566), .ZN(n4652) );
  AND2_X1 U5078 ( .A1(n4569), .A2(n4568), .ZN(n4656) );
  NOR2_X1 U5079 ( .A1(n4656), .A2(n4570), .ZN(n4687) );
  AOI21_X1 U5080 ( .B1(n4571), .B2(n4652), .A(n4687), .ZN(n4572) );
  OAI21_X1 U5081 ( .B1(n4572), .B2(n4691), .A(n4690), .ZN(n4573) );
  AOI21_X1 U5082 ( .B1(n4574), .B2(n4573), .A(n4695), .ZN(n4576) );
  OAI211_X1 U5083 ( .C1(n4576), .C2(n4575), .A(n4693), .B(n4692), .ZN(n4582)
         );
  INV_X1 U5084 ( .A(n5397), .ZN(n5400) );
  INV_X1 U5085 ( .A(n4597), .ZN(n4577) );
  NAND2_X1 U5086 ( .A1(n4717), .A2(n4577), .ZN(n4703) );
  OAI21_X1 U5087 ( .B1(n4718), .B2(n5400), .A(n4703), .ZN(n4618) );
  INV_X1 U5088 ( .A(n4618), .ZN(n4579) );
  NAND2_X1 U5089 ( .A1(n4579), .A2(n4578), .ZN(n4586) );
  NOR3_X1 U5090 ( .A1(n4589), .A2(n4587), .A3(n4586), .ZN(n4580) );
  NAND3_X1 U5091 ( .A1(n4582), .A2(n4581), .A3(n4580), .ZN(n4591) );
  INV_X1 U5092 ( .A(n4583), .ZN(n4585) );
  NOR2_X1 U5093 ( .A1(n4585), .A2(n4584), .ZN(n4588) );
  NAND2_X1 U5094 ( .A1(n4600), .A2(n4588), .ZN(n4698) );
  AOI221_X1 U5095 ( .B1(n4589), .B2(n4588), .C1(n4587), .C2(n4588), .A(n4586), 
        .ZN(n4705) );
  OAI21_X1 U5096 ( .B1(n4803), .B2(n4698), .A(n4705), .ZN(n4590) );
  AOI22_X1 U5097 ( .A1(n4591), .A2(n4590), .B1(n4594), .B2(n5397), .ZN(n4593)
         );
  OR2_X1 U5098 ( .A1(n4593), .A2(n4592), .ZN(n4598) );
  INV_X1 U5099 ( .A(n2864), .ZN(n4708) );
  NAND2_X1 U5100 ( .A1(n4594), .A2(n4597), .ZN(n4596) );
  NAND2_X1 U5101 ( .A1(n4718), .A2(n5400), .ZN(n4595) );
  NAND2_X1 U5102 ( .A1(n4596), .A2(n4595), .ZN(n4704) );
  AOI22_X1 U5103 ( .A1(n4598), .A2(n4708), .B1(n4597), .B2(n4704), .ZN(n4710)
         );
  INV_X1 U5104 ( .A(n4803), .ZN(n4639) );
  NAND2_X1 U5105 ( .A1(n4600), .A2(n4599), .ZN(n4828) );
  INV_X1 U5106 ( .A(n4828), .ZN(n4818) );
  NAND2_X1 U5107 ( .A1(n4601), .A2(n4692), .ZN(n4846) );
  NAND2_X1 U5108 ( .A1(n4603), .A2(n4602), .ZN(n4939) );
  XNOR2_X1 U5109 ( .A(n5331), .B(n4723), .ZN(n5327) );
  NAND2_X1 U5110 ( .A1(n2678), .A2(n4735), .ZN(n4659) );
  NAND2_X1 U5111 ( .A1(n4657), .A2(n4659), .ZN(n5160) );
  NOR4_X1 U5112 ( .A1(n4605), .A2(n4939), .A3(n5327), .A4(n5160), .ZN(n4615)
         );
  INV_X1 U5113 ( .A(n4888), .ZN(n4614) );
  INV_X1 U5114 ( .A(n4606), .ZN(n5182) );
  NOR4_X1 U5115 ( .A1(n4608), .A2(n5182), .A3(n3269), .A4(n4607), .ZN(n4613)
         );
  NOR4_X1 U5116 ( .A1(n4611), .A2(n4978), .A3(n4610), .A4(n4609), .ZN(n4612)
         );
  NAND4_X1 U5117 ( .A1(n4615), .A2(n4614), .A3(n4613), .A4(n4612), .ZN(n4636)
         );
  XNOR2_X1 U5118 ( .A(n4896), .B(n4874), .ZN(n4864) );
  INV_X1 U5119 ( .A(n4864), .ZN(n4635) );
  INV_X1 U5120 ( .A(n4616), .ZN(n4861) );
  NAND2_X1 U5121 ( .A1(n4861), .A2(n4859), .ZN(n4910) );
  INV_X1 U5122 ( .A(n4910), .ZN(n4901) );
  XNOR2_X1 U5123 ( .A(n4943), .B(n4962), .ZN(n4960) );
  INV_X1 U5124 ( .A(n4617), .ZN(n4626) );
  OR2_X1 U5125 ( .A1(n4704), .A2(n5103), .ZN(n4619) );
  NOR2_X1 U5126 ( .A1(n4619), .A2(n4618), .ZN(n4625) );
  INV_X1 U5127 ( .A(n4620), .ZN(n4624) );
  INV_X1 U5128 ( .A(n4621), .ZN(n4623) );
  NAND2_X1 U5129 ( .A1(n4623), .A2(n4622), .ZN(n4997) );
  NAND4_X1 U5130 ( .A1(n4626), .A2(n4625), .A3(n4624), .A4(n4997), .ZN(n4631)
         );
  NAND4_X1 U5131 ( .A1(n4629), .A2(n2597), .A3(n4628), .A4(n5251), .ZN(n4630)
         );
  NOR2_X1 U5132 ( .A1(n4631), .A2(n4630), .ZN(n4632) );
  NAND4_X1 U5133 ( .A1(n4901), .A2(n4633), .A3(n4960), .A4(n4632), .ZN(n4634)
         );
  NOR4_X1 U5134 ( .A1(n4846), .A2(n4636), .A3(n4635), .A4(n4634), .ZN(n4637)
         );
  NAND4_X1 U5135 ( .A1(n4639), .A2(n4638), .A3(n4818), .A4(n4637), .ZN(n4641)
         );
  NOR3_X1 U5136 ( .A1(n4641), .A2(n4775), .A3(n4640), .ZN(n4709) );
  AND2_X1 U5137 ( .A1(n4643), .A2(n4642), .ZN(n4680) );
  INV_X1 U5138 ( .A(n4644), .ZN(n4645) );
  NAND3_X1 U5139 ( .A1(n4680), .A2(n4645), .A3(n4672), .ZN(n4649) );
  NAND3_X1 U5140 ( .A1(n4650), .A2(n4647), .A3(n4646), .ZN(n4682) );
  AOI21_X1 U5141 ( .B1(n4649), .B2(n4648), .A(n4682), .ZN(n4655) );
  OAI211_X1 U5142 ( .C1(n2552), .C2(n4653), .A(n4652), .B(n4651), .ZN(n4654)
         );
  NOR2_X1 U5143 ( .A1(n4655), .A2(n4654), .ZN(n4686) );
  INV_X1 U5144 ( .A(n4656), .ZN(n4685) );
  INV_X1 U5145 ( .A(n4657), .ZN(n4660) );
  OAI211_X1 U5146 ( .C1(n4660), .C2(n5103), .A(n4659), .B(n4658), .ZN(n4663)
         );
  NAND3_X1 U5147 ( .A1(n4663), .A2(n4662), .A3(n4661), .ZN(n4666) );
  NAND3_X1 U5148 ( .A1(n4666), .A2(n4665), .A3(n4664), .ZN(n4669) );
  NAND3_X1 U5149 ( .A1(n4669), .A2(n4668), .A3(n4667), .ZN(n4673) );
  NAND4_X1 U5150 ( .A1(n4673), .A2(n4672), .A3(n4671), .A4(n4670), .ZN(n4675)
         );
  NAND3_X1 U5151 ( .A1(n4675), .A2(n4674), .A3(n3342), .ZN(n4681) );
  NAND2_X1 U5152 ( .A1(n4677), .A2(n4676), .ZN(n4678) );
  AOI22_X1 U5153 ( .A1(n4681), .A2(n4680), .B1(n4679), .B2(n4678), .ZN(n4683)
         );
  OR2_X1 U5154 ( .A1(n4683), .A2(n4682), .ZN(n4684) );
  OAI22_X1 U5155 ( .A1(n4687), .A2(n4686), .B1(n4685), .B2(n4684), .ZN(n4689)
         );
  AOI221_X1 U5156 ( .B1(n4691), .B2(n4690), .C1(n4689), .C2(n4690), .A(n4688), 
        .ZN(n4697) );
  NAND2_X1 U5157 ( .A1(n4693), .A2(n4692), .ZN(n4694) );
  AOI221_X1 U5158 ( .B1(n4697), .B2(n4696), .C1(n4695), .C2(n4696), .A(n4694), 
        .ZN(n4702) );
  INV_X1 U5159 ( .A(n4698), .ZN(n4700) );
  OAI211_X1 U5160 ( .C1(n4702), .C2(n4701), .A(n4700), .B(n4699), .ZN(n4706)
         );
  AOI22_X1 U5161 ( .A1(n4706), .A2(n4705), .B1(n4704), .B2(n4703), .ZN(n4707)
         );
  OAI22_X1 U5162 ( .A1(n4710), .A2(n4709), .B1(n4708), .B2(n4707), .ZN(n4711)
         );
  XNOR2_X1 U5163 ( .A(n4711), .B(n4767), .ZN(n4716) );
  NAND3_X1 U5164 ( .A1(n4712), .A2(n5099), .A3(n5304), .ZN(n4713) );
  OAI211_X1 U5165 ( .C1(n5102), .C2(n4715), .A(n4713), .B(B_REG_SCAN_IN), .ZN(
        n4714) );
  OAI21_X1 U5166 ( .B1(n4716), .B2(n4715), .A(n4714), .ZN(U3239) );
  MUX2_X1 U5167 ( .A(DATAO_REG_31__SCAN_IN), .B(n4717), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U5168 ( .A(n4718), .B(DATAO_REG_30__SCAN_IN), .S(n4734), .Z(U3580)
         );
  INV_X1 U5169 ( .A(n4719), .ZN(n4811) );
  MUX2_X1 U5170 ( .A(DATAO_REG_28__SCAN_IN), .B(n4811), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U5171 ( .A(DATAO_REG_27__SCAN_IN), .B(n4820), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U5172 ( .A(n4720), .B(DATAO_REG_26__SCAN_IN), .S(n4734), .Z(U3576)
         );
  MUX2_X1 U5173 ( .A(DATAO_REG_25__SCAN_IN), .B(n4853), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U5174 ( .A(n4870), .B(DATAO_REG_24__SCAN_IN), .S(n4734), .Z(U3574)
         );
  MUX2_X1 U5175 ( .A(n4896), .B(DATAO_REG_23__SCAN_IN), .S(n4734), .Z(U3573)
         );
  MUX2_X1 U5176 ( .A(n4903), .B(DATAO_REG_22__SCAN_IN), .S(n4734), .Z(U3572)
         );
  MUX2_X1 U5177 ( .A(DATAO_REG_21__SCAN_IN), .B(n4947), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U5178 ( .A(n4905), .B(DATAO_REG_20__SCAN_IN), .S(n4734), .Z(U3570)
         );
  MUX2_X1 U5179 ( .A(n4943), .B(DATAO_REG_19__SCAN_IN), .S(n4734), .Z(U3569)
         );
  MUX2_X1 U5180 ( .A(n4999), .B(DATAO_REG_18__SCAN_IN), .S(n4734), .Z(U3568)
         );
  MUX2_X1 U5181 ( .A(n4721), .B(DATAO_REG_17__SCAN_IN), .S(n4734), .Z(U3567)
         );
  MUX2_X1 U5182 ( .A(n4998), .B(DATAO_REG_16__SCAN_IN), .S(n4734), .Z(U3566)
         );
  MUX2_X1 U5183 ( .A(n4722), .B(DATAO_REG_15__SCAN_IN), .S(n4734), .Z(U3565)
         );
  MUX2_X1 U5184 ( .A(n5303), .B(DATAO_REG_14__SCAN_IN), .S(n4734), .Z(U3564)
         );
  MUX2_X1 U5185 ( .A(n4723), .B(DATAO_REG_13__SCAN_IN), .S(n4734), .Z(U3563)
         );
  MUX2_X1 U5186 ( .A(n5305), .B(DATAO_REG_12__SCAN_IN), .S(n4734), .Z(U3562)
         );
  MUX2_X1 U5187 ( .A(n4724), .B(DATAO_REG_11__SCAN_IN), .S(n4734), .Z(U3561)
         );
  MUX2_X1 U5188 ( .A(n4725), .B(DATAO_REG_10__SCAN_IN), .S(n4734), .Z(U3560)
         );
  MUX2_X1 U5189 ( .A(n4726), .B(DATAO_REG_9__SCAN_IN), .S(n4734), .Z(U3559) );
  MUX2_X1 U5190 ( .A(n4727), .B(DATAO_REG_8__SCAN_IN), .S(n4734), .Z(U3558) );
  MUX2_X1 U5191 ( .A(n4728), .B(DATAO_REG_7__SCAN_IN), .S(n4734), .Z(U3557) );
  MUX2_X1 U5192 ( .A(n4729), .B(DATAO_REG_6__SCAN_IN), .S(n4734), .Z(U3556) );
  MUX2_X1 U5193 ( .A(n4730), .B(DATAO_REG_5__SCAN_IN), .S(n4734), .Z(U3555) );
  MUX2_X1 U5194 ( .A(n4731), .B(DATAO_REG_4__SCAN_IN), .S(n4734), .Z(U3554) );
  MUX2_X1 U5195 ( .A(n4732), .B(DATAO_REG_3__SCAN_IN), .S(n4734), .Z(U3553) );
  MUX2_X1 U5196 ( .A(n4733), .B(DATAO_REG_2__SCAN_IN), .S(n4734), .Z(U3552) );
  MUX2_X1 U5197 ( .A(n2934), .B(DATAO_REG_1__SCAN_IN), .S(n4734), .Z(U3551) );
  MUX2_X1 U5198 ( .A(n4735), .B(DATAO_REG_0__SCAN_IN), .S(n4734), .Z(U3550) );
  AOI21_X1 U5199 ( .B1(n4737), .B2(REG1_REG_16__SCAN_IN), .A(n4736), .ZN(n4745) );
  AOI221_X1 U5200 ( .B1(n4739), .B2(n4738), .C1(n4044), .C2(n4738), .A(n4773), 
        .ZN(n4740) );
  INV_X1 U5201 ( .A(n4740), .ZN(n4744) );
  NOR2_X1 U5202 ( .A1(n4768), .A2(n5379), .ZN(n4741) );
  AOI211_X1 U5203 ( .C1(n5143), .C2(ADDR_REG_16__SCAN_IN), .A(n4742), .B(n4741), .ZN(n4743) );
  OAI211_X1 U5204 ( .C1(n4745), .C2(n4756), .A(n4744), .B(n4743), .ZN(U3256)
         );
  AOI21_X1 U5205 ( .B1(n4747), .B2(n4746), .A(n4305), .ZN(n4757) );
  AOI211_X1 U5206 ( .C1(n4750), .C2(n4749), .A(n4748), .B(n4773), .ZN(n4751)
         );
  AOI211_X1 U5207 ( .C1(n5143), .C2(ADDR_REG_17__SCAN_IN), .A(n4752), .B(n4751), .ZN(n4755) );
  NAND2_X1 U5208 ( .A1(n4753), .A2(n5105), .ZN(n4754) );
  OAI211_X1 U5209 ( .C1(n4757), .C2(n4756), .A(n4755), .B(n4754), .ZN(U3257)
         );
  INV_X1 U5210 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4759) );
  MUX2_X1 U5211 ( .A(REG2_REG_19__SCAN_IN), .B(n4759), .S(n4767), .Z(n4760) );
  XNOR2_X1 U5212 ( .A(n4761), .B(n4760), .ZN(n4774) );
  XNOR2_X1 U5213 ( .A(n4767), .B(REG1_REG_19__SCAN_IN), .ZN(n4763) );
  XNOR2_X1 U5214 ( .A(n4764), .B(n4763), .ZN(n4771) );
  NAND2_X1 U5215 ( .A1(n5143), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4766) );
  OAI211_X1 U5216 ( .C1(n4768), .C2(n4767), .A(n4766), .B(n4765), .ZN(n4769)
         );
  AOI21_X1 U5217 ( .B1(n4771), .B2(n4770), .A(n4769), .ZN(n4772) );
  OAI21_X1 U5218 ( .B1(n4774), .B2(n4773), .A(n4772), .ZN(U3259) );
  XNOR2_X1 U5219 ( .A(n4776), .B(n4775), .ZN(n5055) );
  OAI21_X1 U5220 ( .B1(n4779), .B2(n4778), .A(n4777), .ZN(n4780) );
  NAND2_X1 U5221 ( .A1(n4780), .A2(n5333), .ZN(n4785) );
  OAI22_X1 U5222 ( .A1(n4782), .A2(n5184), .B1(n4781), .B2(n5330), .ZN(n4783)
         );
  INV_X1 U5223 ( .A(n4783), .ZN(n4784) );
  OAI211_X1 U5224 ( .C1(n4786), .C2(n5186), .A(n4785), .B(n4784), .ZN(n5011)
         );
  INV_X1 U5225 ( .A(n4799), .ZN(n4788) );
  INV_X1 U5226 ( .A(n5012), .ZN(n4792) );
  AOI22_X1 U5227 ( .A1(n4790), .A2(n5204), .B1(REG2_REG_28__SCAN_IN), .B2(
        n5402), .ZN(n4791) );
  OAI21_X1 U5228 ( .B1(n4792), .B2(n4877), .A(n4791), .ZN(n4793) );
  AOI21_X1 U5229 ( .B1(n5341), .B2(n5011), .A(n4793), .ZN(n4794) );
  OAI21_X1 U5230 ( .B1(n5055), .B2(n4991), .A(n4794), .ZN(U3262) );
  XNOR2_X1 U5231 ( .A(n4795), .B(n4803), .ZN(n5059) );
  NAND2_X1 U5232 ( .A1(n2486), .A2(n4796), .ZN(n4797) );
  NAND2_X1 U5233 ( .A1(n4797), .A2(n5406), .ZN(n4798) );
  NOR2_X1 U5234 ( .A1(n4799), .A2(n4798), .ZN(n5015) );
  INV_X1 U5235 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4800) );
  OAI22_X1 U5236 ( .A1(n4801), .A2(n5339), .B1(n4800), .B2(n5262), .ZN(n4802)
         );
  AOI21_X1 U5237 ( .B1(n5015), .B2(n4976), .A(n4802), .ZN(n4815) );
  NAND2_X1 U5238 ( .A1(n4804), .A2(n4803), .ZN(n4805) );
  NAND2_X1 U5239 ( .A1(n4806), .A2(n4805), .ZN(n4807) );
  NAND2_X1 U5240 ( .A1(n4807), .A2(n5333), .ZN(n4813) );
  OAI22_X1 U5241 ( .A1(n4809), .A2(n5186), .B1(n5330), .B2(n4808), .ZN(n4810)
         );
  AOI21_X1 U5242 ( .B1(n4811), .B2(n5302), .A(n4810), .ZN(n4812) );
  NAND2_X1 U5243 ( .A1(n4813), .A2(n4812), .ZN(n5016) );
  NAND2_X1 U5244 ( .A1(n5016), .A2(n5262), .ZN(n4814) );
  OAI211_X1 U5245 ( .C1(n5059), .C2(n4991), .A(n4815), .B(n4814), .ZN(U3263)
         );
  NAND2_X1 U5246 ( .A1(n4817), .A2(n4816), .ZN(n4819) );
  XNOR2_X1 U5247 ( .A(n4819), .B(n4818), .ZN(n4826) );
  NAND2_X1 U5248 ( .A1(n4820), .A2(n5302), .ZN(n4823) );
  OR2_X1 U5249 ( .A1(n4821), .A2(n5186), .ZN(n4822) );
  OAI211_X1 U5250 ( .C1(n5330), .C2(n4824), .A(n4823), .B(n4822), .ZN(n4825)
         );
  AOI21_X1 U5251 ( .B1(n4826), .B2(n5333), .A(n4825), .ZN(n5019) );
  XOR2_X1 U5252 ( .A(n4828), .B(n4827), .Z(n5064) );
  INV_X1 U5253 ( .A(n5064), .ZN(n4829) );
  NAND2_X1 U5254 ( .A1(n4829), .A2(n5345), .ZN(n4837) );
  NAND2_X1 U5255 ( .A1(n2505), .A2(n4830), .ZN(n4831) );
  NAND2_X1 U5256 ( .A1(n2486), .A2(n4831), .ZN(n5020) );
  INV_X1 U5257 ( .A(n5020), .ZN(n4835) );
  INV_X1 U5258 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4832) );
  OAI22_X1 U5259 ( .A1(n4833), .A2(n5339), .B1(n4832), .B2(n5341), .ZN(n4834)
         );
  AOI21_X1 U5260 ( .B1(n4835), .B2(n5415), .A(n4834), .ZN(n4836) );
  OAI211_X1 U5261 ( .C1(n5419), .C2(n5019), .A(n4837), .B(n4836), .ZN(U3264)
         );
  XNOR2_X1 U5262 ( .A(n4838), .B(n4846), .ZN(n5068) );
  OAI21_X1 U5263 ( .B1(n4873), .B2(n4851), .A(n5406), .ZN(n4840) );
  NOR2_X1 U5264 ( .A1(n4840), .A2(n4839), .ZN(n5023) );
  INV_X1 U5265 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4841) );
  OAI22_X1 U5266 ( .A1(n4842), .A2(n5339), .B1(n4841), .B2(n5262), .ZN(n4843)
         );
  AOI21_X1 U5267 ( .B1(n5023), .B2(n4976), .A(n4843), .ZN(n4857) );
  NAND2_X1 U5268 ( .A1(n4845), .A2(n4844), .ZN(n4848) );
  INV_X1 U5269 ( .A(n4846), .ZN(n4847) );
  XNOR2_X1 U5270 ( .A(n4848), .B(n4847), .ZN(n4849) );
  NAND2_X1 U5271 ( .A1(n4849), .A2(n5333), .ZN(n4855) );
  NAND2_X1 U5272 ( .A1(n4896), .A2(n5304), .ZN(n4850) );
  OAI21_X1 U5273 ( .B1(n5330), .B2(n4851), .A(n4850), .ZN(n4852) );
  AOI21_X1 U5274 ( .B1(n4853), .B2(n5302), .A(n4852), .ZN(n4854) );
  NAND2_X1 U5275 ( .A1(n4855), .A2(n4854), .ZN(n5024) );
  NAND2_X1 U5276 ( .A1(n5024), .A2(n5262), .ZN(n4856) );
  OAI211_X1 U5277 ( .C1(n5068), .C2(n4991), .A(n4857), .B(n4856), .ZN(U3266)
         );
  XNOR2_X1 U5278 ( .A(n4858), .B(n4864), .ZN(n5072) );
  INV_X1 U5279 ( .A(n4859), .ZN(n4860) );
  OR2_X1 U5280 ( .A1(n4902), .A2(n4860), .ZN(n4862) );
  NAND2_X1 U5281 ( .A1(n4862), .A2(n4861), .ZN(n4889) );
  NAND2_X1 U5282 ( .A1(n4891), .A2(n4863), .ZN(n4865) );
  XNOR2_X1 U5283 ( .A(n4865), .B(n4864), .ZN(n4866) );
  NAND2_X1 U5284 ( .A1(n4866), .A2(n5333), .ZN(n4872) );
  NAND2_X1 U5285 ( .A1(n4903), .A2(n5304), .ZN(n4867) );
  OAI21_X1 U5286 ( .B1(n5330), .B2(n4868), .A(n4867), .ZN(n4869) );
  AOI21_X1 U5287 ( .B1(n4870), .B2(n5302), .A(n4869), .ZN(n4871) );
  NAND2_X1 U5288 ( .A1(n4872), .A2(n4871), .ZN(n5028) );
  AOI211_X1 U5289 ( .C1(n4874), .C2(n4883), .A(n5390), .B(n4873), .ZN(n5027)
         );
  INV_X1 U5290 ( .A(n5027), .ZN(n4878) );
  AOI22_X1 U5291 ( .A1(n4875), .A2(n5204), .B1(REG2_REG_23__SCAN_IN), .B2(
        n5419), .ZN(n4876) );
  OAI21_X1 U5292 ( .B1(n4878), .B2(n4877), .A(n4876), .ZN(n4879) );
  AOI21_X1 U5293 ( .B1(n5341), .B2(n5028), .A(n4879), .ZN(n4880) );
  OAI21_X1 U5294 ( .B1(n5072), .B2(n4991), .A(n4880), .ZN(U3267) );
  XNOR2_X1 U5295 ( .A(n4881), .B(n4888), .ZN(n5076) );
  AOI21_X1 U5296 ( .B1(n4913), .B2(n4882), .A(n5390), .ZN(n4884) );
  AND2_X1 U5297 ( .A1(n4884), .A2(n4883), .ZN(n5031) );
  INV_X1 U5298 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4885) );
  OAI22_X1 U5299 ( .A1(n4886), .A2(n5339), .B1(n4885), .B2(n5341), .ZN(n4887)
         );
  AOI21_X1 U5300 ( .B1(n5031), .B2(n4976), .A(n4887), .ZN(n4900) );
  NAND2_X1 U5301 ( .A1(n4889), .A2(n4888), .ZN(n4890) );
  NAND2_X1 U5302 ( .A1(n4891), .A2(n4890), .ZN(n4892) );
  NAND2_X1 U5303 ( .A1(n4892), .A2(n5333), .ZN(n4898) );
  NAND2_X1 U5304 ( .A1(n4947), .A2(n5304), .ZN(n4893) );
  OAI21_X1 U5305 ( .B1(n5330), .B2(n4894), .A(n4893), .ZN(n4895) );
  AOI21_X1 U5306 ( .B1(n4896), .B2(n5302), .A(n4895), .ZN(n4897) );
  NAND2_X1 U5307 ( .A1(n4898), .A2(n4897), .ZN(n5032) );
  NAND2_X1 U5308 ( .A1(n5032), .A2(n5262), .ZN(n4899) );
  OAI211_X1 U5309 ( .C1(n5076), .C2(n4991), .A(n4900), .B(n4899), .ZN(U3268)
         );
  XNOR2_X1 U5310 ( .A(n4902), .B(n4901), .ZN(n4909) );
  NAND2_X1 U5311 ( .A1(n4903), .A2(n5302), .ZN(n4907) );
  AOI22_X1 U5312 ( .A1(n4905), .A2(n5304), .B1(n4904), .B2(n5396), .ZN(n4906)
         );
  NAND2_X1 U5313 ( .A1(n4907), .A2(n4906), .ZN(n4908) );
  AOI21_X1 U5314 ( .B1(n4909), .B2(n5333), .A(n4908), .ZN(n5036) );
  XNOR2_X1 U5315 ( .A(n4911), .B(n4910), .ZN(n5080) );
  INV_X1 U5316 ( .A(n5080), .ZN(n4912) );
  NAND2_X1 U5317 ( .A1(n4912), .A2(n5345), .ZN(n4920) );
  OAI211_X1 U5318 ( .C1(n4925), .C2(n4914), .A(n5406), .B(n4913), .ZN(n5035)
         );
  INV_X1 U5319 ( .A(n5035), .ZN(n4918) );
  INV_X1 U5320 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4915) );
  OAI22_X1 U5321 ( .A1(n4916), .A2(n5339), .B1(n4915), .B2(n5341), .ZN(n4917)
         );
  AOI21_X1 U5322 ( .B1(n4918), .B2(n4976), .A(n4917), .ZN(n4919) );
  OAI211_X1 U5323 ( .C1(n5419), .C2(n5036), .A(n4920), .B(n4919), .ZN(U3269)
         );
  XNOR2_X1 U5324 ( .A(n4921), .B(n4939), .ZN(n5084) );
  NAND2_X1 U5325 ( .A1(n4963), .A2(n4922), .ZN(n4923) );
  NAND2_X1 U5326 ( .A1(n4923), .A2(n5406), .ZN(n4924) );
  NOR2_X1 U5327 ( .A1(n4925), .A2(n4924), .ZN(n5039) );
  INV_X1 U5328 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4927) );
  OAI22_X1 U5329 ( .A1(n4927), .A2(n5262), .B1(n4926), .B2(n5339), .ZN(n4928)
         );
  AOI21_X1 U5330 ( .B1(n5039), .B2(n4976), .A(n4928), .ZN(n4951) );
  NAND2_X1 U5331 ( .A1(n4930), .A2(n4929), .ZN(n4996) );
  NAND2_X1 U5332 ( .A1(n4996), .A2(n4931), .ZN(n4933) );
  NAND2_X1 U5333 ( .A1(n4933), .A2(n4932), .ZN(n4980) );
  NAND2_X1 U5334 ( .A1(n4980), .A2(n4934), .ZN(n4983) );
  INV_X1 U5335 ( .A(n4935), .ZN(n4936) );
  NAND2_X1 U5336 ( .A1(n4983), .A2(n4936), .ZN(n4938) );
  NAND2_X1 U5337 ( .A1(n4938), .A2(n4937), .ZN(n4941) );
  INV_X1 U5338 ( .A(n4939), .ZN(n4940) );
  XNOR2_X1 U5339 ( .A(n4941), .B(n4940), .ZN(n4942) );
  NAND2_X1 U5340 ( .A1(n4942), .A2(n5333), .ZN(n4949) );
  NAND2_X1 U5341 ( .A1(n4943), .A2(n5304), .ZN(n4944) );
  OAI21_X1 U5342 ( .B1(n5330), .B2(n4945), .A(n4944), .ZN(n4946) );
  AOI21_X1 U5343 ( .B1(n4947), .B2(n5302), .A(n4946), .ZN(n4948) );
  NAND2_X1 U5344 ( .A1(n4949), .A2(n4948), .ZN(n5040) );
  NAND2_X1 U5345 ( .A1(n5040), .A2(n5262), .ZN(n4950) );
  OAI211_X1 U5346 ( .C1(n5084), .C2(n4991), .A(n4951), .B(n4950), .ZN(U3270)
         );
  NAND2_X1 U5347 ( .A1(n4983), .A2(n4977), .ZN(n4953) );
  INV_X1 U5348 ( .A(n4960), .ZN(n4952) );
  XNOR2_X1 U5349 ( .A(n4953), .B(n4952), .ZN(n4958) );
  INV_X1 U5350 ( .A(n4954), .ZN(n4955) );
  OAI21_X1 U5351 ( .B1(n4956), .B2(n5330), .A(n4955), .ZN(n4957) );
  AOI21_X1 U5352 ( .B1(n4958), .B2(n5333), .A(n4957), .ZN(n5044) );
  XOR2_X1 U5353 ( .A(n4960), .B(n4959), .Z(n5088) );
  INV_X1 U5354 ( .A(n5088), .ZN(n4961) );
  NAND2_X1 U5355 ( .A1(n4961), .A2(n5345), .ZN(n4969) );
  AOI21_X1 U5356 ( .B1(n4971), .B2(n4962), .A(n5390), .ZN(n4964) );
  NAND2_X1 U5357 ( .A1(n4964), .A2(n4963), .ZN(n5043) );
  INV_X1 U5358 ( .A(n5043), .ZN(n4967) );
  OAI22_X1 U5359 ( .A1(n5262), .A2(n4759), .B1(n4965), .B2(n5339), .ZN(n4966)
         );
  AOI21_X1 U5360 ( .B1(n4967), .B2(n4976), .A(n4966), .ZN(n4968) );
  OAI211_X1 U5361 ( .C1(n5419), .C2(n5044), .A(n4969), .B(n4968), .ZN(U3271)
         );
  XOR2_X1 U5362 ( .A(n4978), .B(n4970), .Z(n5093) );
  AOI21_X1 U5363 ( .B1(n4994), .B2(n4984), .A(n5390), .ZN(n4972) );
  AND2_X1 U5364 ( .A1(n4972), .A2(n4971), .ZN(n5047) );
  INV_X1 U5365 ( .A(n4973), .ZN(n4974) );
  OAI22_X1 U5366 ( .A1(n5262), .A2(n4319), .B1(n4974), .B2(n5339), .ZN(n4975)
         );
  AOI21_X1 U5367 ( .B1(n5047), .B2(n4976), .A(n4975), .ZN(n4990) );
  INV_X1 U5368 ( .A(n4977), .ZN(n4982) );
  INV_X1 U5369 ( .A(n4978), .ZN(n4979) );
  OR2_X1 U5370 ( .A1(n4980), .A2(n4979), .ZN(n4981) );
  OAI211_X1 U5371 ( .C1(n4983), .C2(n4982), .A(n5333), .B(n4981), .ZN(n4988)
         );
  AND2_X1 U5372 ( .A1(n4984), .A2(n5396), .ZN(n4985) );
  NOR2_X1 U5373 ( .A1(n4986), .A2(n4985), .ZN(n4987) );
  NAND2_X1 U5374 ( .A1(n4988), .A2(n4987), .ZN(n5048) );
  NAND2_X1 U5375 ( .A1(n5048), .A2(n5262), .ZN(n4989) );
  OAI211_X1 U5376 ( .C1(n5093), .C2(n4991), .A(n4990), .B(n4989), .ZN(U3272)
         );
  OR2_X1 U5377 ( .A1(n4992), .A2(n5001), .ZN(n4993) );
  NAND2_X1 U5378 ( .A1(n4994), .A2(n4993), .ZN(n5389) );
  XNOR2_X1 U5379 ( .A(n4995), .B(n4997), .ZN(n5393) );
  NAND2_X1 U5380 ( .A1(n5393), .A2(n5345), .ZN(n5009) );
  XOR2_X1 U5381 ( .A(n4997), .B(n4996), .Z(n5003) );
  AOI22_X1 U5382 ( .A1(n5302), .A2(n4999), .B1(n4998), .B2(n5304), .ZN(n5000)
         );
  OAI21_X1 U5383 ( .B1(n5001), .B2(n5330), .A(n5000), .ZN(n5002) );
  AOI21_X1 U5384 ( .B1(n5003), .B2(n5333), .A(n5002), .ZN(n5388) );
  OAI21_X1 U5385 ( .B1(n5004), .B2(n5339), .A(n5388), .ZN(n5007) );
  INV_X1 U5386 ( .A(REG2_REG_17__SCAN_IN), .ZN(n5005) );
  NOR2_X1 U5387 ( .A1(n5262), .A2(n5005), .ZN(n5006) );
  AOI21_X1 U5388 ( .B1(n5007), .B2(n5262), .A(n5006), .ZN(n5008) );
  OAI211_X1 U5389 ( .C1(n5389), .C2(n5010), .A(n5009), .B(n5008), .ZN(U3273)
         );
  INV_X1 U5390 ( .A(REG1_REG_28__SCAN_IN), .ZN(n5013) );
  NOR2_X1 U5391 ( .A1(n5012), .A2(n5011), .ZN(n5052) );
  MUX2_X1 U5392 ( .A(n5013), .B(n5052), .S(n5410), .Z(n5014) );
  OAI21_X1 U5393 ( .B1(n5055), .B2(n5051), .A(n5014), .ZN(U3546) );
  INV_X1 U5394 ( .A(REG1_REG_27__SCAN_IN), .ZN(n5017) );
  NOR2_X1 U5395 ( .A1(n5016), .A2(n5015), .ZN(n5056) );
  MUX2_X1 U5396 ( .A(n5017), .B(n5056), .S(n5410), .Z(n5018) );
  OAI21_X1 U5397 ( .B1(n5059), .B2(n5051), .A(n5018), .ZN(U3545) );
  OAI21_X1 U5398 ( .B1(n5390), .B2(n5020), .A(n5019), .ZN(n5060) );
  MUX2_X1 U5399 ( .A(REG1_REG_26__SCAN_IN), .B(n5060), .S(n5410), .Z(n5021) );
  INV_X1 U5400 ( .A(n5021), .ZN(n5022) );
  OAI21_X1 U5401 ( .B1(n5064), .B2(n5051), .A(n5022), .ZN(U3544) );
  INV_X1 U5402 ( .A(REG1_REG_24__SCAN_IN), .ZN(n5025) );
  NOR2_X1 U5403 ( .A1(n5024), .A2(n5023), .ZN(n5065) );
  MUX2_X1 U5404 ( .A(n5025), .B(n5065), .S(n5410), .Z(n5026) );
  OAI21_X1 U5405 ( .B1(n5068), .B2(n5051), .A(n5026), .ZN(U3542) );
  INV_X1 U5406 ( .A(REG1_REG_23__SCAN_IN), .ZN(n5029) );
  NOR2_X1 U5407 ( .A1(n5028), .A2(n5027), .ZN(n5069) );
  MUX2_X1 U5408 ( .A(n5029), .B(n5069), .S(n5410), .Z(n5030) );
  OAI21_X1 U5409 ( .B1(n5072), .B2(n5051), .A(n5030), .ZN(U3541) );
  INV_X1 U5410 ( .A(REG1_REG_22__SCAN_IN), .ZN(n5033) );
  NOR2_X1 U5411 ( .A1(n5032), .A2(n5031), .ZN(n5073) );
  MUX2_X1 U5412 ( .A(n5033), .B(n5073), .S(n5410), .Z(n5034) );
  OAI21_X1 U5413 ( .B1(n5076), .B2(n5051), .A(n5034), .ZN(U3540) );
  INV_X1 U5414 ( .A(REG1_REG_21__SCAN_IN), .ZN(n5037) );
  AND2_X1 U5415 ( .A1(n5036), .A2(n5035), .ZN(n5077) );
  MUX2_X1 U5416 ( .A(n5037), .B(n5077), .S(n5410), .Z(n5038) );
  OAI21_X1 U5417 ( .B1(n5080), .B2(n5051), .A(n5038), .ZN(U3539) );
  INV_X1 U5418 ( .A(REG1_REG_20__SCAN_IN), .ZN(n5041) );
  NOR2_X1 U5419 ( .A1(n5040), .A2(n5039), .ZN(n5081) );
  MUX2_X1 U5420 ( .A(n5041), .B(n5081), .S(n5410), .Z(n5042) );
  OAI21_X1 U5421 ( .B1(n5084), .B2(n5051), .A(n5042), .ZN(U3538) );
  INV_X1 U5422 ( .A(REG1_REG_19__SCAN_IN), .ZN(n5045) );
  AND2_X1 U5423 ( .A1(n5044), .A2(n5043), .ZN(n5085) );
  MUX2_X1 U5424 ( .A(n5045), .B(n5085), .S(n5410), .Z(n5046) );
  OAI21_X1 U5425 ( .B1(n5088), .B2(n5051), .A(n5046), .ZN(U3537) );
  INV_X1 U5426 ( .A(REG1_REG_18__SCAN_IN), .ZN(n5049) );
  NOR2_X1 U5427 ( .A1(n5048), .A2(n5047), .ZN(n5089) );
  MUX2_X1 U5428 ( .A(n5049), .B(n5089), .S(n5410), .Z(n5050) );
  OAI21_X1 U5429 ( .B1(n5093), .B2(n5051), .A(n5050), .ZN(U3536) );
  MUX2_X1 U5430 ( .A(n5053), .B(n5052), .S(n5414), .Z(n5054) );
  OAI21_X1 U5431 ( .B1(n5055), .B2(n5092), .A(n5054), .ZN(U3514) );
  MUX2_X1 U5432 ( .A(n5057), .B(n5056), .S(n5414), .Z(n5058) );
  OAI21_X1 U5433 ( .B1(n5059), .B2(n5092), .A(n5058), .ZN(U3513) );
  INV_X1 U5434 ( .A(n5060), .ZN(n5061) );
  MUX2_X1 U5435 ( .A(n5062), .B(n5061), .S(n5414), .Z(n5063) );
  OAI21_X1 U5436 ( .B1(n5064), .B2(n5092), .A(n5063), .ZN(U3512) );
  MUX2_X1 U5437 ( .A(n5066), .B(n5065), .S(n5414), .Z(n5067) );
  OAI21_X1 U5438 ( .B1(n5068), .B2(n5092), .A(n5067), .ZN(U3510) );
  MUX2_X1 U5439 ( .A(n5070), .B(n5069), .S(n5414), .Z(n5071) );
  OAI21_X1 U5440 ( .B1(n5072), .B2(n5092), .A(n5071), .ZN(U3509) );
  MUX2_X1 U5441 ( .A(n5074), .B(n5073), .S(n5414), .Z(n5075) );
  OAI21_X1 U5442 ( .B1(n5076), .B2(n5092), .A(n5075), .ZN(U3508) );
  MUX2_X1 U5443 ( .A(n5078), .B(n5077), .S(n5414), .Z(n5079) );
  OAI21_X1 U5444 ( .B1(n5080), .B2(n5092), .A(n5079), .ZN(U3507) );
  MUX2_X1 U5445 ( .A(n5082), .B(n5081), .S(n5414), .Z(n5083) );
  OAI21_X1 U5446 ( .B1(n5084), .B2(n5092), .A(n5083), .ZN(U3506) );
  MUX2_X1 U5447 ( .A(n5086), .B(n5085), .S(n5414), .Z(n5087) );
  OAI21_X1 U5448 ( .B1(n5088), .B2(n5092), .A(n5087), .ZN(U3505) );
  INV_X1 U5449 ( .A(REG0_REG_18__SCAN_IN), .ZN(n5090) );
  MUX2_X1 U5450 ( .A(n5090), .B(n5089), .S(n5414), .Z(n5091) );
  OAI21_X1 U5451 ( .B1(n5093), .B2(n5092), .A(n5091), .ZN(U3503) );
  NOR3_X1 U5452 ( .A1(n5095), .A2(IR_REG_30__SCAN_IN), .A3(n5094), .ZN(n5096)
         );
  MUX2_X1 U5453 ( .A(n5096), .B(DATAI_31_), .S(U3149), .Z(U3321) );
  MUX2_X1 U5454 ( .A(n5097), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5455 ( .A(n5098), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5456 ( .A(DATAI_27_), .B(n5099), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5457 ( .A(n5100), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5458 ( .A(n5101), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5459 ( .A(n2778), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5460 ( .A(n5102), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5461 ( .A(n5103), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5462 ( .A(DATAI_19_), .B(n5265), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5463 ( .A(DATAI_18_), .B(n5104), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5464 ( .A(n5105), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5465 ( .A(DATAI_14_), .B(n5106), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5466 ( .A(n5107), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  MUX2_X1 U5467 ( .A(n5108), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5468 ( .A(DATAI_8_), .B(n5109), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5469 ( .A(n5110), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5470 ( .A(DATAI_4_), .B(n5111), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5471 ( .A(n5112), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  NOR2_X1 U5472 ( .A1(n5136), .A2(n5113), .ZN(U3320) );
  AND2_X1 U5473 ( .A1(n5130), .A2(D_REG_3__SCAN_IN), .ZN(U3319) );
  NOR2_X1 U5474 ( .A1(n5136), .A2(n5114), .ZN(U3318) );
  AND2_X1 U5475 ( .A1(n5130), .A2(D_REG_5__SCAN_IN), .ZN(U3317) );
  AND2_X1 U5476 ( .A1(n5130), .A2(D_REG_6__SCAN_IN), .ZN(U3316) );
  INV_X1 U5477 ( .A(D_REG_7__SCAN_IN), .ZN(n5115) );
  NOR2_X1 U5478 ( .A1(n5136), .A2(n5115), .ZN(U3315) );
  INV_X1 U5479 ( .A(D_REG_8__SCAN_IN), .ZN(n5116) );
  NOR2_X1 U5480 ( .A1(n5136), .A2(n5116), .ZN(U3314) );
  INV_X1 U5481 ( .A(D_REG_9__SCAN_IN), .ZN(n5117) );
  NOR2_X1 U5482 ( .A1(n5136), .A2(n5117), .ZN(U3313) );
  NOR2_X1 U5483 ( .A1(n5136), .A2(n5118), .ZN(U3312) );
  AND2_X1 U5484 ( .A1(n5130), .A2(D_REG_11__SCAN_IN), .ZN(U3311) );
  NOR2_X1 U5485 ( .A1(n5136), .A2(n5119), .ZN(U3310) );
  INV_X1 U5486 ( .A(D_REG_13__SCAN_IN), .ZN(n5120) );
  NOR2_X1 U5487 ( .A1(n5136), .A2(n5120), .ZN(U3309) );
  NOR2_X1 U5488 ( .A1(n5136), .A2(n5121), .ZN(U3308) );
  NOR2_X1 U5489 ( .A1(n5136), .A2(n5122), .ZN(U3307) );
  INV_X1 U5490 ( .A(D_REG_16__SCAN_IN), .ZN(n5123) );
  NOR2_X1 U5491 ( .A1(n5136), .A2(n5123), .ZN(U3306) );
  AND2_X1 U5492 ( .A1(n5130), .A2(D_REG_17__SCAN_IN), .ZN(U3305) );
  NOR2_X1 U5493 ( .A1(n5136), .A2(n5124), .ZN(U3304) );
  NOR2_X1 U5494 ( .A1(n5136), .A2(n5125), .ZN(U3303) );
  NOR2_X1 U5495 ( .A1(n5136), .A2(n5126), .ZN(U3302) );
  NOR2_X1 U5496 ( .A1(n5136), .A2(n5127), .ZN(U3301) );
  INV_X1 U5497 ( .A(D_REG_22__SCAN_IN), .ZN(n5128) );
  NOR2_X1 U5498 ( .A1(n5136), .A2(n5128), .ZN(U3300) );
  NOR2_X1 U5499 ( .A1(n5136), .A2(n5129), .ZN(U3299) );
  AND2_X1 U5500 ( .A1(n5130), .A2(D_REG_24__SCAN_IN), .ZN(U3298) );
  AND2_X1 U5501 ( .A1(n5130), .A2(D_REG_25__SCAN_IN), .ZN(U3297) );
  AND2_X1 U5502 ( .A1(n5130), .A2(D_REG_26__SCAN_IN), .ZN(U3296) );
  NOR2_X1 U5503 ( .A1(n5136), .A2(n5131), .ZN(U3295) );
  NOR2_X1 U5504 ( .A1(n5136), .A2(n5132), .ZN(U3294) );
  INV_X1 U5505 ( .A(D_REG_29__SCAN_IN), .ZN(n5133) );
  NOR2_X1 U5506 ( .A1(n5136), .A2(n5133), .ZN(U3293) );
  INV_X1 U5507 ( .A(D_REG_30__SCAN_IN), .ZN(n5134) );
  NOR2_X1 U5508 ( .A1(n5136), .A2(n5134), .ZN(U3292) );
  INV_X1 U5509 ( .A(D_REG_31__SCAN_IN), .ZN(n5135) );
  NOR2_X1 U5510 ( .A1(n5136), .A2(n5135), .ZN(U3291) );
  NAND2_X1 U5511 ( .A1(n5137), .A2(n2873), .ZN(n5142) );
  INV_X1 U5512 ( .A(n5138), .ZN(n5141) );
  NAND3_X1 U5513 ( .A1(n5139), .A2(IR_REG_0__SCAN_IN), .A3(n5142), .ZN(n5140)
         );
  OAI211_X1 U5514 ( .C1(IR_REG_0__SCAN_IN), .C2(n5142), .A(n5141), .B(n5140), 
        .ZN(n5145) );
  AOI22_X1 U5515 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n5143), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n5144) );
  OAI21_X1 U5516 ( .B1(n5146), .B2(n5145), .A(n5144), .ZN(U3240) );
  INV_X1 U5517 ( .A(DATAI_0_), .ZN(n5147) );
  AOI22_X1 U5518 ( .A1(STATE_REG_SCAN_IN), .A2(n5148), .B1(n5147), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5519 ( .A(n5228), .ZN(n5198) );
  NOR2_X1 U5520 ( .A1(n2678), .A2(n5149), .ZN(n5157) );
  INV_X1 U5521 ( .A(n3273), .ZN(n5193) );
  OAI21_X1 U5522 ( .B1(n5193), .B2(n5333), .A(n5160), .ZN(n5150) );
  OAI21_X1 U5523 ( .B1(n5151), .B2(n5184), .A(n5150), .ZN(n5155) );
  AOI211_X1 U5524 ( .C1(n5198), .C2(n5160), .A(n5157), .B(n5155), .ZN(n5153)
         );
  AOI22_X1 U5525 ( .A1(n5410), .A2(n5153), .B1(n2873), .B2(n5408), .ZN(U3518)
         );
  INV_X1 U5526 ( .A(REG0_REG_0__SCAN_IN), .ZN(n5152) );
  AOI22_X1 U5527 ( .A1(n5414), .A2(n5153), .B1(n5152), .B2(n5411), .ZN(U3467)
         );
  INV_X1 U5528 ( .A(n5341), .ZN(n5419) );
  INV_X1 U5529 ( .A(n5154), .ZN(n5156) );
  AOI21_X1 U5530 ( .B1(n5157), .B2(n5156), .A(n5155), .ZN(n5162) );
  INV_X1 U5531 ( .A(n5158), .ZN(n5159) );
  AND2_X1 U5532 ( .A1(n5341), .A2(n5159), .ZN(n5206) );
  AOI22_X1 U5533 ( .A1(REG3_REG_0__SCAN_IN), .A2(n5204), .B1(n5206), .B2(n5160), .ZN(n5161) );
  OAI221_X1 U5534 ( .B1(n5419), .B2(n5162), .C1(n5341), .C2(n2877), .A(n5161), 
        .ZN(U3290) );
  AOI22_X1 U5535 ( .A1(STATE_REG_SCAN_IN), .A2(n2840), .B1(n5163), .B2(U3149), 
        .ZN(U3351) );
  INV_X1 U5536 ( .A(n5392), .ZN(n5381) );
  NAND3_X1 U5537 ( .A1(n5165), .A2(n5164), .A3(n5406), .ZN(n5166) );
  OAI211_X1 U5538 ( .C1(n5381), .C2(n5168), .A(n5167), .B(n5166), .ZN(n5169)
         );
  INV_X1 U5539 ( .A(n5169), .ZN(n5172) );
  AOI22_X1 U5540 ( .A1(n5410), .A2(n5172), .B1(n5170), .B2(n5408), .ZN(U3519)
         );
  INV_X1 U5541 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5171) );
  AOI22_X1 U5542 ( .A1(n5414), .A2(n5172), .B1(n5171), .B2(n5411), .ZN(U3469)
         );
  INV_X1 U5543 ( .A(DATAI_2_), .ZN(n5173) );
  AOI22_X1 U5544 ( .A1(STATE_REG_SCAN_IN), .A2(n2838), .B1(n5173), .B2(U3149), 
        .ZN(U3350) );
  OAI22_X1 U5545 ( .A1(n5175), .A2(n5381), .B1(n5390), .B2(n5174), .ZN(n5177)
         );
  NOR2_X1 U5546 ( .A1(n5177), .A2(n5176), .ZN(n5180) );
  AOI22_X1 U5547 ( .A1(n5410), .A2(n5180), .B1(n5178), .B2(n5408), .ZN(U3520)
         );
  INV_X1 U5548 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5179) );
  AOI22_X1 U5549 ( .A1(n5414), .A2(n5180), .B1(n5179), .B2(n5411), .ZN(U3471)
         );
  XNOR2_X1 U5550 ( .A(n5181), .B(n5182), .ZN(n5207) );
  XNOR2_X1 U5551 ( .A(n5183), .B(n5182), .ZN(n5191) );
  OAI22_X1 U5552 ( .A1(n5187), .A2(n5186), .B1(n5185), .B2(n5184), .ZN(n5188)
         );
  AOI21_X1 U5553 ( .B1(n5197), .B2(n5396), .A(n5188), .ZN(n5189) );
  OAI21_X1 U5554 ( .B1(n5191), .B2(n5190), .A(n5189), .ZN(n5192) );
  AOI21_X1 U5555 ( .B1(n5193), .B2(n5207), .A(n5192), .ZN(n5210) );
  INV_X1 U5556 ( .A(n5194), .ZN(n5195) );
  AOI21_X1 U5557 ( .B1(n5197), .B2(n5196), .A(n5195), .ZN(n5205) );
  AOI22_X1 U5558 ( .A1(n5207), .A2(n5198), .B1(n5406), .B2(n5205), .ZN(n5199)
         );
  AND2_X1 U5559 ( .A1(n5210), .A2(n5199), .ZN(n5202) );
  INV_X1 U5560 ( .A(REG1_REG_3__SCAN_IN), .ZN(n5200) );
  AOI22_X1 U5561 ( .A1(n5410), .A2(n5202), .B1(n5200), .B2(n5408), .ZN(U3521)
         );
  INV_X1 U5562 ( .A(REG0_REG_3__SCAN_IN), .ZN(n5201) );
  AOI22_X1 U5563 ( .A1(n5414), .A2(n5202), .B1(n5201), .B2(n5411), .ZN(U3473)
         );
  AOI22_X1 U5564 ( .A1(n5419), .A2(REG2_REG_3__SCAN_IN), .B1(n5204), .B2(n5203), .ZN(n5209) );
  AOI22_X1 U5565 ( .A1(n5207), .A2(n5206), .B1(n5415), .B2(n5205), .ZN(n5208)
         );
  OAI211_X1 U5566 ( .C1(n5419), .C2(n5210), .A(n5209), .B(n5208), .ZN(U3287)
         );
  AOI211_X1 U5567 ( .C1(n5213), .C2(n5392), .A(n5212), .B(n5211), .ZN(n5216)
         );
  AOI22_X1 U5568 ( .A1(n5410), .A2(n5216), .B1(n5214), .B2(n5408), .ZN(U3522)
         );
  INV_X1 U5569 ( .A(REG0_REG_4__SCAN_IN), .ZN(n5215) );
  AOI22_X1 U5570 ( .A1(n5414), .A2(n5216), .B1(n5215), .B2(n5411), .ZN(U3475)
         );
  AOI22_X1 U5571 ( .A1(STATE_REG_SCAN_IN), .A2(n5218), .B1(n5217), .B2(U3149), 
        .ZN(U3347) );
  OAI21_X1 U5572 ( .B1(n5390), .B2(n5220), .A(n5219), .ZN(n5221) );
  AOI21_X1 U5573 ( .B1(n5222), .B2(n5392), .A(n5221), .ZN(n5224) );
  AOI22_X1 U5574 ( .A1(n5410), .A2(n5224), .B1(n2837), .B2(n5408), .ZN(U3523)
         );
  INV_X1 U5575 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5223) );
  AOI22_X1 U5576 ( .A1(n5414), .A2(n5224), .B1(n5223), .B2(n5411), .ZN(U3477)
         );
  OAI22_X1 U5577 ( .A1(U3149), .A2(n5225), .B1(DATAI_6_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5226) );
  INV_X1 U5578 ( .A(n5226), .ZN(U3346) );
  AOI21_X1 U5579 ( .B1(n3273), .B2(n5228), .A(n5227), .ZN(n5229) );
  AOI211_X1 U5580 ( .C1(n5406), .C2(n5231), .A(n5230), .B(n5229), .ZN(n5234)
         );
  INV_X1 U5581 ( .A(REG1_REG_6__SCAN_IN), .ZN(n5232) );
  AOI22_X1 U5582 ( .A1(n5410), .A2(n5234), .B1(n5232), .B2(n5408), .ZN(U3524)
         );
  INV_X1 U5583 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5233) );
  AOI22_X1 U5584 ( .A1(n5414), .A2(n5234), .B1(n5233), .B2(n5411), .ZN(U3479)
         );
  NOR2_X1 U5585 ( .A1(n5235), .A2(n5381), .ZN(n5238) );
  AOI211_X1 U5586 ( .C1(n5238), .C2(n5244), .A(n5237), .B(n5236), .ZN(n5241)
         );
  AOI22_X1 U5587 ( .A1(n5410), .A2(n5241), .B1(n5239), .B2(n5408), .ZN(U3525)
         );
  INV_X1 U5588 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5240) );
  AOI22_X1 U5589 ( .A1(n5414), .A2(n5241), .B1(n5240), .B2(n5411), .ZN(U3481)
         );
  AND2_X1 U5590 ( .A1(n5244), .A2(n5242), .ZN(n5246) );
  NAND2_X1 U5591 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  OAI21_X1 U5592 ( .B1(n5246), .B2(n4627), .A(n5245), .ZN(n5261) );
  INV_X1 U5593 ( .A(n5247), .ZN(n5249) );
  AOI211_X1 U5594 ( .C1(n5250), .C2(n5249), .A(n5390), .B(n5248), .ZN(n5259)
         );
  XNOR2_X1 U5595 ( .A(n5252), .B(n5251), .ZN(n5253) );
  NAND2_X1 U5596 ( .A1(n5253), .A2(n5333), .ZN(n5255) );
  OAI211_X1 U5597 ( .C1(n5330), .C2(n5256), .A(n5255), .B(n5254), .ZN(n5266)
         );
  AOI211_X1 U5598 ( .C1(n5392), .C2(n5261), .A(n5259), .B(n5266), .ZN(n5258)
         );
  AOI22_X1 U5599 ( .A1(n5410), .A2(n5258), .B1(n3232), .B2(n5408), .ZN(U3526)
         );
  INV_X1 U5600 ( .A(REG0_REG_8__SCAN_IN), .ZN(n5257) );
  AOI22_X1 U5601 ( .A1(n5414), .A2(n5258), .B1(n5257), .B2(n5411), .ZN(U3483)
         );
  INV_X1 U5602 ( .A(n5259), .ZN(n5264) );
  NAND2_X1 U5603 ( .A1(n5261), .A2(n5260), .ZN(n5263) );
  OAI211_X1 U5604 ( .C1(n5265), .C2(n5264), .A(n5263), .B(n5262), .ZN(n5267)
         );
  OAI22_X1 U5605 ( .A1(n5267), .A2(n5266), .B1(REG2_REG_8__SCAN_IN), .B2(n5262), .ZN(n5268) );
  OAI21_X1 U5606 ( .B1(n5269), .B2(n5339), .A(n5268), .ZN(U3282) );
  AOI22_X1 U5607 ( .A1(STATE_REG_SCAN_IN), .A2(n5271), .B1(n5270), .B2(U3149), 
        .ZN(U3343) );
  NAND3_X1 U5608 ( .A1(n5273), .A2(n5406), .A3(n5272), .ZN(n5274) );
  OAI211_X1 U5609 ( .C1(n5276), .C2(n5381), .A(n5275), .B(n5274), .ZN(n5277)
         );
  INV_X1 U5610 ( .A(n5277), .ZN(n5280) );
  INV_X1 U5611 ( .A(REG1_REG_9__SCAN_IN), .ZN(n5278) );
  AOI22_X1 U5612 ( .A1(n5410), .A2(n5280), .B1(n5278), .B2(n5408), .ZN(U3527)
         );
  INV_X1 U5613 ( .A(REG0_REG_9__SCAN_IN), .ZN(n5279) );
  AOI22_X1 U5614 ( .A1(n5414), .A2(n5280), .B1(n5279), .B2(n5411), .ZN(U3485)
         );
  AOI22_X1 U5615 ( .A1(STATE_REG_SCAN_IN), .A2(n3428), .B1(n5281), .B2(U3149), 
        .ZN(U3342) );
  OAI22_X1 U5616 ( .A1(n5283), .A2(n5381), .B1(n5282), .B2(n5390), .ZN(n5285)
         );
  NOR2_X1 U5617 ( .A1(n5285), .A2(n5284), .ZN(n5288) );
  INV_X1 U5618 ( .A(REG1_REG_10__SCAN_IN), .ZN(n5286) );
  AOI22_X1 U5619 ( .A1(n5410), .A2(n5288), .B1(n5286), .B2(n5408), .ZN(U3528)
         );
  INV_X1 U5620 ( .A(REG0_REG_10__SCAN_IN), .ZN(n5287) );
  AOI22_X1 U5621 ( .A1(n5414), .A2(n5288), .B1(n5287), .B2(n5411), .ZN(U3487)
         );
  NOR2_X1 U5622 ( .A1(n5289), .A2(n5390), .ZN(n5291) );
  AOI211_X1 U5623 ( .C1(n5292), .C2(n5392), .A(n5291), .B(n5290), .ZN(n5295)
         );
  INV_X1 U5624 ( .A(REG1_REG_11__SCAN_IN), .ZN(n5293) );
  AOI22_X1 U5625 ( .A1(n5410), .A2(n5295), .B1(n5293), .B2(n5408), .ZN(U3529)
         );
  INV_X1 U5626 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5294) );
  AOI22_X1 U5627 ( .A1(n5414), .A2(n5295), .B1(n5294), .B2(n5411), .ZN(U3489)
         );
  AOI211_X1 U5628 ( .C1(n5298), .C2(n5392), .A(n5297), .B(n5296), .ZN(n5301)
         );
  INV_X1 U5629 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5299) );
  AOI22_X1 U5630 ( .A1(n5410), .A2(n5301), .B1(n5299), .B2(n5408), .ZN(U3530)
         );
  INV_X1 U5631 ( .A(REG0_REG_12__SCAN_IN), .ZN(n5300) );
  AOI22_X1 U5632 ( .A1(n5414), .A2(n5301), .B1(n5300), .B2(n5411), .ZN(U3491)
         );
  NAND2_X1 U5633 ( .A1(n5303), .A2(n5302), .ZN(n5307) );
  NAND2_X1 U5634 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  AND2_X1 U5635 ( .A1(n5307), .A2(n5306), .ZN(n5329) );
  INV_X1 U5636 ( .A(n5308), .ZN(n5309) );
  OAI21_X1 U5637 ( .B1(n5329), .B2(n5310), .A(n5309), .ZN(n5319) );
  INV_X1 U5638 ( .A(n5311), .ZN(n5312) );
  NAND3_X1 U5639 ( .A1(n5314), .A2(n5313), .A3(n5312), .ZN(n5316) );
  AOI21_X1 U5640 ( .B1(n5317), .B2(n5316), .A(n5315), .ZN(n5318) );
  AOI211_X1 U5641 ( .C1(n5320), .C2(n5364), .A(n5319), .B(n5318), .ZN(n5321)
         );
  OAI21_X1 U5642 ( .B1(n5340), .B2(n5370), .A(n5321), .ZN(U3231) );
  XOR2_X1 U5643 ( .A(n5327), .B(n5322), .Z(n5346) );
  OAI21_X1 U5644 ( .B1(n5324), .B2(n5331), .A(n5323), .ZN(n5343) );
  NAND2_X1 U5645 ( .A1(n5326), .A2(n5325), .ZN(n5328) );
  XNOR2_X1 U5646 ( .A(n5328), .B(n5327), .ZN(n5334) );
  OAI21_X1 U5647 ( .B1(n5331), .B2(n5330), .A(n5329), .ZN(n5332) );
  AOI21_X1 U5648 ( .B1(n5334), .B2(n5333), .A(n5332), .ZN(n5349) );
  OAI21_X1 U5649 ( .B1(n5390), .B2(n5343), .A(n5349), .ZN(n5335) );
  AOI21_X1 U5650 ( .B1(n5346), .B2(n5392), .A(n5335), .ZN(n5338) );
  INV_X1 U5651 ( .A(REG1_REG_13__SCAN_IN), .ZN(n5336) );
  AOI22_X1 U5652 ( .A1(n5410), .A2(n5338), .B1(n5336), .B2(n5408), .ZN(U3531)
         );
  INV_X1 U5653 ( .A(REG0_REG_13__SCAN_IN), .ZN(n5337) );
  AOI22_X1 U5654 ( .A1(n5414), .A2(n5338), .B1(n5337), .B2(n5411), .ZN(U3493)
         );
  OAI22_X1 U5655 ( .A1(n4140), .A2(n5341), .B1(n5340), .B2(n5339), .ZN(n5342)
         );
  INV_X1 U5656 ( .A(n5342), .ZN(n5348) );
  INV_X1 U5657 ( .A(n5343), .ZN(n5344) );
  AOI22_X1 U5658 ( .A1(n5346), .A2(n5345), .B1(n5415), .B2(n5344), .ZN(n5347)
         );
  OAI211_X1 U5659 ( .C1(n5419), .C2(n5349), .A(n5348), .B(n5347), .ZN(U3277)
         );
  OAI22_X1 U5660 ( .A1(n5351), .A2(n5381), .B1(n5390), .B2(n5350), .ZN(n5352)
         );
  NOR2_X1 U5661 ( .A1(n5353), .A2(n5352), .ZN(n5355) );
  AOI22_X1 U5662 ( .A1(n5410), .A2(n5355), .B1(n4168), .B2(n5408), .ZN(U3532)
         );
  INV_X1 U5663 ( .A(REG0_REG_14__SCAN_IN), .ZN(n5354) );
  AOI22_X1 U5664 ( .A1(n5414), .A2(n5355), .B1(n5354), .B2(n5411), .ZN(U3495)
         );
  AOI22_X1 U5665 ( .A1(STATE_REG_SCAN_IN), .A2(n5357), .B1(n5356), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5666 ( .A1(n5359), .A2(n5358), .B1(REG3_REG_15__SCAN_IN), .B2(
        U3149), .ZN(n5369) );
  NAND2_X1 U5667 ( .A1(n5361), .A2(n5360), .ZN(n5363) );
  XNOR2_X1 U5668 ( .A(n5363), .B(n5362), .ZN(n5367) );
  AOI22_X1 U5669 ( .A1(n5367), .A2(n5366), .B1(n5365), .B2(n5364), .ZN(n5368)
         );
  OAI211_X1 U5670 ( .C1(n5371), .C2(n5370), .A(n5369), .B(n5368), .ZN(U3238)
         );
  AOI211_X1 U5671 ( .C1(n5374), .C2(n5392), .A(n5373), .B(n5372), .ZN(n5377)
         );
  AOI22_X1 U5672 ( .A1(n5410), .A2(n5377), .B1(n5375), .B2(n5408), .ZN(U3533)
         );
  INV_X1 U5673 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5376) );
  AOI22_X1 U5674 ( .A1(n5414), .A2(n5377), .B1(n5376), .B2(n5411), .ZN(U3497)
         );
  AOI22_X1 U5675 ( .A1(STATE_REG_SCAN_IN), .A2(n5379), .B1(n5378), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5676 ( .A1(n5382), .A2(n5381), .B1(n5390), .B2(n5380), .ZN(n5383)
         );
  NOR2_X1 U5677 ( .A1(n5384), .A2(n5383), .ZN(n5387) );
  INV_X1 U5678 ( .A(REG1_REG_16__SCAN_IN), .ZN(n5385) );
  AOI22_X1 U5679 ( .A1(n5410), .A2(n5387), .B1(n5385), .B2(n5408), .ZN(U3534)
         );
  INV_X1 U5680 ( .A(REG0_REG_16__SCAN_IN), .ZN(n5386) );
  AOI22_X1 U5681 ( .A1(n5414), .A2(n5387), .B1(n5386), .B2(n5411), .ZN(U3499)
         );
  OAI21_X1 U5682 ( .B1(n5390), .B2(n5389), .A(n5388), .ZN(n5391) );
  AOI21_X1 U5683 ( .B1(n5393), .B2(n5392), .A(n5391), .ZN(n5395) );
  AOI22_X1 U5684 ( .A1(n5410), .A2(n5395), .B1(n4302), .B2(n5408), .ZN(U3535)
         );
  INV_X1 U5685 ( .A(REG0_REG_17__SCAN_IN), .ZN(n5394) );
  AOI22_X1 U5686 ( .A1(n5414), .A2(n5395), .B1(n5394), .B2(n5411), .ZN(U3501)
         );
  NAND2_X1 U5687 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  AND2_X1 U5688 ( .A1(n5399), .A2(n5398), .ZN(n5404) );
  XNOR2_X1 U5689 ( .A(n5401), .B(n5400), .ZN(n5407) );
  AOI22_X1 U5690 ( .A1(n5407), .A2(n5415), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5402), .ZN(n5403) );
  OAI21_X1 U5691 ( .B1(n5419), .B2(n5404), .A(n5403), .ZN(U3261) );
  INV_X1 U5692 ( .A(n5404), .ZN(n5405) );
  AOI21_X1 U5693 ( .B1(n5407), .B2(n5406), .A(n5405), .ZN(n5413) );
  INV_X1 U5694 ( .A(REG1_REG_30__SCAN_IN), .ZN(n5409) );
  AOI22_X1 U5695 ( .A1(n5410), .A2(n5413), .B1(n5409), .B2(n5408), .ZN(U3548)
         );
  INV_X1 U5696 ( .A(REG0_REG_30__SCAN_IN), .ZN(n5412) );
  AOI22_X1 U5697 ( .A1(n5414), .A2(n5413), .B1(n5412), .B2(n5411), .ZN(U3516)
         );
  AOI22_X1 U5698 ( .A1(n5416), .A2(n5415), .B1(n5419), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5417) );
  OAI21_X1 U5699 ( .B1(n5419), .B2(n5418), .A(n5417), .ZN(U3260) );
endmodule

