

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10980, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11013,
         n11014, n11015, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398;

  NAND2_X1 U11087 ( .A1(n11403), .A2(n12204), .ZN(n16057) );
  BUF_X2 U11088 ( .A(n18768), .Z(n11029) );
  AND2_X1 U11089 ( .A1(n13779), .A2(n13778), .ZN(n21810) );
  NOR2_X1 U11090 ( .A1(n16033), .A2(n16035), .ZN(n13800) );
  AND2_X1 U11091 ( .A1(n13748), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14789)
         );
  INV_X1 U11092 ( .A(n14167), .ZN(n14171) );
  INV_X2 U11093 ( .A(n11028), .ZN(n14857) );
  NAND2_X1 U11094 ( .A1(n14527), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14526) );
  INV_X1 U11095 ( .A(n14081), .ZN(n15510) );
  CLKBUF_X2 U11096 ( .A(n11620), .Z(n10992) );
  INV_X1 U11097 ( .A(n15484), .ZN(n15504) );
  INV_X1 U11098 ( .A(n14462), .ZN(n15512) );
  CLKBUF_X2 U11099 ( .A(n11549), .Z(n17727) );
  CLKBUF_X2 U11100 ( .A(n11621), .Z(n17928) );
  CLKBUF_X2 U11101 ( .A(n11620), .Z(n17803) );
  AND2_X2 U11102 ( .A1(n15520), .A2(n12448), .ZN(n15486) );
  AND2_X2 U11103 ( .A1(n15520), .A2(n14613), .ZN(n15485) );
  BUF_X2 U11104 ( .A(n11644), .Z(n17950) );
  INV_X1 U11105 ( .A(n17690), .ZN(n17940) );
  BUF_X1 U11106 ( .A(n11690), .Z(n17948) );
  CLKBUF_X2 U11108 ( .A(n11991), .Z(n13699) );
  NOR2_X1 U11109 ( .A1(n11944), .A2(n11925), .ZN(n11935) );
  INV_X1 U11110 ( .A(n14193), .ZN(n19720) );
  CLKBUF_X1 U11111 ( .A(n12679), .Z(n19562) );
  BUF_X1 U11112 ( .A(n12628), .Z(n12700) );
  CLKBUF_X1 U11113 ( .A(n11932), .Z(n14689) );
  BUF_X1 U11114 ( .A(n11929), .Z(n11027) );
  AND4_X1 U11115 ( .A1(n11844), .A2(n11843), .A3(n11842), .A4(n11841), .ZN(
        n11845) );
  INV_X1 U11116 ( .A(n11931), .ZN(n10993) );
  OR2_X1 U11117 ( .A1(n11835), .A2(n11836), .ZN(n11931) );
  BUF_X2 U11118 ( .A(n11903), .Z(n11030) );
  AND2_X1 U11119 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14584) );
  NAND2_X1 U11120 ( .A1(n12135), .A2(n21496), .ZN(n10982) );
  NAND2_X1 U11121 ( .A1(n10980), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10983) );
  NAND2_X1 U11122 ( .A1(n10982), .A2(n10983), .ZN(n20153) );
  INV_X1 U11123 ( .A(n12135), .ZN(n10980) );
  BUF_X1 U11125 ( .A(n16105), .Z(n10984) );
  INV_X1 U11127 ( .A(n15026), .ZN(n10986) );
  NOR2_X1 U11128 ( .A1(n14712), .A2(n10993), .ZN(n11915) );
  NAND2_X1 U11129 ( .A1(n11846), .A2(n11845), .ZN(n14712) );
  XNOR2_X1 U11130 ( .A(n11990), .B(n11989), .ZN(n13265) );
  NOR2_X1 U11131 ( .A1(n14195), .A2(n12709), .ZN(n12730) );
  BUF_X1 U11134 ( .A(n11904), .Z(n13636) );
  NOR2_X1 U11136 ( .A1(n11493), .A2(n11492), .ZN(n11691) );
  NAND2_X1 U11137 ( .A1(n12291), .A2(n11027), .ZN(n12381) );
  OAI21_X1 U11138 ( .B1(n17459), .B2(n18604), .A(n16947), .ZN(n16735) );
  NOR2_X1 U11139 ( .A1(n12779), .A2(n12784), .ZN(n12831) );
  CLKBUF_X2 U11140 ( .A(n11690), .Z(n17783) );
  INV_X1 U11141 ( .A(n17649), .ZN(n17927) );
  AND2_X1 U11142 ( .A1(n18011), .A2(n21314), .ZN(n17989) );
  AND2_X1 U11143 ( .A1(n11281), .A2(n10998), .ZN(n11717) );
  AND2_X1 U11144 ( .A1(n21002), .A2(n21010), .ZN(n20988) );
  INV_X2 U11145 ( .A(n20409), .ZN(n11632) );
  OR2_X1 U11146 ( .A1(n15750), .A2(n11458), .ZN(n13728) );
  AND2_X1 U11147 ( .A1(n12064), .A2(n12063), .ZN(n15104) );
  NOR2_X1 U11148 ( .A1(n16694), .A2(n16308), .ZN(n16311) );
  AND2_X1 U11149 ( .A1(n16512), .A2(n11112), .ZN(n16490) );
  AND2_X1 U11150 ( .A1(n12602), .A2(n12601), .ZN(n16730) );
  INV_X2 U11151 ( .A(n18768), .ZN(n18783) );
  NOR3_X2 U11152 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n13191), .A3(
        n13190), .ZN(n13819) );
  INV_X1 U11153 ( .A(n21795), .ZN(n21816) );
  AOI211_X1 U11154 ( .C1(n14694), .C2(n15382), .A(n15007), .B(n15006), .ZN(
        n21828) );
  AND2_X1 U11155 ( .A1(n14444), .A2(n14470), .ZN(n14467) );
  OAI211_X1 U11156 ( .C1(n17459), .C2(n18622), .A(n16711), .B(n16925), .ZN(
        n16713) );
  AOI21_X1 U11157 ( .B1(n16576), .B2(n11331), .A(n11330), .ZN(n11329) );
  NAND2_X1 U11158 ( .A1(n16939), .A2(n16662), .ZN(n16709) );
  AOI221_X1 U11159 ( .B1(n11029), .B2(n18462), .C1(n18783), .C2(n17048), .A(
        n18890), .ZN(n17071) );
  INV_X1 U11160 ( .A(n19220), .ZN(n20779) );
  INV_X1 U11161 ( .A(n20809), .ZN(n20959) );
  NOR2_X1 U11162 ( .A1(n18346), .A2(n18318), .ZN(n18152) );
  NOR2_X2 U11163 ( .A1(n18002), .A2(n21122), .ZN(n21135) );
  XNOR2_X1 U11164 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13860), .ZN(
        n10987) );
  NAND2_X2 U11165 ( .A1(n14454), .A2(n14619), .ZN(n15687) );
  XNOR2_X2 U11166 ( .A(n16325), .B(n16338), .ZN(n16570) );
  OAI211_X2 U11167 ( .C1(n13171), .C2(n13167), .A(n11214), .B(n13170), .ZN(
        n11215) );
  AND2_X1 U11168 ( .A1(n11823), .A2(n11818), .ZN(n10988) );
  AND2_X1 U11169 ( .A1(n11823), .A2(n11818), .ZN(n10989) );
  NOR2_X2 U11170 ( .A1(n20623), .A2(n11802), .ZN(n20658) );
  INV_X2 U11171 ( .A(n15031), .ZN(n14197) );
  NAND2_X2 U11172 ( .A1(n12675), .A2(n12674), .ZN(n15031) );
  OAI21_X2 U11173 ( .B1(n16709), .B2(n16663), .A(n16708), .ZN(n16689) );
  NOR2_X2 U11174 ( .A1(n13836), .A2(n21234), .ZN(n21244) );
  NOR2_X2 U11175 ( .A1(n16414), .A2(n11471), .ZN(n15646) );
  NOR2_X2 U11176 ( .A1(n16413), .A2(n16415), .ZN(n16414) );
  NOR3_X2 U11177 ( .A1(n11039), .A2(n11376), .A3(n16902), .ZN(n11374) );
  BUF_X1 U11178 ( .A(n21284), .Z(n10990) );
  NAND3_X2 U11179 ( .A1(n11587), .A2(n11586), .A3(n11585), .ZN(n20809) );
  NOR2_X2 U11180 ( .A1(n12779), .A2(n12781), .ZN(n12842) );
  NAND2_X1 U11182 ( .A1(n11859), .A2(n11858), .ZN(n11920) );
  AOI21_X4 U11183 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18152), .A(
        n19264), .ZN(n18132) );
  AND2_X1 U11184 ( .A1(n11452), .A2(n11822), .ZN(n10991) );
  AND2_X1 U11185 ( .A1(n11452), .A2(n11822), .ZN(n11904) );
  NOR2_X2 U11186 ( .A1(n18027), .A2(n11286), .ZN(n18221) );
  AND2_X1 U11187 ( .A1(n13183), .A2(n11122), .ZN(n16612) );
  OAI21_X1 U11188 ( .B1(n18143), .B2(n11296), .A(n11295), .ZN(n18124) );
  NOR2_X1 U11189 ( .A1(n11050), .A2(n16451), .ZN(n16452) );
  NOR2_X1 U11190 ( .A1(n11392), .A2(n16155), .ZN(n11391) );
  NOR2_X1 U11191 ( .A1(n20671), .A2(n20670), .ZN(n20697) );
  INV_X1 U11192 ( .A(n18180), .ZN(n18171) );
  INV_X1 U11193 ( .A(n12179), .ZN(n12193) );
  OR2_X1 U11194 ( .A1(n12827), .A2(n12826), .ZN(n11165) );
  NOR2_X1 U11195 ( .A1(n13002), .A2(n13001), .ZN(n13007) );
  INV_X2 U11196 ( .A(n21268), .ZN(n21384) );
  AND2_X1 U11197 ( .A1(n14432), .A2(n14431), .ZN(n14433) );
  OR2_X2 U11198 ( .A1(n14740), .A2(n14749), .ZN(n14807) );
  NAND2_X1 U11199 ( .A1(n21019), .A2(n13195), .ZN(n21321) );
  INV_X2 U11200 ( .A(n16448), .ZN(n16433) );
  OAI21_X1 U11201 ( .B1(n13264), .B2(n12134), .A(n12106), .ZN(n14527) );
  AND2_X1 U11202 ( .A1(n12738), .A2(n12720), .ZN(n12762) );
  OAI211_X1 U11203 ( .C1(n13124), .C2(n16366), .A(n12755), .B(n12754), .ZN(
        n13038) );
  INV_X2 U11204 ( .A(n13892), .ZN(n11350) );
  CLKBUF_X3 U11205 ( .A(n13047), .Z(n14180) );
  NAND2_X1 U11206 ( .A1(n11609), .A2(n20841), .ZN(n20787) );
  NAND2_X2 U11207 ( .A1(n11367), .A2(n11028), .ZN(n14150) );
  NOR2_X1 U11208 ( .A1(n14749), .A2(n11929), .ZN(n11947) );
  NAND3_X1 U11209 ( .A1(n19671), .A2(n12687), .A3(n12700), .ZN(n12706) );
  INV_X1 U11210 ( .A(n12700), .ZN(n12873) );
  CLKBUF_X1 U11211 ( .A(n11924), .Z(n11023) );
  INV_X4 U11212 ( .A(n13931), .ZN(n15667) );
  NAND4_X1 U11213 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11929) );
  INV_X4 U11214 ( .A(n17906), .ZN(n17939) );
  CLKBUF_X2 U11215 ( .A(n17588), .Z(n17943) );
  CLKBUF_X2 U11216 ( .A(n11549), .Z(n17942) );
  CLKBUF_X2 U11217 ( .A(n20053), .Z(n21456) );
  CLKBUF_X2 U11218 ( .A(n11992), .Z(n13680) );
  CLKBUF_X2 U11219 ( .A(n12055), .Z(n13701) );
  INV_X1 U11221 ( .A(n14057), .ZN(n15511) );
  INV_X1 U11222 ( .A(n14078), .ZN(n15508) );
  CLKBUF_X1 U11223 ( .A(n11035), .Z(n11034) );
  BUF_X2 U11224 ( .A(n11958), .Z(n13707) );
  BUF_X2 U11225 ( .A(n11973), .Z(n13709) );
  BUF_X2 U11226 ( .A(n11959), .Z(n13702) );
  CLKBUF_X2 U11227 ( .A(n11998), .Z(n12056) );
  BUF_X2 U11228 ( .A(n11978), .Z(n13502) );
  INV_X1 U11229 ( .A(n17572), .ZN(n21882) );
  INV_X1 U11230 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20991) );
  INV_X2 U11231 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12023) );
  INV_X4 U11232 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12648) );
  AOI21_X1 U11233 ( .B1(n11373), .B2(n18825), .A(n11368), .ZN(n16770) );
  NAND2_X1 U11234 ( .A1(n11172), .A2(n11171), .ZN(n13851) );
  OR2_X1 U11235 ( .A1(n13186), .A2(n16584), .ZN(n16769) );
  NAND2_X1 U11236 ( .A1(n11175), .A2(n11173), .ZN(n11172) );
  OAI21_X1 U11237 ( .B1(n16571), .B2(n17463), .A(n11221), .ZN(n11220) );
  NOR2_X1 U11238 ( .A1(n16605), .A2(n13185), .ZN(n16584) );
  AOI21_X1 U11239 ( .B1(n16689), .B2(n16666), .A(n16665), .ZN(n16668) );
  XNOR2_X1 U11240 ( .A(n13728), .B(n13727), .ZN(n13790) );
  NAND2_X1 U11241 ( .A1(n12200), .A2(n12199), .ZN(n12201) );
  AND2_X1 U11243 ( .A1(n13183), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16734) );
  NAND2_X1 U11244 ( .A1(n11178), .A2(n11176), .ZN(n12992) );
  AND2_X2 U11245 ( .A1(n16739), .A2(n16921), .ZN(n13183) );
  NOR2_X1 U11246 ( .A1(n16112), .A2(n16113), .ZN(n16111) );
  NAND2_X1 U11248 ( .A1(n11341), .A2(n11340), .ZN(n16648) );
  NAND2_X1 U11249 ( .A1(n11149), .A2(n11183), .ZN(n16739) );
  AOI211_X1 U11250 ( .C1(n16289), .C2(n18796), .A(n16343), .B(n16342), .ZN(
        n16344) );
  AOI21_X1 U11251 ( .B1(n11184), .B2(n11186), .A(n11071), .ZN(n11183) );
  AOI21_X1 U11252 ( .B1(n11167), .B2(n11169), .A(n11090), .ZN(n11166) );
  NOR2_X1 U11253 ( .A1(n18124), .A2(n21381), .ZN(n13223) );
  XNOR2_X1 U11254 ( .A(n15702), .B(n14173), .ZN(n16341) );
  AND2_X1 U11255 ( .A1(n12914), .A2(n11089), .ZN(n11169) );
  OAI21_X1 U11256 ( .B1(n15314), .B2(n11186), .A(n17431), .ZN(n11185) );
  AND2_X1 U11257 ( .A1(n11201), .A2(n11076), .ZN(n11203) );
  INV_X1 U11258 ( .A(n13177), .ZN(n11186) );
  AND2_X1 U11259 ( .A1(n11201), .A2(n11060), .ZN(n11205) );
  NOR2_X1 U11260 ( .A1(n13189), .A2(n13192), .ZN(n13818) );
  NAND2_X1 U11261 ( .A1(n20165), .A2(n11397), .ZN(n20174) );
  NAND2_X1 U11262 ( .A1(n20164), .A2(n20166), .ZN(n20165) );
  OAI211_X1 U11263 ( .C1(n11238), .C2(n13859), .A(n11235), .B(n11233), .ZN(
        n12913) );
  NAND2_X1 U11264 ( .A1(n20158), .A2(n12145), .ZN(n20164) );
  NAND2_X1 U11265 ( .A1(n11234), .A2(n16730), .ZN(n11233) );
  NOR2_X1 U11267 ( .A1(n15347), .A2(n15348), .ZN(n16471) );
  OR2_X1 U11268 ( .A1(n10987), .A2(n11336), .ZN(n11335) );
  AOI21_X1 U11269 ( .B1(n15289), .B2(n11020), .A(n11069), .ZN(n11393) );
  NAND2_X1 U11270 ( .A1(n18119), .A2(n21283), .ZN(n18118) );
  OR2_X1 U11271 ( .A1(n13174), .A2(n13173), .ZN(n13178) );
  OR2_X1 U11272 ( .A1(n13014), .A2(n11059), .ZN(n11171) );
  AOI21_X1 U11273 ( .B1(n13161), .B2(n11231), .A(n11236), .ZN(n11235) );
  AND2_X1 U11274 ( .A1(n12177), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11020) );
  INV_X1 U11275 ( .A(n11764), .ZN(n18049) );
  AND2_X1 U11276 ( .A1(n13168), .A2(n16730), .ZN(n11231) );
  OR2_X1 U11277 ( .A1(n11801), .A2(n20586), .ZN(n20623) );
  OR2_X1 U11278 ( .A1(n12906), .A2(n12905), .ZN(n12909) );
  NOR2_X1 U11279 ( .A1(n19440), .A2(n19421), .ZN(n19882) );
  NOR2_X1 U11280 ( .A1(n13250), .A2(n14885), .ZN(n13275) );
  AND2_X1 U11281 ( .A1(n11756), .A2(n21330), .ZN(n11279) );
  AND4_X1 U11282 ( .A1(n12839), .A2(n12838), .A3(n12837), .A4(n12836), .ZN(
        n12856) );
  OR2_X1 U11283 ( .A1(n12815), .A2(n12814), .ZN(n11164) );
  OAI211_X1 U11284 ( .C1(n11747), .C2(n11746), .A(n11745), .B(n11744), .ZN(
        n18249) );
  INV_X1 U11285 ( .A(n12147), .ZN(n11453) );
  AND2_X1 U11286 ( .A1(n13007), .A2(n13006), .ZN(n13853) );
  OAI21_X1 U11287 ( .B1(n15107), .B2(n13373), .A(n13238), .ZN(n14727) );
  CLKBUF_X1 U11288 ( .A(n13750), .Z(n16008) );
  CLKBUF_X1 U11289 ( .A(n15957), .Z(n16010) );
  XNOR2_X1 U11290 ( .A(n12138), .B(n12137), .ZN(n13249) );
  NAND2_X1 U11291 ( .A1(n12138), .A2(n12130), .ZN(n15107) );
  NOR2_X1 U11292 ( .A1(n18026), .A2(n11753), .ZN(n18001) );
  OR2_X1 U11293 ( .A1(n12995), .A2(n12993), .ZN(n13002) );
  INV_X1 U11294 ( .A(n12835), .ZN(n19417) );
  CLKBUF_X1 U11295 ( .A(n12840), .Z(n14852) );
  CLKBUF_X1 U11296 ( .A(n12849), .Z(n17377) );
  CLKBUF_X1 U11297 ( .A(n13251), .Z(n15105) );
  NOR2_X1 U11298 ( .A1(n20968), .A2(n20841), .ZN(n20938) );
  NAND2_X2 U11299 ( .A1(n16015), .A2(n14483), .ZN(n16023) );
  NAND2_X1 U11300 ( .A1(n20136), .A2(n14683), .ZN(n15954) );
  NAND2_X1 U11301 ( .A1(n20778), .A2(n20369), .ZN(n17094) );
  AND2_X1 U11302 ( .A1(n16321), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16323) );
  NAND2_X1 U11303 ( .A1(n12114), .A2(n12113), .ZN(n12115) );
  NAND2_X1 U11304 ( .A1(n18279), .A2(n11742), .ZN(n18272) );
  NOR2_X2 U11305 ( .A1(n21321), .A2(n21386), .ZN(n21285) );
  NOR2_X2 U11306 ( .A1(n16319), .A2(n18740), .ZN(n16321) );
  NOR2_X2 U11307 ( .A1(n21380), .A2(n20322), .ZN(n20369) );
  OR2_X2 U11308 ( .A1(n16317), .A2(n16614), .ZN(n16319) );
  NAND2_X1 U11309 ( .A1(n14428), .A2(n14427), .ZN(n14447) );
  XNOR2_X1 U11310 ( .A(n11741), .B(n11195), .ZN(n18280) );
  OR2_X1 U11311 ( .A1(n12980), .A2(n12979), .ZN(n12985) );
  INV_X1 U11312 ( .A(n12767), .ZN(n12781) );
  NAND2_X1 U11313 ( .A1(n11200), .A2(n11971), .ZN(n12014) );
  NOR2_X2 U11314 ( .A1(n19394), .A2(n19869), .ZN(n14988) );
  NOR2_X2 U11315 ( .A1(n19816), .A2(n19869), .ZN(n17376) );
  NAND2_X1 U11316 ( .A1(n12021), .A2(n12020), .ZN(n12029) );
  NAND2_X1 U11317 ( .A1(n13979), .A2(n13978), .ZN(n15242) );
  XNOR2_X1 U11318 ( .A(n12104), .B(n12103), .ZN(n13264) );
  NAND2_X1 U11319 ( .A1(n12008), .A2(n12007), .ZN(n12104) );
  INV_X1 U11320 ( .A(n12764), .ZN(n12763) );
  AND2_X1 U11321 ( .A1(n12750), .A2(n12749), .ZN(n12756) );
  INV_X2 U11322 ( .A(n20324), .ZN(n20366) );
  OR2_X1 U11323 ( .A1(n12747), .A2(n12748), .ZN(n12750) );
  INV_X1 U11324 ( .A(n18507), .ZN(n11236) );
  XNOR2_X1 U11325 ( .A(n13038), .B(n13039), .ZN(n11230) );
  NAND2_X1 U11326 ( .A1(n18311), .A2(n11735), .ZN(n11737) );
  OR2_X1 U11327 ( .A1(n14920), .A2(n14919), .ZN(n15116) );
  AND2_X1 U11328 ( .A1(n12694), .A2(n11427), .ZN(n11428) );
  AOI21_X1 U11329 ( .B1(n12739), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12751), .ZN(n13039) );
  INV_X2 U11330 ( .A(n10999), .ZN(n13124) );
  AND2_X1 U11331 ( .A1(n11940), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12019) );
  AND3_X1 U11332 ( .A1(n11952), .A2(n11951), .A3(n11479), .ZN(n11953) );
  XNOR2_X1 U11333 ( .A(n13957), .B(n13956), .ZN(n14559) );
  OR2_X1 U11334 ( .A1(n12878), .A2(n12879), .ZN(n12881) );
  AND2_X1 U11335 ( .A1(n14561), .A2(n14560), .ZN(n13957) );
  NOR2_X1 U11336 ( .A1(n14728), .A2(n11318), .ZN(n11317) );
  NAND2_X1 U11337 ( .A1(n16427), .A2(n11440), .ZN(n11439) );
  NAND2_X1 U11338 ( .A1(n11396), .A2(n11395), .ZN(n12875) );
  NOR2_X1 U11339 ( .A1(n20840), .A2(n20841), .ZN(n13212) );
  AND2_X2 U11340 ( .A1(n14453), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13047) );
  AND2_X1 U11341 ( .A1(n14566), .A2(n12693), .ZN(n14453) );
  AND3_X2 U11342 ( .A1(n13899), .A2(n12652), .A3(n14193), .ZN(n12710) );
  CLKBUF_X1 U11343 ( .A(n12215), .Z(n17146) );
  AND2_X1 U11344 ( .A1(n12692), .A2(n12691), .ZN(n14566) );
  AND2_X1 U11345 ( .A1(n12684), .A2(n16279), .ZN(n11212) );
  AND2_X1 U11346 ( .A1(n12689), .A2(n12705), .ZN(n11133) );
  NAND2_X1 U11347 ( .A1(n11922), .A2(n11062), .ZN(n15380) );
  AND2_X1 U11348 ( .A1(n14392), .A2(n11927), .ZN(n12215) );
  OAI211_X1 U11349 ( .C1(n14145), .C2(n14307), .A(n13961), .B(n13947), .ZN(
        n14560) );
  NOR2_X1 U11350 ( .A1(n12388), .A2(n15876), .ZN(n14389) );
  NAND2_X1 U11351 ( .A1(n13861), .A2(n12681), .ZN(n16279) );
  AND2_X1 U11352 ( .A1(n12726), .A2(n19872), .ZN(n12709) );
  CLKBUF_X3 U11353 ( .A(n12873), .Z(n11028) );
  CLKBUF_X1 U11354 ( .A(n11947), .Z(n15876) );
  NOR2_X1 U11355 ( .A1(n17460), .A2(n16300), .ZN(n16303) );
  OR2_X1 U11356 ( .A1(n11554), .A2(n11150), .ZN(n17576) );
  AND2_X1 U11357 ( .A1(n11859), .A2(n13734), .ZN(n14392) );
  NAND2_X1 U11358 ( .A1(n19720), .A2(n14197), .ZN(n13897) );
  NAND2_X1 U11359 ( .A1(n13915), .A2(n12700), .ZN(n14145) );
  AND2_X1 U11360 ( .A1(n14683), .A2(n14689), .ZN(n13752) );
  INV_X1 U11361 ( .A(n13885), .ZN(n16277) );
  INV_X1 U11362 ( .A(n11929), .ZN(n11026) );
  NOR2_X1 U11363 ( .A1(n17441), .A2(n16298), .ZN(n16301) );
  AND2_X1 U11364 ( .A1(n12495), .A2(n12494), .ZN(n13962) );
  NOR2_X1 U11365 ( .A1(n14735), .A2(n11924), .ZN(n11930) );
  NAND2_X1 U11366 ( .A1(n11156), .A2(n11154), .ZN(n14193) );
  NAND2_X1 U11367 ( .A1(n11162), .A2(n11161), .ZN(n12699) );
  NAND2_X2 U11368 ( .A1(n12651), .A2(n12650), .ZN(n12687) );
  INV_X2 U11369 ( .A(n16336), .ZN(n19872) );
  NAND3_X1 U11370 ( .A1(n11826), .A2(n11825), .A3(n11824), .ZN(n11924) );
  NAND3_X1 U11371 ( .A1(n11856), .A2(n11485), .A3(n11053), .ZN(n11932) );
  NAND3_X1 U11372 ( .A1(n11869), .A2(n11487), .A3(n11868), .ZN(n14735) );
  INV_X2 U11373 ( .A(U212), .ZN(n10994) );
  NAND2_X2 U11374 ( .A1(n11914), .A2(n11486), .ZN(n14749) );
  AND4_X1 U11375 ( .A1(n11813), .A2(n11815), .A3(n11814), .A4(n11816), .ZN(
        n11826) );
  AND4_X1 U11376 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n11898) );
  AND4_X1 U11377 ( .A1(n11889), .A2(n11888), .A3(n11887), .A4(n11886), .ZN(
        n11900) );
  AND4_X1 U11378 ( .A1(n11893), .A2(n11892), .A3(n11891), .A4(n11890), .ZN(
        n11899) );
  AND4_X1 U11379 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11837), .ZN(
        n11846) );
  AND4_X1 U11380 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11856) );
  MUX2_X1 U11381 ( .A(n12473), .B(n12472), .S(n12648), .Z(n16336) );
  NAND2_X2 U11382 ( .A1(U214), .A2(n20243), .ZN(n20309) );
  AND4_X1 U11383 ( .A1(n11913), .A2(n11912), .A3(n11911), .A4(n11910), .ZN(
        n11914) );
  AND4_X1 U11384 ( .A1(n11885), .A2(n11884), .A3(n11883), .A4(n11882), .ZN(
        n11901) );
  INV_X2 U11385 ( .A(n14082), .ZN(n15509) );
  AND2_X1 U11386 ( .A1(n12613), .A2(n12612), .ZN(n12617) );
  AND2_X1 U11387 ( .A1(n12620), .A2(n12619), .ZN(n12624) );
  CLKBUF_X2 U11388 ( .A(n11972), .Z(n12054) );
  INV_X2 U11389 ( .A(n17690), .ZN(n17914) );
  BUF_X4 U11390 ( .A(n11547), .Z(n17907) );
  CLKBUF_X2 U11391 ( .A(n11903), .Z(n11031) );
  CLKBUF_X2 U11392 ( .A(n13637), .Z(n11037) );
  AND2_X2 U11393 ( .A1(n11002), .A2(n11817), .ZN(n11997) );
  AND2_X2 U11394 ( .A1(n11002), .A2(n14584), .ZN(n11992) );
  AND2_X2 U11395 ( .A1(n11002), .A2(n11015), .ZN(n12055) );
  CLKBUF_X1 U11396 ( .A(n11909), .Z(n13681) );
  INV_X2 U11397 ( .A(n21329), .ZN(n10995) );
  CLKBUF_X1 U11398 ( .A(n14361), .Z(n15697) );
  INV_X2 U11399 ( .A(n17816), .ZN(n17881) );
  NAND2_X1 U11400 ( .A1(n11197), .A2(n11196), .ZN(n17649) );
  NOR2_X1 U11401 ( .A1(n11493), .A2(n21005), .ZN(n11620) );
  BUF_X4 U11402 ( .A(n11537), .Z(n10996) );
  OR2_X2 U11403 ( .A1(n21004), .A2(n20368), .ZN(n17816) );
  OR2_X2 U11404 ( .A1(n21004), .A2(n11493), .ZN(n17690) );
  AND2_X2 U11405 ( .A1(n11817), .A2(n11822), .ZN(n11991) );
  AND2_X1 U11406 ( .A1(n12023), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11002) );
  AND2_X2 U11407 ( .A1(n11817), .A2(n15009), .ZN(n11958) );
  INV_X2 U11408 ( .A(n19986), .ZN(n20029) );
  NAND2_X1 U11409 ( .A1(n14604), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12441) );
  NAND2_X1 U11410 ( .A1(n21003), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11493) );
  NAND2_X1 U11411 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21029), .ZN(
        n11495) );
  AND2_X1 U11412 ( .A1(n15385), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11015) );
  AND2_X1 U11413 ( .A1(n15008), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11005) );
  AND2_X1 U11414 ( .A1(n15008), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11198) );
  AND2_X2 U11415 ( .A1(n14594), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11817) );
  AND2_X1 U11416 ( .A1(n15008), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11004) );
  AND2_X1 U11417 ( .A1(n15385), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11452) );
  NAND2_X1 U11418 ( .A1(n21029), .A2(n21394), .ZN(n21005) );
  NOR2_X1 U11419 ( .A1(n21872), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22398) );
  OR2_X2 U11420 ( .A1(n21862), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U11421 ( .A1(n20991), .A2(n21003), .ZN(n20368) );
  NAND2_X2 U11422 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20991), .ZN(
        n11494) );
  AND2_X1 U11423 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21013) );
  INV_X2 U11424 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21394) );
  NAND2_X1 U11425 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21004) );
  AND2_X2 U11426 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12447) );
  NOR2_X2 U11427 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11822) );
  AND2_X1 U11428 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15009) );
  OAI211_X1 U11429 ( .C1(n13171), .C2(n13167), .A(n11214), .B(n13170), .ZN(
        n10997) );
  NAND2_X1 U11430 ( .A1(n11391), .A2(n11394), .ZN(n11201) );
  AND2_X1 U11431 ( .A1(n14450), .A2(n14331), .ZN(n12782) );
  OR2_X1 U11432 ( .A1(n14450), .A2(n14426), .ZN(n12785) );
  OR2_X2 U11433 ( .A1(n14450), .A2(n14331), .ZN(n12779) );
  AND2_X1 U11434 ( .A1(n12782), .A2(n12775), .ZN(n19462) );
  AND2_X1 U11435 ( .A1(n12782), .A2(n12780), .ZN(n14985) );
  AND2_X1 U11436 ( .A1(n12782), .A2(n12767), .ZN(n19478) );
  AND2_X1 U11437 ( .A1(n12782), .A2(n12766), .ZN(n19446) );
  NOR2_X1 U11438 ( .A1(n12785), .A2(n12781), .ZN(n15170) );
  NOR2_X1 U11439 ( .A1(n12779), .A2(n12783), .ZN(n12829) );
  AND2_X1 U11440 ( .A1(n11484), .A2(n12767), .ZN(n12841) );
  AND2_X1 U11441 ( .A1(n11484), .A2(n12780), .ZN(n12843) );
  NAND2_X1 U11442 ( .A1(n11484), .A2(n12775), .ZN(n12835) );
  NAND2_X1 U11443 ( .A1(n11358), .A2(n12750), .ZN(n11320) );
  CLKBUF_X1 U11444 ( .A(n13642), .Z(n13708) );
  NAND2_X1 U11445 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11716), .ZN(
        n10998) );
  INV_X2 U11446 ( .A(n21311), .ZN(n21192) );
  NOR2_X1 U11447 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15008), .ZN(
        n11818) );
  AND2_X1 U11448 ( .A1(n11409), .A2(n12648), .ZN(n15520) );
  NAND2_X2 U11449 ( .A1(n12447), .A2(n11409), .ZN(n15650) );
  INV_X1 U11450 ( .A(n12743), .ZN(n10999) );
  NAND2_X4 U11451 ( .A1(n11350), .A2(n11064), .ZN(n12743) );
  NAND2_X1 U11452 ( .A1(n14405), .A2(n14404), .ZN(n14429) );
  NOR2_X2 U11453 ( .A1(n12985), .A2(n12984), .ZN(n12989) );
  NAND2_X1 U11454 ( .A1(n14449), .A2(n14448), .ZN(n11000) );
  AND2_X4 U11455 ( .A1(n12447), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11001) );
  AND2_X1 U11456 ( .A1(n14749), .A2(n14735), .ZN(n12388) );
  AND4_X1 U11457 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(
        n11869) );
  AND2_X1 U11458 ( .A1(n14450), .A2(n14426), .ZN(n11484) );
  NAND2_X1 U11459 ( .A1(n14449), .A2(n14448), .ZN(n14466) );
  INV_X1 U11460 ( .A(n12763), .ZN(n11003) );
  NOR2_X2 U11461 ( .A1(n18247), .A2(n21322), .ZN(n18184) );
  INV_X2 U11462 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15008) );
  AND2_X1 U11463 ( .A1(n11764), .A2(n11763), .ZN(n18119) );
  AND2_X2 U11464 ( .A1(n11452), .A2(n11198), .ZN(n11903) );
  CLKBUF_X1 U11465 ( .A(n12697), .Z(n11006) );
  CLKBUF_X1 U11466 ( .A(n13899), .Z(n11007) );
  NAND2_X1 U11467 ( .A1(n13895), .A2(n19671), .ZN(n13899) );
  INV_X1 U11468 ( .A(n15385), .ZN(n11008) );
  NAND2_X1 U11469 ( .A1(n20143), .A2(n12128), .ZN(n11009) );
  INV_X2 U11471 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U11472 ( .A1(n20143), .A2(n12128), .ZN(n12135) );
  NAND2_X1 U11473 ( .A1(n20151), .A2(n12136), .ZN(n12144) );
  AND2_X2 U11475 ( .A1(n11933), .A2(n12395), .ZN(n12208) );
  CLKBUF_X1 U11476 ( .A(n13893), .Z(n11013) );
  NAND2_X1 U11477 ( .A1(n12758), .A2(n12738), .ZN(n12757) );
  NAND2_X1 U11478 ( .A1(n12762), .A2(n12764), .ZN(n12758) );
  AND2_X1 U11479 ( .A1(n12696), .A2(n13892), .ZN(n12697) );
  NOR2_X1 U11480 ( .A1(n18470), .A2(n18452), .ZN(n12767) );
  NAND2_X1 U11481 ( .A1(n11939), .A2(n11935), .ZN(n11014) );
  NAND2_X1 U11482 ( .A1(n11935), .A2(n11939), .ZN(n11936) );
  OAI21_X2 U11483 ( .B1(n11754), .B2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18258), .ZN(n11759) );
  AOI22_X2 U11484 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18168), .B1(
        n18169), .B2(n18178), .ZN(n13820) );
  NAND3_X1 U11485 ( .A1(n18112), .A2(n18050), .A3(n18118), .ZN(n18108) );
  INV_X2 U11487 ( .A(n15104), .ZN(n11129) );
  NAND2_X2 U11488 ( .A1(n12734), .A2(n12713), .ZN(n12739) );
  CLKBUF_X1 U11490 ( .A(n20139), .Z(n11017) );
  XNOR2_X1 U11491 ( .A(n14526), .B(n12115), .ZN(n11018) );
  XNOR2_X1 U11492 ( .A(n11010), .B(n21492), .ZN(n11019) );
  XNOR2_X1 U11493 ( .A(n14526), .B(n12115), .ZN(n20138) );
  XNOR2_X1 U11494 ( .A(n12144), .B(n21492), .ZN(n20160) );
  INV_X1 U11495 ( .A(n11020), .ZN(n12178) );
  AND2_X2 U11496 ( .A1(n15906), .A2(n15909), .ZN(n15799) );
  NAND2_X2 U11497 ( .A1(n14668), .A2(n11955), .ZN(n12021) );
  XNOR2_X1 U11498 ( .A(n11941), .B(n12019), .ZN(n11957) );
  AND2_X2 U11499 ( .A1(n16323), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16324) );
  NOR2_X2 U11500 ( .A1(n16745), .A2(n16302), .ZN(n16305) );
  NOR2_X2 U11501 ( .A1(n14596), .A2(n15181), .ZN(n14597) );
  NAND2_X2 U11502 ( .A1(n15428), .A2(n11451), .ZN(n14596) );
  NAND2_X2 U11503 ( .A1(n16460), .A2(n16462), .ZN(n16454) );
  NOR2_X4 U11504 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14604) );
  CLKBUF_X1 U11505 ( .A(n20151), .Z(n11021) );
  XNOR2_X1 U11506 ( .A(n11009), .B(n21496), .ZN(n11022) );
  BUF_X1 U11507 ( .A(n16119), .Z(n11024) );
  INV_X1 U11508 ( .A(n14938), .ZN(n11025) );
  OAI211_X2 U11509 ( .C1(n16393), .C2(n16405), .A(n16395), .B(n16402), .ZN(
        n15665) );
  NOR2_X2 U11510 ( .A1(n15646), .A2(n15645), .ZN(n16393) );
  AND2_X2 U11511 ( .A1(n15775), .A2(n13613), .ZN(n15761) );
  NOR2_X2 U11512 ( .A1(n15784), .A2(n15786), .ZN(n15775) );
  OR2_X2 U11513 ( .A1(n20178), .A2(n20179), .ZN(n20177) );
  NOR2_X2 U11515 ( .A1(n15084), .A2(n15083), .ZN(n15143) );
  NOR2_X2 U11516 ( .A1(n18783), .A2(n16371), .ZN(n17063) );
  NOR2_X2 U11517 ( .A1(n15188), .A2(n15230), .ZN(n15202) );
  XNOR2_X1 U11518 ( .A(n12127), .B(n21479), .ZN(n20145) );
  NOR2_X2 U11519 ( .A1(n14884), .A2(n14910), .ZN(n14908) );
  OAI21_X4 U11520 ( .B1(n15253), .B2(n15254), .A(n13358), .ZN(n15329) );
  XNOR2_X2 U11521 ( .A(n15147), .B(n13357), .ZN(n15253) );
  NAND3_X2 U11522 ( .A1(n13298), .A2(n13297), .A3(n11094), .ZN(n15147) );
  NOR2_X2 U11523 ( .A1(n15283), .A2(n11446), .ZN(n16460) );
  AOI22_X2 U11524 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14221), .B1(n16570), 
        .B2(n14841), .ZN(n18768) );
  INV_X2 U11525 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11409) );
  NAND2_X2 U11526 ( .A1(n12208), .A2(n14741), .ZN(n12287) );
  OAI21_X2 U11527 ( .B1(n16119), .B2(n11408), .A(n11405), .ZN(n16105) );
  NAND2_X2 U11528 ( .A1(n16097), .A2(n12202), .ZN(n16044) );
  NOR2_X4 U11529 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11823) );
  AND2_X1 U11530 ( .A1(n11817), .A2(n11005), .ZN(n11035) );
  AND2_X1 U11531 ( .A1(n11817), .A2(n11004), .ZN(n11036) );
  AND2_X2 U11532 ( .A1(n11005), .A2(n11823), .ZN(n13637) );
  AND2_X2 U11533 ( .A1(n15520), .A2(n11182), .ZN(n15498) );
  NAND2_X1 U11534 ( .A1(n15667), .A2(n16277), .ZN(n11351) );
  AND2_X1 U11535 ( .A1(n15667), .A2(n11074), .ZN(n11367) );
  NAND2_X1 U11536 ( .A1(n14185), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12714) );
  NAND2_X1 U11537 ( .A1(n12699), .A2(n12687), .ZN(n12682) );
  NAND2_X1 U11538 ( .A1(n12859), .A2(n13168), .ZN(n11237) );
  AND2_X1 U11539 ( .A1(n12828), .A2(n12825), .ZN(n11163) );
  NOR2_X1 U11540 ( .A1(n13897), .A2(n14841), .ZN(n11211) );
  NAND2_X1 U11541 ( .A1(n15738), .A2(n11461), .ZN(n11460) );
  INV_X1 U11542 ( .A(n15751), .ZN(n11461) );
  AND2_X1 U11543 ( .A1(n11093), .A2(n15328), .ZN(n11128) );
  INV_X1 U11544 ( .A(n11455), .ZN(n11454) );
  NAND2_X1 U11545 ( .A1(n11391), .A2(n20177), .ZN(n11204) );
  INV_X1 U11546 ( .A(n15380), .ZN(n13422) );
  OAI21_X1 U11547 ( .B1(n13256), .B2(n13257), .A(n12016), .ZN(n12120) );
  NAND2_X1 U11548 ( .A1(n15284), .A2(n11450), .ZN(n11449) );
  INV_X1 U11549 ( .A(n15364), .ZN(n11450) );
  INV_X1 U11550 ( .A(n15627), .ZN(n15582) );
  NAND2_X1 U11551 ( .A1(n13179), .A2(n13859), .ZN(n13180) );
  AOI21_X1 U11552 ( .B1(n11179), .B2(n11181), .A(n11177), .ZN(n11176) );
  NAND2_X1 U11553 ( .A1(n16648), .A2(n11179), .ZN(n11178) );
  INV_X1 U11554 ( .A(n16631), .ZN(n11177) );
  AND2_X1 U11555 ( .A1(n12921), .A2(n11348), .ZN(n11347) );
  INV_X1 U11556 ( .A(n17031), .ZN(n11348) );
  NAND2_X1 U11557 ( .A1(n15212), .A2(n15210), .ZN(n13171) );
  AND2_X1 U11558 ( .A1(n15209), .A2(n13164), .ZN(n11187) );
  AND2_X1 U11559 ( .A1(n14841), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14438) );
  OAI211_X1 U11560 ( .C1(n18138), .C2(n18108), .A(n11765), .B(n18158), .ZN(
        n11766) );
  AND2_X1 U11561 ( .A1(n11715), .A2(n20816), .ZN(n11688) );
  AOI21_X1 U11562 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17090), .A(
        n11509), .ZN(n11616) );
  INV_X1 U11563 ( .A(n14520), .ZN(n13766) );
  AND2_X1 U11564 ( .A1(n15748), .A2(n15736), .ZN(n15734) );
  NOR2_X1 U11565 ( .A1(n16477), .A2(n15703), .ZN(n15702) );
  NAND2_X1 U11566 ( .A1(n16490), .A2(n16475), .ZN(n16477) );
  AND2_X1 U11567 ( .A1(n14127), .A2(n14126), .ZN(n16970) );
  INV_X1 U11568 ( .A(n11339), .ZN(n11336) );
  NAND2_X1 U11569 ( .A1(n16613), .A2(n14232), .ZN(n16583) );
  NAND2_X1 U11570 ( .A1(n12967), .A2(n12968), .ZN(n11344) );
  AND2_X1 U11571 ( .A1(n14148), .A2(n14147), .ZN(n16945) );
  OR2_X1 U11572 ( .A1(n16984), .A2(n16970), .ZN(n11039) );
  AND2_X1 U11573 ( .A1(n17010), .A2(n17007), .ZN(n12932) );
  NAND2_X1 U11574 ( .A1(n13912), .A2(n18907), .ZN(n14234) );
  AND4_X1 U11575 ( .A1(n13909), .A2(n14286), .A3(n13908), .A4(n13907), .ZN(
        n13910) );
  AND2_X1 U11576 ( .A1(n18471), .A2(n17481), .ZN(n19492) );
  NOR2_X1 U11577 ( .A1(n13836), .A2(n18137), .ZN(n21245) );
  NAND2_X1 U11578 ( .A1(n11293), .A2(n11290), .ZN(n11289) );
  INV_X1 U11579 ( .A(n18315), .ZN(n11290) );
  NAND2_X1 U11580 ( .A1(n21029), .A2(n21013), .ZN(n21012) );
  NAND2_X1 U11581 ( .A1(n20988), .A2(n11794), .ZN(n15373) );
  NAND2_X1 U11582 ( .A1(n14659), .A2(n18907), .ZN(n18911) );
  XNOR2_X1 U11583 ( .A(n16583), .B(n14221), .ZN(n16571) );
  NOR2_X1 U11584 ( .A1(n21263), .A2(n21381), .ZN(n21110) );
  AND2_X1 U11585 ( .A1(n11472), .A2(n14683), .ZN(n12209) );
  CLKBUF_X1 U11586 ( .A(n11031), .Z(n13700) );
  AOI21_X1 U11587 ( .B1(n20214), .B2(n21585), .A(n11209), .ZN(n11408) );
  NAND2_X1 U11588 ( .A1(n12076), .A2(n12075), .ZN(n12137) );
  INV_X1 U11589 ( .A(n12108), .ZN(n11987) );
  OR2_X1 U11590 ( .A1(n11027), .A2(n21832), .ZN(n12031) );
  NAND2_X1 U11591 ( .A1(n12688), .A2(n12699), .ZN(n13893) );
  NAND2_X1 U11592 ( .A1(n12746), .A2(n12745), .ZN(n12748) );
  NAND2_X1 U11593 ( .A1(n12753), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12746) );
  INV_X1 U11594 ( .A(n12866), .ZN(n11239) );
  AOI22_X1 U11595 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19417), .B1(
        n19462), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12822) );
  NAND2_X1 U11596 ( .A1(n12753), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11430) );
  OR2_X1 U11597 ( .A1(n12685), .A2(n14193), .ZN(n11213) );
  OR2_X1 U11598 ( .A1(n12683), .A2(n19720), .ZN(n12684) );
  AND2_X1 U11599 ( .A1(n12698), .A2(n12687), .ZN(n12703) );
  NAND2_X1 U11600 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21394), .ZN(
        n11492) );
  AOI21_X1 U11601 ( .B1(n21388), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11503), .ZN(n11513) );
  NOR2_X1 U11602 ( .A1(n11615), .A2(n11502), .ZN(n11503) );
  OAI22_X1 U11603 ( .A1(n21394), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n21398), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11512) );
  NOR2_X1 U11604 ( .A1(n11228), .A2(n11226), .ZN(n11225) );
  NAND2_X1 U11605 ( .A1(n11575), .A2(n11227), .ZN(n11226) );
  INV_X1 U11606 ( .A(n11571), .ZN(n11228) );
  NAND2_X1 U11607 ( .A1(n11620), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11227) );
  OR2_X1 U11608 ( .A1(n12235), .A2(n12234), .ZN(n12274) );
  NOR2_X1 U11609 ( .A1(n11931), .A2(n14712), .ZN(n13734) );
  NAND2_X1 U11610 ( .A1(n13565), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13606) );
  NAND2_X1 U11611 ( .A1(n13234), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13344) );
  AND2_X1 U11612 ( .A1(n13242), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13277) );
  NOR2_X2 U11613 ( .A1(n14689), .A2(n13234), .ZN(n13417) );
  INV_X1 U11614 ( .A(n15758), .ZN(n11306) );
  NAND2_X1 U11615 ( .A1(n16096), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12202) );
  NOR2_X1 U11616 ( .A1(n16132), .A2(n20215), .ZN(n12195) );
  NAND2_X1 U11617 ( .A1(n11209), .A2(n11121), .ZN(n11407) );
  NAND2_X1 U11618 ( .A1(n11408), .A2(n11405), .ZN(n11404) );
  INV_X1 U11619 ( .A(n11393), .ZN(n11392) );
  AND2_X1 U11620 ( .A1(n15126), .A2(n11092), .ZN(n15154) );
  INV_X1 U11621 ( .A(n15155), .ZN(n11297) );
  INV_X1 U11622 ( .A(n14706), .ZN(n11315) );
  NAND2_X1 U11623 ( .A1(n11319), .A2(n14888), .ZN(n11318) );
  INV_X1 U11624 ( .A(n14705), .ZN(n11319) );
  NAND2_X1 U11625 ( .A1(n12009), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12032) );
  OR2_X1 U11626 ( .A1(n11984), .A2(n11983), .ZN(n12181) );
  INV_X1 U11627 ( .A(n12248), .ZN(n12263) );
  AND3_X1 U11628 ( .A1(n14712), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n11027), 
        .ZN(n12248) );
  OR2_X1 U11629 ( .A1(n11915), .A2(n11926), .ZN(n11880) );
  AND2_X1 U11630 ( .A1(n11991), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11867) );
  OAI21_X1 U11631 ( .B1(n21838), .B2(n21834), .A(n21825), .ZN(n14673) );
  INV_X1 U11632 ( .A(n16540), .ZN(n11390) );
  OR2_X1 U11633 ( .A1(n11051), .A2(n12943), .ZN(n12958) );
  OR2_X1 U11634 ( .A1(n11421), .A2(n11420), .ZN(n11419) );
  INV_X1 U11635 ( .A(n12948), .ZN(n11420) );
  INV_X1 U11636 ( .A(n12951), .ZN(n11421) );
  AND2_X1 U11637 ( .A1(n12911), .A2(n11411), .ZN(n12924) );
  AND2_X1 U11638 ( .A1(n11057), .A2(n11412), .ZN(n11411) );
  INV_X1 U11639 ( .A(n11107), .ZN(n11412) );
  NOR2_X1 U11640 ( .A1(n15582), .A2(n19761), .ZN(n14442) );
  NOR2_X1 U11641 ( .A1(n12875), .A2(n12876), .ZN(n12868) );
  OR2_X1 U11642 ( .A1(n15649), .A2(n12648), .ZN(n14082) );
  OR2_X1 U11643 ( .A1(n15543), .A2(n12648), .ZN(n14057) );
  NAND2_X1 U11644 ( .A1(n11001), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14081) );
  INV_X1 U11645 ( .A(n16500), .ZN(n11385) );
  AND2_X1 U11646 ( .A1(n11444), .A2(n15495), .ZN(n11443) );
  INV_X1 U11647 ( .A(n16456), .ZN(n11444) );
  INV_X1 U11648 ( .A(n16429), .ZN(n11360) );
  AND2_X1 U11649 ( .A1(n16444), .A2(n16436), .ZN(n11361) );
  AND2_X1 U11650 ( .A1(n11366), .A2(n11365), .ZN(n11364) );
  INV_X1 U11651 ( .A(n15205), .ZN(n11365) );
  INV_X1 U11652 ( .A(n14865), .ZN(n11355) );
  NOR2_X1 U11653 ( .A1(n11357), .A2(n14507), .ZN(n11356) );
  INV_X1 U11654 ( .A(n14595), .ZN(n11357) );
  NAND2_X1 U11655 ( .A1(n13005), .A2(n13004), .ZN(n11175) );
  NAND2_X1 U11656 ( .A1(n11410), .A2(n13859), .ZN(n12986) );
  NOR2_X1 U11657 ( .A1(n16661), .A2(n11244), .ZN(n11243) );
  INV_X1 U11658 ( .A(n11246), .ZN(n11244) );
  NOR2_X1 U11659 ( .A1(n16995), .A2(n17002), .ZN(n11247) );
  NOR2_X1 U11660 ( .A1(n14926), .A2(n14925), .ZN(n14924) );
  NAND2_X1 U11661 ( .A1(n14402), .A2(n19472), .ZN(n14440) );
  NOR2_X1 U11662 ( .A1(n11492), .A2(n20368), .ZN(n11690) );
  NOR2_X1 U11663 ( .A1(n11493), .A2(n11495), .ZN(n11644) );
  INV_X1 U11664 ( .A(n20840), .ZN(n11609) );
  NOR2_X1 U11665 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n11259), .ZN(
        n11258) );
  NOR2_X1 U11666 ( .A1(n20609), .A2(n11268), .ZN(n11267) );
  INV_X1 U11667 ( .A(n18096), .ZN(n11760) );
  NAND2_X1 U11668 ( .A1(n11280), .A2(n18258), .ZN(n11764) );
  NOR2_X1 U11669 ( .A1(n18271), .A2(n21116), .ZN(n11743) );
  NAND2_X1 U11670 ( .A1(n18291), .A2(n11739), .ZN(n11741) );
  NOR2_X1 U11671 ( .A1(n20959), .A2(n19135), .ZN(n13206) );
  INV_X1 U11672 ( .A(n20368), .ZN(n11196) );
  INV_X1 U11673 ( .A(n21005), .ZN(n11197) );
  NOR2_X1 U11674 ( .A1(n13420), .A2(n15839), .ZN(n13438) );
  NOR2_X1 U11675 ( .A1(n13313), .A2(n13312), .ZN(n13329) );
  NOR2_X1 U11676 ( .A1(n13769), .A2(n21639), .ZN(n21720) );
  INV_X1 U11677 ( .A(n13752), .ZN(n13749) );
  OAI21_X1 U11678 ( .B1(n12287), .B2(n13733), .A(n13732), .ZN(n14554) );
  INV_X1 U11679 ( .A(n21844), .ZN(n15390) );
  INV_X1 U11680 ( .A(n13344), .ZN(n13724) );
  NAND2_X1 U11681 ( .A1(n15714), .A2(n11459), .ZN(n11458) );
  OR2_X1 U11682 ( .A1(n13760), .A2(n15717), .ZN(n13761) );
  INV_X1 U11683 ( .A(n11459), .ZN(n11457) );
  NAND2_X1 U11684 ( .A1(n13612), .A2(n13611), .ZN(n15777) );
  OR2_X1 U11685 ( .A1(n16076), .A2(n11099), .ZN(n13611) );
  AND2_X1 U11686 ( .A1(n11128), .A2(n11127), .ZN(n11126) );
  INV_X1 U11687 ( .A(n15942), .ZN(n11127) );
  NAND2_X1 U11688 ( .A1(n13808), .A2(n13807), .ZN(n17133) );
  AND2_X1 U11689 ( .A1(n15389), .A2(n10985), .ZN(n13807) );
  INV_X1 U11690 ( .A(n12380), .ZN(n14512) );
  AND2_X1 U11691 ( .A1(n15944), .A2(n11096), .ZN(n15930) );
  INV_X1 U11692 ( .A(n15931), .ZN(n11309) );
  NAND2_X1 U11693 ( .A1(n15944), .A2(n11081), .ZN(n15937) );
  NAND2_X1 U11694 ( .A1(n15944), .A2(n11311), .ZN(n15935) );
  AND2_X1 U11695 ( .A1(n15944), .A2(n15943), .ZN(n15946) );
  NOR2_X1 U11696 ( .A1(n20171), .A2(n11398), .ZN(n11397) );
  INV_X1 U11697 ( .A(n12155), .ZN(n11398) );
  NAND2_X1 U11698 ( .A1(n11315), .A2(n11317), .ZN(n14912) );
  INV_X1 U11699 ( .A(n12129), .ZN(n11130) );
  NAND2_X1 U11700 ( .A1(n15108), .A2(n15107), .ZN(n21953) );
  OR2_X1 U11701 ( .A1(n14667), .A2(n14938), .ZN(n21977) );
  NOR2_X1 U11702 ( .A1(n22044), .A2(n21924), .ZN(n22002) );
  NAND2_X1 U11703 ( .A1(n21832), .A2(n14673), .ZN(n21924) );
  NOR2_X1 U11704 ( .A1(n21999), .A2(n21924), .ZN(n22057) );
  AND2_X1 U11705 ( .A1(n14667), .A2(n11025), .ZN(n22041) );
  NOR2_X1 U11706 ( .A1(n16336), .A2(n13931), .ZN(n14564) );
  NOR2_X1 U11707 ( .A1(n14190), .A2(n13900), .ZN(n14640) );
  NAND2_X1 U11708 ( .A1(n13000), .A2(n12998), .ZN(n12995) );
  AND2_X1 U11709 ( .A1(n12989), .A2(n12987), .ZN(n13000) );
  AND2_X1 U11710 ( .A1(n16877), .A2(n11387), .ZN(n16529) );
  AND2_X1 U11711 ( .A1(n11106), .A2(n11388), .ZN(n11387) );
  INV_X1 U11712 ( .A(n16527), .ZN(n11388) );
  NOR2_X1 U11713 ( .A1(n12958), .A2(n12957), .ZN(n12959) );
  NOR3_X1 U11714 ( .A1(n12934), .A2(n12933), .A3(n11421), .ZN(n12954) );
  OR2_X1 U11715 ( .A1(n12926), .A2(n12925), .ZN(n12934) );
  AND2_X1 U11716 ( .A1(n13109), .A2(n13108), .ZN(n16451) );
  NOR2_X1 U11717 ( .A1(n11437), .A2(n11435), .ZN(n11434) );
  AND2_X1 U11718 ( .A1(n13052), .A2(n13051), .ZN(n14476) );
  NAND2_X1 U11719 ( .A1(n11445), .A2(n11443), .ZN(n11442) );
  INV_X1 U11720 ( .A(n16435), .ZN(n11445) );
  NAND2_X1 U11721 ( .A1(n11447), .A2(n16469), .ZN(n11446) );
  INV_X1 U11722 ( .A(n11449), .ZN(n11447) );
  NOR2_X1 U11723 ( .A1(n13968), .A2(n11380), .ZN(n18479) );
  NAND2_X1 U11724 ( .A1(n11383), .A2(n11382), .ZN(n11380) );
  AND2_X1 U11725 ( .A1(n13942), .A2(n13941), .ZN(n18478) );
  NAND2_X1 U11726 ( .A1(n15081), .A2(n11362), .ZN(n15347) );
  AND2_X1 U11727 ( .A1(n11364), .A2(n11363), .ZN(n11362) );
  INV_X1 U11728 ( .A(n15266), .ZN(n11363) );
  NAND2_X1 U11729 ( .A1(n15081), .A2(n11364), .ZN(n15267) );
  NAND2_X1 U11730 ( .A1(n15081), .A2(n11366), .ZN(n15227) );
  AND2_X1 U11731 ( .A1(n15081), .A2(n15138), .ZN(n15229) );
  AND2_X1 U11732 ( .A1(n13079), .A2(n13078), .ZN(n15079) );
  NAND2_X1 U11733 ( .A1(n11352), .A2(n11356), .ZN(n14864) );
  INV_X1 U11734 ( .A(n11185), .ZN(n11184) );
  NAND2_X1 U11735 ( .A1(n12887), .A2(n11467), .ZN(n15214) );
  AND2_X1 U11736 ( .A1(n15431), .A2(n15430), .ZN(n15433) );
  NOR2_X1 U11737 ( .A1(n11343), .A2(n16651), .ZN(n11340) );
  INV_X1 U11738 ( .A(n11377), .ZN(n11375) );
  OAI21_X1 U11739 ( .B1(n15234), .B2(n11168), .A(n11166), .ZN(n17008) );
  INV_X1 U11740 ( .A(n11169), .ZN(n11168) );
  NAND2_X1 U11741 ( .A1(n11055), .A2(n13167), .ZN(n11214) );
  NAND2_X1 U11742 ( .A1(n14260), .A2(n14292), .ZN(n14639) );
  NAND2_X1 U11743 ( .A1(n15683), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15484) );
  NAND2_X1 U11744 ( .A1(n13890), .A2(n13887), .ZN(n14647) );
  NAND2_X1 U11745 ( .A1(n16277), .A2(n13886), .ZN(n13887) );
  INV_X1 U11746 ( .A(n14985), .ZN(n14981) );
  AND2_X1 U11747 ( .A1(n19475), .A2(n19508), .ZN(n19511) );
  NAND2_X1 U11748 ( .A1(n14844), .A2(n14843), .ZN(n19475) );
  INV_X1 U11749 ( .A(n14842), .ZN(n14843) );
  NAND2_X1 U11750 ( .A1(n18897), .A2(n14841), .ZN(n14844) );
  OR2_X1 U11751 ( .A1(n19613), .A2(n19611), .ZN(n19421) );
  AND3_X1 U11752 ( .A1(n18890), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18907) );
  OAI21_X1 U11753 ( .B1(n17578), .B2(n17577), .A(n21440), .ZN(n20777) );
  NAND2_X1 U11754 ( .A1(n15373), .A2(n11795), .ZN(n20781) );
  NAND3_X1 U11755 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n21013), .ZN(n20409) );
  NOR2_X1 U11756 ( .A1(n21414), .A2(n13200), .ZN(n17092) );
  NOR2_X1 U11757 ( .A1(n21900), .A2(n20322), .ZN(n20782) );
  OR2_X1 U11758 ( .A1(n18125), .A2(n18258), .ZN(n11296) );
  OR2_X1 U11759 ( .A1(n13190), .A2(n18125), .ZN(n11295) );
  NOR2_X2 U11760 ( .A1(n18088), .A2(n18087), .ZN(n18103) );
  NAND2_X1 U11761 ( .A1(n20812), .A2(n21440), .ZN(n11229) );
  XNOR2_X1 U11762 ( .A(n11737), .B(n11194), .ZN(n18302) );
  INV_X1 U11763 ( .A(n11736), .ZN(n11194) );
  NAND2_X1 U11764 ( .A1(n18302), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18301) );
  OR2_X1 U11765 ( .A1(n11749), .A2(n21039), .ZN(n21272) );
  OR2_X1 U11766 ( .A1(n21038), .A2(n11749), .ZN(n18091) );
  NAND2_X1 U11767 ( .A1(n18048), .A2(n21177), .ZN(n21039) );
  NAND2_X1 U11768 ( .A1(n21192), .A2(n18048), .ZN(n21038) );
  INV_X1 U11769 ( .A(n11755), .ZN(n11756) );
  OAI22_X1 U11770 ( .A1(n11757), .A2(n21338), .B1(n18258), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11755) );
  NAND2_X1 U11771 ( .A1(n21132), .A2(n21163), .ZN(n18197) );
  NOR2_X1 U11772 ( .A1(n18273), .A2(n18272), .ZN(n18271) );
  OR2_X1 U11773 ( .A1(n18316), .A2(n18315), .ZN(n11292) );
  NOR2_X2 U11774 ( .A1(n11535), .A2(n11534), .ZN(n20370) );
  NAND2_X1 U11775 ( .A1(n21412), .A2(n21402), .ZN(n11148) );
  OR2_X1 U11776 ( .A1(n21412), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11147) );
  NAND2_X1 U11777 ( .A1(n11145), .A2(n11143), .ZN(n11142) );
  INV_X1 U11778 ( .A(n21409), .ZN(n11145) );
  AND2_X1 U11779 ( .A1(n21442), .A2(n11144), .ZN(n11143) );
  XNOR2_X1 U11780 ( .A(n12389), .B(n13765), .ZN(n15718) );
  INV_X1 U11781 ( .A(n16015), .ZN(n16019) );
  AND2_X1 U11782 ( .A1(n12415), .A2(n12290), .ZN(n21624) );
  AND2_X1 U11783 ( .A1(n12415), .A2(n12392), .ZN(n21625) );
  INV_X1 U11784 ( .A(n21624), .ZN(n21635) );
  OR2_X1 U11785 ( .A1(n21953), .A2(n15043), .ZN(n22326) );
  AND2_X1 U11786 ( .A1(n15427), .A2(n11468), .ZN(n11451) );
  INV_X1 U11787 ( .A(n16474), .ZN(n16457) );
  OR2_X1 U11788 ( .A1(n16433), .A2(n14575), .ZN(n16474) );
  INV_X1 U11789 ( .A(n16564), .ZN(n19763) );
  AOI21_X1 U11790 ( .B1(n16289), .B2(n17474), .A(n16572), .ZN(n11221) );
  OR2_X1 U11791 ( .A1(n16576), .A2(n11335), .ZN(n11322) );
  INV_X1 U11792 ( .A(n16390), .ZN(n18775) );
  NAND2_X1 U11793 ( .A1(n18911), .A2(n13139), .ZN(n17459) );
  AND2_X1 U11794 ( .A1(n10987), .A2(n16578), .ZN(n11331) );
  INV_X1 U11795 ( .A(n11332), .ZN(n11330) );
  OAI21_X1 U11796 ( .B1(n10987), .B2(n11065), .A(n11333), .ZN(n11332) );
  OAI21_X1 U11797 ( .B1(n16571), .B2(n18881), .A(n14235), .ZN(n11338) );
  INV_X1 U11798 ( .A(n11335), .ZN(n11326) );
  OAI21_X1 U11799 ( .B1(n11335), .B2(n11325), .A(n18856), .ZN(n11324) );
  INV_X1 U11800 ( .A(n11370), .ZN(n11369) );
  OAI21_X1 U11801 ( .B1(n18781), .B2(n18870), .A(n11371), .ZN(n11370) );
  NOR2_X1 U11802 ( .A1(n16763), .A2(n11372), .ZN(n11371) );
  OR2_X1 U11803 ( .A1(n14429), .A2(n14407), .ZN(n17481) );
  NOR2_X2 U11804 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19508) );
  INV_X1 U11805 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19432) );
  NAND2_X1 U11806 ( .A1(n14432), .A2(n14418), .ZN(n18471) );
  AND2_X1 U11807 ( .A1(n14449), .A2(n14435), .ZN(n17488) );
  OR2_X1 U11808 ( .A1(n14434), .A2(n14433), .ZN(n14435) );
  INV_X1 U11809 ( .A(n19939), .ZN(n19743) );
  INV_X1 U11810 ( .A(n17092), .ZN(n20322) );
  INV_X1 U11811 ( .A(n20755), .ZN(n11255) );
  INV_X1 U11812 ( .A(n20757), .ZN(n11254) );
  NAND2_X1 U11813 ( .A1(n20760), .A2(n20759), .ZN(n11249) );
  NOR2_X1 U11814 ( .A1(n11252), .A2(n11251), .ZN(n11250) );
  NOR2_X1 U11815 ( .A1(n20762), .A2(n20763), .ZN(n11251) );
  INV_X1 U11816 ( .A(n20761), .ZN(n11252) );
  NAND2_X1 U11817 ( .A1(n20742), .A2(n20743), .ZN(n20756) );
  NOR2_X1 U11818 ( .A1(n11642), .A2(n11641), .ZN(n20830) );
  INV_X1 U11819 ( .A(n13829), .ZN(n11193) );
  XNOR2_X1 U11820 ( .A(n13822), .B(n20983), .ZN(n13844) );
  NOR3_X1 U11821 ( .A1(n18157), .A2(n21206), .A3(n18138), .ZN(n18166) );
  NAND2_X1 U11822 ( .A1(n18184), .A2(n18048), .ZN(n18157) );
  INV_X1 U11823 ( .A(n18187), .ZN(n18261) );
  AOI22_X1 U11824 ( .A1(n21251), .A2(n21384), .B1(n21252), .B2(n21293), .ZN(
        n11191) );
  AND2_X1 U11825 ( .A1(n21253), .A2(n11190), .ZN(n11189) );
  OR2_X1 U11826 ( .A1(n21285), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11190) );
  INV_X1 U11827 ( .A(n21219), .ZN(n21293) );
  INV_X1 U11828 ( .A(n21238), .ZN(n21275) );
  OAI21_X2 U11829 ( .B1(n13217), .B2(n13216), .A(n21440), .ZN(n21263) );
  OAI21_X1 U11830 ( .B1(n12850), .B2(n12773), .A(n16334), .ZN(n12778) );
  AOI22_X1 U11831 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12831), .B1(
        n12842), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12816) );
  INV_X1 U11832 ( .A(n12715), .ZN(n12677) );
  NAND2_X1 U11833 ( .A1(n11008), .A2(n22029), .ZN(n12243) );
  NAND2_X1 U11834 ( .A1(n11923), .A2(n15380), .ZN(n11945) );
  INV_X1 U11835 ( .A(n12137), .ZN(n11210) );
  NAND2_X1 U11836 ( .A1(n12088), .A2(n12087), .ZN(n12146) );
  OR2_X1 U11837 ( .A1(n12098), .A2(n12097), .ZN(n12172) );
  INV_X1 U11838 ( .A(n12181), .ZN(n12013) );
  OR2_X1 U11839 ( .A1(n12042), .A2(n12041), .ZN(n12121) );
  AOI22_X1 U11840 ( .A1(n11991), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n11903), .ZN(n11834) );
  NAND2_X1 U11841 ( .A1(n13637), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U11842 ( .A1(n12055), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11854) );
  AOI22_X1 U11843 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11851) );
  INV_X1 U11844 ( .A(n11237), .ZN(n11234) );
  NAND2_X1 U11845 ( .A1(n12861), .A2(n12860), .ZN(n13174) );
  NOR2_X1 U11846 ( .A1(n12687), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13949) );
  AOI22_X1 U11847 ( .A1(n15683), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12667), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12460) );
  AOI21_X1 U11848 ( .B1(n12668), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12648), .ZN(n12620) );
  NAND2_X1 U11849 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12612) );
  AOI21_X1 U11850 ( .B1(n12668), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12613) );
  NOR2_X1 U11851 ( .A1(n20830), .A2(n11729), .ZN(n11707) );
  AOI21_X1 U11852 ( .B1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B2(n17783), .A(
        n11152), .ZN(n11151) );
  INV_X1 U11853 ( .A(n11557), .ZN(n11152) );
  INV_X1 U11854 ( .A(n11555), .ZN(n11153) );
  NOR2_X1 U11855 ( .A1(n15385), .A2(n21832), .ZN(n11400) );
  NAND2_X1 U11856 ( .A1(n13274), .A2(n13273), .ZN(n14726) );
  NOR2_X1 U11857 ( .A1(n11460), .A2(n15726), .ZN(n11459) );
  AND2_X1 U11858 ( .A1(n11113), .A2(n11463), .ZN(n11462) );
  NOR2_X1 U11859 ( .A1(n15929), .A2(n11464), .ZN(n11463) );
  INV_X1 U11860 ( .A(n15933), .ZN(n11464) );
  NAND2_X1 U11861 ( .A1(n11456), .A2(n13389), .ZN(n11455) );
  INV_X1 U11862 ( .A(n15846), .ZN(n11456) );
  XNOR2_X1 U11863 ( .A(n12170), .B(n12169), .ZN(n13296) );
  AND2_X1 U11864 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13231), .ZN(
        n13242) );
  NOR2_X1 U11865 ( .A1(n15771), .A2(n11308), .ZN(n11307) );
  INV_X1 U11866 ( .A(n15789), .ZN(n11308) );
  INV_X1 U11867 ( .A(n15934), .ZN(n11310) );
  NOR2_X1 U11868 ( .A1(n11313), .A2(n11312), .ZN(n11311) );
  INV_X1 U11869 ( .A(n15818), .ZN(n11313) );
  INV_X1 U11870 ( .A(n15943), .ZN(n11312) );
  NAND2_X1 U11871 ( .A1(n16122), .A2(n12194), .ZN(n20214) );
  NOR2_X1 U11872 ( .A1(n15134), .A2(n11299), .ZN(n11298) );
  INV_X1 U11873 ( .A(n15125), .ZN(n11299) );
  OR2_X1 U11874 ( .A1(n12074), .A2(n12073), .ZN(n12148) );
  NAND2_X1 U11875 ( .A1(n13764), .A2(n12380), .ZN(n12378) );
  AND2_X1 U11876 ( .A1(n14749), .A2(n11858), .ZN(n12246) );
  AND3_X1 U11877 ( .A1(n12394), .A2(n12110), .A3(n12211), .ZN(n13808) );
  NOR2_X1 U11878 ( .A1(n14532), .A2(n11858), .ZN(n14537) );
  OR2_X1 U11879 ( .A1(n12032), .A2(n11987), .ZN(n11971) );
  NOR2_X1 U11880 ( .A1(n12032), .A2(n12013), .ZN(n12100) );
  OR2_X1 U11881 ( .A1(n12062), .A2(n12061), .ZN(n12139) );
  NAND2_X1 U11882 ( .A1(n12032), .A2(n12031), .ZN(n12250) );
  AND2_X1 U11883 ( .A1(n12248), .A2(n12246), .ZN(n12265) );
  AND2_X1 U11884 ( .A1(n11915), .A2(n11026), .ZN(n12395) );
  AOI22_X1 U11885 ( .A1(n12055), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13637), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U11886 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11958), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U11887 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11991), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U11888 ( .A1(n11031), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11991), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11844) );
  INV_X1 U11889 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22018) );
  OR2_X1 U11890 ( .A1(n13022), .A2(n13023), .ZN(n13880) );
  NAND2_X1 U11891 ( .A1(n13024), .A2(n13023), .ZN(n13029) );
  INV_X1 U11892 ( .A(n16841), .ZN(n11389) );
  INV_X1 U11893 ( .A(n12915), .ZN(n11413) );
  NOR2_X1 U11894 ( .A1(n11415), .A2(n12918), .ZN(n11414) );
  INV_X1 U11895 ( .A(n12910), .ZN(n11415) );
  NAND2_X1 U11896 ( .A1(n12911), .A2(n12910), .ZN(n12920) );
  NAND2_X1 U11897 ( .A1(n11028), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11395) );
  NAND2_X1 U11898 ( .A1(n13019), .A2(n14857), .ZN(n11396) );
  INV_X1 U11899 ( .A(n13861), .ZN(n16287) );
  CLKBUF_X1 U11900 ( .A(n15588), .Z(n15677) );
  AND2_X1 U11901 ( .A1(n16511), .A2(n16505), .ZN(n11386) );
  INV_X1 U11902 ( .A(n13949), .ZN(n14167) );
  AND2_X1 U11903 ( .A1(n11382), .A2(n15218), .ZN(n11381) );
  AND2_X1 U11904 ( .A1(n12564), .A2(n12563), .ZN(n13976) );
  INV_X1 U11905 ( .A(n18478), .ZN(n11382) );
  NAND2_X1 U11906 ( .A1(n16336), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13885) );
  NOR2_X1 U11907 ( .A1(n16312), .A2(n18688), .ZN(n16314) );
  AND2_X1 U11908 ( .A1(n15138), .A2(n15228), .ZN(n11366) );
  NAND2_X1 U11909 ( .A1(n12757), .A2(n12756), .ZN(n11358) );
  NOR2_X1 U11910 ( .A1(n11059), .A2(n11174), .ZN(n11173) );
  INV_X1 U11911 ( .A(n13009), .ZN(n11174) );
  NOR2_X1 U11912 ( .A1(n11068), .A2(n11346), .ZN(n11345) );
  INV_X1 U11913 ( .A(n16632), .ZN(n11346) );
  NOR2_X1 U11914 ( .A1(n14216), .A2(n11278), .ZN(n11277) );
  INV_X1 U11915 ( .A(n11476), .ZN(n11278) );
  NOR2_X1 U11916 ( .A1(n11378), .A2(n16945), .ZN(n11377) );
  NAND2_X1 U11917 ( .A1(n16995), .A2(n17002), .ZN(n11246) );
  AND2_X1 U11918 ( .A1(n18576), .A2(n13859), .ZN(n12955) );
  NAND2_X1 U11919 ( .A1(n13168), .A2(n13161), .ZN(n11232) );
  NAND2_X1 U11920 ( .A1(n13174), .A2(n12862), .ZN(n13165) );
  INV_X1 U11921 ( .A(n12865), .ZN(n11269) );
  NAND2_X1 U11922 ( .A1(n12868), .A2(n12867), .ZN(n12879) );
  NAND2_X1 U11923 ( .A1(n11164), .A2(n12813), .ZN(n12866) );
  NAND2_X1 U11924 ( .A1(n11429), .A2(n12717), .ZN(n12719) );
  INV_X1 U11925 ( .A(n14150), .ZN(n13948) );
  OAI21_X1 U11926 ( .B1(n12687), .B2(n17514), .A(n19472), .ZN(n13943) );
  NAND4_X1 U11927 ( .A1(n12811), .A2(n12810), .A3(n12809), .A4(n12808), .ZN(
        n13148) );
  NAND2_X1 U11928 ( .A1(n12652), .A2(n13899), .ZN(n11426) );
  CLKBUF_X1 U11929 ( .A(n12447), .Z(n12448) );
  NOR2_X2 U11930 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14613) );
  NAND2_X1 U11931 ( .A1(n11134), .A2(n14292), .ZN(n14185) );
  AND2_X1 U11932 ( .A1(n19872), .A2(n14468), .ZN(n11135) );
  NAND2_X1 U11933 ( .A1(n14426), .A2(n14438), .ZN(n14428) );
  CLKBUF_X1 U11934 ( .A(n14454), .Z(n14603) );
  INV_X1 U11935 ( .A(n13029), .ZN(n13886) );
  NAND2_X1 U11936 ( .A1(n11157), .A2(n12648), .ZN(n11156) );
  NAND2_X1 U11937 ( .A1(n11155), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11154) );
  NAND2_X1 U11938 ( .A1(n12637), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11162) );
  NAND2_X1 U11939 ( .A1(n12638), .A2(n12648), .ZN(n11161) );
  AND2_X1 U11940 ( .A1(n14840), .A2(n18900), .ZN(n14842) );
  NOR2_X1 U11941 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20995), .ZN(
        n11549) );
  NOR2_X1 U11942 ( .A1(n18035), .A2(n11265), .ZN(n11264) );
  NAND2_X1 U11943 ( .A1(n18221), .A2(n11750), .ZN(n18026) );
  INV_X1 U11944 ( .A(n18304), .ZN(n11293) );
  NAND2_X1 U11945 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20379) );
  NAND2_X1 U11946 ( .A1(n11598), .A2(n11040), .ZN(n17574) );
  INV_X1 U11947 ( .A(n20988), .ZN(n21011) );
  NOR3_X1 U11948 ( .A1(n13203), .A2(n11600), .A3(n11040), .ZN(n11608) );
  NAND2_X1 U11949 ( .A1(n21379), .A2(n11136), .ZN(n15375) );
  NAND2_X1 U11950 ( .A1(n11138), .A2(n11137), .ZN(n11136) );
  INV_X1 U11951 ( .A(n11613), .ZN(n11137) );
  NOR2_X1 U11952 ( .A1(n21029), .A2(n20995), .ZN(n17588) );
  NOR3_X1 U11953 ( .A1(n17576), .A2(n11599), .A3(n11601), .ZN(n11794) );
  NAND3_X1 U11954 ( .A1(n11546), .A2(n11545), .A3(n11544), .ZN(n11611) );
  AOI211_X1 U11955 ( .C1(n10992), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n11543), .B(n11542), .ZN(n11544) );
  OR2_X1 U11956 ( .A1(n21412), .A2(n21413), .ZN(n11144) );
  NOR2_X1 U11957 ( .A1(n12279), .A2(n12278), .ZN(n14396) );
  AND2_X1 U11958 ( .A1(n12277), .A2(n12276), .ZN(n12278) );
  INV_X1 U11959 ( .A(n15878), .ZN(n15875) );
  OR2_X1 U11960 ( .A1(n21720), .A2(n21721), .ZN(n21781) );
  AOI22_X1 U11961 ( .A1(n13672), .A2(n13671), .B1(n13757), .B2(n15739), .ZN(
        n15738) );
  AOI22_X1 U11962 ( .A1(n13630), .A2(n13629), .B1(n13757), .B2(n15763), .ZN(
        n15762) );
  AND2_X1 U11963 ( .A1(n15392), .A2(n21447), .ZN(n20035) );
  NAND2_X1 U11964 ( .A1(n15391), .A2(n14807), .ZN(n15392) );
  AOI21_X1 U11965 ( .B1(n13723), .B2(n13722), .A(n13721), .ZN(n15714) );
  OR2_X1 U11966 ( .A1(n13676), .A2(n13675), .ZN(n13760) );
  OR2_X1 U11967 ( .A1(n13609), .A2(n13608), .ZN(n13631) );
  INV_X1 U11968 ( .A(n15777), .ZN(n13613) );
  AND2_X1 U11969 ( .A1(n13570), .A2(n13569), .ZN(n15800) );
  AND2_X1 U11970 ( .A1(n13538), .A2(n13537), .ZN(n15909) );
  NOR2_X1 U11971 ( .A1(n13518), .A2(n13517), .ZN(n13519) );
  NOR2_X1 U11972 ( .A1(n13481), .A2(n21756), .ZN(n13482) );
  NAND2_X1 U11973 ( .A1(n13482), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13518) );
  OR2_X1 U11974 ( .A1(n13453), .A2(n15826), .ZN(n13481) );
  NAND2_X1 U11975 ( .A1(n13438), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13453) );
  AOI21_X1 U11976 ( .B1(n15821), .B2(n13757), .A(n13451), .ZN(n15817) );
  AND2_X1 U11977 ( .A1(n13437), .A2(n13436), .ZN(n15942) );
  NAND2_X1 U11978 ( .A1(n13405), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13420) );
  NOR2_X1 U11979 ( .A1(n13369), .A2(n15262), .ZN(n13374) );
  OR2_X1 U11980 ( .A1(n15147), .A2(n13357), .ZN(n13358) );
  AND2_X1 U11981 ( .A1(n13329), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13343) );
  AND3_X1 U11982 ( .A1(n13326), .A2(n13325), .A3(n13324), .ZN(n13327) );
  INV_X1 U11983 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13312) );
  NAND2_X1 U11984 ( .A1(n13292), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13313) );
  NAND2_X1 U11985 ( .A1(n13287), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13291) );
  AND2_X1 U11986 ( .A1(n13277), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13287) );
  CLKBUF_X1 U11987 ( .A(n14884), .Z(n14909) );
  NAND2_X1 U11988 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U11989 ( .A1(n12204), .A2(n11086), .ZN(n11402) );
  AND2_X1 U11990 ( .A1(n15803), .A2(n11114), .ZN(n15748) );
  INV_X1 U11991 ( .A(n15747), .ZN(n11305) );
  NAND2_X1 U11992 ( .A1(n15803), .A2(n11104), .ZN(n15760) );
  NAND2_X1 U11993 ( .A1(n15803), .A2(n11307), .ZN(n15772) );
  NAND2_X1 U11994 ( .A1(n15803), .A2(n15789), .ZN(n15788) );
  NOR2_X1 U11995 ( .A1(n15912), .A2(n15801), .ZN(n15803) );
  OR2_X1 U11996 ( .A1(n15920), .A2(n15910), .ZN(n15912) );
  NAND2_X1 U11997 ( .A1(n11404), .A2(n11044), .ZN(n11207) );
  NAND2_X1 U11998 ( .A1(n15924), .A2(n15918), .ZN(n15920) );
  AND2_X1 U11999 ( .A1(n15930), .A2(n15922), .ZN(n15924) );
  NOR2_X1 U12000 ( .A1(n15867), .A2(n12342), .ZN(n15944) );
  OR2_X1 U12001 ( .A1(n15865), .A2(n15864), .ZN(n15867) );
  NAND2_X1 U12002 ( .A1(n20231), .A2(n21556), .ZN(n11199) );
  NAND2_X1 U12003 ( .A1(n15257), .A2(n15331), .ZN(n15865) );
  AND2_X1 U12004 ( .A1(n15154), .A2(n15256), .ZN(n15257) );
  AND2_X1 U12005 ( .A1(n12327), .A2(n12326), .ZN(n15155) );
  INV_X1 U12006 ( .A(n21633), .ZN(n21534) );
  NAND2_X1 U12007 ( .A1(n15126), .A2(n11298), .ZN(n15156) );
  NAND2_X1 U12008 ( .A1(n15126), .A2(n15125), .ZN(n15135) );
  NOR2_X1 U12009 ( .A1(n15116), .A2(n15115), .ZN(n15126) );
  INV_X1 U12010 ( .A(n14913), .ZN(n11314) );
  NAND2_X1 U12011 ( .A1(n20153), .A2(n20152), .ZN(n20151) );
  OR2_X1 U12012 ( .A1(n14706), .A2(n14705), .ZN(n14730) );
  AND2_X1 U12013 ( .A1(n12417), .A2(n16266), .ZN(n21554) );
  NAND2_X1 U12014 ( .A1(n12415), .A2(n14397), .ZN(n21501) );
  OR2_X1 U12015 ( .A1(n21551), .A2(n21575), .ZN(n21633) );
  AND2_X1 U12016 ( .A1(n13764), .A2(n12381), .ZN(n14520) );
  NAND2_X1 U12017 ( .A1(n12415), .A2(n17118), .ZN(n21608) );
  OAI211_X1 U12018 ( .C1(n12263), .C2(n12012), .A(n12011), .B(n12010), .ZN(
        n12103) );
  AOI21_X1 U12019 ( .B1(n12104), .B2(n12103), .A(n12100), .ZN(n13257) );
  OAI21_X1 U12020 ( .B1(n12022), .B2(n12023), .A(n12027), .ZN(n12028) );
  NAND2_X1 U12021 ( .A1(n12120), .A2(n12118), .ZN(n12129) );
  INV_X1 U12022 ( .A(n14749), .ZN(n14741) );
  OR2_X1 U12023 ( .A1(n21953), .A2(n21977), .ZN(n21930) );
  NAND2_X1 U12024 ( .A1(n14693), .A2(n15108), .ZN(n21993) );
  AOI21_X1 U12025 ( .B1(n11031), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n11867), .ZN(n11868) );
  AND3_X1 U12026 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21832), .A3(n14673), 
        .ZN(n14750) );
  NAND2_X1 U12027 ( .A1(n20236), .A2(n14732), .ZN(n14747) );
  NAND2_X1 U12028 ( .A1(n20236), .A2(n14789), .ZN(n14748) );
  NAND2_X1 U12029 ( .A1(n17154), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17148) );
  NAND2_X2 U12030 ( .A1(n13931), .A2(n16336), .ZN(n13861) );
  NAND2_X1 U12031 ( .A1(n16877), .A2(n11102), .ZN(n16842) );
  NAND2_X1 U12032 ( .A1(n16877), .A2(n11106), .ZN(n16844) );
  NOR2_X1 U12033 ( .A1(n11425), .A2(n11423), .ZN(n11422) );
  OR2_X1 U12034 ( .A1(n12941), .A2(n11108), .ZN(n11425) );
  NAND2_X1 U12035 ( .A1(n11424), .A2(n12936), .ZN(n11423) );
  NAND2_X1 U12036 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16307), .ZN(
        n16306) );
  NAND2_X1 U12037 ( .A1(n11418), .A2(n11417), .ZN(n11416) );
  NOR2_X1 U12038 ( .A1(n12961), .A2(n11419), .ZN(n11417) );
  AND2_X1 U12039 ( .A1(n14106), .A2(n14105), .ZN(n16999) );
  NAND2_X1 U12040 ( .A1(n12911), .A2(n11414), .ZN(n13858) );
  INV_X1 U12041 ( .A(n14441), .ZN(n11431) );
  AND2_X1 U12042 ( .A1(n13104), .A2(n13103), .ZN(n16464) );
  AND2_X1 U12043 ( .A1(n13089), .A2(n13088), .ZN(n15205) );
  NAND2_X1 U12044 ( .A1(n14863), .A2(n11087), .ZN(n11437) );
  INV_X1 U12045 ( .A(n16491), .ZN(n11384) );
  AND2_X1 U12046 ( .A1(n16512), .A2(n16511), .ZN(n16514) );
  NAND2_X1 U12047 ( .A1(n16418), .A2(n16420), .ZN(n16419) );
  INV_X1 U12048 ( .A(n11443), .ZN(n11441) );
  NAND2_X1 U12049 ( .A1(n16554), .A2(n11377), .ZN(n11376) );
  AND2_X1 U12050 ( .A1(n15362), .A2(n15361), .ZN(n15364) );
  OR2_X1 U12051 ( .A1(n15201), .A2(n15200), .ZN(n15204) );
  CLKBUF_X1 U12052 ( .A(n15283), .Z(n15203) );
  NOR2_X1 U12053 ( .A1(n15582), .A2(n19711), .ZN(n15427) );
  AND2_X1 U12054 ( .A1(n19556), .A2(n14574), .ZN(n15698) );
  NOR2_X1 U12055 ( .A1(n14424), .A2(n21893), .ZN(n17512) );
  AOI21_X1 U12056 ( .B1(n14423), .B2(n14422), .A(n14369), .ZN(n14424) );
  INV_X1 U12057 ( .A(n14361), .ZN(n15695) );
  AND2_X1 U12058 ( .A1(n16452), .A2(n11116), .ZN(n16422) );
  INV_X1 U12059 ( .A(n16421), .ZN(n11359) );
  AND2_X1 U12060 ( .A1(n13117), .A2(n13116), .ZN(n16429) );
  NAND2_X1 U12061 ( .A1(n16452), .A2(n11105), .ZN(n16431) );
  NAND2_X1 U12062 ( .A1(n16452), .A2(n11361), .ZN(n16438) );
  AND2_X1 U12063 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13142), .ZN(
        n16313) );
  NAND2_X1 U12064 ( .A1(n16313), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16312) );
  NAND2_X1 U12065 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16311), .ZN(
        n16310) );
  NOR2_X1 U12066 ( .A1(n18622), .A2(n16306), .ZN(n16309) );
  NAND2_X1 U12067 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16309), .ZN(
        n16308) );
  AND2_X1 U12068 ( .A1(n13098), .A2(n13097), .ZN(n15348) );
  NOR2_X1 U12069 ( .A1(n18604), .A2(n16304), .ZN(n16307) );
  INV_X1 U12070 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18604) );
  INV_X1 U12071 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16745) );
  INV_X1 U12072 ( .A(n15079), .ZN(n13080) );
  NAND2_X1 U12073 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16301), .ZN(
        n16300) );
  NOR2_X1 U12074 ( .A1(n11054), .A2(n11354), .ZN(n11353) );
  INV_X1 U12075 ( .A(n14873), .ZN(n11354) );
  AND2_X1 U12076 ( .A1(n13064), .A2(n13063), .ZN(n14865) );
  NOR2_X1 U12077 ( .A1(n15320), .A2(n16296), .ZN(n16299) );
  NAND2_X1 U12078 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16297), .ZN(
        n16296) );
  NOR2_X1 U12079 ( .A1(n17414), .A2(n16294), .ZN(n16297) );
  NAND2_X1 U12080 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16295), .ZN(
        n16294) );
  NAND2_X1 U12081 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16293) );
  NOR2_X1 U12082 ( .A1(n17400), .A2(n16293), .ZN(n16295) );
  NAND2_X1 U12083 ( .A1(n10987), .A2(n11339), .ZN(n11333) );
  INV_X1 U12084 ( .A(n16578), .ZN(n11334) );
  NAND2_X1 U12085 ( .A1(n16768), .A2(n16761), .ZN(n11372) );
  AND3_X1 U12086 ( .A1(n18777), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13859), .ZN(n16575) );
  AND2_X1 U12087 ( .A1(n13012), .A2(n16798), .ZN(n16619) );
  NAND2_X1 U12088 ( .A1(n12992), .A2(n16632), .ZN(n16621) );
  AOI21_X1 U12089 ( .B1(n16644), .B2(n11180), .A(n11070), .ZN(n11179) );
  INV_X1 U12090 ( .A(n12983), .ZN(n11180) );
  INV_X1 U12091 ( .A(n16644), .ZN(n11181) );
  AND2_X1 U12092 ( .A1(n16452), .A2(n16444), .ZN(n16445) );
  AND2_X1 U12093 ( .A1(n16662), .A2(n12947), .ZN(n16715) );
  NAND2_X1 U12094 ( .A1(n11242), .A2(n11240), .ZN(n16716) );
  AOI21_X1 U12095 ( .B1(n11243), .B2(n11247), .A(n11241), .ZN(n11240) );
  INV_X1 U12096 ( .A(n16660), .ZN(n11241) );
  INV_X1 U12097 ( .A(n13183), .ZN(n16959) );
  NAND2_X1 U12098 ( .A1(n11245), .A2(n11246), .ZN(n16744) );
  OR2_X1 U12099 ( .A1(n16659), .A2(n11247), .ZN(n11245) );
  INV_X1 U12100 ( .A(n12955), .ZN(n16995) );
  AND2_X1 U12101 ( .A1(n12928), .A2(n17016), .ZN(n17009) );
  AND2_X1 U12102 ( .A1(n14053), .A2(n14052), .ZN(n18556) );
  INV_X1 U12103 ( .A(n14476), .ZN(n13053) );
  NAND2_X1 U12104 ( .A1(n15213), .A2(n15214), .ZN(n11321) );
  OR2_X1 U12105 ( .A1(n14234), .A2(n14206), .ZN(n16917) );
  NAND2_X1 U12106 ( .A1(n18452), .A2(n14438), .ZN(n14405) );
  AOI21_X1 U12107 ( .B1(n18470), .B2(n14438), .A(n14414), .ZN(n14416) );
  XNOR2_X1 U12108 ( .A(n14447), .B(n14445), .ZN(n14434) );
  NAND2_X1 U12109 ( .A1(n11001), .A2(n12648), .ZN(n14462) );
  BUF_X1 U12110 ( .A(n12834), .Z(n19534) );
  INV_X1 U12111 ( .A(n19414), .ZN(n19452) );
  INV_X1 U12112 ( .A(n19462), .ZN(n19458) );
  INV_X1 U12113 ( .A(n19440), .ZN(n19498) );
  INV_X1 U12114 ( .A(n19446), .ZN(n19443) );
  NAND3_X1 U12115 ( .A1(n15697), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19511), 
        .ZN(n19559) );
  NAND3_X1 U12116 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n15695), .A3(n19511), 
        .ZN(n19560) );
  NAND2_X1 U12117 ( .A1(n19420), .A2(n19865), .ZN(n19440) );
  NAND2_X1 U12118 ( .A1(n12666), .A2(n12648), .ZN(n12675) );
  INV_X1 U12119 ( .A(n19559), .ZN(n19875) );
  INV_X1 U12120 ( .A(n19560), .ZN(n19876) );
  NAND2_X1 U12121 ( .A1(n18471), .A2(n19865), .ZN(n19467) );
  AND2_X1 U12122 ( .A1(n11140), .A2(n11139), .ZN(n11612) );
  NOR2_X1 U12123 ( .A1(n11610), .A2(n11609), .ZN(n11139) );
  INV_X1 U12124 ( .A(n11608), .ZN(n11140) );
  NOR2_X1 U12125 ( .A1(n15375), .A2(n20781), .ZN(n21380) );
  NAND2_X1 U12126 ( .A1(n20580), .A2(n11473), .ZN(n14254) );
  NAND2_X1 U12127 ( .A1(n14254), .A2(n18195), .ZN(n14253) );
  NAND2_X1 U12128 ( .A1(n11661), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11662) );
  AND2_X1 U12129 ( .A1(n20312), .A2(n15375), .ZN(n17091) );
  INV_X1 U12130 ( .A(n18398), .ZN(n18399) );
  NOR2_X1 U12131 ( .A1(n21379), .A2(n20322), .ZN(n20324) );
  NOR2_X1 U12132 ( .A1(n20763), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11257) );
  NOR2_X1 U12133 ( .A1(n13823), .A2(n20374), .ZN(n11778) );
  AND2_X1 U12134 ( .A1(n18103), .A2(n11115), .ZN(n11771) );
  NAND2_X1 U12135 ( .A1(n18103), .A2(n11038), .ZN(n18131) );
  NOR2_X1 U12136 ( .A1(n18091), .A2(n21283), .ZN(n18101) );
  NAND2_X1 U12137 ( .A1(n17976), .A2(n11266), .ZN(n18088) );
  AND2_X1 U12138 ( .A1(n11049), .A2(n11098), .ZN(n11266) );
  NAND2_X1 U12139 ( .A1(n17976), .A2(n11267), .ZN(n18076) );
  NAND2_X1 U12140 ( .A1(n17976), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17991) );
  NOR2_X1 U12141 ( .A1(n18183), .A2(n18182), .ZN(n17976) );
  NAND2_X1 U12142 ( .A1(n18213), .A2(n11082), .ZN(n17997) );
  AND2_X1 U12143 ( .A1(n18213), .A2(n11264), .ZN(n18199) );
  NAND2_X1 U12144 ( .A1(n18213), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18029) );
  NOR2_X1 U12145 ( .A1(n18269), .A2(n11719), .ZN(n18260) );
  NAND2_X1 U12146 ( .A1(n18285), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20482) );
  NOR2_X1 U12147 ( .A1(n20406), .A2(n18297), .ZN(n18285) );
  AOI22_X2 U12148 ( .A1(n13213), .A2(n21384), .B1(n21382), .B2(n21084), .ZN(
        n21407) );
  NOR2_X1 U12149 ( .A1(n21283), .A2(n21272), .ZN(n18107) );
  NOR2_X1 U12150 ( .A1(n11760), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11761) );
  NAND2_X1 U12151 ( .A1(n18196), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21311) );
  AND2_X1 U12152 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21188), .ZN(
        n21177) );
  NOR2_X1 U12153 ( .A1(n13191), .A2(n21122), .ZN(n11286) );
  NOR2_X1 U12154 ( .A1(n18260), .A2(n11287), .ZN(n18027) );
  AND2_X1 U12155 ( .A1(n13191), .A2(n21122), .ZN(n11287) );
  NAND2_X1 U12156 ( .A1(n18248), .A2(n11748), .ZN(n21132) );
  INV_X1 U12157 ( .A(n11740), .ZN(n11195) );
  NAND2_X1 U12158 ( .A1(n18280), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18279) );
  INV_X1 U12159 ( .A(n11712), .ZN(n11711) );
  NAND2_X1 U12160 ( .A1(n18301), .A2(n11738), .ZN(n18292) );
  AND2_X1 U12161 ( .A1(n18290), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18296) );
  NAND2_X1 U12162 ( .A1(n20779), .A2(n21285), .ZN(n21381) );
  OAI21_X1 U12163 ( .B1(n11617), .B2(n11619), .A(n11616), .ZN(n13200) );
  NOR2_X1 U12164 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20379), .ZN(
        n20380) );
  NOR2_X1 U12165 ( .A1(n21011), .A2(n11794), .ZN(n21019) );
  NOR2_X1 U12166 ( .A1(n15375), .A2(n11222), .ZN(n21002) );
  NAND2_X1 U12167 ( .A1(n11795), .A2(n11083), .ZN(n11222) );
  NOR2_X1 U12168 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18941), .ZN(n19265) );
  INV_X1 U12169 ( .A(n11606), .ZN(n19135) );
  INV_X1 U12170 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18980) );
  INV_X1 U12171 ( .A(n17576), .ZN(n19095) );
  NOR2_X1 U12172 ( .A1(n11567), .A2(n11566), .ZN(n20840) );
  NOR2_X1 U12173 ( .A1(n11573), .A2(n11224), .ZN(n11223) );
  INV_X1 U12174 ( .A(n19265), .ZN(n19176) );
  AOI211_X1 U12175 ( .C1(n17914), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n11584), .B(n11583), .ZN(n11585) );
  NOR2_X1 U12176 ( .A1(n11303), .A2(n11302), .ZN(n11301) );
  INV_X1 U12177 ( .A(n15720), .ZN(n11302) );
  INV_X1 U12178 ( .A(n15721), .ZN(n11303) );
  OR2_X1 U12179 ( .A1(n15718), .A2(n21812), .ZN(n11304) );
  INV_X1 U12180 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15826) );
  INV_X1 U12181 ( .A(n21781), .ZN(n21804) );
  INV_X1 U12182 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15839) );
  INV_X1 U12183 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15863) );
  INV_X1 U12184 ( .A(n21732), .ZN(n21721) );
  INV_X1 U12185 ( .A(n21820), .ZN(n21792) );
  OR2_X1 U12186 ( .A1(n21720), .A2(n15151), .ZN(n21795) );
  INV_X1 U12187 ( .A(n21690), .ZN(n21679) );
  INV_X1 U12188 ( .A(n20136), .ZN(n15949) );
  AND2_X2 U12189 ( .A1(n14515), .A2(n15390), .ZN(n20136) );
  NAND2_X1 U12190 ( .A1(n14551), .A2(n14514), .ZN(n14515) );
  INV_X1 U12191 ( .A(n16030), .ZN(n15960) );
  INV_X1 U12192 ( .A(n15955), .ZN(n16007) );
  INV_X1 U12193 ( .A(n16014), .ZN(n16021) );
  AND2_X1 U12194 ( .A1(n13737), .A2(n15390), .ZN(n16015) );
  OR2_X1 U12195 ( .A1(n14554), .A2(n13736), .ZN(n13737) );
  OR2_X1 U12196 ( .A1(n16019), .A2(n14483), .ZN(n16014) );
  NOR2_X1 U12197 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17152), .ZN(n20053) );
  INV_X1 U12198 ( .A(n20230), .ZN(n16114) );
  INV_X1 U12199 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n21756) );
  NAND2_X1 U12200 ( .A1(n15290), .A2(n15289), .ZN(n15288) );
  NAND2_X1 U12201 ( .A1(n20177), .A2(n12178), .ZN(n15290) );
  AND2_X2 U12202 ( .A1(n21822), .A2(n13811), .ZN(n20230) );
  NAND2_X1 U12203 ( .A1(n11401), .A2(n12204), .ZN(n16064) );
  AOI21_X1 U12204 ( .B1(n21500), .B2(n21575), .A(n21555), .ZN(n21549) );
  NAND2_X1 U12205 ( .A1(n20165), .A2(n12155), .ZN(n20172) );
  NOR2_X1 U12206 ( .A1(n14706), .A2(n11316), .ZN(n14889) );
  OR2_X1 U12207 ( .A1(n14728), .A2(n14705), .ZN(n11316) );
  AND2_X1 U12208 ( .A1(n21551), .A2(n21631), .ZN(n21573) );
  INV_X1 U12209 ( .A(n22077), .ZN(n22043) );
  INV_X1 U12210 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21944) );
  OAI21_X1 U12211 ( .B1(n15023), .B2(n21835), .A(n21924), .ZN(n17155) );
  AND2_X1 U12212 ( .A1(n12208), .A2(n14749), .ZN(n17118) );
  NOR2_X1 U12213 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n17081) );
  OAI21_X1 U12214 ( .B1(n15047), .B2(n15048), .A(n22057), .ZN(n15072) );
  OAI211_X1 U12215 ( .C1(n22341), .C2(n22021), .A(n21985), .B(n22002), .ZN(
        n22344) );
  NOR2_X2 U12216 ( .A1(n21993), .A2(n22037), .ZN(n22355) );
  OAI21_X1 U12217 ( .B1(n22009), .B2(n22008), .A(n22007), .ZN(n22356) );
  OR2_X1 U12218 ( .A1(n21993), .A2(n15043), .ZN(n14812) );
  NOR2_X1 U12219 ( .A1(n21924), .A2(n14771), .ZN(n22048) );
  INV_X1 U12220 ( .A(n22113), .ZN(n22107) );
  NOR2_X1 U12221 ( .A1(n21924), .A2(n14769), .ZN(n22106) );
  INV_X1 U12222 ( .A(n22150), .ZN(n22144) );
  NOR2_X1 U12223 ( .A1(n21924), .A2(n14811), .ZN(n22143) );
  INV_X1 U12224 ( .A(n22187), .ZN(n22181) );
  NOR2_X1 U12225 ( .A1(n21924), .A2(n14838), .ZN(n22180) );
  INV_X1 U12226 ( .A(n22225), .ZN(n22219) );
  NOR2_X1 U12227 ( .A1(n21924), .A2(n14893), .ZN(n22218) );
  NOR2_X1 U12228 ( .A1(n21924), .A2(n14915), .ZN(n22255) );
  INV_X1 U12229 ( .A(n22299), .ZN(n22293) );
  NOR2_X1 U12230 ( .A1(n21924), .A2(n14978), .ZN(n22292) );
  INV_X1 U12231 ( .A(n22386), .ZN(n22376) );
  NOR2_X1 U12232 ( .A1(n21924), .A2(n15130), .ZN(n22374) );
  OAI211_X1 U12233 ( .C1(n22375), .C2(n22058), .A(n22057), .B(n22056), .ZN(
        n22379) );
  AND2_X1 U12234 ( .A1(n22042), .A2(n22038), .ZN(n22378) );
  INV_X1 U12235 ( .A(n22048), .ZN(n22069) );
  INV_X1 U12236 ( .A(n22106), .ZN(n22112) );
  INV_X1 U12237 ( .A(n22143), .ZN(n22149) );
  INV_X1 U12238 ( .A(n22218), .ZN(n22224) );
  INV_X1 U12239 ( .A(n22255), .ZN(n22261) );
  INV_X1 U12240 ( .A(n22292), .ZN(n22298) );
  INV_X1 U12241 ( .A(n22374), .ZN(n22383) );
  OR2_X1 U12242 ( .A1(n17148), .A2(n21832), .ZN(n21844) );
  INV_X1 U12243 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n17154) );
  INV_X1 U12244 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21873) );
  NAND2_X1 U12245 ( .A1(n18791), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18765) );
  XNOR2_X1 U12246 ( .A(n12995), .B(n12994), .ZN(n18734) );
  AOI21_X1 U12247 ( .B1(n12984), .B2(n12985), .A(n12989), .ZN(n11410) );
  NOR2_X1 U12248 ( .A1(n12934), .A2(n12933), .ZN(n12952) );
  INV_X1 U12249 ( .A(n18788), .ZN(n18774) );
  INV_X1 U12250 ( .A(n18795), .ZN(n18780) );
  AND2_X1 U12251 ( .A1(n16290), .A2(n16332), .ZN(n18796) );
  INV_X1 U12252 ( .A(n18765), .ZN(n18794) );
  AND2_X1 U12253 ( .A1(n14142), .A2(n14141), .ZN(n15230) );
  CLKBUF_X1 U12254 ( .A(n15188), .Z(n15144) );
  AND2_X1 U12255 ( .A1(n13930), .A2(n13929), .ZN(n15083) );
  CLKBUF_X1 U12256 ( .A(n15084), .Z(n14929) );
  AND2_X1 U12257 ( .A1(n14410), .A2(n18907), .ZN(n16448) );
  OAI21_X1 U12258 ( .B1(n16454), .B2(n11442), .A(n15542), .ZN(n16428) );
  INV_X1 U12259 ( .A(n19860), .ZN(n19549) );
  NAND2_X1 U12260 ( .A1(n19556), .A2(n14573), .ZN(n16564) );
  AND2_X1 U12261 ( .A1(n15698), .A2(n15697), .ZN(n19764) );
  NAND2_X1 U12262 ( .A1(n14571), .A2(n14570), .ZN(n19556) );
  NAND2_X1 U12263 ( .A1(n14569), .A2(n18907), .ZN(n14571) );
  NAND2_X1 U12264 ( .A1(n11379), .A2(n11383), .ZN(n18477) );
  NAND2_X1 U12265 ( .A1(n19556), .A2(n14572), .ZN(n19812) );
  INV_X1 U12266 ( .A(n17481), .ZN(n19865) );
  AND2_X1 U12267 ( .A1(n19556), .A2(n14575), .ZN(n19860) );
  INV_X1 U12268 ( .A(n19556), .ZN(n19859) );
  CLKBUF_X1 U12269 ( .A(n17529), .Z(n17537) );
  NOR2_X1 U12271 ( .A1(n17512), .A2(n17538), .ZN(n17529) );
  NAND2_X1 U12272 ( .A1(n16583), .A2(n11273), .ZN(n11272) );
  NOR2_X1 U12273 ( .A1(n17463), .A2(n11275), .ZN(n11273) );
  NAND2_X1 U12274 ( .A1(n16734), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16920) );
  INV_X1 U12275 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17460) );
  NAND2_X1 U12276 ( .A1(n15316), .A2(n13177), .ZN(n17432) );
  INV_X1 U12277 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17400) );
  INV_X1 U12278 ( .A(n17461), .ZN(n17475) );
  AND2_X1 U12279 ( .A1(n17459), .A2(n14301), .ZN(n17453) );
  NAND2_X1 U12280 ( .A1(n16645), .A2(n16644), .ZN(n16643) );
  NAND2_X1 U12281 ( .A1(n16648), .A2(n12983), .ZN(n16645) );
  NAND2_X1 U12282 ( .A1(n11341), .A2(n11342), .ZN(n16650) );
  NOR2_X1 U12283 ( .A1(n11039), .A2(n16945), .ZN(n16349) );
  NAND2_X1 U12284 ( .A1(n11349), .A2(n12921), .ZN(n17030) );
  NAND2_X1 U12285 ( .A1(n11215), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17415) );
  INV_X1 U12286 ( .A(n10997), .ZN(n15236) );
  OR2_X1 U12287 ( .A1(n14234), .A2(n14176), .ZN(n18870) );
  NAND2_X1 U12288 ( .A1(n16912), .A2(n16917), .ZN(n18808) );
  INV_X1 U12289 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19488) );
  INV_X1 U12290 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n17490) );
  INV_X1 U12291 ( .A(n18471), .ZN(n19420) );
  AND2_X1 U12292 ( .A1(n14647), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18897) );
  INV_X1 U12293 ( .A(n19965), .ZN(n19846) );
  OAI21_X1 U12294 ( .B1(n19505), .B2(n19504), .A(n19503), .ZN(n19934) );
  INV_X1 U12295 ( .A(n19913), .ZN(n19915) );
  OAI21_X1 U12296 ( .B1(n19449), .B2(n19448), .A(n19447), .ZN(n19909) );
  OR2_X1 U12297 ( .A1(n14984), .A2(n14983), .ZN(n19903) );
  INV_X1 U12298 ( .A(n19889), .ZN(n19899) );
  INV_X1 U12299 ( .A(n19958), .ZN(n19976) );
  INV_X1 U12300 ( .A(n19842), .ZN(n19854) );
  INV_X1 U12301 ( .A(n19791), .ZN(n19803) );
  INV_X1 U12302 ( .A(n19749), .ZN(n19756) );
  AOI22_X1 U12303 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19875), .ZN(n19655) );
  INV_X1 U12304 ( .A(n19635), .ZN(n19652) );
  INV_X1 U12305 ( .A(n19426), .ZN(n19543) );
  AND2_X1 U12306 ( .A1(n15031), .A2(n15030), .ZN(n19802) );
  AND2_X1 U12307 ( .A1(n14857), .A2(n15030), .ZN(n19650) );
  NOR2_X2 U12308 ( .A1(n19421), .A2(n19467), .ZN(n19975) );
  AND2_X1 U12309 ( .A1(n12687), .A2(n15030), .ZN(n19531) );
  NAND2_X1 U12310 ( .A1(n19492), .A2(n19397), .ZN(n19886) );
  XNOR2_X1 U12311 ( .A(n20779), .B(n20370), .ZN(n20314) );
  INV_X1 U12312 ( .A(n21907), .ZN(n21900) );
  NAND2_X1 U12313 ( .A1(n20725), .A2(n20726), .ZN(n20724) );
  NAND2_X1 U12314 ( .A1(n20713), .A2(n20714), .ZN(n20712) );
  NAND2_X1 U12315 ( .A1(n20625), .A2(n20580), .ZN(n20640) );
  NAND2_X1 U12316 ( .A1(n20640), .A2(n20641), .ZN(n20639) );
  NAND2_X1 U12317 ( .A1(n20615), .A2(n20580), .ZN(n20626) );
  NAND2_X1 U12318 ( .A1(n20626), .A2(n20627), .ZN(n20625) );
  NAND2_X1 U12319 ( .A1(n20616), .A2(n20617), .ZN(n20615) );
  NOR2_X1 U12320 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n20591), .ZN(n20597) );
  NOR2_X1 U12321 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n20539), .ZN(n20563) );
  INV_X1 U12322 ( .A(n21422), .ZN(n20741) );
  INV_X1 U12323 ( .A(n20456), .ZN(n20492) );
  INV_X1 U12324 ( .A(n20764), .ZN(n20727) );
  INV_X1 U12325 ( .A(n20749), .ZN(n20765) );
  INV_X1 U12326 ( .A(n20430), .ZN(n20768) );
  NOR2_X1 U12327 ( .A1(n20677), .A2(n17865), .ZN(n17870) );
  NOR2_X1 U12328 ( .A1(n17962), .A2(n17958), .ZN(n17918) );
  INV_X1 U12329 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17815) );
  INV_X1 U12330 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17891) );
  INV_X1 U12331 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17905) );
  NOR2_X1 U12332 ( .A1(n20914), .A2(n20915), .ZN(n20913) );
  NAND2_X1 U12333 ( .A1(n20891), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n20914) );
  NOR2_X1 U12334 ( .A1(n20923), .A2(n20885), .ZN(n20891) );
  OR2_X1 U12335 ( .A1(n20921), .A2(n20922), .ZN(n20923) );
  NOR2_X1 U12336 ( .A1(n20931), .A2(n20930), .ZN(n20929) );
  NOR2_X1 U12337 ( .A1(n20878), .A2(n20877), .ZN(n20873) );
  INV_X1 U12338 ( .A(n20873), .ZN(n20879) );
  NOR2_X1 U12339 ( .A1(n20952), .A2(n20941), .ZN(n20940) );
  INV_X1 U12340 ( .A(n20933), .ZN(n20939) );
  NAND2_X1 U12341 ( .A1(n20953), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n20952) );
  NOR2_X1 U12342 ( .A1(n20948), .A2(n20947), .ZN(n20953) );
  NOR2_X1 U12343 ( .A1(n20785), .A2(n20801), .ZN(n20798) );
  INV_X1 U12344 ( .A(n20814), .ZN(n20964) );
  AOI21_X1 U12345 ( .B1(n20782), .B2(n20781), .A(n20780), .ZN(n20966) );
  NOR2_X1 U12346 ( .A1(n11501), .A2(n11500), .ZN(n20812) );
  NOR2_X1 U12347 ( .A1(n20958), .A2(n20975), .ZN(n20814) );
  INV_X1 U12348 ( .A(n20823), .ZN(n20832) );
  AND2_X1 U12349 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n20834), .ZN(n20838) );
  AOI211_X1 U12350 ( .C1(n11661), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n11697), .B(n11696), .ZN(n11698) );
  INV_X1 U12351 ( .A(n20839), .ZN(n20973) );
  NOR2_X1 U12352 ( .A1(n20364), .A2(n20324), .ZN(n20357) );
  CLKBUF_X1 U12353 ( .A(n20357), .Z(n20363) );
  INV_X1 U12354 ( .A(n11294), .ZN(n18126) );
  OAI21_X1 U12355 ( .B1(n18143), .B2(n18258), .A(n13190), .ZN(n11294) );
  NAND2_X1 U12356 ( .A1(n18103), .A2(n11047), .ZN(n18151) );
  NAND2_X1 U12357 ( .A1(n18213), .A2(n11262), .ZN(n18183) );
  AND2_X1 U12358 ( .A1(n11082), .A2(n11263), .ZN(n11262) );
  INV_X1 U12359 ( .A(n18015), .ZN(n11263) );
  INV_X1 U12360 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20496) );
  AOI22_X1 U12361 ( .A1(n21135), .A2(n18262), .B1(n18275), .B2(n21132), .ZN(
        n18247) );
  NAND2_X1 U12362 ( .A1(n18307), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20406) );
  AND2_X1 U12363 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18307) );
  INV_X1 U12364 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20401) );
  NAND2_X1 U12365 ( .A1(n18181), .A2(n18180), .ZN(n18321) );
  INV_X1 U12366 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20378) );
  INV_X1 U12367 ( .A(n18321), .ZN(n18342) );
  NAND2_X1 U12368 ( .A1(n11191), .A2(n21260), .ZN(n21262) );
  INV_X1 U12369 ( .A(n18091), .ZN(n21269) );
  INV_X1 U12370 ( .A(n11280), .ZN(n18185) );
  NAND2_X1 U12371 ( .A1(n11759), .A2(n11756), .ZN(n18186) );
  NOR2_X1 U12372 ( .A1(n18205), .A2(n18204), .ZN(n21188) );
  INV_X1 U12373 ( .A(n21075), .ZN(n21363) );
  NOR2_X1 U12374 ( .A1(n21112), .A2(n21111), .ZN(n21140) );
  INV_X1 U12375 ( .A(n21381), .ZN(n21084) );
  INV_X1 U12376 ( .A(n11706), .ZN(n11291) );
  INV_X1 U12377 ( .A(n11292), .ZN(n18314) );
  INV_X1 U12378 ( .A(n21367), .ZN(n21162) );
  INV_X1 U12379 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21398) );
  INV_X1 U12380 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17090) );
  INV_X1 U12381 ( .A(n20380), .ZN(n20995) );
  INV_X2 U12382 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21029) );
  NAND2_X1 U12383 ( .A1(n11146), .A2(n11141), .ZN(n21434) );
  AOI21_X1 U12384 ( .B1(n21410), .B2(n21411), .A(n11142), .ZN(n11141) );
  NOR2_X1 U12385 ( .A1(n21438), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n21419) );
  CLKBUF_X1 U12386 ( .A(n18937), .Z(n19261) );
  NAND2_X1 U12387 ( .A1(n11132), .A2(n11131), .ZN(P1_U2810) );
  AND2_X1 U12388 ( .A1(n11300), .A2(n11304), .ZN(n11131) );
  NAND2_X1 U12389 ( .A1(n16030), .A2(n21771), .ZN(n11132) );
  NOR2_X1 U12390 ( .A1(n15719), .A2(n11301), .ZN(n11300) );
  AND2_X1 U12391 ( .A1(n12425), .A2(n12424), .ZN(n12426) );
  CLKBUF_X1 U12392 ( .A(n14861), .Z(n14598) );
  INV_X1 U12393 ( .A(n11220), .ZN(n16573) );
  OAI211_X1 U12394 ( .C1(n16760), .C2(n17461), .A(n11271), .B(n11270), .ZN(
        P2_U2984) );
  AND2_X1 U12395 ( .A1(n11274), .A2(n11272), .ZN(n11271) );
  NAND2_X1 U12396 ( .A1(n11072), .A2(n16584), .ZN(n11270) );
  AOI21_X1 U12397 ( .B1(n18797), .B2(n17474), .A(n16585), .ZN(n11274) );
  AOI21_X1 U12398 ( .B1(n18775), .B2(n17474), .A(n13146), .ZN(n13147) );
  INV_X1 U12399 ( .A(n11323), .ZN(n11328) );
  INV_X1 U12400 ( .A(n11338), .ZN(n11337) );
  INV_X1 U12401 ( .A(n11329), .ZN(n11327) );
  NOR2_X1 U12402 ( .A1(n11159), .A2(n11158), .ZN(n16759) );
  OAI21_X1 U12403 ( .B1(n16758), .B2(n18849), .A(n16757), .ZN(n11158) );
  NOR2_X1 U12404 ( .A1(n16756), .A2(n18881), .ZN(n11159) );
  OAI21_X1 U12405 ( .B1(n16390), .B2(n18849), .A(n11369), .ZN(n11368) );
  INV_X1 U12406 ( .A(n16769), .ZN(n11373) );
  OR2_X1 U12407 ( .A1(n20758), .A2(n11248), .ZN(P3_U2640) );
  OAI211_X1 U12408 ( .C1(n20756), .C2(n11253), .A(n11250), .B(n11249), .ZN(
        n11248) );
  NAND2_X1 U12409 ( .A1(n11255), .A2(n11254), .ZN(n11253) );
  AOI21_X1 U12410 ( .B1(n13838), .B2(n18262), .A(n11193), .ZN(n11192) );
  NAND2_X1 U12411 ( .A1(n18166), .A2(n18167), .ZN(n18179) );
  OR2_X1 U12412 ( .A1(n11777), .A2(n11776), .ZN(P3_U2801) );
  OAI21_X1 U12413 ( .B1(n11775), .B2(n20743), .A(n11774), .ZN(n11776) );
  AOI21_X1 U12414 ( .B1(n13824), .B2(n11773), .A(n21249), .ZN(n11774) );
  AOI21_X1 U12415 ( .B1(n13847), .B2(n21369), .A(n13846), .ZN(n13848) );
  NAND2_X1 U12416 ( .A1(n11191), .A2(n11189), .ZN(n21254) );
  NOR2_X1 U12417 ( .A1(n13225), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13229) );
  OAI21_X1 U12418 ( .B1(n13220), .B2(n13219), .A(n21329), .ZN(n13230) );
  OR2_X1 U12419 ( .A1(n20243), .A2(n20296), .ZN(U212) );
  NAND2_X1 U12420 ( .A1(n15329), .A2(n11128), .ZN(n15831) );
  AND2_X1 U12421 ( .A1(n11048), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11038) );
  AND2_X1 U12422 ( .A1(n20841), .A2(n17576), .ZN(n11040) );
  OR3_X1 U12423 ( .A1(n21407), .A2(n19220), .A3(n11229), .ZN(n11041) );
  AND2_X1 U12424 ( .A1(n15815), .A2(n11463), .ZN(n11042) );
  AND3_X1 U12425 ( .A1(n13297), .A2(n11011), .A3(n11084), .ZN(n11043) );
  OR2_X1 U12426 ( .A1(n15327), .A2(n15855), .ZN(n15845) );
  INV_X1 U12427 ( .A(n11448), .ZN(n15363) );
  INV_X1 U12428 ( .A(n11125), .ZN(n15814) );
  AND2_X1 U12429 ( .A1(n11406), .A2(n12196), .ZN(n11044) );
  NAND2_X1 U12430 ( .A1(n11206), .A2(n15289), .ZN(n11208) );
  INV_X1 U12431 ( .A(n11795), .ZN(n20323) );
  AND2_X1 U12432 ( .A1(n16334), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11045) );
  AND2_X1 U12433 ( .A1(n11383), .A2(n11381), .ZN(n11046) );
  NAND2_X1 U12434 ( .A1(n11436), .A2(n14863), .ZN(n14900) );
  NAND2_X1 U12435 ( .A1(n12021), .A2(n21933), .ZN(n14582) );
  AND2_X1 U12436 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11047) );
  AND2_X1 U12437 ( .A1(n11047), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11048) );
  AND2_X1 U12438 ( .A1(n11267), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11049) );
  NOR2_X1 U12439 ( .A1(n13967), .A2(n11118), .ZN(n11383) );
  INV_X1 U12440 ( .A(n20580), .ZN(n20523) );
  NAND2_X2 U12441 ( .A1(n11260), .A2(n11256), .ZN(n20580) );
  AND2_X2 U12442 ( .A1(n12446), .A2(n15520), .ZN(n12479) );
  OR2_X1 U12443 ( .A1(n16463), .A2(n16464), .ZN(n11050) );
  INV_X1 U12444 ( .A(n12802), .ZN(n12536) );
  OR2_X1 U12445 ( .A1(n12934), .A2(n11416), .ZN(n11051) );
  NOR2_X1 U12446 ( .A1(n21004), .A2(n11494), .ZN(n11525) );
  INV_X1 U12447 ( .A(n20231), .ZN(n11209) );
  XNOR2_X1 U12448 ( .A(n14184), .B(n14183), .ZN(n16289) );
  NAND2_X1 U12449 ( .A1(n11208), .A2(n11391), .ZN(n11483) );
  NAND2_X1 U12450 ( .A1(n15815), .A2(n15933), .ZN(n15928) );
  NAND2_X1 U12451 ( .A1(n16877), .A2(n16876), .ZN(n16538) );
  AND2_X1 U12452 ( .A1(n11349), .A2(n11347), .ZN(n17028) );
  NAND2_X1 U12453 ( .A1(n15315), .A2(n15314), .ZN(n15316) );
  AND2_X1 U12454 ( .A1(n13183), .A2(n11476), .ZN(n11052) );
  INV_X2 U12455 ( .A(n13042), .ZN(n14179) );
  INV_X1 U12456 ( .A(n12753), .ZN(n13042) );
  AND3_X1 U12457 ( .A1(n11855), .A2(n11854), .A3(n11853), .ZN(n11053) );
  AND2_X2 U12458 ( .A1(n11823), .A2(n11818), .ZN(n11909) );
  NAND2_X1 U12459 ( .A1(n11356), .A2(n11355), .ZN(n11054) );
  NAND2_X1 U12460 ( .A1(n16512), .A2(n11386), .ZN(n16497) );
  NAND2_X1 U12461 ( .A1(n11170), .A2(n12914), .ZN(n15299) );
  AND2_X1 U12462 ( .A1(n11188), .A2(n11187), .ZN(n11055) );
  NAND2_X1 U12463 ( .A1(n15815), .A2(n11462), .ZN(n11056) );
  AND2_X1 U12464 ( .A1(n11414), .A2(n11413), .ZN(n11057) );
  OR3_X1 U12465 ( .A1(n12934), .A2(n12933), .A3(n11419), .ZN(n11058) );
  OAI21_X1 U12466 ( .B1(n16648), .B2(n11181), .A(n11179), .ZN(n16630) );
  OR2_X1 U12467 ( .A1(n13013), .A2(n16620), .ZN(n11059) );
  NAND2_X1 U12468 ( .A1(n20231), .A2(n12407), .ZN(n11060) );
  NAND2_X1 U12469 ( .A1(n11204), .A2(n11205), .ZN(n16119) );
  INV_X1 U12470 ( .A(n11924), .ZN(n11926) );
  INV_X1 U12471 ( .A(n21386), .ZN(n21312) );
  NOR2_X2 U12472 ( .A1(n20314), .A2(n17574), .ZN(n21386) );
  XNOR2_X1 U12473 ( .A(n15606), .B(n11465), .ZN(n16413) );
  OR2_X1 U12474 ( .A1(n12938), .A2(n12935), .ZN(n11061) );
  AND2_X1 U12475 ( .A1(n14683), .A2(n14712), .ZN(n11062) );
  NAND2_X1 U12476 ( .A1(n11570), .A2(n11223), .ZN(n19017) );
  INV_X1 U12477 ( .A(n19017), .ZN(n20841) );
  AND2_X1 U12478 ( .A1(n13183), .A2(n11277), .ZN(n11063) );
  AND2_X1 U12479 ( .A1(n16334), .A2(n16277), .ZN(n11064) );
  AND2_X1 U12480 ( .A1(n11334), .A2(n11339), .ZN(n11065) );
  OR2_X1 U12481 ( .A1(n15586), .A2(n16426), .ZN(n11066) );
  NOR2_X1 U12482 ( .A1(n16412), .A2(n16407), .ZN(n16397) );
  OR2_X1 U12483 ( .A1(n13850), .A2(n16575), .ZN(n11067) );
  INV_X1 U12484 ( .A(n11276), .ZN(n16640) );
  NAND2_X1 U12485 ( .A1(n13183), .A2(n11120), .ZN(n11276) );
  OR2_X1 U12486 ( .A1(n16611), .A2(n16619), .ZN(n11068) );
  INV_X1 U12487 ( .A(n13161), .ZN(n12861) );
  NAND2_X1 U12488 ( .A1(n12203), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11403) );
  INV_X1 U12489 ( .A(n11403), .ZN(n11401) );
  INV_X1 U12490 ( .A(n11343), .ZN(n11342) );
  NAND2_X1 U12491 ( .A1(n12978), .A2(n11344), .ZN(n11343) );
  AND2_X1 U12492 ( .A1(n12184), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11069) );
  AND2_X1 U12493 ( .A1(n12986), .A2(n16833), .ZN(n11070) );
  NAND2_X1 U12494 ( .A1(n12209), .A2(n12009), .ZN(n11919) );
  AND2_X1 U12495 ( .A1(n13181), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11071) );
  AND2_X1 U12496 ( .A1(n12909), .A2(n12908), .ZN(n13168) );
  INV_X1 U12497 ( .A(n13168), .ZN(n13173) );
  AND2_X1 U12498 ( .A1(n16583), .A2(n17473), .ZN(n11072) );
  AND2_X1 U12499 ( .A1(n12858), .A2(n12857), .ZN(n12860) );
  INV_X1 U12500 ( .A(n11406), .ZN(n11405) );
  NAND2_X1 U12501 ( .A1(n12195), .A2(n11407), .ZN(n11406) );
  NOR3_X1 U12502 ( .A1(n12938), .A2(n12935), .A3(n12941), .ZN(n11073) );
  AND2_X1 U12503 ( .A1(n12687), .A2(n19472), .ZN(n11074) );
  AND2_X1 U12504 ( .A1(n12204), .A2(n12203), .ZN(n11075) );
  NAND2_X1 U12505 ( .A1(n16419), .A2(n11066), .ZN(n15606) );
  AND2_X1 U12506 ( .A1(n11060), .A2(n12196), .ZN(n11076) );
  OR2_X1 U12507 ( .A1(n13844), .A2(n18351), .ZN(n11077) );
  NOR2_X1 U12508 ( .A1(n14442), .A2(n11431), .ZN(n11078) );
  INV_X1 U12509 ( .A(n15289), .ZN(n11394) );
  INV_X1 U12510 ( .A(n14155), .ZN(n14152) );
  AND2_X2 U12511 ( .A1(n13931), .A2(n19472), .ZN(n14155) );
  INV_X1 U12512 ( .A(n12933), .ZN(n11418) );
  INV_X1 U12513 ( .A(n12935), .ZN(n11424) );
  OR2_X1 U12514 ( .A1(n16454), .A2(n11441), .ZN(n11079) );
  NOR2_X1 U12515 ( .A1(n11039), .A2(n11375), .ZN(n16347) );
  NOR2_X1 U12516 ( .A1(n16454), .A2(n16456), .ZN(n16441) );
  NOR2_X1 U12517 ( .A1(n15283), .A2(n11449), .ZN(n15449) );
  NOR2_X1 U12518 ( .A1(n15327), .A2(n11455), .ZN(n15830) );
  AND2_X1 U12519 ( .A1(n12911), .A2(n11057), .ZN(n11080) );
  AND2_X1 U12520 ( .A1(n14924), .A2(n13080), .ZN(n15081) );
  AND2_X1 U12521 ( .A1(n11311), .A2(n11310), .ZN(n11081) );
  OR2_X1 U12522 ( .A1(n21720), .A2(n13763), .ZN(n21813) );
  INV_X1 U12523 ( .A(n11011), .ZN(n14916) );
  NOR2_X1 U12524 ( .A1(n16998), .A2(n16999), .ZN(n16981) );
  NAND2_X1 U12525 ( .A1(n15329), .A2(n15328), .ZN(n15327) );
  XNOR2_X1 U12526 ( .A(n12888), .B(n15215), .ZN(n15213) );
  AND2_X1 U12527 ( .A1(n11264), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11082) );
  OR3_X1 U12528 ( .A1(n20779), .A2(n11607), .A3(n17575), .ZN(n11083) );
  AND2_X1 U12529 ( .A1(n15122), .A2(n15131), .ZN(n11084) );
  AND3_X1 U12530 ( .A1(n13297), .A2(n11011), .A3(n15122), .ZN(n11085) );
  XNOR2_X1 U12531 ( .A(n16426), .B(n15585), .ZN(n16418) );
  OR2_X1 U12532 ( .A1(n12179), .A2(n16183), .ZN(n11086) );
  INV_X1 U12533 ( .A(n20177), .ZN(n11206) );
  NAND2_X1 U12534 ( .A1(n15329), .A2(n11126), .ZN(n11125) );
  AND2_X1 U12535 ( .A1(n14899), .A2(n14898), .ZN(n11087) );
  AND2_X1 U12536 ( .A1(n12146), .A2(n12099), .ZN(n11088) );
  NOR2_X1 U12537 ( .A1(n17426), .A2(n17423), .ZN(n11089) );
  NOR2_X1 U12538 ( .A1(n15283), .A2(n15285), .ZN(n11448) );
  INV_X1 U12539 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21832) );
  NAND2_X1 U12540 ( .A1(n11347), .A2(n17445), .ZN(n11090) );
  OR2_X1 U12541 ( .A1(n11039), .A2(n11376), .ZN(n11091) );
  AND2_X1 U12542 ( .A1(n11298), .A2(n11297), .ZN(n11092) );
  AND2_X1 U12543 ( .A1(n11454), .A2(n15832), .ZN(n11093) );
  AND2_X1 U12544 ( .A1(n11084), .A2(n15148), .ZN(n11094) );
  AND2_X1 U12545 ( .A1(n12813), .A2(n11163), .ZN(n11095) );
  AND2_X1 U12546 ( .A1(n11081), .A2(n11309), .ZN(n11096) );
  AND2_X1 U12547 ( .A1(n13523), .A2(n11462), .ZN(n11097) );
  AND2_X1 U12548 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11098) );
  OR2_X1 U12549 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n11099) );
  INV_X1 U12550 ( .A(n14150), .ZN(n14170) );
  INV_X1 U12551 ( .A(n17463), .ZN(n17473) );
  INV_X1 U12552 ( .A(n18881), .ZN(n18825) );
  NAND2_X1 U12553 ( .A1(n15428), .A2(n15427), .ZN(n14473) );
  AND2_X1 U12554 ( .A1(n17976), .A2(n11049), .ZN(n11100) );
  AND2_X1 U12555 ( .A1(n18103), .A2(n11048), .ZN(n11101) );
  NOR2_X2 U12556 ( .A1(n11524), .A2(n11523), .ZN(n19220) );
  NOR2_X1 U12557 ( .A1(n14506), .A2(n14507), .ZN(n14505) );
  NOR2_X1 U12558 ( .A1(n14861), .A2(n11437), .ZN(n14928) );
  NOR2_X1 U12559 ( .A1(n14506), .A2(n11054), .ZN(n14866) );
  AND2_X1 U12560 ( .A1(n16876), .A2(n11390), .ZN(n11102) );
  AND2_X1 U12561 ( .A1(n12215), .A2(n11027), .ZN(n11103) );
  AND2_X1 U12562 ( .A1(n11307), .A2(n11306), .ZN(n11104) );
  AND2_X1 U12563 ( .A1(n11361), .A2(n11360), .ZN(n11105) );
  NOR2_X1 U12564 ( .A1(n18555), .A2(n18556), .ZN(n17017) );
  INV_X1 U12565 ( .A(n14930), .ZN(n11435) );
  AND2_X1 U12566 ( .A1(n11102), .A2(n11389), .ZN(n11106) );
  NOR2_X1 U12567 ( .A1(n13968), .A2(n13967), .ZN(n16362) );
  AND2_X1 U12568 ( .A1(n11028), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11107) );
  AND2_X1 U12569 ( .A1(n11028), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11108) );
  AND2_X1 U12570 ( .A1(n13134), .A2(n13138), .ZN(n11109) );
  AND2_X1 U12571 ( .A1(n11386), .A2(n11385), .ZN(n11110) );
  NAND2_X1 U12572 ( .A1(n11213), .A2(n11212), .ZN(n14174) );
  NOR2_X1 U12573 ( .A1(n18296), .A2(n11714), .ZN(n11111) );
  AND2_X1 U12574 ( .A1(n11110), .A2(n11384), .ZN(n11112) );
  AND2_X1 U12575 ( .A1(n13501), .A2(n13500), .ZN(n11113) );
  INV_X1 U12576 ( .A(n14861), .ZN(n11436) );
  INV_X1 U12577 ( .A(n11138), .ZN(n21403) );
  OR2_X1 U12578 ( .A1(n11612), .A2(n13204), .ZN(n11138) );
  AND2_X1 U12579 ( .A1(n11104), .A2(n11305), .ZN(n11114) );
  AND2_X1 U12580 ( .A1(n11038), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11115) );
  AND2_X1 U12581 ( .A1(n11105), .A2(n11359), .ZN(n11116) );
  AND2_X1 U12582 ( .A1(n11109), .A2(n15706), .ZN(n11117) );
  AND2_X2 U12583 ( .A1(n13789), .A2(n22077), .ZN(n20236) );
  CLKBUF_X3 U12584 ( .A(n17588), .Z(n21008) );
  INV_X1 U12585 ( .A(n13583), .ZN(n13725) );
  AND3_X1 U12586 ( .A1(n13973), .A2(n13972), .A3(n13971), .ZN(n11118) );
  INV_X1 U12587 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11268) );
  AND2_X1 U12588 ( .A1(n11292), .A2(n11291), .ZN(n11119) );
  INV_X1 U12589 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11261) );
  AND2_X1 U12590 ( .A1(n11277), .A2(n14223), .ZN(n11120) );
  OR2_X1 U12591 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11121) );
  AND2_X1 U12592 ( .A1(n11120), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11122) );
  INV_X1 U12593 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11259) );
  INV_X1 U12594 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11283) );
  INV_X1 U12595 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11265) );
  INV_X1 U12596 ( .A(n18869), .ZN(n18856) );
  NOR2_X4 U12597 ( .A1(n21873), .A2(n22395), .ZN(n20104) );
  AOI221_X2 U12598 ( .B1(n21424), .B2(n15368), .C1(n21424), .C2(
        P3_FLUSH_REG_SCAN_IN), .A(n19265), .ZN(n18356) );
  NOR2_X1 U12599 ( .A1(n19671), .A2(n19871), .ZN(n11123) );
  NOR2_X1 U12600 ( .A1(n19671), .A2(n19871), .ZN(n11124) );
  NAND2_X1 U12601 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19475), .ZN(n19871) );
  NAND2_X1 U12602 ( .A1(n11930), .A2(n11947), .ZN(n14532) );
  NAND2_X1 U12603 ( .A1(n14537), .A2(n13752), .ZN(n12391) );
  NOR2_X2 U12604 ( .A1(n15750), .A2(n11457), .ZN(n15725) );
  NAND2_X2 U12605 ( .A1(n15761), .A2(n15762), .ZN(n15750) );
  AND2_X2 U12606 ( .A1(n14908), .A2(n14917), .ZN(n13298) );
  OR2_X2 U12607 ( .A1(n12138), .A2(n11210), .ZN(n12147) );
  NAND2_X2 U12608 ( .A1(n11130), .A2(n11129), .ZN(n12138) );
  OAI211_X2 U12609 ( .C1(n11351), .C2(n13892), .A(n12723), .B(n12714), .ZN(
        n12753) );
  NAND2_X2 U12610 ( .A1(n11133), .A2(n14199), .ZN(n14292) );
  NAND3_X1 U12611 ( .A1(n14565), .A2(n13914), .A3(n11135), .ZN(n11134) );
  NAND3_X1 U12612 ( .A1(n21401), .A2(n11148), .A3(n11147), .ZN(n11146) );
  NAND2_X1 U12613 ( .A1(n15315), .A2(n11184), .ZN(n11149) );
  NAND3_X1 U12614 ( .A1(n11153), .A2(n11556), .A3(n11151), .ZN(n11150) );
  NAND4_X1 U12615 ( .A1(n12653), .A2(n12654), .A3(n12655), .A4(n12656), .ZN(
        n11155) );
  NAND4_X1 U12616 ( .A1(n12658), .A2(n12659), .A3(n12660), .A4(n12661), .ZN(
        n11157) );
  NAND3_X1 U12617 ( .A1(n13174), .A2(n12862), .A3(n16730), .ZN(n11160) );
  NAND2_X1 U12618 ( .A1(n11160), .A2(n18497), .ZN(n12888) );
  INV_X2 U12619 ( .A(n12699), .ZN(n19671) );
  INV_X1 U12620 ( .A(n12706), .ZN(n12705) );
  NAND2_X1 U12621 ( .A1(n11165), .A2(n12825), .ZN(n12865) );
  NAND3_X1 U12622 ( .A1(n11164), .A2(n11165), .A3(n11095), .ZN(n13161) );
  INV_X1 U12623 ( .A(n15235), .ZN(n11167) );
  NAND2_X1 U12624 ( .A1(n11170), .A2(n11169), .ZN(n11349) );
  NAND2_X1 U12625 ( .A1(n15234), .A2(n15235), .ZN(n11170) );
  XNOR2_X1 U12626 ( .A(n13851), .B(n11067), .ZN(n16771) );
  AND2_X4 U12627 ( .A1(n11182), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15683) );
  NOR2_X2 U12628 ( .A1(n12428), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11182) );
  NAND2_X2 U12629 ( .A1(n12710), .A2(n12676), .ZN(n13892) );
  AND2_X2 U12630 ( .A1(n13893), .A2(n12687), .ZN(n12652) );
  NAND2_X1 U12631 ( .A1(n12690), .A2(n12688), .ZN(n13895) );
  OAI21_X1 U12632 ( .B1(n15315), .B2(n11186), .A(n11184), .ZN(n17430) );
  NAND2_X1 U12633 ( .A1(n11188), .A2(n13164), .ZN(n15212) );
  OR2_X2 U12634 ( .A1(n17405), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11188) );
  NAND3_X1 U12635 ( .A1(n13830), .A2(n11192), .A3(n11077), .ZN(P3_U2799) );
  NOR2_X2 U12636 ( .A1(n18197), .A2(n18205), .ZN(n18196) );
  INV_X2 U12637 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21003) );
  AND2_X2 U12638 ( .A1(n11005), .A2(n14584), .ZN(n11972) );
  AND2_X4 U12639 ( .A1(n11817), .A2(n11004), .ZN(n11964) );
  AND2_X1 U12640 ( .A1(n11199), .A2(n16147), .ZN(n20199) );
  NAND2_X1 U12641 ( .A1(n16146), .A2(n11199), .ZN(n12187) );
  NAND2_X1 U12642 ( .A1(n20198), .A2(n11199), .ZN(n16149) );
  NAND3_X1 U12643 ( .A1(n12021), .A2(n21832), .A3(n21933), .ZN(n11200) );
  NAND2_X1 U12644 ( .A1(n11957), .A2(n11956), .ZN(n21933) );
  INV_X1 U12645 ( .A(n11957), .ZN(n14668) );
  NAND3_X1 U12646 ( .A1(n11207), .A2(n11202), .A3(n20231), .ZN(n16096) );
  NAND3_X1 U12647 ( .A1(n11204), .A2(n11404), .A3(n11203), .ZN(n11202) );
  NAND2_X2 U12648 ( .A1(n11453), .A2(n11088), .ZN(n12170) );
  NAND3_X1 U12649 ( .A1(n11213), .A2(n11212), .A3(n11211), .ZN(n12723) );
  NOR2_X1 U12650 ( .A1(n14174), .A2(n13897), .ZN(n14187) );
  NAND2_X1 U12651 ( .A1(n11216), .A2(n12648), .ZN(n11219) );
  NAND4_X1 U12652 ( .A1(n12458), .A2(n12459), .A3(n12457), .A4(n12456), .ZN(
        n11216) );
  NAND2_X1 U12653 ( .A1(n11217), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11218) );
  NAND4_X1 U12654 ( .A1(n12462), .A2(n12460), .A3(n12461), .A4(n12463), .ZN(
        n11217) );
  NAND2_X2 U12655 ( .A1(n11219), .A2(n11218), .ZN(n13931) );
  INV_X1 U12656 ( .A(n21321), .ZN(n21362) );
  INV_X1 U12657 ( .A(n21285), .ZN(n21336) );
  NAND2_X2 U12658 ( .A1(n21285), .A2(n19220), .ZN(n21268) );
  NOR2_X2 U12659 ( .A1(n21012), .A2(n21003), .ZN(n11661) );
  NAND4_X1 U12660 ( .A1(n11574), .A2(n11225), .A3(n11569), .A4(n11572), .ZN(
        n11224) );
  NOR3_X2 U12661 ( .A1(n21407), .A2(n19220), .A3(n21414), .ZN(n18339) );
  NOR2_X2 U12662 ( .A1(n21407), .A2(n21414), .ZN(n21443) );
  INV_X1 U12663 ( .A(n18339), .ZN(n18350) );
  AOI21_X1 U12664 ( .B1(n11320), .B2(n11230), .A(n13041), .ZN(n15431) );
  XNOR2_X2 U12665 ( .A(n11320), .B(n11230), .ZN(n14450) );
  NAND3_X1 U12666 ( .A1(n11238), .A2(n11232), .A3(n11237), .ZN(n13166) );
  NAND3_X1 U12667 ( .A1(n12861), .A2(n12860), .A3(n13173), .ZN(n11238) );
  NAND2_X1 U12668 ( .A1(n11239), .A2(n11269), .ZN(n13159) );
  OAI21_X2 U12669 ( .B1(n17008), .B2(n17009), .A(n12932), .ZN(n16659) );
  NAND2_X1 U12670 ( .A1(n16659), .A2(n11243), .ZN(n11242) );
  NAND2_X1 U12671 ( .A1(n11350), .A2(n16277), .ZN(n12715) );
  INV_X1 U12672 ( .A(n12743), .ZN(n12752) );
  AOI21_X1 U12673 ( .B1(n11778), .B2(n11258), .A(n11257), .ZN(n11256) );
  OR2_X1 U12674 ( .A1(n11778), .A2(n20763), .ZN(n11260) );
  OAI21_X1 U12675 ( .B1(n16584), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16583), .ZN(n16756) );
  INV_X1 U12676 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11275) );
  NAND2_X1 U12677 ( .A1(n11279), .A2(n11759), .ZN(n11280) );
  INV_X1 U12678 ( .A(n11281), .ZN(n18281) );
  OAI211_X1 U12679 ( .C1(n11714), .C2(n18290), .A(n11282), .B(n11285), .ZN(
        n11281) );
  NAND2_X1 U12680 ( .A1(n11284), .A2(n11283), .ZN(n11282) );
  XNOR2_X1 U12681 ( .A(n11713), .B(n11711), .ZN(n18290) );
  INV_X1 U12682 ( .A(n11714), .ZN(n11284) );
  INV_X1 U12683 ( .A(n18282), .ZN(n11285) );
  NAND2_X1 U12684 ( .A1(n11293), .A2(n11706), .ZN(n11288) );
  OAI21_X2 U12685 ( .B1(n18316), .B2(n11289), .A(n11288), .ZN(n18303) );
  XNOR2_X1 U12686 ( .A(n11705), .B(n11704), .ZN(n18316) );
  INV_X1 U12687 ( .A(n13190), .ZN(n13227) );
  INV_X2 U12688 ( .A(n12388), .ZN(n13764) );
  NAND2_X1 U12689 ( .A1(n11026), .A2(n14749), .ZN(n21448) );
  NAND3_X1 U12690 ( .A1(n11315), .A2(n11317), .A3(n11314), .ZN(n14920) );
  NAND2_X1 U12691 ( .A1(n11321), .A2(n12889), .ZN(n15234) );
  NAND2_X1 U12692 ( .A1(n11329), .A2(n11322), .ZN(n16574) );
  AOI21_X1 U12693 ( .B1(n13851), .B2(n11326), .A(n11324), .ZN(n11323) );
  INV_X1 U12694 ( .A(n13850), .ZN(n11325) );
  NOR2_X2 U12695 ( .A1(n13851), .A2(n13850), .ZN(n16576) );
  OAI21_X1 U12696 ( .B1(n11328), .B2(n11327), .A(n11337), .ZN(P2_U3015) );
  NOR2_X1 U12697 ( .A1(n16575), .A2(n16577), .ZN(n11339) );
  NAND4_X1 U12698 ( .A1(n11428), .A2(n11429), .A3(n12717), .A4(n11430), .ZN(
        n12738) );
  NAND2_X1 U12699 ( .A1(n16659), .A2(n12967), .ZN(n11341) );
  NAND2_X1 U12700 ( .A1(n12992), .A2(n11345), .ZN(n16586) );
  INV_X1 U12701 ( .A(n16586), .ZN(n13005) );
  INV_X1 U12702 ( .A(n14506), .ZN(n11352) );
  NAND2_X1 U12703 ( .A1(n11352), .A2(n11353), .ZN(n14872) );
  AND2_X1 U12704 ( .A1(n16397), .A2(n13134), .ZN(n13137) );
  NAND2_X1 U12705 ( .A1(n16397), .A2(n11109), .ZN(n15707) );
  NAND2_X1 U12706 ( .A1(n16397), .A2(n11117), .ZN(n14184) );
  AND3_X1 U12707 ( .A1(n12873), .A2(n15667), .A3(n12687), .ZN(n13914) );
  INV_X1 U12708 ( .A(n11374), .ZN(n16901) );
  INV_X1 U12709 ( .A(n16348), .ZN(n11378) );
  INV_X1 U12710 ( .A(n13968), .ZN(n11379) );
  NAND2_X1 U12711 ( .A1(n11379), .A2(n11046), .ZN(n13979) );
  NAND2_X1 U12712 ( .A1(n16512), .A2(n11110), .ZN(n16498) );
  NAND2_X1 U12713 ( .A1(n11208), .A2(n11393), .ZN(n16154) );
  NAND2_X1 U12714 ( .A1(n11014), .A2(n11400), .ZN(n11399) );
  NAND2_X1 U12715 ( .A1(n11399), .A2(n11943), .ZN(n11990) );
  NAND2_X1 U12716 ( .A1(n11936), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12022) );
  NAND2_X1 U12717 ( .A1(n13265), .A2(n21832), .ZN(n12008) );
  OAI21_X2 U12718 ( .B1(n11402), .B2(n11401), .A(n13791), .ZN(n16033) );
  INV_X1 U12719 ( .A(n11410), .ZN(n18699) );
  NAND2_X1 U12720 ( .A1(n12959), .A2(n11422), .ZN(n12980) );
  NAND2_X1 U12721 ( .A1(n12959), .A2(n12936), .ZN(n12938) );
  NOR2_X1 U12722 ( .A1(n14174), .A2(n11006), .ZN(n14648) );
  NAND2_X1 U12723 ( .A1(n11426), .A2(n16334), .ZN(n14614) );
  NAND2_X1 U12724 ( .A1(n12677), .A2(n11045), .ZN(n11427) );
  NAND2_X1 U12725 ( .A1(n11428), .A2(n11430), .ZN(n12718) );
  NAND2_X1 U12726 ( .A1(n12739), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11429) );
  NAND2_X1 U12727 ( .A1(n14450), .A2(n14438), .ZN(n11432) );
  NAND2_X1 U12728 ( .A1(n11432), .A2(n14441), .ZN(n14443) );
  NAND2_X1 U12729 ( .A1(n11432), .A2(n11078), .ZN(n14444) );
  INV_X1 U12730 ( .A(n14861), .ZN(n11433) );
  NAND2_X1 U12731 ( .A1(n11433), .A2(n11434), .ZN(n15084) );
  INV_X1 U12732 ( .A(n11438), .ZN(n16426) );
  AOI21_X2 U12733 ( .B1(n16454), .B2(n15542), .A(n11439), .ZN(n11438) );
  NAND2_X1 U12734 ( .A1(n11442), .A2(n15542), .ZN(n11440) );
  NAND2_X2 U12735 ( .A1(n14472), .A2(n14471), .ZN(n15428) );
  AND2_X2 U12736 ( .A1(n11015), .A2(n15009), .ZN(n11973) );
  NAND2_X1 U12737 ( .A1(n11453), .A2(n12146), .ZN(n12157) );
  NAND2_X1 U12738 ( .A1(n13297), .A2(n11011), .ZN(n15112) );
  NOR2_X1 U12739 ( .A1(n15750), .A2(n15751), .ZN(n15737) );
  OR2_X2 U12740 ( .A1(n15750), .A2(n11460), .ZN(n15724) );
  AND2_X2 U12741 ( .A1(n15815), .A2(n11097), .ZN(n15906) );
  NAND2_X1 U12742 ( .A1(n20145), .A2(n20144), .ZN(n20143) );
  XNOR2_X1 U12743 ( .A(n11702), .B(n11701), .ZN(n18325) );
  NAND2_X1 U12744 ( .A1(n13054), .A2(n13053), .ZN(n14506) );
  XNOR2_X2 U12745 ( .A(n16605), .B(n16595), .ZN(n16776) );
  AND2_X1 U12746 ( .A1(n17485), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12871) );
  INV_X1 U12747 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12427) );
  CLKBUF_X1 U12748 ( .A(n16454), .Z(n16461) );
  NOR2_X1 U12749 ( .A1(n19671), .A2(n19871), .ZN(n19705) );
  INV_X1 U12750 ( .A(n14475), .ZN(n13054) );
  NAND2_X1 U12751 ( .A1(n20160), .A2(n20159), .ZN(n20158) );
  AND2_X1 U12752 ( .A1(n11926), .A2(n14735), .ZN(n12110) );
  OR2_X1 U12753 ( .A1(n14417), .A2(n14416), .ZN(n14418) );
  NAND2_X1 U12754 ( .A1(n14416), .A2(n14417), .ZN(n14432) );
  CLKBUF_X1 U12755 ( .A(n14450), .Z(n17397) );
  AND2_X1 U12756 ( .A1(n15605), .A2(n15627), .ZN(n11465) );
  INV_X1 U12757 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n14841) );
  OR2_X1 U12758 ( .A1(n14234), .A2(n14188), .ZN(n18849) );
  OR2_X1 U12759 ( .A1(n17133), .A2(n21844), .ZN(n21822) );
  INV_X1 U12760 ( .A(n21822), .ZN(n20237) );
  NOR3_X1 U12761 ( .A1(n16787), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16752), .ZN(n11466) );
  AND2_X1 U12762 ( .A1(n12886), .A2(n12885), .ZN(n11467) );
  AND2_X1 U12763 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11468) );
  NOR2_X1 U12764 ( .A1(n21980), .A2(n21998), .ZN(n11469) );
  AND2_X1 U12765 ( .A1(n13228), .A2(n11475), .ZN(n11470) );
  AND2_X1 U12766 ( .A1(n15606), .A2(n11465), .ZN(n11471) );
  NAND2_X1 U12767 ( .A1(n10993), .A2(n11932), .ZN(n11472) );
  NAND2_X1 U12768 ( .A1(n18470), .A2(n18805), .ZN(n12772) );
  OR2_X1 U12769 ( .A1(n18183), .A2(n20521), .ZN(n11473) );
  OR2_X1 U12770 ( .A1(n19176), .A2(n18976), .ZN(n18333) );
  AND2_X1 U12771 ( .A1(n14197), .A2(n12700), .ZN(n11474) );
  OR2_X1 U12772 ( .A1(n21329), .A2(n20720), .ZN(n11475) );
  AND2_X1 U12773 ( .A1(n16923), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11476) );
  AND4_X1 U12774 ( .A1(n11658), .A2(n11657), .A3(n11656), .A4(n11655), .ZN(
        n11477) );
  INV_X1 U12775 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17084) );
  INV_X1 U12776 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11751) );
  INV_X1 U12777 ( .A(n12784), .ZN(n12775) );
  NAND2_X2 U12778 ( .A1(n13226), .A2(n11688), .ZN(n18258) );
  OR2_X1 U12779 ( .A1(n14749), .A2(n12217), .ZN(n11478) );
  INV_X1 U12780 ( .A(n11920), .ZN(n11922) );
  INV_X2 U12781 ( .A(n17965), .ZN(n17935) );
  INV_X1 U12782 ( .A(n15143), .ZN(n15140) );
  AND2_X1 U12783 ( .A1(n12405), .A2(n11950), .ZN(n11479) );
  NOR2_X1 U12784 ( .A1(n14278), .A2(n16334), .ZN(n14369) );
  OR2_X1 U12785 ( .A1(n13766), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11480) );
  OR2_X1 U12786 ( .A1(n13766), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11481) );
  OR2_X1 U12787 ( .A1(n13766), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11482) );
  AND2_X1 U12788 ( .A1(n18520), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17423) );
  INV_X1 U12789 ( .A(n16328), .ZN(n18848) );
  AND2_X1 U12790 ( .A1(n14025), .A2(n14024), .ZN(n14862) );
  AND2_X1 U12791 ( .A1(n14122), .A2(n14121), .ZN(n15141) );
  INV_X1 U12792 ( .A(n18152), .ZN(n18181) );
  INV_X1 U12793 ( .A(n15562), .ZN(n15541) );
  INV_X1 U12794 ( .A(n16730), .ZN(n13859) );
  INV_X1 U12795 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n18890) );
  AND2_X2 U12796 ( .A1(n15009), .A2(n14584), .ZN(n11998) );
  AND2_X1 U12797 ( .A1(n11852), .A2(n11851), .ZN(n11485) );
  AND4_X1 U12798 ( .A1(n11908), .A2(n11907), .A3(n11906), .A4(n11905), .ZN(
        n11486) );
  AND3_X1 U12799 ( .A1(n11866), .A2(n11865), .A3(n11864), .ZN(n11487) );
  OAI21_X1 U12800 ( .B1(n10993), .B2(n14749), .A(n13735), .ZN(n12260) );
  OR2_X1 U12801 ( .A1(n12245), .A2(n12243), .ZN(n12222) );
  AOI22_X1 U12802 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19406), .B1(
        n19478), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12819) );
  NAND2_X1 U12803 ( .A1(n11474), .A2(n14468), .ZN(n12701) );
  AND2_X1 U12804 ( .A1(n12224), .A2(n12223), .ZN(n12237) );
  OR2_X1 U12805 ( .A1(n11970), .A2(n11969), .ZN(n12108) );
  AND4_X1 U12806 ( .A1(n12532), .A2(n12531), .A3(n12530), .A4(n12529), .ZN(
        n12539) );
  NAND2_X1 U12807 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12619) );
  OR2_X1 U12808 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12225), .ZN(
        n12229) );
  INV_X1 U12809 ( .A(n13563), .ZN(n13564) );
  OR2_X1 U12810 ( .A1(n12086), .A2(n12085), .ZN(n12159) );
  AND3_X1 U12811 ( .A1(n11821), .A2(n11820), .A3(n11819), .ZN(n11825) );
  INV_X1 U12812 ( .A(n12744), .ZN(n12745) );
  OR2_X1 U12813 ( .A1(n11512), .A2(n11513), .ZN(n11504) );
  INV_X1 U12814 ( .A(n13606), .ZN(n13607) );
  AND2_X1 U12815 ( .A1(n13564), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13565) );
  INV_X1 U12816 ( .A(n15855), .ZN(n13389) );
  INV_X1 U12817 ( .A(n12156), .ZN(n12099) );
  INV_X1 U12818 ( .A(n14712), .ZN(n12009) );
  INV_X1 U12819 ( .A(n15676), .ZN(n15649) );
  AND2_X1 U12820 ( .A1(n16334), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14415) );
  AOI22_X1 U12821 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12665) );
  OAI21_X1 U12822 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21394), .A(
        n11504), .ZN(n11505) );
  AOI21_X1 U12823 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21832), .A(
        n12267), .ZN(n12268) );
  AND2_X1 U12824 ( .A1(n16025), .A2(n13757), .ZN(n13721) );
  NAND2_X1 U12825 ( .A1(n13607), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13609) );
  INV_X1 U12826 ( .A(n13276), .ZN(n13583) );
  NAND2_X1 U12827 ( .A1(n13374), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13390) );
  NOR2_X1 U12828 ( .A1(n12101), .A2(n12134), .ZN(n12102) );
  OR2_X1 U12829 ( .A1(n12004), .A2(n12003), .ZN(n12109) );
  OR2_X1 U12830 ( .A1(n16316), .A2(n16625), .ZN(n16317) );
  OR2_X1 U12831 ( .A1(n13022), .A2(n13021), .ZN(n13024) );
  INV_X1 U12832 ( .A(n15141), .ZN(n15142) );
  AND2_X1 U12833 ( .A1(n14415), .A2(n19562), .ZN(n15627) );
  OR2_X1 U12834 ( .A1(n16589), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13004) );
  OR2_X1 U12835 ( .A1(n18564), .A2(n16730), .ZN(n12928) );
  NOR2_X1 U12836 ( .A1(n12785), .A2(n12772), .ZN(n12849) );
  NOR2_X1 U12837 ( .A1(n12779), .A2(n12772), .ZN(n12830) );
  OAI21_X1 U12838 ( .B1(n11577), .B2(n13203), .A(n11576), .ZN(n11604) );
  NOR2_X1 U12839 ( .A1(n11609), .A2(n20841), .ZN(n13203) );
  NOR2_X1 U12840 ( .A1(n20820), .A2(n11710), .ZN(n11715) );
  AND2_X1 U12841 ( .A1(n12227), .A2(n12233), .ZN(n12279) );
  AND2_X1 U12842 ( .A1(n21805), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15778) );
  NAND2_X1 U12843 ( .A1(n13769), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15878) );
  INV_X1 U12844 ( .A(n11988), .ZN(n11989) );
  AOI22_X1 U12845 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11998), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11874) );
  NAND2_X1 U12846 ( .A1(n13422), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13694) );
  OR2_X1 U12847 ( .A1(n13634), .A2(n13633), .ZN(n13673) );
  INV_X1 U12848 ( .A(n13694), .ZN(n13718) );
  NOR2_X1 U12849 ( .A1(n13390), .A2(n15863), .ZN(n13405) );
  NAND2_X1 U12850 ( .A1(n13343), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13369) );
  OAI21_X1 U12851 ( .B1(n13794), .B2(n12179), .A(n13793), .ZN(n13795) );
  AND2_X1 U12852 ( .A1(n12348), .A2(n11480), .ZN(n15818) );
  NAND2_X1 U12853 ( .A1(n12049), .A2(n12048), .ZN(n15010) );
  INV_X1 U12854 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12225) );
  INV_X1 U12855 ( .A(n14172), .ZN(n14173) );
  INV_X1 U12856 ( .A(n16310), .ZN(n13142) );
  AND2_X1 U12857 ( .A1(n13121), .A2(n13120), .ZN(n16421) );
  INV_X1 U12858 ( .A(n16442), .ZN(n15495) );
  NAND2_X1 U12859 ( .A1(n16324), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16325) );
  AND2_X1 U12860 ( .A1(n13094), .A2(n13093), .ZN(n15266) );
  NAND2_X1 U12861 ( .A1(n16289), .A2(n14189), .ZN(n14230) );
  AND2_X1 U12862 ( .A1(n13074), .A2(n13073), .ZN(n14925) );
  INV_X1 U12863 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14616) );
  AND2_X1 U12864 ( .A1(n12698), .A2(n14468), .ZN(n12689) );
  INV_X1 U12865 ( .A(n12850), .ZN(n19406) );
  INV_X1 U12866 ( .A(n18258), .ZN(n13191) );
  INV_X1 U12867 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11701) );
  AOI21_X1 U12868 ( .B1(n11762), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11761), .ZN(n11763) );
  AND3_X1 U12869 ( .A1(n13191), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17989), .ZN(n18071) );
  INV_X1 U12870 ( .A(n21160), .ZN(n21163) );
  INV_X1 U12871 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11704) );
  NAND2_X1 U12872 ( .A1(n12270), .A2(n12269), .ZN(n12271) );
  AND2_X1 U12873 ( .A1(n15778), .A2(n13770), .ZN(n15752) );
  INV_X1 U12874 ( .A(n20221), .ZN(n15821) );
  AND2_X1 U12875 ( .A1(n11027), .A2(n15875), .ZN(n13775) );
  INV_X1 U12876 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15262) );
  NAND2_X1 U12877 ( .A1(n13774), .A2(n13775), .ZN(n21732) );
  OR2_X1 U12878 ( .A1(n21453), .A2(n13759), .ZN(n13769) );
  OR2_X1 U12879 ( .A1(n14511), .A2(n15389), .ZN(n14551) );
  XNOR2_X1 U12880 ( .A(n13761), .B(n13780), .ZN(n15150) );
  INV_X1 U12881 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13517) );
  AND3_X1 U12882 ( .A1(n21832), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n13789) );
  AND2_X1 U12883 ( .A1(n12285), .A2(n15390), .ZN(n12415) );
  OR2_X1 U12884 ( .A1(n21953), .A2(n21941), .ZN(n22318) );
  INV_X1 U12885 ( .A(n13264), .ZN(n14938) );
  OR2_X1 U12886 ( .A1(n14939), .A2(n22037), .ZN(n22334) );
  INV_X1 U12887 ( .A(n15105), .ZN(n15108) );
  AOI21_X1 U12888 ( .B1(n22029), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n21924), 
        .ZN(n22035) );
  AND2_X1 U12889 ( .A1(n14667), .A2(n14938), .ZN(n21919) );
  OR2_X1 U12890 ( .A1(n13892), .A2(n19872), .ZN(n14260) );
  NAND2_X1 U12891 ( .A1(n15667), .A2(n15541), .ZN(n15542) );
  NAND2_X1 U12892 ( .A1(n13983), .A2(n13982), .ZN(n15305) );
  INV_X1 U12893 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15320) );
  AND2_X1 U12894 ( .A1(n16755), .A2(n16754), .ZN(n16757) );
  OR2_X1 U12895 ( .A1(n16848), .A2(n14224), .ZN(n16809) );
  NAND2_X1 U12896 ( .A1(n18829), .A2(n14211), .ZN(n17037) );
  INV_X1 U12897 ( .A(n14924), .ZN(n15080) );
  INV_X1 U12898 ( .A(n18808), .ZN(n17047) );
  OR2_X1 U12899 ( .A1(n14234), .A2(n14191), .ZN(n16912) );
  INV_X1 U12900 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19472) );
  OR2_X1 U12901 ( .A1(n19613), .A2(n17488), .ZN(n19455) );
  NAND2_X1 U12902 ( .A1(n19420), .A2(n17481), .ZN(n19414) );
  INV_X1 U12903 ( .A(n19508), .ZN(n19532) );
  OAI211_X1 U12904 ( .C1(n11513), .C2(n11512), .A(n11511), .B(n11510), .ZN(
        n11619) );
  NOR2_X1 U12905 ( .A1(n11666), .A2(n11665), .ZN(n11667) );
  NOR3_X1 U12906 ( .A1(n20779), .A2(n20778), .A3(n20777), .ZN(n20780) );
  INV_X1 U12907 ( .A(n18211), .ZN(n18002) );
  INV_X1 U12908 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18297) );
  NAND3_X1 U12909 ( .A1(n21855), .A2(n18345), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18180) );
  INV_X1 U12910 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21388) );
  AND2_X1 U12911 ( .A1(n12272), .A2(n12271), .ZN(n15389) );
  NAND2_X1 U12912 ( .A1(n14295), .A2(n14740), .ZN(n21453) );
  AND3_X1 U12913 ( .A1(n13776), .A2(n13775), .A3(n17143), .ZN(n21801) );
  NOR2_X1 U12914 ( .A1(n15255), .A2(n21732), .ZN(n15857) );
  INV_X1 U12915 ( .A(n21813), .ZN(n21771) );
  INV_X1 U12916 ( .A(n15954), .ZN(n20132) );
  INV_X1 U12917 ( .A(n15952), .ZN(n20131) );
  INV_X1 U12918 ( .A(n14745), .ZN(n14808) );
  OR2_X1 U12919 ( .A1(n14740), .A2(n14739), .ZN(n14804) );
  NAND2_X1 U12920 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13519), .ZN(
        n13563) );
  INV_X1 U12921 ( .A(n20240), .ZN(n20222) );
  INV_X1 U12922 ( .A(n13291), .ZN(n13292) );
  OR2_X1 U12923 ( .A1(n13803), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13804) );
  INV_X1 U12924 ( .A(n21501), .ZN(n21575) );
  NAND2_X1 U12925 ( .A1(n21608), .A2(n16268), .ZN(n21551) );
  NAND2_X1 U12926 ( .A1(n15389), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21825) );
  INV_X1 U12927 ( .A(n21930), .ZN(n22312) );
  INV_X1 U12928 ( .A(n22316), .ZN(n22320) );
  INV_X1 U12929 ( .A(n22318), .ZN(n22328) );
  INV_X1 U12930 ( .A(n22326), .ZN(n22201) );
  INV_X1 U12931 ( .A(n15078), .ZN(n14974) );
  INV_X1 U12932 ( .A(n14757), .ZN(n22336) );
  INV_X1 U12933 ( .A(n14725), .ZN(n22343) );
  INV_X1 U12934 ( .A(n21993), .ZN(n21978) );
  INV_X1 U12935 ( .A(n21919), .ZN(n15043) );
  AND2_X1 U12936 ( .A1(n21978), .A2(n22041), .ZN(n22354) );
  INV_X1 U12937 ( .A(n14812), .ZN(n22362) );
  INV_X1 U12938 ( .A(n21977), .ZN(n22012) );
  INV_X1 U12939 ( .A(n22070), .ZN(n22049) );
  INV_X1 U12940 ( .A(n22262), .ZN(n22256) );
  AND2_X1 U12941 ( .A1(n22042), .A2(n21919), .ZN(n22389) );
  AND2_X1 U12942 ( .A1(n15105), .A2(n11129), .ZN(n22042) );
  INV_X1 U12943 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21872) );
  NOR2_X1 U12944 ( .A1(n14638), .A2(n18904), .ZN(n14264) );
  AND2_X1 U12945 ( .A1(n16290), .A2(n16288), .ZN(n18776) );
  NOR2_X2 U12946 ( .A1(n17388), .A2(n16330), .ZN(n18755) );
  AND2_X1 U12947 ( .A1(n17388), .A2(n16327), .ZN(n18795) );
  AND2_X1 U12948 ( .A1(n15698), .A2(n15695), .ZN(n19765) );
  INV_X1 U12949 ( .A(n19812), .ZN(n19862) );
  INV_X1 U12950 ( .A(n14319), .ZN(n14382) );
  INV_X1 U12951 ( .A(n16623), .ZN(n18720) );
  NAND2_X1 U12952 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16305), .ZN(
        n16304) );
  NAND2_X1 U12953 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16303), .ZN(
        n16302) );
  NAND2_X1 U12954 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16299), .ZN(
        n16298) );
  INV_X1 U12955 ( .A(n17459), .ZN(n17470) );
  NOR2_X1 U12956 ( .A1(n17037), .A2(n14217), .ZN(n16908) );
  NOR2_X1 U12957 ( .A1(n15249), .A2(n15237), .ZN(n18829) );
  AOI21_X1 U12958 ( .B1(n16912), .B2(n14213), .A(n17047), .ZN(n18847) );
  INV_X1 U12959 ( .A(n18870), .ZN(n18852) );
  INV_X1 U12960 ( .A(n13148), .ZN(n14307) );
  INV_X1 U12961 ( .A(n19475), .ZN(n19869) );
  NOR2_X1 U12962 ( .A1(n19440), .A2(n19539), .ZN(n19961) );
  NAND2_X1 U12963 ( .A1(n19613), .A2(n19611), .ZN(n19539) );
  INV_X1 U12964 ( .A(n19849), .ZN(n19953) );
  INV_X1 U12965 ( .A(n19944), .ZN(n19946) );
  AND2_X1 U12966 ( .A1(n19499), .A2(n19498), .ZN(n19939) );
  AND2_X1 U12967 ( .A1(n19613), .A2(n17488), .ZN(n19499) );
  INV_X1 U12968 ( .A(n19837), .ZN(n19928) );
  INV_X1 U12969 ( .A(n19906), .ZN(n19908) );
  INV_X1 U12970 ( .A(n19455), .ZN(n19453) );
  NOR2_X1 U12971 ( .A1(n19414), .A2(n19421), .ZN(n19889) );
  INV_X1 U12972 ( .A(n19699), .ZN(n19706) );
  INV_X1 U12973 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n13888) );
  OAI211_X1 U12974 ( .C1(n11618), .C2(n11514), .A(n11616), .B(n11619), .ZN(
        n21385) );
  INV_X1 U12975 ( .A(n20754), .ZN(n11810) );
  NAND4_X1 U12976 ( .A1(n11804), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n20779), 
        .A4(n11803), .ZN(n20764) );
  NOR2_X1 U12977 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n20571), .ZN(n20593) );
  NOR2_X1 U12978 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n20509), .ZN(n20531) );
  INV_X1 U12979 ( .A(n20762), .ZN(n20718) );
  NOR2_X1 U12980 ( .A1(n20652), .A2(n17889), .ZN(n17871) );
  NOR2_X1 U12981 ( .A1(n20530), .A2(n17687), .ZN(n17637) );
  INV_X1 U12982 ( .A(n17968), .ZN(n17962) );
  INV_X1 U12983 ( .A(n20910), .ZN(n20905) );
  NOR2_X1 U12984 ( .A1(n20859), .A2(n20879), .ZN(n20867) );
  INV_X1 U12985 ( .A(n20966), .ZN(n20843) );
  INV_X1 U12986 ( .A(n20370), .ZN(n20778) );
  NAND2_X1 U12987 ( .A1(n13226), .A2(n18339), .ZN(n18187) );
  INV_X2 U12988 ( .A(n18351), .ZN(n18275) );
  INV_X1 U12989 ( .A(n20812), .ZN(n13226) );
  INV_X1 U12990 ( .A(n21333), .ZN(n21373) );
  INV_X1 U12991 ( .A(n21263), .ZN(n21369) );
  NOR2_X1 U12992 ( .A1(n10995), .A2(n21369), .ZN(n21238) );
  NAND2_X1 U12993 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21419), .ZN(n21414) );
  INV_X1 U12994 ( .A(n21429), .ZN(n21026) );
  INV_X1 U12995 ( .A(n19244), .ZN(n19341) );
  INV_X1 U12996 ( .A(n21414), .ZN(n21440) );
  INV_X1 U12997 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21862) );
  INV_X1 U12998 ( .A(n18444), .ZN(n18438) );
  OAI21_X1 U12999 ( .B1(n14246), .B2(n14245), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14361) );
  NOR2_X1 U13000 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14249), .ZN(n18937)
         );
  NAND3_X1 U13001 ( .A1(n11103), .A2(n15390), .A3(n15389), .ZN(n14740) );
  OR2_X1 U13002 ( .A1(n21720), .A2(n22021), .ZN(n21820) );
  INV_X1 U13003 ( .A(n21801), .ZN(n21812) );
  INV_X1 U13004 ( .A(n21810), .ZN(n21765) );
  AND2_X1 U13005 ( .A1(n21813), .A2(n15877), .ZN(n21690) );
  NAND2_X1 U13006 ( .A1(n20136), .A2(n15956), .ZN(n15952) );
  INV_X1 U13007 ( .A(n20195), .ZN(n15297) );
  INV_X1 U13008 ( .A(n20035), .ZN(n20066) );
  INV_X1 U13009 ( .A(n14804), .ZN(n14745) );
  INV_X1 U13010 ( .A(n20236), .ZN(n16118) );
  NAND2_X2 U13011 ( .A1(n16114), .A2(n14528), .ZN(n20240) );
  OR2_X1 U13012 ( .A1(n13810), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21596) );
  INV_X1 U13013 ( .A(n21625), .ZN(n21642) );
  INV_X1 U13014 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22029) );
  INV_X2 U13015 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14594) );
  AOI22_X1 U13016 ( .A1(n21928), .A2(n21925), .B1(n11469), .B2(n21999), .ZN(
        n22309) );
  OR2_X1 U13017 ( .A1(n21953), .A2(n22037), .ZN(n22316) );
  AOI22_X1 U13018 ( .A1(n21943), .A2(n21947), .B1(n21999), .B2(n21967), .ZN(
        n22324) );
  INV_X1 U13019 ( .A(n21956), .ZN(n22332) );
  OR2_X1 U13020 ( .A1(n14939), .A2(n21977), .ZN(n15078) );
  AOI22_X1 U13021 ( .A1(n21968), .A2(n21973), .B1(n22044), .B2(n21967), .ZN(
        n22340) );
  OR2_X1 U13022 ( .A1(n14939), .A2(n21941), .ZN(n14757) );
  NAND2_X1 U13023 ( .A1(n21978), .A2(n22012), .ZN(n22352) );
  AOI22_X1 U13024 ( .A1(n22000), .A2(n22008), .B1(n21999), .B2(n22045), .ZN(
        n22359) );
  INV_X1 U13025 ( .A(n22354), .ZN(n14837) );
  INV_X1 U13026 ( .A(n22180), .ZN(n22186) );
  AOI22_X1 U13027 ( .A1(n22017), .A2(n22025), .B1(n22044), .B2(n22016), .ZN(
        n22366) );
  NAND2_X1 U13028 ( .A1(n22042), .A2(n22012), .ZN(n22372) );
  NAND2_X1 U13029 ( .A1(n22042), .A2(n22041), .ZN(n22393) );
  NOR2_X1 U13030 ( .A1(n17154), .A2(n13234), .ZN(n21834) );
  CLKBUF_X1 U13031 ( .A(n17117), .Z(n21848) );
  OR2_X1 U13032 ( .A1(n22395), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20092) );
  NAND2_X1 U13033 ( .A1(n14261), .A2(n14264), .ZN(n14278) );
  AND2_X1 U13034 ( .A1(n14639), .A2(n14264), .ZN(n17388) );
  INV_X1 U13035 ( .A(n18776), .ZN(n18800) );
  INV_X1 U13036 ( .A(n18755), .ZN(n18791) );
  INV_X1 U13037 ( .A(n18796), .ZN(n18737) );
  XNOR2_X1 U13038 ( .A(n14467), .B(n11000), .ZN(n19613) );
  INV_X1 U13039 ( .A(n17488), .ZN(n19611) );
  AND2_X1 U13040 ( .A1(n19549), .A2(n19812), .ZN(n19620) );
  INV_X1 U13041 ( .A(n19606), .ZN(n19868) );
  INV_X1 U13042 ( .A(n17512), .ZN(n17540) );
  INV_X1 U13043 ( .A(n14369), .ZN(n14319) );
  OR2_X1 U13044 ( .A1(n18911), .A2(n16334), .ZN(n17463) );
  INV_X1 U13045 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17441) );
  INV_X1 U13046 ( .A(n17453), .ZN(n17479) );
  OR2_X1 U13047 ( .A1(n14234), .A2(n13913), .ZN(n18869) );
  OR2_X1 U13048 ( .A1(n14234), .A2(n14644), .ZN(n18881) );
  INV_X1 U13049 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17485) );
  INV_X1 U13050 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14656) );
  AOI22_X1 U13051 ( .A1(n15174), .A2(n15173), .B1(n15172), .B2(n15171), .ZN(
        n19984) );
  INV_X1 U13052 ( .A(n19961), .ZN(n19971) );
  OR2_X1 U13053 ( .A1(n19539), .A2(n19467), .ZN(n19849) );
  OR2_X1 U13054 ( .A1(n19539), .A2(n14856), .ZN(n19965) );
  AOI21_X1 U13055 ( .B1(n15093), .B2(n15098), .A(n15092), .ZN(n19951) );
  NAND2_X1 U13056 ( .A1(n19499), .A2(n19452), .ZN(n19944) );
  NAND2_X1 U13057 ( .A1(n19499), .A2(n19492), .ZN(n19937) );
  NAND2_X1 U13058 ( .A1(n19499), .A2(n19468), .ZN(n19837) );
  NAND2_X1 U13059 ( .A1(n19453), .A2(n19452), .ZN(n19925) );
  NAND2_X1 U13060 ( .A1(n19453), .A2(n19498), .ZN(n19913) );
  NAND2_X1 U13061 ( .A1(n19453), .A2(n19492), .ZN(n19906) );
  INV_X1 U13062 ( .A(n19882), .ZN(n19893) );
  AOI22_X1 U13063 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19875), .ZN(n19546) );
  INV_X1 U13064 ( .A(n19600), .ZN(n19593) );
  INV_X1 U13065 ( .A(n21853), .ZN(n17098) );
  INV_X1 U13066 ( .A(n21888), .ZN(n17567) );
  AOI211_X1 U13067 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n20751), .A(n11810), 
        .B(n11809), .ZN(n11811) );
  NAND2_X1 U13068 ( .A1(n11793), .A2(n20741), .ZN(n11812) );
  INV_X1 U13069 ( .A(n20766), .ZN(n20719) );
  NAND2_X1 U13070 ( .A1(n20768), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20762) );
  NOR2_X1 U13071 ( .A1(n20701), .A2(n17855), .ZN(n17860) );
  NOR2_X1 U13072 ( .A1(n20608), .A2(n17921), .ZN(n17937) );
  NOR2_X1 U13073 ( .A1(n20493), .A2(n17714), .ZN(n17702) );
  INV_X1 U13074 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17782) );
  NOR2_X2 U13075 ( .A1(n17962), .A2(n20959), .ZN(n17965) );
  INV_X1 U13076 ( .A(n20968), .ZN(n20946) );
  NOR3_X1 U13077 ( .A1(n20963), .A2(n20783), .A3(n20964), .ZN(n20807) );
  NOR2_X1 U13078 ( .A1(n11631), .A2(n11630), .ZN(n20820) );
  INV_X1 U13079 ( .A(n20972), .ZN(n20956) );
  NAND2_X1 U13080 ( .A1(n18399), .A2(n20778), .ZN(n18417) );
  NAND2_X1 U13081 ( .A1(n17092), .A2(n17091), .ZN(n18398) );
  INV_X1 U13082 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20374) );
  NAND2_X1 U13083 ( .A1(n13226), .A2(n21110), .ZN(n21333) );
  INV_X1 U13084 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21376) );
  INV_X1 U13085 ( .A(n21172), .ZN(n21246) );
  INV_X1 U13086 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18975) );
  INV_X1 U13087 ( .A(n19359), .ZN(n19339) );
  INV_X1 U13088 ( .A(n19329), .ZN(n19321) );
  INV_X1 U13089 ( .A(n19306), .ZN(n19298) );
  INV_X1 U13090 ( .A(n19122), .ZN(n19133) );
  INV_X1 U13091 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21438) );
  INV_X1 U13092 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21426) );
  INV_X1 U13093 ( .A(n21858), .ZN(n17086) );
  INV_X1 U13094 ( .A(n18436), .ZN(n18443) );
  NAND2_X1 U13095 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21864), .ZN(n18444) );
  NAND2_X1 U13096 ( .A1(n11812), .A2(n11811), .ZN(P3_U2641) );
  OAI21_X1 U13097 ( .B1(n13230), .B2(n13229), .A(n11470), .ZN(P3_U2834) );
  NOR2_X2 U13098 ( .A1(n21005), .A2(n11494), .ZN(n11621) );
  NOR2_X2 U13099 ( .A1(n11492), .A2(n11494), .ZN(n11547) );
  AOI22_X1 U13100 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11547), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U13101 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11490) );
  CLKBUF_X3 U13102 ( .A(n11661), .Z(n17941) );
  AOI22_X1 U13103 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U13104 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17942), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11488) );
  NAND4_X1 U13105 ( .A1(n11491), .A2(n11490), .A3(n11489), .A4(n11488), .ZN(
        n11501) );
  AOI22_X1 U13106 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17927), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11499) );
  INV_X2 U13107 ( .A(n11525), .ZN(n17906) );
  BUF_X4 U13108 ( .A(n11691), .Z(n17949) );
  AOI22_X1 U13109 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U13110 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17803), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11497) );
  NOR2_X2 U13111 ( .A1(n11494), .A2(n11495), .ZN(n11537) );
  NOR2_X2 U13112 ( .A1(n20368), .A2(n11495), .ZN(n11654) );
  CLKBUF_X3 U13113 ( .A(n11654), .Z(n17938) );
  AOI22_X1 U13114 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11496) );
  NAND4_X1 U13115 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11500) );
  NAND2_X1 U13116 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18980), .ZN(
        n11615) );
  OAI21_X1 U13117 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18980), .A(
        n11615), .ZN(n11618) );
  AOI22_X1 U13118 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21388), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20991), .ZN(n11614) );
  INV_X1 U13119 ( .A(n11614), .ZN(n11502) );
  OAI22_X1 U13120 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17090), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11505), .ZN(n11507) );
  NOR2_X1 U13121 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17090), .ZN(
        n11506) );
  NAND2_X1 U13122 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11505), .ZN(
        n11508) );
  AOI22_X1 U13123 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11507), .B1(
        n11506), .B2(n11508), .ZN(n11511) );
  NAND2_X1 U13124 ( .A1(n11614), .A2(n11511), .ZN(n11514) );
  AOI21_X1 U13125 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11508), .A(
        n11507), .ZN(n11509) );
  NAND2_X1 U13126 ( .A1(n11513), .A2(n11512), .ZN(n11510) );
  INV_X1 U13127 ( .A(n21385), .ZN(n13213) );
  INV_X2 U13128 ( .A(n17649), .ZN(n17732) );
  AOI22_X1 U13129 ( .A1(n17949), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U13130 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U13131 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U13132 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11515) );
  NAND4_X1 U13133 ( .A1(n11518), .A2(n11517), .A3(n11516), .A4(n11515), .ZN(
        n11524) );
  AOI22_X1 U13134 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U13135 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17783), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U13136 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U13137 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11519) );
  NAND4_X1 U13138 ( .A1(n11522), .A2(n11521), .A3(n11520), .A4(n11519), .ZN(
        n11523) );
  AOI22_X1 U13139 ( .A1(n17949), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U13140 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U13141 ( .A1(n11661), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U13142 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11526) );
  NAND4_X1 U13143 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11535) );
  AOI22_X1 U13144 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U13145 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11654), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U13146 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U13147 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U13148 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11534) );
  INV_X2 U13149 ( .A(n17816), .ZN(n17951) );
  AOI22_X1 U13150 ( .A1(n17951), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U13151 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U13152 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11536) );
  OAI21_X1 U13153 ( .B1(n17649), .B2(n17905), .A(n11536), .ZN(n11543) );
  AOI22_X1 U13154 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U13155 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11547), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U13156 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17943), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U13157 ( .A1(n11661), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17942), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11538) );
  NAND4_X1 U13158 ( .A1(n11541), .A2(n11540), .A3(n11539), .A4(n11538), .ZN(
        n11542) );
  AOI22_X1 U13159 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U13160 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U13161 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11548) );
  OAI21_X1 U13162 ( .B1(n17649), .B2(n17891), .A(n11548), .ZN(n11555) );
  AOI22_X1 U13163 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11691), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U13164 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U13165 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U13166 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11550) );
  NAND4_X1 U13167 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11554) );
  NOR2_X1 U13168 ( .A1(n11611), .A2(n17576), .ZN(n13210) );
  INV_X1 U13169 ( .A(n13210), .ZN(n11577) );
  AOI22_X1 U13170 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17927), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U13171 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10992), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U13172 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U13173 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11558) );
  NAND4_X1 U13174 ( .A1(n11561), .A2(n11560), .A3(n11559), .A4(n11558), .ZN(
        n11567) );
  AOI22_X1 U13175 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U13176 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U13177 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U13178 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11562) );
  NAND4_X1 U13179 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11566) );
  AOI22_X1 U13180 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U13181 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17783), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U13182 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11568) );
  OAI21_X1 U13183 ( .B1(n17649), .B2(n17815), .A(n11568), .ZN(n11573) );
  AOI22_X1 U13184 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11691), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U13185 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11621), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U13186 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U13187 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11569) );
  NOR2_X1 U13188 ( .A1(n20840), .A2(n11611), .ZN(n13201) );
  INV_X1 U13189 ( .A(n13201), .ZN(n11576) );
  AOI22_X1 U13190 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U13191 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U13192 ( .A1(n11620), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11691), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11578) );
  OAI21_X1 U13193 ( .B1(n17649), .B2(n17782), .A(n11578), .ZN(n11584) );
  AOI22_X1 U13194 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U13195 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U13196 ( .A1(n11661), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U13197 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11579) );
  NAND4_X1 U13198 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11583) );
  AOI22_X1 U13199 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U13200 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11596) );
  INV_X1 U13201 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17582) );
  AOI22_X1 U13202 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11588) );
  OAI21_X1 U13203 ( .B1(n17649), .B2(n17582), .A(n11588), .ZN(n11594) );
  AOI22_X1 U13204 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U13205 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U13206 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U13207 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11589) );
  NAND4_X1 U13208 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n11593) );
  AOI211_X1 U13209 ( .C1(n17914), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n11594), .B(n11593), .ZN(n11595) );
  NAND3_X1 U13210 ( .A1(n11597), .A2(n11596), .A3(n11595), .ZN(n11606) );
  NAND2_X1 U13211 ( .A1(n11604), .A2(n13206), .ZN(n11610) );
  INV_X1 U13212 ( .A(n11610), .ZN(n11598) );
  NAND2_X1 U13213 ( .A1(n20809), .A2(n20370), .ZN(n11607) );
  OR2_X1 U13214 ( .A1(n11606), .A2(n11607), .ZN(n11599) );
  INV_X1 U13215 ( .A(n13212), .ZN(n11601) );
  INV_X1 U13216 ( .A(n11611), .ZN(n19177) );
  NAND2_X1 U13217 ( .A1(n20370), .A2(n20779), .ZN(n11613) );
  NAND2_X1 U13218 ( .A1(n19177), .A2(n11613), .ZN(n13202) );
  INV_X1 U13219 ( .A(n20787), .ZN(n20978) );
  NOR2_X1 U13220 ( .A1(n20959), .A2(n20978), .ZN(n20786) );
  NOR3_X1 U13221 ( .A1(n20370), .A2(n20786), .A3(n20779), .ZN(n13208) );
  OAI21_X1 U13222 ( .B1(n20778), .B2(n11611), .A(n20787), .ZN(n13209) );
  INV_X1 U13223 ( .A(n13209), .ZN(n11600) );
  AOI211_X1 U13224 ( .C1(n11601), .C2(n13202), .A(n13208), .B(n11608), .ZN(
        n11603) );
  NAND2_X1 U13225 ( .A1(n19135), .A2(n11607), .ZN(n11602) );
  OAI211_X1 U13226 ( .C1(n11604), .C2(n19135), .A(n11603), .B(n11602), .ZN(
        n11605) );
  AOI221_X2 U13227 ( .B1(n20959), .B2(n17576), .C1(n13212), .C2(n17576), .A(
        n11605), .ZN(n21010) );
  NOR2_X1 U13228 ( .A1(n11611), .A2(n11606), .ZN(n20989) );
  NAND2_X1 U13229 ( .A1(n13203), .A2(n20989), .ZN(n17575) );
  NAND2_X1 U13230 ( .A1(n20779), .A2(n11612), .ZN(n11795) );
  AND2_X1 U13231 ( .A1(n11611), .A2(n11794), .ZN(n13204) );
  NAND2_X1 U13232 ( .A1(n19220), .A2(n11612), .ZN(n21379) );
  NOR2_X1 U13233 ( .A1(n19220), .A2(n13206), .ZN(n20987) );
  NOR2_X1 U13234 ( .A1(n20989), .A2(n20987), .ZN(n13195) );
  XOR2_X1 U13235 ( .A(n11615), .B(n11614), .Z(n11617) );
  INV_X1 U13236 ( .A(n13200), .ZN(n21405) );
  OAI21_X1 U13237 ( .B1(n11619), .B2(n11618), .A(n21405), .ZN(n13211) );
  INV_X1 U13238 ( .A(n13211), .ZN(n21382) );
  INV_X2 U13239 ( .A(n11041), .ZN(n18262) );
  INV_X1 U13240 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21205) );
  INV_X1 U13241 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21229) );
  NOR2_X1 U13242 ( .A1(n21205), .A2(n21229), .ZN(n13194) );
  INV_X1 U13243 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21283) );
  INV_X1 U13244 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18095) );
  INV_X1 U13245 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21280) );
  NOR2_X1 U13246 ( .A1(n18095), .A2(n21280), .ZN(n18112) );
  INV_X1 U13247 ( .A(n18112), .ZN(n11749) );
  INV_X1 U13248 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21338) );
  INV_X1 U13249 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21330) );
  NOR2_X1 U13250 ( .A1(n21338), .A2(n21330), .ZN(n21314) );
  NAND2_X1 U13251 ( .A1(n21314), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17987) );
  INV_X1 U13252 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18082) );
  INV_X1 U13253 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21300) );
  NOR2_X1 U13254 ( .A1(n18082), .A2(n21300), .ZN(n21042) );
  NAND2_X1 U13255 ( .A1(n21042), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13833) );
  NOR2_X1 U13256 ( .A1(n17987), .A2(n13833), .ZN(n18048) );
  INV_X1 U13257 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18205) );
  INV_X1 U13258 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21351) );
  NOR2_X1 U13259 ( .A1(n21376), .A2(n21351), .ZN(n21130) );
  NAND3_X1 U13260 ( .A1(n21130), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18041) );
  INV_X1 U13261 ( .A(n18041), .ZN(n21152) );
  NAND2_X1 U13262 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21152), .ZN(
        n21160) );
  AOI22_X1 U13263 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U13264 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11547), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U13265 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17943), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U13266 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17942), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11622) );
  NAND4_X1 U13267 ( .A1(n11625), .A2(n11624), .A3(n11623), .A4(n11622), .ZN(
        n11631) );
  AOI22_X1 U13268 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U13269 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17927), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U13270 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U13271 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11626) );
  NAND4_X1 U13272 ( .A1(n11629), .A2(n11628), .A3(n11627), .A4(n11626), .ZN(
        n11630) );
  AOI22_X1 U13273 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U13274 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17803), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U13275 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17942), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U13276 ( .A1(n11661), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17943), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11633) );
  NAND4_X1 U13277 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n11642) );
  AOI22_X1 U13278 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17927), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U13279 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U13280 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U13281 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11547), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11637) );
  NAND4_X1 U13282 ( .A1(n11640), .A2(n11639), .A3(n11638), .A4(n11637), .ZN(
        n11641) );
  AOI22_X1 U13283 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U13284 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17927), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U13285 ( .A1(n17588), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11549), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11643) );
  OAI21_X1 U13286 ( .B1(n20409), .B2(n17905), .A(n11643), .ZN(n11650) );
  AOI22_X1 U13287 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11621), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U13288 ( .A1(n11620), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11644), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U13289 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11547), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U13290 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11654), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11645) );
  NAND4_X1 U13291 ( .A1(n11648), .A2(n11647), .A3(n11646), .A4(n11645), .ZN(
        n11649) );
  AOI211_X1 U13292 ( .C1(n11661), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n11650), .B(n11649), .ZN(n11651) );
  NAND3_X1 U13293 ( .A1(n11653), .A2(n11652), .A3(n11651), .ZN(n20835) );
  AOI22_X1 U13294 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11654), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11658) );
  INV_X1 U13295 ( .A(n17906), .ZN(n17771) );
  AOI22_X1 U13296 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17771), .B1(
        n11547), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U13297 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17927), .ZN(n11656) );
  AOI22_X1 U13298 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n11621), .ZN(n11655) );
  INV_X1 U13299 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U13300 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17943), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17942), .ZN(n11659) );
  OAI21_X1 U13301 ( .B1(n11660), .B2(n20409), .A(n11659), .ZN(n11666) );
  AOI22_X1 U13302 ( .A1(n11620), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11644), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U13303 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11691), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11663) );
  NAND3_X1 U13304 ( .A1(n11664), .A2(n11663), .A3(n11662), .ZN(n11665) );
  NAND2_X2 U13305 ( .A1(n11477), .A2(n11667), .ZN(n20965) );
  NAND2_X1 U13306 ( .A1(n20835), .A2(n20965), .ZN(n11729) );
  AOI22_X1 U13307 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U13308 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17927), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U13309 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17942), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11668) );
  OAI21_X1 U13310 ( .B1(n20409), .B2(n17891), .A(n11668), .ZN(n11674) );
  AOI22_X1 U13311 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U13312 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U13313 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U13314 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U13315 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  AOI211_X1 U13316 ( .C1(n11661), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n11674), .B(n11673), .ZN(n11675) );
  NAND3_X1 U13317 ( .A1(n11677), .A2(n11676), .A3(n11675), .ZN(n20825) );
  NAND2_X1 U13318 ( .A1(n11707), .A2(n20825), .ZN(n11710) );
  AOI22_X1 U13319 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U13320 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U13321 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17942), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11678) );
  OAI21_X1 U13322 ( .B1(n20409), .B2(n17815), .A(n11678), .ZN(n11684) );
  AOI22_X1 U13323 ( .A1(n11547), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U13324 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17803), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U13325 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U13326 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17927), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11679) );
  NAND4_X1 U13327 ( .A1(n11682), .A2(n11681), .A3(n11680), .A4(n11679), .ZN(
        n11683) );
  AOI211_X1 U13328 ( .C1(n11661), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n11684), .B(n11683), .ZN(n11685) );
  NAND3_X1 U13329 ( .A1(n11687), .A2(n11686), .A3(n11685), .ZN(n20816) );
  INV_X1 U13330 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21116) );
  OAI21_X1 U13331 ( .B1(n11688), .B2(n13226), .A(n18258), .ZN(n11718) );
  INV_X1 U13332 ( .A(n20965), .ZN(n11720) );
  INV_X1 U13333 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20982) );
  XNOR2_X1 U13334 ( .A(n20965), .B(n20982), .ZN(n18335) );
  AOI22_X1 U13335 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U13336 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11699) );
  INV_X1 U13337 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17770) );
  AOI22_X1 U13338 ( .A1(n17588), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11549), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11689) );
  OAI21_X1 U13339 ( .B1(n20409), .B2(n17770), .A(n11689), .ZN(n11697) );
  AOI22_X1 U13340 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11620), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U13341 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11621), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U13342 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11691), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U13343 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11692) );
  NAND4_X1 U13344 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n11696) );
  NAND3_X1 U13345 ( .A1(n11700), .A2(n11699), .A3(n11698), .ZN(n20971) );
  NAND2_X1 U13346 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20971), .ZN(
        n18344) );
  NOR2_X1 U13347 ( .A1(n18335), .A2(n18344), .ZN(n18334) );
  AOI21_X1 U13348 ( .B1(n11720), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18334), .ZN(n18326) );
  XNOR2_X1 U13349 ( .A(n20835), .B(n20965), .ZN(n11702) );
  NOR2_X1 U13350 ( .A1(n18326), .A2(n18325), .ZN(n18324) );
  NOR2_X1 U13351 ( .A1(n11701), .A2(n11702), .ZN(n11703) );
  NOR2_X1 U13352 ( .A1(n18324), .A2(n11703), .ZN(n11705) );
  XNOR2_X1 U13353 ( .A(n20830), .B(n11729), .ZN(n18315) );
  NOR2_X1 U13354 ( .A1(n11705), .A2(n11704), .ZN(n11706) );
  XNOR2_X1 U13355 ( .A(n20825), .B(n11707), .ZN(n11708) );
  XOR2_X1 U13356 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11708), .Z(
        n18304) );
  INV_X1 U13357 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21095) );
  NOR2_X1 U13358 ( .A1(n21095), .A2(n11708), .ZN(n11709) );
  NOR2_X2 U13359 ( .A1(n18303), .A2(n11709), .ZN(n11713) );
  XNOR2_X1 U13360 ( .A(n20820), .B(n11710), .ZN(n11712) );
  NOR2_X1 U13361 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  INV_X1 U13362 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21112) );
  XOR2_X1 U13363 ( .A(n20816), .B(n11715), .Z(n11716) );
  XOR2_X1 U13364 ( .A(n21112), .B(n11716), .Z(n18282) );
  XNOR2_X1 U13365 ( .A(n11718), .B(n11717), .ZN(n18270) );
  NOR2_X1 U13366 ( .A1(n21116), .A2(n18270), .ZN(n18269) );
  NOR2_X1 U13367 ( .A1(n11717), .A2(n11718), .ZN(n11719) );
  NAND2_X1 U13368 ( .A1(n18258), .A2(n18260), .ZN(n18211) );
  INV_X1 U13369 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21122) );
  NAND2_X1 U13370 ( .A1(n21163), .A2(n21135), .ZN(n18204) );
  NAND2_X1 U13371 ( .A1(n13194), .A2(n18107), .ZN(n21234) );
  INV_X1 U13372 ( .A(n21234), .ZN(n21220) );
  NAND2_X1 U13373 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13836) );
  INV_X1 U13374 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21250) );
  NOR2_X1 U13375 ( .A1(n13836), .A2(n21250), .ZN(n18167) );
  NAND2_X1 U13376 ( .A1(n21220), .A2(n18167), .ZN(n21252) );
  NAND2_X2 U13377 ( .A1(n19220), .A2(n21443), .ZN(n18351) );
  INV_X1 U13378 ( .A(n20971), .ZN(n11731) );
  NOR2_X1 U13379 ( .A1(n11720), .A2(n11731), .ZN(n11732) );
  NOR2_X1 U13380 ( .A1(n11732), .A2(n20835), .ZN(n11726) );
  NOR2_X1 U13381 ( .A1(n20830), .A2(n11726), .ZN(n11725) );
  NAND2_X1 U13382 ( .A1(n11725), .A2(n20825), .ZN(n11723) );
  NOR2_X1 U13383 ( .A1(n20820), .A2(n11723), .ZN(n11722) );
  NAND2_X1 U13384 ( .A1(n11722), .A2(n20816), .ZN(n11721) );
  NOR2_X1 U13385 ( .A1(n20812), .A2(n11721), .ZN(n11747) );
  XOR2_X1 U13386 ( .A(n20812), .B(n11721), .Z(n18273) );
  XOR2_X1 U13387 ( .A(n20816), .B(n11722), .Z(n11740) );
  XOR2_X1 U13388 ( .A(n20820), .B(n11723), .Z(n11724) );
  NAND2_X1 U13389 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11724), .ZN(
        n11739) );
  XOR2_X1 U13390 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11724), .Z(
        n18293) );
  XOR2_X1 U13391 ( .A(n20825), .B(n11725), .Z(n11736) );
  INV_X1 U13392 ( .A(n11726), .ZN(n11728) );
  XNOR2_X1 U13393 ( .A(n20830), .B(n11728), .ZN(n11727) );
  NAND2_X1 U13394 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11727), .ZN(
        n11735) );
  XOR2_X1 U13395 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11727), .Z(
        n18313) );
  OAI21_X1 U13396 ( .B1(n11731), .B2(n11729), .A(n11728), .ZN(n11730) );
  NAND2_X1 U13397 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11730), .ZN(
        n11734) );
  XNOR2_X1 U13398 ( .A(n11701), .B(n11730), .ZN(n18330) );
  NOR2_X1 U13399 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20965), .ZN(
        n11733) );
  INV_X1 U13400 ( .A(n18335), .ZN(n18337) );
  INV_X1 U13401 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21137) );
  NAND2_X1 U13402 ( .A1(n11731), .A2(n21137), .ZN(n18343) );
  NOR2_X1 U13403 ( .A1(n18337), .A2(n18343), .ZN(n18336) );
  NOR3_X1 U13404 ( .A1(n11733), .A2(n11732), .A3(n18336), .ZN(n18329) );
  NAND2_X1 U13405 ( .A1(n18330), .A2(n18329), .ZN(n18328) );
  NAND2_X1 U13406 ( .A1(n11734), .A2(n18328), .ZN(n18312) );
  NAND2_X1 U13407 ( .A1(n18313), .A2(n18312), .ZN(n18311) );
  NAND2_X1 U13408 ( .A1(n11736), .A2(n11737), .ZN(n11738) );
  NAND2_X1 U13409 ( .A1(n18293), .A2(n18292), .ZN(n18291) );
  NAND2_X1 U13410 ( .A1(n11740), .A2(n11741), .ZN(n11742) );
  NAND2_X1 U13411 ( .A1(n11747), .A2(n11743), .ZN(n11748) );
  INV_X1 U13412 ( .A(n11743), .ZN(n11746) );
  NAND2_X1 U13413 ( .A1(n18273), .A2(n18272), .ZN(n11745) );
  NAND2_X1 U13414 ( .A1(n11747), .A2(n11746), .ZN(n11744) );
  NAND2_X1 U13415 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18249), .ZN(
        n18248) );
  NAND2_X1 U13416 ( .A1(n13194), .A2(n18101), .ZN(n18137) );
  INV_X1 U13417 ( .A(n18137), .ZN(n21236) );
  NAND2_X1 U13418 ( .A1(n21236), .A2(n18167), .ZN(n21251) );
  AOI22_X1 U13419 ( .A1(n18262), .A2(n21252), .B1(n18275), .B2(n21251), .ZN(
        n18177) );
  AOI211_X1 U13420 ( .C1(n21245), .C2(n18275), .A(n21244), .B(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11768) );
  INV_X1 U13421 ( .A(n13194), .ZN(n18138) );
  NOR2_X1 U13422 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18226) );
  INV_X1 U13423 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18220) );
  AND2_X1 U13424 ( .A1(n18226), .A2(n18220), .ZN(n11750) );
  INV_X1 U13425 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U13426 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  NAND2_X1 U13427 ( .A1(n18001), .A2(n18205), .ZN(n11754) );
  NAND2_X1 U13428 ( .A1(n21163), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18006) );
  INV_X1 U13429 ( .A(n18006), .ZN(n21183) );
  NAND2_X1 U13430 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21183), .ZN(
        n21322) );
  NOR2_X1 U13431 ( .A1(n18221), .A2(n21322), .ZN(n11757) );
  INV_X1 U13432 ( .A(n11757), .ZN(n11758) );
  NAND2_X1 U13433 ( .A1(n11759), .A2(n11758), .ZN(n18011) );
  INV_X1 U13434 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17985) );
  NOR3_X1 U13435 ( .A1(n17988), .A2(n13833), .A3(n17985), .ZN(n18050) );
  NAND2_X1 U13436 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18048), .ZN(
        n13197) );
  INV_X1 U13437 ( .A(n13197), .ZN(n13193) );
  NAND2_X1 U13438 ( .A1(n13193), .A2(n18011), .ZN(n11762) );
  NOR2_X1 U13439 ( .A1(n13191), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18072) );
  INV_X1 U13440 ( .A(n18072), .ZN(n17981) );
  NOR4_X1 U13441 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n17981), .ZN(n18051) );
  NAND2_X1 U13442 ( .A1(n18051), .A2(n18095), .ZN(n18096) );
  OAI21_X1 U13443 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n18258), .ZN(n11765) );
  NAND2_X1 U13444 ( .A1(n18258), .A2(n18118), .ZN(n18158) );
  OR2_X2 U13445 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11766), .ZN(
        n13190) );
  NAND2_X1 U13446 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11766), .ZN(
        n13189) );
  NAND2_X1 U13447 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n13191), .ZN(
        n13192) );
  NOR2_X1 U13448 ( .A1(n13819), .A2(n13818), .ZN(n11767) );
  XOR2_X1 U13449 ( .A(n11767), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n21257) );
  OAI22_X1 U13450 ( .A1(n18177), .A2(n11768), .B1(n21257), .B2(n18187), .ZN(
        n11777) );
  NAND2_X1 U13451 ( .A1(n21438), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18346) );
  NAND2_X1 U13452 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n15367) );
  INV_X1 U13453 ( .A(n15367), .ZN(n17972) );
  NOR2_X1 U13454 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17972), .ZN(n20319) );
  AOI21_X4 U13455 ( .B1(n20319), .B2(n21438), .A(n21443), .ZN(n18318) );
  NOR2_X1 U13456 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18181), .ZN(
        n13825) );
  INV_X1 U13457 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21855) );
  INV_X2 U13458 ( .A(n18318), .ZN(n18345) );
  NOR2_X1 U13459 ( .A1(n13825), .A2(n18171), .ZN(n11775) );
  INV_X1 U13460 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20738) );
  NAND3_X1 U13461 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20481) );
  NOR3_X2 U13462 ( .A1(n20482), .A2(n20481), .A3(n20496), .ZN(n18213) );
  NAND2_X1 U13463 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18035) );
  NAND2_X1 U13464 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18015) );
  INV_X1 U13465 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18182) );
  INV_X1 U13466 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20609) );
  INV_X1 U13467 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18075) );
  INV_X1 U13468 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18087) );
  INV_X1 U13469 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18150) );
  INV_X1 U13470 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18130) );
  NAND2_X1 U13471 ( .A1(n11771), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11790) );
  NAND2_X1 U13472 ( .A1(n11771), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13823) );
  AOI21_X1 U13473 ( .B1(n20738), .B2(n11790), .A(n11778), .ZN(n11769) );
  INV_X1 U13474 ( .A(n11769), .ZN(n20743) );
  INV_X1 U13475 ( .A(n18346), .ZN(n18086) );
  INV_X1 U13476 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18347) );
  INV_X1 U13477 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21417) );
  NAND2_X1 U13478 ( .A1(n18347), .A2(n21417), .ZN(n21430) );
  INV_X1 U13479 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21413) );
  NAND2_X1 U13480 ( .A1(n21413), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21429) );
  AOI21_X1 U13481 ( .B1(n21430), .B2(n15367), .A(n21026), .ZN(n18941) );
  NAND3_X1 U13482 ( .A1(n21417), .A2(n21426), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18976) );
  INV_X2 U13483 ( .A(n18333), .ZN(n19264) );
  AOI22_X1 U13484 ( .A1(n18086), .A2(n11790), .B1(n19264), .B2(n13823), .ZN(
        n11770) );
  NAND2_X1 U13485 ( .A1(n11770), .A2(n18345), .ZN(n13824) );
  INV_X1 U13486 ( .A(n11771), .ZN(n11772) );
  OAI21_X1 U13487 ( .B1(n11772), .B2(n18333), .A(n20738), .ZN(n11773) );
  NOR2_X1 U13488 ( .A1(n21430), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17969) );
  NAND2_X2 U13489 ( .A1(n21438), .A2(n17969), .ZN(n21329) );
  INV_X1 U13490 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18442) );
  NOR2_X1 U13491 ( .A1(n21329), .A2(n18442), .ZN(n21249) );
  XNOR2_X1 U13492 ( .A(n11778), .B(n11259), .ZN(n20757) );
  INV_X1 U13493 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20763) );
  INV_X1 U13494 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18104) );
  NAND2_X1 U13495 ( .A1(n18103), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11781) );
  NOR2_X1 U13496 ( .A1(n18104), .A2(n11781), .ZN(n11780) );
  NOR2_X1 U13497 ( .A1(n18151), .A2(n20374), .ZN(n18127) );
  INV_X1 U13498 ( .A(n18127), .ZN(n11779) );
  OAI21_X1 U13499 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n11780), .A(
        n11779), .ZN(n20692) );
  XNOR2_X1 U13500 ( .A(n18104), .B(n11781), .ZN(n20676) );
  NOR2_X1 U13501 ( .A1(n18088), .A2(n20374), .ZN(n11782) );
  OAI21_X1 U13502 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n11782), .A(
        n11781), .ZN(n20666) );
  INV_X1 U13503 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20636) );
  NAND2_X1 U13504 ( .A1(n11100), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11787) );
  NOR2_X1 U13505 ( .A1(n20636), .A2(n11787), .ZN(n11783) );
  INV_X1 U13506 ( .A(n11782), .ZN(n18085) );
  OAI21_X1 U13507 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11783), .A(
        n18085), .ZN(n20651) );
  NOR2_X1 U13508 ( .A1(n18076), .A2(n20374), .ZN(n11784) );
  OAI21_X1 U13509 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11784), .A(
        n11787), .ZN(n20627) );
  NOR2_X1 U13510 ( .A1(n17991), .A2(n20374), .ZN(n11785) );
  INV_X1 U13511 ( .A(n11784), .ZN(n18054) );
  OAI21_X1 U13512 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11785), .A(
        n18054), .ZN(n20617) );
  NAND2_X1 U13513 ( .A1(n17976), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17977) );
  AOI21_X1 U13514 ( .B1(n11268), .B2(n17977), .A(n11785), .ZN(n11786) );
  INV_X1 U13515 ( .A(n11786), .ZN(n20603) );
  NOR2_X1 U13516 ( .A1(n20374), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20384) );
  INV_X1 U13517 ( .A(n20384), .ZN(n20521) );
  NOR2_X1 U13518 ( .A1(n18183), .A2(n20374), .ZN(n18012) );
  OAI21_X1 U13519 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18012), .A(
        n17977), .ZN(n18195) );
  NAND2_X1 U13520 ( .A1(n20580), .A2(n14253), .ZN(n20602) );
  NAND2_X1 U13521 ( .A1(n20603), .A2(n20602), .ZN(n20601) );
  NAND2_X1 U13522 ( .A1(n20580), .A2(n20601), .ZN(n20616) );
  XOR2_X1 U13523 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n11787), .Z(
        n20641) );
  NAND2_X1 U13524 ( .A1(n20580), .A2(n20639), .ZN(n20650) );
  NAND2_X1 U13525 ( .A1(n20651), .A2(n20650), .ZN(n20649) );
  NAND2_X1 U13526 ( .A1(n20580), .A2(n20649), .ZN(n20665) );
  NAND2_X1 U13527 ( .A1(n20666), .A2(n20665), .ZN(n20664) );
  NAND2_X1 U13528 ( .A1(n20580), .A2(n20664), .ZN(n20675) );
  NAND2_X1 U13529 ( .A1(n20676), .A2(n20675), .ZN(n20674) );
  NAND2_X1 U13530 ( .A1(n20580), .A2(n20674), .ZN(n20691) );
  NAND2_X1 U13531 ( .A1(n20692), .A2(n20691), .ZN(n20690) );
  NAND2_X1 U13532 ( .A1(n20580), .A2(n20690), .ZN(n20700) );
  NAND2_X1 U13533 ( .A1(n11101), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11788) );
  OAI21_X1 U13534 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18127), .A(
        n11788), .ZN(n20699) );
  NAND2_X1 U13535 ( .A1(n20700), .A2(n20699), .ZN(n20698) );
  NAND2_X1 U13536 ( .A1(n20580), .A2(n20698), .ZN(n20713) );
  NOR2_X1 U13537 ( .A1(n18131), .A2(n20374), .ZN(n11791) );
  AOI21_X1 U13538 ( .B1(n11261), .B2(n11788), .A(n11791), .ZN(n11789) );
  INV_X1 U13539 ( .A(n11789), .ZN(n20714) );
  NAND2_X1 U13540 ( .A1(n20580), .A2(n20712), .ZN(n20725) );
  OAI21_X1 U13541 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11791), .A(
        n11790), .ZN(n20726) );
  NAND2_X1 U13542 ( .A1(n20580), .A2(n20724), .ZN(n20742) );
  NAND2_X1 U13543 ( .A1(n20580), .A2(n20756), .ZN(n11792) );
  XNOR2_X1 U13544 ( .A(n20757), .B(n11792), .ZN(n11793) );
  NAND4_X1 U13545 ( .A1(n21438), .A2(n21417), .A3(n21855), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n21422) );
  INV_X1 U13546 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20720) );
  NAND2_X1 U13547 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n11797) );
  NAND3_X1 U13548 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .ZN(n11796) );
  INV_X1 U13549 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n21342) );
  INV_X1 U13550 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18431) );
  NAND2_X1 U13551 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n20554) );
  NOR2_X1 U13552 ( .A1(n18431), .A2(n20554), .ZN(n20577) );
  NAND2_X1 U13553 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n20577), .ZN(n20587) );
  NOR2_X1 U13554 ( .A1(n21342), .A2(n20587), .ZN(n14251) );
  NAND2_X1 U13555 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n14251), .ZN(n11801) );
  INV_X1 U13556 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18428) );
  INV_X1 U13557 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20484) );
  INV_X1 U13558 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n21102) );
  INV_X1 U13559 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20408) );
  NAND3_X1 U13560 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20407) );
  NOR2_X1 U13561 ( .A1(n20408), .A2(n20407), .ZN(n20432) );
  NAND2_X1 U13562 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20432), .ZN(n20429) );
  NOR2_X1 U13563 ( .A1(n21102), .A2(n20429), .ZN(n20455) );
  NAND2_X1 U13564 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20455), .ZN(n20483) );
  NOR2_X1 U13565 ( .A1(n20484), .A2(n20483), .ZN(n20472) );
  NAND2_X1 U13566 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20472), .ZN(n20491) );
  NOR2_X1 U13567 ( .A1(n18428), .A2(n20491), .ZN(n11800) );
  NOR2_X1 U13568 ( .A1(n21426), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18992) );
  AND2_X1 U13569 ( .A1(n21419), .A2(n18992), .ZN(n21433) );
  NOR4_X2 U13570 ( .A1(n10995), .A2(n20369), .A3(n21433), .A4(n20741), .ZN(
        n20430) );
  NAND3_X1 U13571 ( .A1(n11800), .A2(P3_REIP_REG_11__SCAN_IN), .A3(n20768), 
        .ZN(n20552) );
  NOR2_X1 U13572 ( .A1(n11801), .A2(n20552), .ZN(n14252) );
  NAND4_X1 U13573 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(P3_REIP_REG_19__SCAN_IN), .A4(n14252), .ZN(n20621) );
  NOR2_X1 U13574 ( .A1(n11796), .A2(n20621), .ZN(n20659) );
  NAND2_X1 U13575 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20659), .ZN(n20683) );
  NOR2_X1 U13576 ( .A1(n11797), .A2(n20683), .ZN(n20696) );
  NAND2_X1 U13577 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n20696), .ZN(n20722) );
  NOR2_X1 U13578 ( .A1(n20720), .A2(n20722), .ZN(n11799) );
  INV_X1 U13579 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21861) );
  NAND2_X1 U13580 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21861), .ZN(n21905) );
  INV_X2 U13581 ( .A(n11798), .ZN(n21864) );
  AOI21_X1 U13582 ( .B1(n11798), .B2(n21905), .A(n18438), .ZN(n20312) );
  NAND2_X1 U13583 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21907) );
  OAI211_X1 U13584 ( .C1(n20312), .C2(n20779), .A(n21907), .B(n21855), .ZN(
        n11805) );
  NOR2_X2 U13585 ( .A1(n11805), .A2(n17094), .ZN(n20456) );
  NAND2_X1 U13586 ( .A1(n20492), .A2(n20768), .ZN(n20766) );
  AOI21_X1 U13587 ( .B1(n11799), .B2(P3_REIP_REG_29__SCAN_IN), .A(n20719), 
        .ZN(n20751) );
  INV_X1 U13588 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18441) );
  INV_X1 U13589 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20671) );
  INV_X1 U13590 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n21146) );
  NAND2_X1 U13591 ( .A1(n20456), .A2(n11800), .ZN(n20519) );
  NOR2_X2 U13592 ( .A1(n21146), .A2(n20519), .ZN(n20576) );
  INV_X1 U13593 ( .A(n20576), .ZN(n20586) );
  NAND3_X1 U13594 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(P3_REIP_REG_19__SCAN_IN), .ZN(n11802) );
  NAND4_X1 U13595 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .A4(n20658), .ZN(n20670) );
  NAND3_X1 U13596 ( .A1(n20697), .A2(P3_REIP_REG_26__SCAN_IN), .A3(
        P3_REIP_REG_25__SCAN_IN), .ZN(n20717) );
  NOR2_X1 U13597 ( .A1(n18441), .A2(n20717), .ZN(n20721) );
  NAND2_X1 U13598 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n20721), .ZN(n20746) );
  NOR2_X1 U13599 ( .A1(n18442), .A2(n20746), .ZN(n20760) );
  INV_X1 U13600 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20750) );
  NAND2_X1 U13601 ( .A1(n20760), .A2(n20750), .ZN(n20754) );
  NOR2_X1 U13602 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20389) );
  INV_X1 U13603 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20388) );
  NAND2_X1 U13604 ( .A1(n20389), .A2(n20388), .ZN(n20396) );
  NOR2_X1 U13605 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n20396), .ZN(n20421) );
  INV_X1 U13606 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20420) );
  NAND2_X1 U13607 ( .A1(n20421), .A2(n20420), .ZN(n20427) );
  NOR2_X1 U13608 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n20427), .ZN(n20447) );
  INV_X1 U13609 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20446) );
  NAND2_X1 U13610 ( .A1(n20447), .A2(n20446), .ZN(n20453) );
  NOR2_X1 U13611 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n20453), .ZN(n20468) );
  INV_X1 U13612 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20470) );
  NAND2_X1 U13613 ( .A1(n20468), .A2(n20470), .ZN(n20477) );
  NOR2_X1 U13614 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n20477), .ZN(n20494) );
  INV_X1 U13615 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20493) );
  NAND2_X1 U13616 ( .A1(n20494), .A2(n20493), .ZN(n20509) );
  INV_X1 U13617 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n20530) );
  NAND2_X1 U13618 ( .A1(n20531), .A2(n20530), .ZN(n20539) );
  INV_X1 U13619 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20562) );
  NAND2_X1 U13620 ( .A1(n20563), .A2(n20562), .ZN(n20571) );
  INV_X1 U13621 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n20592) );
  NAND2_X1 U13622 ( .A1(n20593), .A2(n20592), .ZN(n20591) );
  INV_X1 U13623 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20599) );
  NAND2_X1 U13624 ( .A1(n20597), .A2(n20599), .ZN(n20607) );
  NOR2_X1 U13625 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n20607), .ZN(n20629) );
  INV_X1 U13626 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n20628) );
  NAND2_X1 U13627 ( .A1(n20629), .A2(n20628), .ZN(n20634) );
  NOR2_X1 U13628 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n20634), .ZN(n20653) );
  INV_X1 U13629 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n20652) );
  NAND2_X1 U13630 ( .A1(n20653), .A2(n20652), .ZN(n20660) );
  NOR2_X1 U13631 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n20660), .ZN(n20678) );
  INV_X1 U13632 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20677) );
  NAND2_X1 U13633 ( .A1(n20678), .A2(n20677), .ZN(n20684) );
  NOR2_X1 U13634 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n20684), .ZN(n20702) );
  INV_X1 U13635 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n20701) );
  NAND2_X1 U13636 ( .A1(n20702), .A2(n20701), .ZN(n20707) );
  NOR2_X1 U13637 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n20707), .ZN(n20729) );
  INV_X1 U13638 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n20728) );
  NAND2_X1 U13639 ( .A1(n20729), .A2(n20728), .ZN(n20736) );
  NOR2_X1 U13640 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n20736), .ZN(n11806) );
  INV_X1 U13641 ( .A(n17094), .ZN(n11804) );
  NAND2_X1 U13642 ( .A1(n21907), .A2(n21855), .ZN(n11803) );
  NOR2_X1 U13643 ( .A1(n11806), .A2(n20764), .ZN(n20734) );
  INV_X1 U13644 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20747) );
  AOI22_X1 U13645 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20718), .B1(
        n20734), .B2(n20747), .ZN(n11808) );
  INV_X1 U13646 ( .A(n11805), .ZN(n21416) );
  AOI211_X4 U13647 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20779), .A(n21416), .B(
        n17094), .ZN(n20749) );
  AND2_X1 U13648 ( .A1(n20727), .A2(n11806), .ZN(n20748) );
  OAI21_X1 U13649 ( .B1(n20749), .B2(n20748), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n11807) );
  NAND2_X1 U13650 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  AOI22_X1 U13651 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11909), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11815) );
  AND2_X4 U13652 ( .A1(n11823), .A2(n11822), .ZN(n13642) );
  AOI22_X1 U13653 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U13654 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11998), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11820) );
  AND2_X2 U13655 ( .A1(n11822), .A2(n14584), .ZN(n11959) );
  AOI22_X1 U13656 ( .A1(n11992), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11819) );
  AND2_X2 U13657 ( .A1(n11823), .A2(n15009), .ZN(n11978) );
  AOI22_X1 U13658 ( .A1(n13636), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11978), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U13659 ( .A1(n12055), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13637), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U13660 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U13661 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U13662 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11827) );
  NAND4_X1 U13663 ( .A1(n11830), .A2(n11829), .A3(n11828), .A4(n11827), .ZN(
        n11836) );
  AOI22_X1 U13664 ( .A1(n11992), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11978), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U13665 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10991), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U13666 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11998), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11831) );
  NAND4_X1 U13667 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n11835) );
  NAND2_X1 U13668 ( .A1(n11926), .A2(n11931), .ZN(n11857) );
  AOI22_X1 U13669 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11909), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U13670 ( .A1(n12055), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13637), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U13671 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U13672 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11998), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U13673 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11904), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U13674 ( .A1(n11992), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U13675 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11978), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U13676 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11991), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U13677 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11904), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U13678 ( .A1(n11992), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U13679 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11978), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U13680 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11909), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U13681 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11998), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11853) );
  INV_X2 U13682 ( .A(n11932), .ZN(n11859) );
  MUX2_X1 U13683 ( .A(n11857), .B(n14712), .S(n11859), .Z(n11881) );
  AOI22_X1 U13684 ( .A1(n12055), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13637), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U13685 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U13686 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U13687 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11998), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U13688 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11978), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U13689 ( .A1(n11992), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U13690 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11904), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11864) );
  NAND2_X1 U13691 ( .A1(n11920), .A2(n14735), .ZN(n11948) );
  AOI22_X1 U13692 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13636), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U13693 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11991), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U13694 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11978), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U13695 ( .A1(n11992), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11870) );
  NAND4_X1 U13696 ( .A1(n11873), .A2(n11872), .A3(n11871), .A4(n11870), .ZN(
        n11879) );
  AOI22_X1 U13697 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11909), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U13698 ( .A1(n12055), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13637), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U13699 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11875) );
  NAND4_X1 U13700 ( .A1(n11877), .A2(n11876), .A3(n11875), .A4(n11874), .ZN(
        n11878) );
  AND4_X2 U13702 ( .A1(n11881), .A2(n11880), .A3(n11948), .A4(n14683), .ZN(
        n11933) );
  INV_X1 U13703 ( .A(n11933), .ZN(n11902) );
  NAND2_X1 U13704 ( .A1(n11904), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11885) );
  NAND2_X1 U13705 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11884) );
  NAND2_X1 U13706 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11883) );
  NAND2_X1 U13707 ( .A1(n11978), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11882) );
  NAND2_X1 U13708 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U13709 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11888) );
  NAND2_X1 U13710 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11887) );
  NAND2_X1 U13711 ( .A1(n11998), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11886) );
  NAND2_X1 U13712 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11893) );
  NAND2_X1 U13713 ( .A1(n11909), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11892) );
  NAND2_X1 U13714 ( .A1(n12055), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11891) );
  NAND2_X1 U13715 ( .A1(n13637), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11890) );
  NAND2_X1 U13716 ( .A1(n11992), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11897) );
  NAND2_X1 U13717 ( .A1(n11991), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11896) );
  NAND2_X1 U13718 ( .A1(n11031), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11895) );
  NAND2_X1 U13719 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11894) );
  NAND2_X1 U13720 ( .A1(n11902), .A2(n11026), .ZN(n12402) );
  AOI22_X1 U13721 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13637), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U13722 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U13723 ( .A1(n11991), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U13724 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11904), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U13725 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11978), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U13726 ( .A1(n11997), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11992), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U13727 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11998), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U13728 ( .A1(n11909), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11910) );
  AND2_X2 U13729 ( .A1(n14741), .A2(n11027), .ZN(n17144) );
  NAND2_X1 U13730 ( .A1(n11919), .A2(n17144), .ZN(n11918) );
  NAND2_X1 U13731 ( .A1(n11023), .A2(n11027), .ZN(n11916) );
  NAND2_X1 U13732 ( .A1(n21448), .A2(n11916), .ZN(n12396) );
  AOI21_X1 U13733 ( .B1(n10985), .B2(n12388), .A(n12396), .ZN(n11917) );
  NAND3_X1 U13734 ( .A1(n12402), .A2(n11918), .A3(n11917), .ZN(n11944) );
  INV_X1 U13735 ( .A(n11919), .ZN(n11921) );
  NAND2_X1 U13736 ( .A1(n11921), .A2(n11920), .ZN(n11923) );
  INV_X1 U13737 ( .A(n11930), .ZN(n11949) );
  NAND2_X1 U13738 ( .A1(n11945), .A2(n11949), .ZN(n11925) );
  AND2_X1 U13739 ( .A1(n12110), .A2(n14683), .ZN(n11927) );
  NAND2_X1 U13740 ( .A1(n21873), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21865) );
  NAND2_X1 U13741 ( .A1(n21872), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U13742 ( .A1(n21865), .A2(n11928), .ZN(n12217) );
  INV_X1 U13743 ( .A(n12391), .ZN(n12288) );
  AOI21_X1 U13744 ( .B1(n11103), .B2(n11478), .A(n12288), .ZN(n11934) );
  AND2_X2 U13745 ( .A1(n11934), .A2(n12287), .ZN(n11939) );
  NAND2_X1 U13746 ( .A1(n17081), .A2(n21832), .ZN(n13810) );
  XNOR2_X1 U13747 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21979) );
  NAND2_X1 U13748 ( .A1(n17148), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12017) );
  OAI21_X1 U13749 ( .B1(n13810), .B2(n21979), .A(n12017), .ZN(n11937) );
  INV_X1 U13750 ( .A(n11937), .ZN(n11938) );
  OAI21_X2 U13751 ( .B1(n12022), .B2(n14594), .A(n11938), .ZN(n11941) );
  INV_X1 U13752 ( .A(n11939), .ZN(n11940) );
  INV_X1 U13753 ( .A(n17148), .ZN(n11942) );
  MUX2_X1 U13754 ( .A(n11942), .B(n13810), .S(n22029), .Z(n11943) );
  INV_X1 U13755 ( .A(n11944), .ZN(n11954) );
  INV_X1 U13756 ( .A(n11945), .ZN(n11946) );
  NAND2_X1 U13757 ( .A1(n11946), .A2(n14749), .ZN(n11952) );
  INV_X1 U13758 ( .A(n15876), .ZN(n13735) );
  NAND2_X1 U13759 ( .A1(n14389), .A2(n11948), .ZN(n11951) );
  NAND2_X1 U13760 ( .A1(n11930), .A2(n11859), .ZN(n12405) );
  AND2_X1 U13761 ( .A1(n17081), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11950) );
  NAND2_X1 U13762 ( .A1(n11954), .A2(n11953), .ZN(n11988) );
  NAND2_X1 U13763 ( .A1(n11990), .A2(n11988), .ZN(n11956) );
  INV_X1 U13764 ( .A(n11956), .ZN(n11955) );
  AOI22_X1 U13765 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U13766 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U13767 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U13768 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11960) );
  NAND4_X1 U13769 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11970) );
  AOI22_X1 U13770 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U13771 ( .A1(n11031), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U13772 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U13773 ( .A1(n10989), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11965) );
  NAND4_X1 U13774 ( .A1(n11968), .A2(n11967), .A3(n11966), .A4(n11965), .ZN(
        n11969) );
  AOI22_X1 U13775 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U13776 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11909), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U13777 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U13778 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11974) );
  NAND4_X1 U13779 ( .A1(n11977), .A2(n11976), .A3(n11975), .A4(n11974), .ZN(
        n11984) );
  AOI22_X1 U13780 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U13781 ( .A1(n11031), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U13782 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U13783 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11979) );
  NAND4_X1 U13784 ( .A1(n11982), .A2(n11981), .A3(n11980), .A4(n11979), .ZN(
        n11983) );
  OR2_X1 U13785 ( .A1(n12032), .A2(n12181), .ZN(n11986) );
  NAND2_X1 U13786 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11985) );
  OAI211_X1 U13787 ( .C1(n11987), .C2(n12031), .A(n11986), .B(n11985), .ZN(
        n12015) );
  XNOR2_X1 U13788 ( .A(n12014), .B(n12015), .ZN(n13256) );
  INV_X1 U13789 ( .A(n12032), .ZN(n12006) );
  AOI22_X1 U13790 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U13791 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n13699), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U13792 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n10989), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U13793 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11993) );
  NAND4_X1 U13794 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n12004) );
  AOI22_X1 U13795 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U13796 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13701), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U13797 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U13798 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11999) );
  NAND4_X1 U13799 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n12003) );
  XNOR2_X1 U13800 ( .A(n12013), .B(n12109), .ZN(n12005) );
  NAND2_X1 U13801 ( .A1(n12006), .A2(n12005), .ZN(n12007) );
  INV_X1 U13802 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12012) );
  AOI21_X1 U13803 ( .B1(n12009), .B2(n12181), .A(n21832), .ZN(n12011) );
  NAND2_X1 U13804 ( .A1(n11026), .A2(n12109), .ZN(n12010) );
  INV_X1 U13805 ( .A(n12014), .ZN(n12107) );
  NAND2_X1 U13806 ( .A1(n12014), .A2(n12015), .ZN(n12016) );
  NAND2_X1 U13807 ( .A1(n12017), .A2(n14594), .ZN(n12018) );
  NAND2_X1 U13808 ( .A1(n12019), .A2(n12018), .ZN(n12020) );
  INV_X1 U13809 ( .A(n13810), .ZN(n12047) );
  NAND2_X1 U13810 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12024) );
  NAND2_X1 U13811 ( .A1(n22018), .A2(n12024), .ZN(n12026) );
  NAND2_X1 U13812 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22067) );
  INV_X1 U13813 ( .A(n22067), .ZN(n12025) );
  NAND2_X1 U13814 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12025), .ZN(
        n12045) );
  AND2_X1 U13815 ( .A1(n12026), .A2(n12045), .ZN(n15049) );
  AOI22_X1 U13816 ( .A1(n12047), .A2(n15049), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17148), .ZN(n12027) );
  OR2_X2 U13817 ( .A1(n12029), .A2(n12028), .ZN(n12030) );
  NAND2_X2 U13818 ( .A1(n12029), .A2(n12028), .ZN(n15011) );
  NAND2_X2 U13819 ( .A1(n12030), .A2(n15011), .ZN(n14536) );
  AOI22_X1 U13820 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U13821 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U13822 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U13823 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12033) );
  NAND4_X1 U13824 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n12042) );
  AOI22_X1 U13825 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U13826 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11909), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U13827 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U13828 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12037) );
  NAND4_X1 U13829 ( .A1(n12040), .A2(n12039), .A3(n12038), .A4(n12037), .ZN(
        n12041) );
  AOI22_X1 U13830 ( .A1(n12250), .A2(n12121), .B1(n12248), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12043) );
  OAI21_X2 U13831 ( .B1(n14536), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12043), 
        .ZN(n12118) );
  INV_X1 U13832 ( .A(n12022), .ZN(n12044) );
  NAND2_X1 U13833 ( .A1(n12044), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12049) );
  INV_X1 U13834 ( .A(n12045), .ZN(n22063) );
  NAND2_X1 U13835 ( .A1(n22063), .A2(n12225), .ZN(n14751) );
  NAND2_X1 U13836 ( .A1(n12045), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12046) );
  NAND2_X1 U13837 ( .A1(n14751), .A2(n12046), .ZN(n21980) );
  AOI22_X1 U13838 ( .A1(n12047), .A2(n21980), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17148), .ZN(n12048) );
  XNOR2_X2 U13839 ( .A(n15011), .B(n15010), .ZN(n14694) );
  NAND2_X1 U13840 ( .A1(n14694), .A2(n21832), .ZN(n12064) );
  AOI22_X1 U13841 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U13842 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U13843 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U13844 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12050) );
  NAND4_X1 U13845 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n12062) );
  AOI22_X1 U13846 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U13847 ( .A1(n12055), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U13848 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U13849 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12057) );
  NAND4_X1 U13850 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(
        n12061) );
  AOI22_X1 U13851 ( .A1(n12250), .A2(n12139), .B1(n12248), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U13852 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U13853 ( .A1(n11031), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U13854 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U13855 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12065) );
  NAND4_X1 U13856 ( .A1(n12068), .A2(n12067), .A3(n12066), .A4(n12065), .ZN(
        n12074) );
  AOI22_X1 U13857 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10989), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U13858 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U13859 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U13860 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12069) );
  NAND4_X1 U13861 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(
        n12073) );
  NAND2_X1 U13862 ( .A1(n12250), .A2(n12148), .ZN(n12076) );
  NAND2_X1 U13863 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12075) );
  AOI22_X1 U13864 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U13865 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U13866 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U13867 ( .A1(n11031), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U13868 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12086) );
  AOI22_X1 U13869 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U13870 ( .A1(n11909), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U13871 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U13872 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U13873 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12085) );
  NAND2_X1 U13874 ( .A1(n12250), .A2(n12159), .ZN(n12088) );
  NAND2_X1 U13875 ( .A1(n12248), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12087) );
  AOI22_X1 U13876 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U13877 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U13878 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U13879 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12089) );
  NAND4_X1 U13880 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12089), .ZN(
        n12098) );
  AOI22_X1 U13881 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11909), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U13882 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U13883 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U13884 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12093) );
  NAND4_X1 U13885 ( .A1(n12096), .A2(n12095), .A3(n12094), .A4(n12093), .ZN(
        n12097) );
  AOI22_X1 U13886 ( .A1(n12250), .A2(n12172), .B1(n12248), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12156) );
  INV_X1 U13887 ( .A(n12100), .ZN(n12101) );
  INV_X1 U13888 ( .A(n12246), .ZN(n12134) );
  NAND2_X4 U13889 ( .A1(n12170), .A2(n12102), .ZN(n12179) );
  NOR2_X1 U13890 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16183) );
  NAND2_X1 U13891 ( .A1(n11209), .A2(n16183), .ZN(n12205) );
  NAND2_X1 U13892 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16174) );
  INV_X1 U13893 ( .A(n16174), .ZN(n16184) );
  NAND2_X1 U13894 ( .A1(n16184), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12414) );
  INV_X1 U13895 ( .A(n17144), .ZN(n21446) );
  NAND2_X1 U13896 ( .A1(n11026), .A2(n14735), .ZN(n12122) );
  OAI21_X1 U13897 ( .B1(n21446), .B2(n12109), .A(n12122), .ZN(n12105) );
  INV_X1 U13898 ( .A(n12105), .ZN(n12106) );
  NAND2_X1 U13899 ( .A1(n12107), .A2(n12246), .ZN(n12114) );
  NAND2_X1 U13900 ( .A1(n12109), .A2(n12108), .ZN(n12132) );
  OAI21_X1 U13901 ( .B1(n12109), .B2(n12108), .A(n12132), .ZN(n12111) );
  OAI211_X1 U13902 ( .C1(n12111), .C2(n21446), .A(n12110), .B(n11858), .ZN(
        n12112) );
  INV_X1 U13903 ( .A(n12112), .ZN(n12113) );
  NAND2_X1 U13904 ( .A1(n20138), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20139) );
  INV_X1 U13905 ( .A(n12115), .ZN(n12116) );
  OR2_X1 U13906 ( .A1(n14526), .A2(n12116), .ZN(n12117) );
  NAND2_X1 U13907 ( .A1(n20139), .A2(n12117), .ZN(n12127) );
  INV_X1 U13908 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21479) );
  INV_X1 U13909 ( .A(n12118), .ZN(n12119) );
  XNOR2_X1 U13910 ( .A(n12120), .B(n12119), .ZN(n13251) );
  NAND2_X1 U13911 ( .A1(n13251), .A2(n12246), .ZN(n12126) );
  INV_X1 U13912 ( .A(n12121), .ZN(n12131) );
  XNOR2_X1 U13913 ( .A(n12132), .B(n12131), .ZN(n12124) );
  INV_X1 U13914 ( .A(n12122), .ZN(n12123) );
  AOI21_X1 U13915 ( .B1(n12124), .B2(n17144), .A(n12123), .ZN(n12125) );
  NAND2_X1 U13916 ( .A1(n12126), .A2(n12125), .ZN(n20144) );
  NAND2_X1 U13917 ( .A1(n12127), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12128) );
  INV_X1 U13918 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21496) );
  NAND2_X1 U13919 ( .A1(n12129), .A2(n15104), .ZN(n12130) );
  NAND2_X1 U13920 ( .A1(n12132), .A2(n12131), .ZN(n12140) );
  XNOR2_X1 U13921 ( .A(n12140), .B(n12139), .ZN(n12133) );
  OAI22_X1 U13922 ( .A1(n15107), .A2(n12134), .B1(n21446), .B2(n12133), .ZN(
        n20152) );
  NAND2_X1 U13923 ( .A1(n11009), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12136) );
  INV_X1 U13924 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21492) );
  NAND2_X1 U13925 ( .A1(n13249), .A2(n12246), .ZN(n12143) );
  NAND2_X1 U13926 ( .A1(n12140), .A2(n12139), .ZN(n12150) );
  XNOR2_X1 U13927 ( .A(n12150), .B(n12148), .ZN(n12141) );
  NAND2_X1 U13928 ( .A1(n12141), .A2(n17144), .ZN(n12142) );
  NAND2_X1 U13929 ( .A1(n12143), .A2(n12142), .ZN(n20159) );
  NAND2_X1 U13930 ( .A1(n11010), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12145) );
  XNOR2_X1 U13931 ( .A(n12147), .B(n12146), .ZN(n13285) );
  NAND2_X1 U13932 ( .A1(n13285), .A2(n12246), .ZN(n12153) );
  INV_X1 U13933 ( .A(n12148), .ZN(n12149) );
  OR2_X1 U13934 ( .A1(n12150), .A2(n12149), .ZN(n12158) );
  XNOR2_X1 U13935 ( .A(n12158), .B(n12159), .ZN(n12151) );
  NAND2_X1 U13936 ( .A1(n12151), .A2(n17144), .ZN(n12152) );
  NAND2_X1 U13937 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  INV_X1 U13938 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21462) );
  XNOR2_X1 U13939 ( .A(n12154), .B(n21462), .ZN(n20166) );
  NAND2_X1 U13940 ( .A1(n12154), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12155) );
  NAND2_X1 U13941 ( .A1(n12157), .A2(n12156), .ZN(n13286) );
  NAND3_X1 U13942 ( .A1(n12170), .A2(n13286), .A3(n12246), .ZN(n12163) );
  INV_X1 U13943 ( .A(n12158), .ZN(n12160) );
  NAND2_X1 U13944 ( .A1(n12160), .A2(n12159), .ZN(n12171) );
  XNOR2_X1 U13945 ( .A(n12171), .B(n12172), .ZN(n12161) );
  NAND2_X1 U13946 ( .A1(n12161), .A2(n17144), .ZN(n12162) );
  NAND2_X1 U13947 ( .A1(n12163), .A2(n12162), .ZN(n12164) );
  XNOR2_X1 U13948 ( .A(n12164), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20171) );
  INV_X1 U13949 ( .A(n12164), .ZN(n12165) );
  INV_X1 U13950 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21521) );
  NAND2_X1 U13951 ( .A1(n12165), .A2(n21521), .ZN(n12166) );
  NAND2_X1 U13952 ( .A1(n20174), .A2(n12166), .ZN(n20178) );
  INV_X1 U13953 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12168) );
  NAND2_X1 U13954 ( .A1(n12250), .A2(n12181), .ZN(n12167) );
  OAI21_X1 U13955 ( .B1(n12168), .B2(n12263), .A(n12167), .ZN(n12169) );
  NAND2_X1 U13956 ( .A1(n13296), .A2(n12246), .ZN(n12176) );
  INV_X1 U13957 ( .A(n12171), .ZN(n12173) );
  NAND2_X1 U13958 ( .A1(n12173), .A2(n12172), .ZN(n12180) );
  XNOR2_X1 U13959 ( .A(n12180), .B(n12181), .ZN(n12174) );
  NAND2_X1 U13960 ( .A1(n12174), .A2(n17144), .ZN(n12175) );
  NAND2_X1 U13961 ( .A1(n12176), .A2(n12175), .ZN(n12177) );
  XNOR2_X1 U13962 ( .A(n12177), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n20179) );
  INV_X1 U13963 ( .A(n12180), .ZN(n12182) );
  NAND3_X1 U13964 ( .A1(n12182), .A2(n17144), .A3(n12181), .ZN(n12183) );
  NAND2_X1 U13965 ( .A1(n12179), .A2(n12183), .ZN(n12184) );
  INV_X1 U13966 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21523) );
  XNOR2_X1 U13967 ( .A(n12184), .B(n21523), .ZN(n15289) );
  INV_X1 U13968 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12407) );
  XNOR2_X1 U13969 ( .A(n20231), .B(n12407), .ZN(n16155) );
  INV_X4 U13970 ( .A(n12193), .ZN(n20231) );
  NAND2_X1 U13971 ( .A1(n12193), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16120) );
  INV_X1 U13972 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12189) );
  NAND2_X1 U13973 ( .A1(n20231), .A2(n12189), .ZN(n12185) );
  NAND2_X1 U13974 ( .A1(n16120), .A2(n12185), .ZN(n16148) );
  INV_X1 U13975 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21556) );
  NAND2_X1 U13976 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12186) );
  NAND2_X1 U13977 ( .A1(n20231), .A2(n12186), .ZN(n16146) );
  NOR2_X1 U13978 ( .A1(n16148), .A2(n12187), .ZN(n16135) );
  INV_X1 U13979 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21464) );
  NAND2_X1 U13980 ( .A1(n20231), .A2(n21464), .ZN(n12188) );
  NAND2_X1 U13981 ( .A1(n16135), .A2(n12188), .ZN(n16122) );
  INV_X1 U13982 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21597) );
  NAND3_X1 U13983 ( .A1(n21597), .A2(n12189), .A3(n21464), .ZN(n12190) );
  NAND2_X1 U13984 ( .A1(n12193), .A2(n12190), .ZN(n12194) );
  NAND2_X1 U13985 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21589) );
  INV_X1 U13986 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21588) );
  NOR2_X1 U13987 ( .A1(n21589), .A2(n21588), .ZN(n21585) );
  INV_X1 U13988 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12323) );
  INV_X1 U13989 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12191) );
  NAND2_X1 U13990 ( .A1(n12323), .A2(n12191), .ZN(n12192) );
  NAND2_X1 U13991 ( .A1(n12193), .A2(n12192), .ZN(n16144) );
  NAND2_X1 U13992 ( .A1(n12193), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16147) );
  NAND2_X1 U13993 ( .A1(n16144), .A2(n16147), .ZN(n16132) );
  INV_X1 U13994 ( .A(n12194), .ZN(n20215) );
  NAND3_X1 U13995 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16247) );
  INV_X1 U13996 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12349) );
  NOR2_X1 U13997 ( .A1(n16247), .A2(n12349), .ZN(n12196) );
  INV_X1 U13998 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12355) );
  INV_X1 U13999 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U14000 ( .A1(n21629), .A2(n12355), .A3(n12197), .A4(n12349), .ZN(
        n12198) );
  OAI21_X1 U14001 ( .B1(n16105), .B2(n12198), .A(n11209), .ZN(n16097) );
  INV_X1 U14002 ( .A(n16044), .ZN(n12200) );
  INV_X1 U14003 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16223) );
  INV_X1 U14004 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16073) );
  INV_X1 U14005 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16228) );
  NAND3_X1 U14006 ( .A1(n16223), .A2(n16073), .A3(n16228), .ZN(n16046) );
  INV_X1 U14007 ( .A(n16046), .ZN(n12199) );
  NAND2_X1 U14008 ( .A1(n12202), .A2(n20231), .ZN(n16071) );
  AND2_X1 U14009 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16214) );
  NAND2_X1 U14010 ( .A1(n16214), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16204) );
  NAND2_X1 U14011 ( .A1(n12179), .A2(n16204), .ZN(n16045) );
  AND2_X1 U14012 ( .A1(n16071), .A2(n16045), .ZN(n12203) );
  MUX2_X1 U14013 ( .A(n12205), .B(n12414), .S(n16057), .Z(n12206) );
  AND2_X1 U14014 ( .A1(n11209), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16034) );
  NOR2_X2 U14015 ( .A1(n12206), .A2(n16034), .ZN(n12207) );
  XNOR2_X1 U14016 ( .A(n12207), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16032) );
  INV_X1 U14017 ( .A(n12208), .ZN(n12214) );
  NAND2_X1 U14018 ( .A1(n10985), .A2(n11859), .ZN(n12210) );
  AND2_X1 U14019 ( .A1(n12210), .A2(n12209), .ZN(n12394) );
  NAND2_X1 U14020 ( .A1(n15380), .A2(n11026), .ZN(n12211) );
  INV_X1 U14021 ( .A(n13808), .ZN(n12213) );
  MUX2_X1 U14022 ( .A(n11919), .B(n14741), .S(n11922), .Z(n12212) );
  AND2_X1 U14023 ( .A1(n12212), .A2(n11027), .ZN(n12403) );
  AOI21_X1 U14024 ( .B1(n12214), .B2(n12213), .A(n12403), .ZN(n14552) );
  INV_X1 U14025 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12216) );
  NAND2_X1 U14026 ( .A1(n12217), .A2(n12216), .ZN(n21875) );
  INV_X1 U14027 ( .A(n21875), .ZN(n21447) );
  NAND2_X1 U14028 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21455) );
  OAI21_X1 U14029 ( .B1(n14749), .B2(n21447), .A(n21455), .ZN(n13773) );
  INV_X1 U14030 ( .A(n13773), .ZN(n12218) );
  NAND2_X1 U14031 ( .A1(n17146), .A2(n12218), .ZN(n12219) );
  NAND3_X1 U14032 ( .A1(n12219), .A2(n11027), .A3(n13749), .ZN(n12273) );
  NAND2_X1 U14033 ( .A1(n21944), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12221) );
  NAND2_X1 U14034 ( .A1(n14594), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12220) );
  NAND2_X1 U14035 ( .A1(n12221), .A2(n12220), .ZN(n12245) );
  NAND2_X1 U14036 ( .A1(n12222), .A2(n12221), .ZN(n12238) );
  NAND2_X1 U14037 ( .A1(n22018), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12224) );
  NAND2_X1 U14038 ( .A1(n12023), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12223) );
  NAND2_X1 U14039 ( .A1(n12238), .A2(n12237), .ZN(n12236) );
  NAND2_X1 U14040 ( .A1(n12236), .A2(n12224), .ZN(n12228) );
  NAND2_X1 U14041 ( .A1(n12228), .A2(n12229), .ZN(n12232) );
  INV_X1 U14042 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17156) );
  NAND2_X1 U14043 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17156), .ZN(
        n12226) );
  NAND2_X1 U14044 ( .A1(n12225), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12230) );
  NAND3_X1 U14045 ( .A1(n12232), .A2(n12226), .A3(n12230), .ZN(n12227) );
  NAND2_X1 U14046 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17084), .ZN(
        n12233) );
  NAND2_X1 U14047 ( .A1(n12250), .A2(n12279), .ZN(n12272) );
  NAND2_X1 U14048 ( .A1(n12265), .A2(n12279), .ZN(n12270) );
  AOI21_X1 U14049 ( .B1(n12229), .B2(n12230), .A(n12228), .ZN(n12235) );
  INV_X1 U14050 ( .A(n12230), .ZN(n12231) );
  AOI21_X1 U14051 ( .B1(n12233), .B2(n12232), .A(n12231), .ZN(n12234) );
  OAI21_X1 U14052 ( .B1(n12238), .B2(n12237), .A(n12236), .ZN(n12275) );
  INV_X1 U14053 ( .A(n12275), .ZN(n12257) );
  NAND2_X1 U14054 ( .A1(n12257), .A2(n12250), .ZN(n12255) );
  INV_X1 U14055 ( .A(n12255), .ZN(n12261) );
  OAI21_X1 U14056 ( .B1(n11008), .B2(n22029), .A(n12243), .ZN(n12239) );
  AOI211_X1 U14057 ( .C1(n10985), .C2(n11027), .A(n12239), .B(n12260), .ZN(
        n12242) );
  INV_X1 U14058 ( .A(n12239), .ZN(n12240) );
  AOI21_X1 U14059 ( .B1(n12250), .B2(n12240), .A(n12265), .ZN(n12241) );
  NOR2_X1 U14060 ( .A1(n12242), .A2(n12241), .ZN(n12249) );
  INV_X1 U14061 ( .A(n12243), .ZN(n12244) );
  XNOR2_X1 U14062 ( .A(n12245), .B(n12244), .ZN(n12277) );
  NOR3_X1 U14063 ( .A1(n12246), .A2(n12249), .A3(n12277), .ZN(n12254) );
  INV_X1 U14064 ( .A(n12277), .ZN(n12247) );
  AOI22_X1 U14065 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n10993), .B1(n12248), 
        .B2(n12247), .ZN(n12253) );
  OAI21_X1 U14066 ( .B1(n14749), .B2(n12277), .A(n12249), .ZN(n12252) );
  NAND3_X1 U14067 ( .A1(n12250), .A2(n14749), .A3(n12277), .ZN(n12251) );
  OAI211_X1 U14068 ( .C1(n12254), .C2(n12253), .A(n12252), .B(n12251), .ZN(
        n12259) );
  INV_X1 U14069 ( .A(n12260), .ZN(n12256) );
  OAI211_X1 U14070 ( .C1(n12257), .C2(n12263), .A(n12256), .B(n12255), .ZN(
        n12258) );
  AOI22_X1 U14071 ( .A1(n12261), .A2(n12260), .B1(n12259), .B2(n12258), .ZN(
        n12262) );
  AOI21_X1 U14072 ( .B1(n12263), .B2(n12274), .A(n12262), .ZN(n12264) );
  AOI21_X1 U14073 ( .B1(n12265), .B2(n12274), .A(n12264), .ZN(n12266) );
  INV_X1 U14074 ( .A(n12266), .ZN(n12267) );
  INV_X1 U14075 ( .A(n12268), .ZN(n12269) );
  NAND2_X1 U14076 ( .A1(n12273), .A2(n15389), .ZN(n12282) );
  NOR2_X1 U14077 ( .A1(n12275), .A2(n12274), .ZN(n12276) );
  NAND2_X1 U14078 ( .A1(n14396), .A2(n21455), .ZN(n13733) );
  AND2_X1 U14079 ( .A1(n14749), .A2(n21875), .ZN(n12280) );
  OR2_X1 U14080 ( .A1(n13733), .A2(n12280), .ZN(n12281) );
  MUX2_X1 U14081 ( .A(n12282), .B(n12281), .S(n11023), .Z(n12284) );
  INV_X1 U14082 ( .A(n15389), .ZN(n14548) );
  NAND3_X1 U14083 ( .A1(n14548), .A2(n13422), .A3(n14749), .ZN(n12283) );
  NAND3_X1 U14084 ( .A1(n14552), .A2(n12284), .A3(n12283), .ZN(n12285) );
  NAND2_X1 U14085 ( .A1(n13808), .A2(n10985), .ZN(n12286) );
  INV_X1 U14086 ( .A(n12110), .ZN(n12398) );
  NOR2_X1 U14087 ( .A1(n12398), .A2(n15380), .ZN(n14533) );
  NAND2_X1 U14088 ( .A1(n14533), .A2(n15876), .ZN(n13729) );
  AND2_X1 U14089 ( .A1(n12286), .A2(n13729), .ZN(n14394) );
  AND2_X2 U14090 ( .A1(n14749), .A2(n11929), .ZN(n12380) );
  NAND2_X1 U14091 ( .A1(n17146), .A2(n12380), .ZN(n13730) );
  NAND2_X1 U14092 ( .A1(n12288), .A2(n14712), .ZN(n12289) );
  NAND4_X1 U14093 ( .A1(n14394), .A2(n12287), .A3(n13730), .A4(n12289), .ZN(
        n12290) );
  AND2_X2 U14094 ( .A1(n12388), .A2(n12380), .ZN(n12373) );
  INV_X1 U14095 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21649) );
  NAND2_X1 U14096 ( .A1(n12373), .A2(n21649), .ZN(n12295) );
  INV_X1 U14097 ( .A(n14735), .ZN(n12291) );
  INV_X1 U14098 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21632) );
  NAND2_X1 U14099 ( .A1(n12381), .A2(n21632), .ZN(n12293) );
  NAND2_X1 U14100 ( .A1(n12380), .A2(n21649), .ZN(n12292) );
  NAND3_X1 U14101 ( .A1(n12293), .A2(n13764), .A3(n12292), .ZN(n12294) );
  NAND2_X1 U14102 ( .A1(n12295), .A2(n12294), .ZN(n12297) );
  NAND2_X1 U14103 ( .A1(n12381), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12296) );
  OAI21_X1 U14104 ( .B1(n12388), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12296), .ZN(
        n14521) );
  XNOR2_X1 U14105 ( .A(n12297), .B(n14521), .ZN(n21648) );
  NAND2_X1 U14106 ( .A1(n21648), .A2(n12380), .ZN(n14517) );
  NAND2_X1 U14107 ( .A1(n14517), .A2(n12297), .ZN(n14706) );
  INV_X1 U14108 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12298) );
  NAND2_X1 U14109 ( .A1(n12373), .A2(n12298), .ZN(n12302) );
  NAND2_X1 U14110 ( .A1(n12381), .A2(n21479), .ZN(n12300) );
  NAND2_X1 U14111 ( .A1(n12380), .A2(n12298), .ZN(n12299) );
  NAND3_X1 U14112 ( .A1(n12300), .A2(n13764), .A3(n12299), .ZN(n12301) );
  AND2_X1 U14113 ( .A1(n12302), .A2(n12301), .ZN(n14705) );
  MUX2_X1 U14114 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12304) );
  NAND2_X1 U14115 ( .A1(n14520), .A2(n21496), .ZN(n12303) );
  NAND2_X1 U14116 ( .A1(n12304), .A2(n12303), .ZN(n14728) );
  INV_X1 U14117 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21683) );
  NAND2_X1 U14118 ( .A1(n12373), .A2(n21683), .ZN(n12308) );
  NAND2_X1 U14119 ( .A1(n12381), .A2(n21492), .ZN(n12306) );
  NAND2_X1 U14120 ( .A1(n12380), .A2(n21683), .ZN(n12305) );
  NAND3_X1 U14121 ( .A1(n12306), .A2(n13764), .A3(n12305), .ZN(n12307) );
  NAND2_X1 U14122 ( .A1(n12308), .A2(n12307), .ZN(n14888) );
  MUX2_X1 U14123 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12309) );
  NAND2_X1 U14124 ( .A1(n11481), .A2(n12309), .ZN(n14913) );
  INV_X1 U14125 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21700) );
  NAND2_X1 U14126 ( .A1(n12373), .A2(n21700), .ZN(n12313) );
  NAND2_X1 U14127 ( .A1(n12381), .A2(n21521), .ZN(n12311) );
  NAND2_X1 U14128 ( .A1(n12380), .A2(n21700), .ZN(n12310) );
  NAND3_X1 U14129 ( .A1(n12311), .A2(n13764), .A3(n12310), .ZN(n12312) );
  AND2_X1 U14130 ( .A1(n12313), .A2(n12312), .ZN(n14919) );
  INV_X1 U14131 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21522) );
  INV_X1 U14132 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n15119) );
  NAND2_X1 U14133 ( .A1(n12380), .A2(n15119), .ZN(n12314) );
  OAI211_X1 U14134 ( .C1(n12388), .C2(n21522), .A(n12314), .B(n12381), .ZN(
        n12315) );
  OAI21_X1 U14135 ( .B1(n12378), .B2(P1_EBX_REG_7__SCAN_IN), .A(n12315), .ZN(
        n15115) );
  INV_X1 U14136 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21723) );
  NAND2_X1 U14137 ( .A1(n12373), .A2(n21723), .ZN(n12319) );
  NAND2_X1 U14138 ( .A1(n12381), .A2(n21523), .ZN(n12317) );
  NAND2_X1 U14139 ( .A1(n12380), .A2(n21723), .ZN(n12316) );
  NAND3_X1 U14140 ( .A1(n12317), .A2(n13764), .A3(n12316), .ZN(n12318) );
  NAND2_X1 U14141 ( .A1(n12319), .A2(n12318), .ZN(n15125) );
  INV_X1 U14142 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U14143 ( .A1(n12380), .A2(n12320), .ZN(n12321) );
  OAI211_X1 U14144 ( .C1(n12388), .C2(n12407), .A(n12321), .B(n12381), .ZN(
        n12322) );
  OAI21_X1 U14145 ( .B1(n12378), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12322), .ZN(
        n15134) );
  INV_X1 U14146 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15185) );
  NAND2_X1 U14147 ( .A1(n12373), .A2(n15185), .ZN(n12327) );
  NAND2_X1 U14148 ( .A1(n12381), .A2(n12323), .ZN(n12325) );
  NAND2_X1 U14149 ( .A1(n12380), .A2(n15185), .ZN(n12324) );
  NAND3_X1 U14150 ( .A1(n12325), .A2(n13764), .A3(n12324), .ZN(n12326) );
  NAND2_X1 U14151 ( .A1(n14520), .A2(n12191), .ZN(n12329) );
  MUX2_X1 U14152 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12328) );
  AND2_X1 U14153 ( .A1(n12329), .A2(n12328), .ZN(n15256) );
  INV_X1 U14154 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15337) );
  NAND2_X1 U14155 ( .A1(n12373), .A2(n15337), .ZN(n12333) );
  NAND2_X1 U14156 ( .A1(n12381), .A2(n21556), .ZN(n12331) );
  NAND2_X1 U14157 ( .A1(n12380), .A2(n15337), .ZN(n12330) );
  NAND3_X1 U14158 ( .A1(n12331), .A2(n13764), .A3(n12330), .ZN(n12332) );
  NAND2_X1 U14159 ( .A1(n12333), .A2(n12332), .ZN(n15331) );
  INV_X1 U14160 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n20135) );
  NAND2_X1 U14161 ( .A1(n12380), .A2(n20135), .ZN(n12334) );
  OAI211_X1 U14162 ( .C1(n12388), .C2(n12189), .A(n12334), .B(n12381), .ZN(
        n12335) );
  OAI21_X1 U14163 ( .B1(n12378), .B2(P1_EBX_REG_13__SCAN_IN), .A(n12335), .ZN(
        n15864) );
  NAND2_X1 U14164 ( .A1(n14520), .A2(n21597), .ZN(n12337) );
  MUX2_X1 U14165 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12336) );
  AND2_X1 U14166 ( .A1(n12337), .A2(n12336), .ZN(n15833) );
  OAI21_X1 U14167 ( .B1(n12388), .B2(n21464), .A(n12381), .ZN(n12339) );
  INV_X1 U14168 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15953) );
  NAND2_X1 U14169 ( .A1(n12380), .A2(n15953), .ZN(n12338) );
  NAND2_X1 U14170 ( .A1(n12339), .A2(n12338), .ZN(n12341) );
  NAND2_X1 U14171 ( .A1(n12373), .A2(n15953), .ZN(n12340) );
  NAND2_X1 U14172 ( .A1(n12341), .A2(n12340), .ZN(n15847) );
  NAND2_X1 U14173 ( .A1(n15833), .A2(n15847), .ZN(n12342) );
  INV_X1 U14174 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21754) );
  NAND2_X1 U14175 ( .A1(n12373), .A2(n21754), .ZN(n12347) );
  INV_X1 U14176 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12343) );
  NAND2_X1 U14177 ( .A1(n12381), .A2(n12343), .ZN(n12345) );
  NAND2_X1 U14178 ( .A1(n12380), .A2(n21754), .ZN(n12344) );
  NAND3_X1 U14179 ( .A1(n12345), .A2(n13764), .A3(n12344), .ZN(n12346) );
  NAND2_X1 U14180 ( .A1(n12347), .A2(n12346), .ZN(n15943) );
  MUX2_X1 U14181 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12348) );
  INV_X1 U14182 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15938) );
  NAND2_X1 U14183 ( .A1(n12373), .A2(n15938), .ZN(n12353) );
  NAND2_X1 U14184 ( .A1(n12381), .A2(n12349), .ZN(n12351) );
  NAND2_X1 U14185 ( .A1(n12380), .A2(n15938), .ZN(n12350) );
  NAND3_X1 U14186 ( .A1(n12351), .A2(n13764), .A3(n12350), .ZN(n12352) );
  AND2_X1 U14187 ( .A1(n12353), .A2(n12352), .ZN(n15934) );
  MUX2_X1 U14188 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12354) );
  NAND2_X1 U14189 ( .A1(n11482), .A2(n12354), .ZN(n15931) );
  INV_X1 U14190 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15925) );
  NAND2_X1 U14191 ( .A1(n12373), .A2(n15925), .ZN(n12359) );
  NAND2_X1 U14192 ( .A1(n12381), .A2(n12355), .ZN(n12357) );
  NAND2_X1 U14193 ( .A1(n12380), .A2(n15925), .ZN(n12356) );
  NAND3_X1 U14194 ( .A1(n12357), .A2(n13764), .A3(n12356), .ZN(n12358) );
  NAND2_X1 U14195 ( .A1(n12359), .A2(n12358), .ZN(n15922) );
  INV_X1 U14196 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21629) );
  NAND2_X1 U14197 ( .A1(n14520), .A2(n21629), .ZN(n12361) );
  MUX2_X1 U14198 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12360) );
  AND2_X1 U14199 ( .A1(n12361), .A2(n12360), .ZN(n15918) );
  INV_X1 U14200 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15913) );
  NAND2_X1 U14201 ( .A1(n12373), .A2(n15913), .ZN(n12365) );
  INV_X1 U14202 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16098) );
  NAND2_X1 U14203 ( .A1(n12381), .A2(n16098), .ZN(n12363) );
  NAND2_X1 U14204 ( .A1(n12380), .A2(n15913), .ZN(n12362) );
  NAND3_X1 U14205 ( .A1(n12363), .A2(n13764), .A3(n12362), .ZN(n12364) );
  AND2_X1 U14206 ( .A1(n12365), .A2(n12364), .ZN(n15910) );
  MUX2_X1 U14207 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12367) );
  NAND2_X1 U14208 ( .A1(n14520), .A2(n16223), .ZN(n12366) );
  NAND2_X1 U14209 ( .A1(n12367), .A2(n12366), .ZN(n15801) );
  INV_X1 U14210 ( .A(n12373), .ZN(n12383) );
  OAI21_X1 U14211 ( .B1(n12388), .B2(n16228), .A(n12381), .ZN(n12369) );
  INV_X1 U14212 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15791) );
  NAND2_X1 U14213 ( .A1(n12380), .A2(n15791), .ZN(n12368) );
  NAND2_X1 U14214 ( .A1(n12369), .A2(n12368), .ZN(n12370) );
  OAI21_X1 U14215 ( .B1(n12383), .B2(P1_EBX_REG_24__SCAN_IN), .A(n12370), .ZN(
        n15789) );
  MUX2_X1 U14216 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12372) );
  NAND2_X1 U14217 ( .A1(n14520), .A2(n16073), .ZN(n12371) );
  NAND2_X1 U14218 ( .A1(n12372), .A2(n12371), .ZN(n15771) );
  INV_X1 U14219 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15902) );
  NAND2_X1 U14220 ( .A1(n12373), .A2(n15902), .ZN(n12377) );
  INV_X1 U14221 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U14222 ( .A1(n12381), .A2(n12412), .ZN(n12375) );
  NAND2_X1 U14223 ( .A1(n12380), .A2(n15902), .ZN(n12374) );
  NAND3_X1 U14224 ( .A1(n12375), .A2(n13764), .A3(n12374), .ZN(n12376) );
  AND2_X1 U14225 ( .A1(n12377), .A2(n12376), .ZN(n15758) );
  MUX2_X1 U14226 ( .A(n12378), .B(n13764), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12379) );
  OAI21_X1 U14227 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13766), .A(
        n12379), .ZN(n15747) );
  OAI21_X1 U14228 ( .B1(n14512), .B2(P1_EBX_REG_28__SCAN_IN), .A(n13764), .ZN(
        n12385) );
  INV_X1 U14229 ( .A(n12381), .ZN(n12382) );
  NOR2_X1 U14230 ( .A1(n12382), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12384) );
  OAI22_X1 U14231 ( .A1(n12385), .A2(n12384), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n12383), .ZN(n15736) );
  NOR2_X1 U14232 ( .A1(n14512), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12386) );
  INV_X1 U14233 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13792) );
  AOI21_X1 U14234 ( .B1(n14520), .B2(n13792), .A(n12386), .ZN(n12387) );
  MUX2_X1 U14235 ( .A(n12386), .B(n12387), .S(n13764), .Z(n15723) );
  NAND2_X1 U14236 ( .A1(n15734), .A2(n15723), .ZN(n15722) );
  AOI22_X1 U14237 ( .A1(n15722), .A2(n12388), .B1(n12387), .B2(n15734), .ZN(
        n12389) );
  OAI22_X1 U14238 ( .A1(n13766), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n14512), .ZN(n13765) );
  INV_X1 U14239 ( .A(n15718), .ZN(n12393) );
  NAND2_X1 U14240 ( .A1(n17146), .A2(n17144), .ZN(n12390) );
  OAI21_X1 U14241 ( .B1(n12391), .B2(n14712), .A(n12390), .ZN(n12392) );
  NAND2_X1 U14242 ( .A1(n12393), .A2(n21625), .ZN(n12425) );
  OR2_X1 U14243 ( .A1(n12394), .A2(n14741), .ZN(n12401) );
  INV_X1 U14244 ( .A(n12395), .ZN(n12397) );
  NAND2_X1 U14245 ( .A1(n12397), .A2(n12396), .ZN(n12400) );
  NAND2_X1 U14246 ( .A1(n13766), .A2(n12398), .ZN(n12399) );
  NAND4_X1 U14247 ( .A1(n12402), .A2(n12401), .A3(n12400), .A4(n12399), .ZN(
        n12404) );
  NOR2_X1 U14248 ( .A1(n12404), .A2(n12403), .ZN(n14539) );
  NAND2_X1 U14249 ( .A1(n14539), .A2(n12405), .ZN(n12406) );
  NAND2_X1 U14250 ( .A1(n12415), .A2(n12406), .ZN(n16268) );
  INV_X1 U14251 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21472) );
  NAND2_X1 U14252 ( .A1(n21472), .A2(n21608), .ZN(n21631) );
  NOR3_X1 U14253 ( .A1(n21523), .A2(n21522), .A3(n21521), .ZN(n21533) );
  INV_X1 U14254 ( .A(n21533), .ZN(n21536) );
  NOR2_X1 U14255 ( .A1(n12407), .A2(n21536), .ZN(n21540) );
  NAND2_X1 U14256 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n21540), .ZN(
        n21463) );
  NOR2_X1 U14257 ( .A1(n21479), .A2(n21632), .ZN(n21484) );
  NOR2_X1 U14258 ( .A1(n21492), .A2(n21496), .ZN(n21486) );
  NAND2_X1 U14259 ( .A1(n21484), .A2(n21486), .ZN(n21461) );
  NOR3_X1 U14260 ( .A1(n21462), .A2(n21463), .A3(n21461), .ZN(n16261) );
  INV_X1 U14261 ( .A(n16261), .ZN(n21550) );
  NOR3_X1 U14262 ( .A1(n12191), .A2(n21556), .A3(n21550), .ZN(n16264) );
  NOR2_X1 U14263 ( .A1(n21464), .A2(n12189), .ZN(n16252) );
  AND3_X1 U14264 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21585), .A3(
        n16252), .ZN(n16245) );
  NAND2_X1 U14265 ( .A1(n16264), .A2(n16245), .ZN(n21616) );
  NOR2_X1 U14266 ( .A1(n16098), .A2(n16247), .ZN(n12409) );
  INV_X1 U14267 ( .A(n12409), .ZN(n12408) );
  NOR2_X1 U14268 ( .A1(n21616), .A2(n12408), .ZN(n12420) );
  NAND2_X1 U14269 ( .A1(n21573), .A2(n12420), .ZN(n12411) );
  NAND2_X1 U14270 ( .A1(n14533), .A2(n12380), .ZN(n14511) );
  INV_X1 U14271 ( .A(n14511), .ZN(n14397) );
  NOR2_X1 U14272 ( .A1(n12191), .A2(n21463), .ZN(n21560) );
  OAI21_X1 U14273 ( .B1(n21472), .B2(n21632), .A(n21479), .ZN(n21485) );
  NAND2_X1 U14274 ( .A1(n21486), .A2(n21485), .ZN(n21509) );
  NOR2_X1 U14275 ( .A1(n21462), .A2(n21509), .ZN(n21500) );
  NAND2_X1 U14276 ( .A1(n21560), .A2(n21500), .ZN(n21552) );
  NOR2_X1 U14277 ( .A1(n21556), .A2(n21552), .ZN(n16273) );
  NAND3_X1 U14278 ( .A1(n16245), .A2(n12409), .A3(n16273), .ZN(n12418) );
  OR2_X1 U14279 ( .A1(n21501), .A2(n12418), .ZN(n12410) );
  NAND2_X1 U14280 ( .A1(n12411), .A2(n12410), .ZN(n16225) );
  NOR2_X1 U14281 ( .A1(n16204), .A2(n12412), .ZN(n12413) );
  NAND2_X1 U14282 ( .A1(n16225), .A2(n12413), .ZN(n16194) );
  NOR2_X1 U14283 ( .A1(n16194), .A2(n12414), .ZN(n16165) );
  INV_X1 U14284 ( .A(n21551), .ZN(n21503) );
  OR2_X1 U14285 ( .A1(n16268), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12417) );
  INV_X1 U14286 ( .A(n12415), .ZN(n12416) );
  NAND2_X1 U14287 ( .A1(n12416), .A2(n21596), .ZN(n16266) );
  OAI21_X1 U14288 ( .B1(n16223), .B2(n12418), .A(n21575), .ZN(n12419) );
  OAI211_X1 U14289 ( .C1(n21503), .C2(n12420), .A(n21554), .B(n12419), .ZN(
        n16235) );
  AOI21_X1 U14290 ( .B1(n16204), .B2(n21633), .A(n16235), .ZN(n16216) );
  NAND2_X1 U14291 ( .A1(n16216), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12421) );
  NAND2_X1 U14292 ( .A1(n21534), .A2(n21554), .ZN(n21515) );
  NAND2_X1 U14293 ( .A1(n12421), .A2(n21515), .ZN(n16199) );
  NAND2_X1 U14294 ( .A1(n21633), .A2(n13792), .ZN(n12422) );
  NAND3_X1 U14295 ( .A1(n16199), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12422), .ZN(n16162) );
  INV_X1 U14296 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n17357) );
  NOR2_X1 U14297 ( .A1(n21596), .A2(n17357), .ZN(n16026) );
  OAI21_X1 U14298 ( .B1(n12421), .B2(n16174), .A(n21515), .ZN(n16173) );
  INV_X1 U14299 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13798) );
  AOI21_X1 U14300 ( .B1(n16173), .B2(n12422), .A(n13798), .ZN(n12423) );
  AOI211_X1 U14301 ( .C1(n16165), .C2(n16162), .A(n16026), .B(n12423), .ZN(
        n12424) );
  OAI21_X1 U14302 ( .B1(n16032), .B2(n21635), .A(n12426), .ZN(P1_U3001) );
  INV_X4 U14303 ( .A(n12441), .ZN(n15588) );
  AND2_X2 U14304 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14454) );
  INV_X2 U14305 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14619) );
  INV_X2 U14306 ( .A(n15687), .ZN(n12618) );
  AOI22_X1 U14307 ( .A1(n15588), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12618), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12432) );
  AND2_X2 U14308 ( .A1(n12427), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12446) );
  AND2_X4 U14309 ( .A1(n12446), .A2(n11409), .ZN(n12667) );
  INV_X1 U14310 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U14311 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12431) );
  NAND2_X2 U14312 ( .A1(n14604), .A2(n14619), .ZN(n15543) );
  INV_X4 U14313 ( .A(n15543), .ZN(n15566) );
  AND2_X4 U14314 ( .A1(n14613), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15676) );
  AOI22_X1 U14315 ( .A1(n15566), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15676), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U14316 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12429) );
  NAND4_X1 U14317 ( .A1(n12432), .A2(n12431), .A3(n12430), .A4(n12429), .ZN(
        n12433) );
  NAND2_X1 U14318 ( .A1(n12433), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12440) );
  AOI22_X1 U14319 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U14320 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U14321 ( .A1(n15566), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12435) );
  INV_X2 U14322 ( .A(n15687), .ZN(n12657) );
  AOI22_X1 U14323 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12434) );
  NAND4_X1 U14324 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n12434), .ZN(
        n12438) );
  NAND2_X1 U14325 ( .A1(n12438), .A2(n12648), .ZN(n12439) );
  NAND2_X2 U14326 ( .A1(n12439), .A2(n12440), .ZN(n12628) );
  NAND2_X1 U14327 ( .A1(n11028), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13852) );
  AND2_X2 U14328 ( .A1(n15683), .A2(n12648), .ZN(n12793) );
  AOI22_X1 U14329 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15512), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12445) );
  OR2_X1 U14330 ( .A1(n12441), .A2(n12648), .ZN(n14078) );
  NAND3_X1 U14331 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13033) );
  NOR2_X1 U14332 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n13033), .ZN(
        n12803) );
  AOI22_X1 U14333 ( .A1(n15508), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n15513), .ZN(n12444) );
  AND2_X2 U14334 ( .A1(n12618), .A2(n12648), .ZN(n12802) );
  AOI22_X1 U14335 ( .A1(n15510), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12443) );
  AND2_X2 U14336 ( .A1(n15676), .A2(n12648), .ZN(n15499) );
  AOI22_X1 U14337 ( .A1(n15504), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15499), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12442) );
  NAND4_X1 U14338 ( .A1(n12445), .A2(n12444), .A3(n12443), .A4(n12442), .ZN(
        n12454) );
  AOI22_X1 U14339 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12479), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U14340 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n15498), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12451) );
  AND2_X2 U14341 ( .A1(n12667), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14086) );
  AOI22_X1 U14342 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n14086), .B1(
        n15511), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12450) );
  INV_X2 U14343 ( .A(n15650), .ZN(n15681) );
  AND2_X2 U14344 ( .A1(n15681), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12500) );
  AOI22_X1 U14345 ( .A1(n15509), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12449) );
  NAND4_X1 U14346 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        n12453) );
  NOR2_X1 U14347 ( .A1(n12454), .A2(n12453), .ZN(n13952) );
  OR2_X1 U14348 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(
        n12455) );
  MUX2_X1 U14349 ( .A(n13952), .B(n12455), .S(n11028), .Z(n12876) );
  AOI22_X1 U14350 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12457) );
  INV_X2 U14351 ( .A(n15650), .ZN(n12668) );
  AOI22_X1 U14352 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U14353 ( .A1(n15566), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U14354 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U14355 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U14356 ( .A1(n15566), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U14357 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12461) );
  AOI22_X1 U14358 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U14359 ( .A1(n15566), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U14360 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U14361 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12464) );
  NAND4_X1 U14362 ( .A1(n12467), .A2(n12466), .A3(n12465), .A4(n12464), .ZN(
        n12473) );
  AOI22_X1 U14363 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U14364 ( .A1(n15566), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U14365 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U14366 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12468) );
  NAND4_X1 U14367 ( .A1(n12471), .A2(n12470), .A3(n12469), .A4(n12468), .ZN(
        n12472) );
  XNOR2_X1 U14368 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13028) );
  NAND2_X1 U14369 ( .A1(n13028), .A2(n12871), .ZN(n12475) );
  NAND2_X1 U14370 ( .A1(n19488), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12474) );
  NAND2_X1 U14371 ( .A1(n12475), .A2(n12474), .ZN(n12517) );
  XNOR2_X1 U14372 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12516) );
  INV_X1 U14373 ( .A(n12516), .ZN(n12476) );
  XNOR2_X1 U14374 ( .A(n12517), .B(n12476), .ZN(n13863) );
  AND2_X1 U14375 ( .A1(n13861), .A2(n13863), .ZN(n13875) );
  INV_X1 U14376 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14029) );
  NAND2_X1 U14377 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12478) );
  NAND2_X1 U14378 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12477) );
  OAI211_X1 U14379 ( .C1(n14029), .C2(n15484), .A(n12478), .B(n12477), .ZN(
        n12485) );
  NAND2_X1 U14380 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12483) );
  AOI22_X1 U14381 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U14382 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12481) );
  NAND2_X1 U14383 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12480) );
  NAND4_X1 U14384 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n12480), .ZN(
        n12484) );
  NOR2_X1 U14385 ( .A1(n12485), .A2(n12484), .ZN(n12495) );
  INV_X1 U14386 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12486) );
  INV_X1 U14387 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14031) );
  OAI22_X1 U14388 ( .A1(n14082), .A2(n12486), .B1(n14078), .B2(n14031), .ZN(
        n12488) );
  INV_X1 U14389 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15574) );
  INV_X1 U14390 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19808) );
  OAI22_X1 U14391 ( .A1(n14057), .A2(n15574), .B1(n14081), .B2(n19808), .ZN(
        n12487) );
  OR2_X1 U14392 ( .A1(n12488), .A2(n12487), .ZN(n12493) );
  INV_X1 U14393 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12491) );
  NAND2_X1 U14394 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12490) );
  NAND2_X1 U14395 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12489) );
  OAI211_X1 U14396 ( .C1(n12491), .C2(n14462), .A(n12490), .B(n12489), .ZN(
        n12492) );
  NOR2_X1 U14397 ( .A1(n12493), .A2(n12492), .ZN(n12494) );
  NOR2_X1 U14398 ( .A1(n13861), .A2(n13962), .ZN(n12496) );
  NOR2_X1 U14399 ( .A1(n13875), .A2(n12496), .ZN(n13019) );
  INV_X1 U14400 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12497) );
  INV_X1 U14401 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14056) );
  OAI22_X1 U14402 ( .A1(n14082), .A2(n12497), .B1(n14078), .B2(n14056), .ZN(
        n12499) );
  INV_X1 U14403 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15597) );
  INV_X1 U14404 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19761) );
  OAI22_X1 U14405 ( .A1(n14057), .A2(n15597), .B1(n14081), .B2(n19761), .ZN(
        n12498) );
  NOR2_X1 U14406 ( .A1(n12499), .A2(n12498), .ZN(n12515) );
  INV_X1 U14407 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14055) );
  NAND2_X1 U14408 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12502) );
  NAND2_X1 U14409 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12501) );
  OAI211_X1 U14410 ( .C1(n14055), .C2(n15484), .A(n12502), .B(n12501), .ZN(
        n12503) );
  INV_X1 U14411 ( .A(n12503), .ZN(n12514) );
  NAND2_X1 U14412 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12507) );
  AOI22_X1 U14413 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U14414 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12505) );
  NAND2_X1 U14415 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12504) );
  AND4_X1 U14416 ( .A1(n12507), .A2(n12506), .A3(n12505), .A4(n12504), .ZN(
        n12513) );
  INV_X1 U14417 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12510) );
  NAND2_X1 U14418 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12509) );
  NAND2_X1 U14419 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12508) );
  OAI211_X1 U14420 ( .C1(n12510), .C2(n14462), .A(n12509), .B(n12508), .ZN(
        n12511) );
  INV_X1 U14421 ( .A(n12511), .ZN(n12512) );
  NAND4_X1 U14422 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n13969) );
  NAND2_X1 U14423 ( .A1(n12517), .A2(n12516), .ZN(n12519) );
  NAND2_X1 U14424 ( .A1(n17490), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12518) );
  NAND2_X1 U14425 ( .A1(n12519), .A2(n12518), .ZN(n12543) );
  XNOR2_X1 U14426 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12542) );
  INV_X1 U14427 ( .A(n12542), .ZN(n12520) );
  XNOR2_X1 U14428 ( .A(n12543), .B(n12520), .ZN(n13876) );
  MUX2_X1 U14429 ( .A(n13969), .B(n13876), .S(n13861), .Z(n13018) );
  INV_X1 U14430 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12521) );
  MUX2_X1 U14431 ( .A(n13018), .B(n12521), .S(n11028), .Z(n12867) );
  INV_X1 U14432 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12523) );
  INV_X1 U14433 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12522) );
  OAI22_X1 U14434 ( .A1(n12523), .A2(n14082), .B1(n14078), .B2(n12522), .ZN(
        n12525) );
  INV_X1 U14435 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15618) );
  INV_X1 U14436 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19711) );
  OAI22_X1 U14437 ( .A1(n15618), .A2(n14057), .B1(n14081), .B2(n19711), .ZN(
        n12524) );
  NOR2_X1 U14438 ( .A1(n12525), .A2(n12524), .ZN(n12541) );
  INV_X1 U14439 ( .A(n12793), .ZN(n14017) );
  INV_X1 U14440 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14080) );
  NAND2_X1 U14441 ( .A1(n15504), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12527) );
  NAND2_X1 U14442 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12526) );
  OAI211_X1 U14443 ( .C1(n14017), .C2(n14080), .A(n12527), .B(n12526), .ZN(
        n12528) );
  INV_X1 U14444 ( .A(n12528), .ZN(n12540) );
  NAND2_X1 U14445 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12532) );
  AOI22_X1 U14446 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12479), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U14447 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n15498), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12530) );
  NAND2_X1 U14448 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12529) );
  INV_X1 U14449 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12535) );
  NAND2_X1 U14450 ( .A1(n15512), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12534) );
  NAND2_X1 U14451 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12533) );
  OAI211_X1 U14452 ( .C1(n12536), .C2(n12535), .A(n12534), .B(n12533), .ZN(
        n12537) );
  INV_X1 U14453 ( .A(n12537), .ZN(n12538) );
  NAND4_X1 U14454 ( .A1(n12541), .A2(n12540), .A3(n12539), .A4(n12538), .ZN(
        n12828) );
  NAND2_X1 U14455 ( .A1(n12543), .A2(n12542), .ZN(n12545) );
  NAND2_X1 U14456 ( .A1(n19432), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12544) );
  NAND2_X1 U14457 ( .A1(n12545), .A2(n12544), .ZN(n13022) );
  NAND2_X1 U14458 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14656), .ZN(
        n13023) );
  MUX2_X1 U14459 ( .A(n12828), .B(n13880), .S(n13861), .Z(n13017) );
  INV_X1 U14460 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n15434) );
  MUX2_X1 U14461 ( .A(n13017), .B(n15434), .S(n11028), .Z(n12546) );
  INV_X1 U14462 ( .A(n12546), .ZN(n12878) );
  INV_X1 U14463 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12549) );
  NAND2_X1 U14464 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12548) );
  NAND2_X1 U14465 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12547) );
  OAI211_X1 U14466 ( .C1(n12549), .C2(n15484), .A(n12548), .B(n12547), .ZN(
        n12555) );
  NAND2_X1 U14467 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12553) );
  AOI22_X1 U14468 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U14469 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12551) );
  NAND2_X1 U14470 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12550) );
  NAND4_X1 U14471 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12554) );
  NOR2_X1 U14472 ( .A1(n12555), .A2(n12554), .ZN(n12564) );
  INV_X1 U14473 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12556) );
  INV_X1 U14474 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15640) );
  OAI22_X1 U14475 ( .A1(n14082), .A2(n12556), .B1(n14078), .B2(n15640), .ZN(
        n12558) );
  INV_X1 U14476 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12846) );
  INV_X1 U14477 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15469) );
  OAI22_X1 U14478 ( .A1(n14057), .A2(n12846), .B1(n14081), .B2(n15469), .ZN(
        n12557) );
  OR2_X1 U14479 ( .A1(n12558), .A2(n12557), .ZN(n12562) );
  INV_X1 U14480 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U14481 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12560) );
  NAND2_X1 U14482 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12559) );
  OAI211_X1 U14483 ( .C1(n12832), .C2(n14462), .A(n12560), .B(n12559), .ZN(
        n12561) );
  NOR2_X1 U14484 ( .A1(n12562), .A2(n12561), .ZN(n12563) );
  MUX2_X1 U14485 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n13976), .S(n14857), .Z(
        n12863) );
  NOR2_X2 U14486 ( .A1(n12881), .A2(n12863), .ZN(n12911) );
  INV_X1 U14487 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18506) );
  INV_X1 U14488 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12565) );
  INV_X1 U14489 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12897) );
  OAI22_X1 U14490 ( .A1(n12565), .A2(n14082), .B1(n14078), .B2(n12897), .ZN(
        n12567) );
  INV_X1 U14491 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12890) );
  INV_X1 U14492 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19605) );
  OAI22_X1 U14493 ( .A1(n12890), .A2(n14057), .B1(n14081), .B2(n19605), .ZN(
        n12566) );
  NOR2_X1 U14494 ( .A1(n12567), .A2(n12566), .ZN(n12582) );
  INV_X1 U14495 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12570) );
  NAND2_X1 U14496 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12569) );
  NAND2_X1 U14497 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12568) );
  OAI211_X1 U14498 ( .C1(n15484), .C2(n12570), .A(n12569), .B(n12568), .ZN(
        n12571) );
  INV_X1 U14499 ( .A(n12571), .ZN(n12581) );
  NAND2_X1 U14500 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12575) );
  AOI22_X1 U14501 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12479), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U14502 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n15498), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12573) );
  NAND2_X1 U14503 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12572) );
  AND4_X1 U14504 ( .A1(n12575), .A2(n12574), .A3(n12573), .A4(n12572), .ZN(
        n12580) );
  INV_X1 U14505 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12899) );
  NAND2_X1 U14506 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12577) );
  NAND2_X1 U14507 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12576) );
  OAI211_X1 U14508 ( .C1(n14462), .C2(n12899), .A(n12577), .B(n12576), .ZN(
        n12578) );
  INV_X1 U14509 ( .A(n12578), .ZN(n12579) );
  NAND4_X1 U14510 ( .A1(n12582), .A2(n12581), .A3(n12580), .A4(n12579), .ZN(
        n12907) );
  MUX2_X1 U14511 ( .A(n18506), .B(n12907), .S(n14857), .Z(n12910) );
  INV_X1 U14512 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U14513 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12584) );
  NAND2_X1 U14514 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12583) );
  OAI211_X1 U14515 ( .C1(n15484), .C2(n12585), .A(n12584), .B(n12583), .ZN(
        n12591) );
  NAND2_X1 U14516 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12589) );
  AOI22_X1 U14517 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U14518 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12587) );
  NAND2_X1 U14519 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12586) );
  NAND4_X1 U14520 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n12586), .ZN(
        n12590) );
  NOR2_X1 U14521 ( .A1(n12591), .A2(n12590), .ZN(n12602) );
  INV_X1 U14522 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12592) );
  INV_X1 U14523 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15686) );
  OAI22_X1 U14524 ( .A1(n12592), .A2(n14082), .B1(n14078), .B2(n15686), .ZN(
        n12595) );
  INV_X1 U14525 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12593) );
  INV_X1 U14526 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15181) );
  OAI22_X1 U14527 ( .A1(n14057), .A2(n12593), .B1(n14081), .B2(n15181), .ZN(
        n12594) );
  OR2_X1 U14528 ( .A1(n12595), .A2(n12594), .ZN(n12600) );
  INV_X1 U14529 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12598) );
  NAND2_X1 U14530 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12597) );
  NAND2_X1 U14531 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12596) );
  OAI211_X1 U14532 ( .C1(n14462), .C2(n12598), .A(n12597), .B(n12596), .ZN(
        n12599) );
  NOR2_X1 U14533 ( .A1(n12600), .A2(n12599), .ZN(n12601) );
  MUX2_X1 U14534 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n16730), .S(n14857), .Z(
        n12918) );
  INV_X1 U14535 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12603) );
  NOR2_X1 U14536 ( .A1(n14857), .A2(n12603), .ZN(n12915) );
  NAND2_X1 U14537 ( .A1(n11028), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12922) );
  NAND2_X1 U14538 ( .A1(n12924), .A2(n12922), .ZN(n12926) );
  INV_X1 U14539 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12604) );
  NOR2_X1 U14540 ( .A1(n14857), .A2(n12604), .ZN(n12925) );
  INV_X1 U14541 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12605) );
  NOR2_X1 U14542 ( .A1(n14857), .A2(n12605), .ZN(n12933) );
  NAND2_X1 U14543 ( .A1(n11028), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12951) );
  NAND2_X1 U14544 ( .A1(n11028), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12948) );
  INV_X1 U14545 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n18605) );
  NOR2_X1 U14546 ( .A1(n14857), .A2(n18605), .ZN(n12961) );
  INV_X1 U14547 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12606) );
  NOR2_X1 U14548 ( .A1(n14857), .A2(n12606), .ZN(n12943) );
  INV_X1 U14549 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12607) );
  NOR2_X1 U14550 ( .A1(n14857), .A2(n12607), .ZN(n12957) );
  NAND2_X1 U14551 ( .A1(n11028), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12936) );
  INV_X1 U14552 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12608) );
  NOR2_X1 U14553 ( .A1(n14857), .A2(n12608), .ZN(n12935) );
  INV_X1 U14554 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n12609) );
  NOR2_X1 U14555 ( .A1(n14857), .A2(n12609), .ZN(n12941) );
  INV_X1 U14556 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n18680) );
  NOR2_X1 U14557 ( .A1(n14857), .A2(n18680), .ZN(n12979) );
  INV_X1 U14558 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12610) );
  NOR2_X1 U14559 ( .A1(n14857), .A2(n12610), .ZN(n12984) );
  NAND2_X1 U14560 ( .A1(n11028), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12987) );
  NAND2_X1 U14561 ( .A1(n11028), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12998) );
  INV_X1 U14562 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n18730) );
  NOR2_X1 U14563 ( .A1(n14857), .A2(n18730), .ZN(n12993) );
  INV_X1 U14564 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12611) );
  NOR2_X1 U14565 ( .A1(n14857), .A2(n12611), .ZN(n13001) );
  NAND2_X1 U14566 ( .A1(n11028), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13006) );
  XOR2_X1 U14567 ( .A(n13852), .B(n13853), .Z(n18777) );
  AOI21_X1 U14568 ( .B1(n18777), .B2(n13859), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13850) );
  INV_X1 U14569 ( .A(n12628), .ZN(n12627) );
  AOI22_X1 U14570 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U14571 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U14572 ( .A1(n15566), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12614) );
  NAND4_X1 U14573 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n12626) );
  AOI22_X1 U14574 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U14575 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U14576 ( .A1(n15566), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12621) );
  NAND4_X1 U14577 ( .A1(n12624), .A2(n12623), .A3(n12622), .A4(n12621), .ZN(
        n12625) );
  NAND2_X1 U14578 ( .A1(n12626), .A2(n12625), .ZN(n12679) );
  INV_X1 U14579 ( .A(n12679), .ZN(n12686) );
  NAND2_X1 U14580 ( .A1(n12627), .A2(n12686), .ZN(n12690) );
  NAND2_X2 U14581 ( .A1(n12628), .A2(n12679), .ZN(n12688) );
  INV_X2 U14582 ( .A(n15543), .ZN(n15678) );
  AOI22_X1 U14583 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U14584 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U14585 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U14586 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12629) );
  NAND4_X1 U14587 ( .A1(n12632), .A2(n12631), .A3(n12630), .A4(n12629), .ZN(
        n12638) );
  AOI22_X1 U14588 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U14589 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U14590 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U14591 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12633) );
  NAND4_X1 U14592 ( .A1(n12636), .A2(n12635), .A3(n12634), .A4(n12633), .ZN(
        n12637) );
  AOI22_X1 U14593 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U14594 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U14595 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U14596 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12639) );
  NAND4_X1 U14597 ( .A1(n12642), .A2(n12641), .A3(n12640), .A4(n12639), .ZN(
        n12643) );
  NAND2_X1 U14598 ( .A1(n12643), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12651) );
  AOI22_X1 U14599 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U14600 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U14601 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12645) );
  AOI22_X1 U14602 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12644) );
  NAND4_X1 U14603 ( .A1(n12647), .A2(n12646), .A3(n12645), .A4(n12644), .ZN(
        n12649) );
  NAND2_X1 U14604 ( .A1(n12649), .A2(n12648), .ZN(n12650) );
  AOI22_X1 U14605 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U14606 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U14607 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U14608 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U14609 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U14610 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U14611 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U14612 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12658) );
  AOI22_X1 U14613 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U14614 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U14615 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12662) );
  NAND4_X1 U14616 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12666) );
  AOI22_X1 U14617 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15683), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U14618 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U14619 ( .A1(n15676), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12670) );
  AOI22_X1 U14620 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12669) );
  NAND4_X1 U14621 ( .A1(n12672), .A2(n12671), .A3(n12670), .A4(n12669), .ZN(
        n12673) );
  NAND2_X1 U14622 ( .A1(n12673), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12674) );
  NOR2_X1 U14623 ( .A1(n15031), .A2(n12700), .ZN(n12676) );
  INV_X4 U14624 ( .A(n15667), .ZN(n16334) );
  INV_X1 U14625 ( .A(n12682), .ZN(n12678) );
  NAND2_X1 U14626 ( .A1(n12678), .A2(n15667), .ZN(n13900) );
  NAND2_X1 U14627 ( .A1(n19562), .A2(n12873), .ZN(n12680) );
  NOR2_X1 U14628 ( .A1(n13900), .A2(n12680), .ZN(n12685) );
  INV_X1 U14629 ( .A(n14564), .ZN(n12681) );
  NOR2_X1 U14630 ( .A1(n12688), .A2(n12682), .ZN(n12683) );
  INV_X1 U14631 ( .A(n13897), .ZN(n14565) );
  AND2_X2 U14632 ( .A1(n19872), .A2(n15031), .ZN(n14199) );
  NAND2_X1 U14633 ( .A1(n12688), .A2(n14193), .ZN(n12698) );
  INV_X1 U14634 ( .A(n12690), .ZN(n12692) );
  NOR2_X1 U14635 ( .A1(n12687), .A2(n12699), .ZN(n12691) );
  NOR2_X1 U14636 ( .A1(n13897), .A2(n13861), .ZN(n12693) );
  AOI22_X1 U14637 ( .A1(n13047), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12694) );
  AND2_X1 U14638 ( .A1(n14197), .A2(n14468), .ZN(n12695) );
  NAND2_X2 U14639 ( .A1(n12710), .A2(n12695), .ZN(n13015) );
  NAND3_X1 U14640 ( .A1(n13015), .A2(n14197), .A3(n16334), .ZN(n12696) );
  NAND2_X1 U14641 ( .A1(n12697), .A2(n16277), .ZN(n12734) );
  NAND2_X1 U14642 ( .A1(n19562), .A2(n19671), .ZN(n12702) );
  NAND3_X1 U14643 ( .A1(n12703), .A2(n12702), .A3(n12701), .ZN(n12704) );
  NAND2_X1 U14644 ( .A1(n12704), .A2(n19872), .ZN(n12708) );
  NAND2_X1 U14645 ( .A1(n14199), .A2(n12706), .ZN(n12707) );
  NAND2_X1 U14646 ( .A1(n12708), .A2(n12707), .ZN(n14195) );
  NAND2_X1 U14647 ( .A1(n12688), .A2(n15667), .ZN(n12726) );
  INV_X1 U14648 ( .A(n14566), .ZN(n12727) );
  INV_X1 U14649 ( .A(n12710), .ZN(n12728) );
  OAI211_X1 U14650 ( .C1(n14193), .C2(n12727), .A(n12728), .B(n16287), .ZN(
        n12711) );
  NAND2_X1 U14651 ( .A1(n12730), .A2(n12711), .ZN(n12712) );
  NAND2_X1 U14652 ( .A1(n12712), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12713) );
  NAND2_X1 U14653 ( .A1(n14841), .A2(n18890), .ZN(n18882) );
  OAI211_X1 U14654 ( .C1(n18882), .C2(n19488), .A(n12715), .B(n12714), .ZN(
        n12716) );
  INV_X1 U14655 ( .A(n12716), .ZN(n12717) );
  NAND2_X1 U14656 ( .A1(n12719), .A2(n12718), .ZN(n12720) );
  AND3_X1 U14657 ( .A1(n14565), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n16287), 
        .ZN(n12721) );
  OAI22_X1 U14658 ( .A1(n12739), .A2(n12721), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13047), .ZN(n12725) );
  INV_X1 U14659 ( .A(n18882), .ZN(n13144) );
  NAND2_X1 U14660 ( .A1(n13144), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12722) );
  AND2_X1 U14661 ( .A1(n12723), .A2(n12722), .ZN(n12724) );
  NAND2_X1 U14662 ( .A1(n12725), .A2(n12724), .ZN(n12760) );
  NAND2_X1 U14663 ( .A1(n12753), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12737) );
  AND2_X1 U14664 ( .A1(n12727), .A2(n12726), .ZN(n14196) );
  OAI21_X1 U14665 ( .B1(n14196), .B2(n14193), .A(n12728), .ZN(n12729) );
  AOI21_X1 U14666 ( .B1(n12730), .B2(n12729), .A(n14841), .ZN(n12731) );
  AOI21_X1 U14667 ( .B1(n12752), .B2(P2_REIP_REG_0__SCAN_IN), .A(n12731), .ZN(
        n12736) );
  NAND2_X1 U14668 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12732) );
  NAND2_X1 U14669 ( .A1(n18882), .A2(n12732), .ZN(n12733) );
  AOI21_X1 U14670 ( .B1(n13047), .B2(P2_EBX_REG_0__SCAN_IN), .A(n12733), .ZN(
        n12735) );
  NAND4_X1 U14671 ( .A1(n12737), .A2(n12736), .A3(n12735), .A4(n12734), .ZN(
        n12759) );
  NAND2_X1 U14672 ( .A1(n12760), .A2(n12759), .ZN(n12764) );
  NAND2_X1 U14673 ( .A1(n12739), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12741) );
  AOI21_X1 U14674 ( .B1(n14841), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12740) );
  NAND2_X1 U14675 ( .A1(n12741), .A2(n12740), .ZN(n12747) );
  INV_X1 U14676 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n14336) );
  AOI22_X1 U14677 ( .A1(n13047), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12742) );
  OAI21_X1 U14678 ( .B1(n12743), .B2(n14336), .A(n12742), .ZN(n12744) );
  NAND2_X1 U14679 ( .A1(n12748), .A2(n12747), .ZN(n12749) );
  NOR2_X1 U14680 ( .A1(n18882), .A2(n19432), .ZN(n12751) );
  NAND2_X1 U14681 ( .A1(n12753), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12755) );
  AOI22_X1 U14682 ( .A1(n14180), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12754) );
  XNOR2_X2 U14683 ( .A(n12757), .B(n12756), .ZN(n14426) );
  INV_X1 U14684 ( .A(n12758), .ZN(n12761) );
  OR2_X1 U14685 ( .A1(n12760), .A2(n12759), .ZN(n12765) );
  NAND2_X1 U14686 ( .A1(n12761), .A2(n12765), .ZN(n12783) );
  INV_X1 U14687 ( .A(n12762), .ZN(n12774) );
  XNOR2_X2 U14688 ( .A(n12774), .B(n12763), .ZN(n18470) );
  AND2_X2 U14689 ( .A1(n12765), .A2(n11003), .ZN(n18452) );
  AOI22_X1 U14690 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12829), .B1(
        n12842), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12771) );
  INV_X1 U14691 ( .A(n18452), .ZN(n18805) );
  INV_X1 U14692 ( .A(n14426), .ZN(n14331) );
  INV_X1 U14693 ( .A(n12772), .ZN(n12766) );
  AOI22_X1 U14694 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12849), .B1(
        n19446), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12770) );
  INV_X1 U14695 ( .A(n12783), .ZN(n12780) );
  AOI22_X1 U14696 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19478), .B1(
        n12843), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U14697 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12830), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12768) );
  NAND4_X1 U14698 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n12768), .ZN(
        n12815) );
  NAND2_X1 U14699 ( .A1(n11484), .A2(n12766), .ZN(n12850) );
  INV_X1 U14700 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12773) );
  NAND2_X1 U14701 ( .A1(n18452), .A2(n12774), .ZN(n12784) );
  INV_X1 U14702 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12776) );
  NOR2_X1 U14703 ( .A1(n12835), .A2(n12776), .ZN(n12777) );
  NOR2_X1 U14704 ( .A1(n12778), .A2(n12777), .ZN(n12789) );
  AOI22_X1 U14705 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12831), .B1(
        n14985), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U14706 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n15170), .B1(
        n19462), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12787) );
  NOR2_X1 U14707 ( .A1(n12785), .A2(n12783), .ZN(n12840) );
  NOR2_X1 U14708 ( .A1(n12785), .A2(n12784), .ZN(n12834) );
  AOI22_X1 U14709 ( .A1(n12840), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12786) );
  NAND4_X1 U14710 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12814) );
  INV_X1 U14711 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12790) );
  INV_X1 U14712 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13988) );
  OAI22_X1 U14713 ( .A1(n14082), .A2(n12790), .B1(n14078), .B2(n13988), .ZN(
        n12792) );
  INV_X1 U14714 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15531) );
  INV_X1 U14715 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19983) );
  OAI22_X1 U14716 ( .A1(n14057), .A2(n15531), .B1(n14081), .B2(n19983), .ZN(
        n12791) );
  NOR2_X1 U14717 ( .A1(n12792), .A2(n12791), .ZN(n12811) );
  INV_X1 U14718 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12796) );
  NAND2_X1 U14719 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12795) );
  NAND2_X1 U14720 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12794) );
  OAI211_X1 U14721 ( .C1(n12796), .C2(n15484), .A(n12795), .B(n12794), .ZN(
        n12797) );
  INV_X1 U14722 ( .A(n12797), .ZN(n12810) );
  NAND2_X1 U14723 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12801) );
  AOI22_X1 U14724 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U14725 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U14726 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12798) );
  AND4_X1 U14727 ( .A1(n12801), .A2(n12800), .A3(n12799), .A4(n12798), .ZN(
        n12809) );
  INV_X1 U14728 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12806) );
  NAND2_X1 U14729 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12805) );
  NAND2_X1 U14730 ( .A1(n12803), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12804) );
  OAI211_X1 U14731 ( .C1(n12806), .C2(n14462), .A(n12805), .B(n12804), .ZN(
        n12807) );
  INV_X1 U14732 ( .A(n12807), .ZN(n12808) );
  NOR2_X1 U14733 ( .A1(n14307), .A2(n13952), .ZN(n12812) );
  NAND2_X1 U14734 ( .A1(n15667), .A2(n12812), .ZN(n13153) );
  NAND2_X1 U14735 ( .A1(n13153), .A2(n13962), .ZN(n12813) );
  AOI22_X1 U14736 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12830), .B1(
        n12843), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U14737 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12829), .B1(
        n19446), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12817) );
  NAND4_X1 U14738 ( .A1(n12819), .A2(n12818), .A3(n12817), .A4(n12816), .ZN(
        n12827) );
  AOI22_X1 U14739 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n15170), .B1(
        n12834), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U14740 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12849), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U14741 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12840), .B1(
        n14985), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12820) );
  NAND4_X1 U14742 ( .A1(n12823), .A2(n12822), .A3(n12821), .A4(n12820), .ZN(
        n12826) );
  INV_X1 U14743 ( .A(n13969), .ZN(n12824) );
  NAND2_X1 U14744 ( .A1(n12824), .A2(n15667), .ZN(n12825) );
  INV_X1 U14745 ( .A(n12828), .ZN(n13939) );
  AOI22_X1 U14746 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n12829), .B1(
        n12830), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U14747 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n15170), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12838) );
  INV_X1 U14748 ( .A(n19478), .ZN(n12898) );
  OAI22_X1 U14749 ( .A1(n12832), .A2(n12898), .B1(n19443), .B2(n15640), .ZN(
        n12833) );
  INV_X1 U14750 ( .A(n12833), .ZN(n12837) );
  AOI22_X1 U14751 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19534), .B1(
        n19417), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U14752 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14852), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U14753 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n12842), .B1(
        n12843), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12844) );
  NAND2_X1 U14754 ( .A1(n12845), .A2(n12844), .ZN(n12854) );
  INV_X1 U14755 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12847) );
  OAI22_X1 U14756 ( .A1(n12847), .A2(n14981), .B1(n19458), .B2(n12846), .ZN(
        n12848) );
  INV_X1 U14757 ( .A(n12848), .ZN(n12852) );
  AOI22_X1 U14758 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n17377), .B1(
        n19406), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12851) );
  NAND2_X1 U14759 ( .A1(n12852), .A2(n12851), .ZN(n12853) );
  NOR2_X1 U14760 ( .A1(n12854), .A2(n12853), .ZN(n12855) );
  NAND2_X1 U14761 ( .A1(n12856), .A2(n12855), .ZN(n12858) );
  NAND2_X1 U14762 ( .A1(n15667), .A2(n13976), .ZN(n12857) );
  INV_X1 U14763 ( .A(n12860), .ZN(n12859) );
  NAND2_X1 U14764 ( .A1(n13161), .A2(n12859), .ZN(n12862) );
  AND2_X1 U14765 ( .A1(n12881), .A2(n12863), .ZN(n12864) );
  OR2_X1 U14766 ( .A1(n12864), .A2(n12911), .ZN(n18497) );
  INV_X1 U14767 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15215) );
  XNOR2_X1 U14768 ( .A(n12866), .B(n12865), .ZN(n17392) );
  OR2_X1 U14769 ( .A1(n17392), .A2(n13859), .ZN(n12869) );
  OAI21_X1 U14770 ( .B1(n12868), .B2(n12867), .A(n12879), .ZN(n16363) );
  NAND2_X1 U14771 ( .A1(n12869), .A2(n16363), .ZN(n17390) );
  NAND3_X1 U14772 ( .A1(n11028), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n12870) );
  AND2_X1 U14773 ( .A1(n12876), .A2(n12870), .ZN(n18466) );
  INV_X1 U14774 ( .A(n12871), .ZN(n13027) );
  NAND2_X1 U14775 ( .A1(n14619), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12872) );
  AND2_X1 U14776 ( .A1(n13027), .A2(n12872), .ZN(n13865) );
  INV_X1 U14777 ( .A(n13865), .ZN(n13869) );
  MUX2_X1 U14778 ( .A(n14307), .B(n13869), .S(n13861), .Z(n13020) );
  INV_X1 U14779 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14411) );
  MUX2_X1 U14780 ( .A(n13020), .B(n14411), .S(n11028), .Z(n18453) );
  INV_X1 U14781 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17048) );
  NOR2_X1 U14782 ( .A1(n18453), .A2(n17048), .ZN(n14303) );
  NAND2_X1 U14783 ( .A1(n18466), .A2(n14303), .ZN(n12874) );
  XOR2_X1 U14784 ( .A(n18466), .B(n14303), .Z(n14270) );
  NAND2_X1 U14785 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14270), .ZN(
        n14269) );
  NAND2_X1 U14786 ( .A1(n12874), .A2(n14269), .ZN(n14330) );
  XNOR2_X1 U14787 ( .A(n12876), .B(n12875), .ZN(n16378) );
  XNOR2_X1 U14788 ( .A(n16378), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14329) );
  INV_X1 U14789 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13154) );
  NOR2_X1 U14790 ( .A1(n16378), .A2(n13154), .ZN(n12877) );
  AOI21_X1 U14791 ( .B1(n14330), .B2(n14329), .A(n12877), .ZN(n17391) );
  INV_X1 U14792 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18860) );
  NAND2_X1 U14793 ( .A1(n12879), .A2(n12878), .ZN(n12880) );
  NAND2_X1 U14794 ( .A1(n12881), .A2(n12880), .ZN(n18482) );
  INV_X1 U14795 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18844) );
  AND2_X1 U14796 ( .A1(n18482), .A2(n18844), .ZN(n12883) );
  AOI21_X1 U14797 ( .B1(n17391), .B2(n18860), .A(n12883), .ZN(n12882) );
  NAND2_X1 U14798 ( .A1(n17390), .A2(n12882), .ZN(n12887) );
  INV_X1 U14799 ( .A(n17391), .ZN(n17401) );
  INV_X1 U14800 ( .A(n12883), .ZN(n12884) );
  NAND3_X1 U14801 ( .A1(n17401), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n12884), .ZN(n12886) );
  OR2_X1 U14802 ( .A1(n18482), .A2(n18844), .ZN(n12885) );
  NAND2_X1 U14803 ( .A1(n12888), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12889) );
  AOI22_X1 U14804 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12830), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U14805 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12829), .B1(
        n12843), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U14806 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14852), .B1(
        n12841), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12894) );
  INV_X1 U14807 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12891) );
  OAI22_X1 U14808 ( .A1(n12891), .A2(n14981), .B1(n19458), .B2(n12890), .ZN(
        n12892) );
  INV_X1 U14809 ( .A(n12892), .ZN(n12893) );
  NAND4_X1 U14810 ( .A1(n12896), .A2(n12895), .A3(n12894), .A4(n12893), .ZN(
        n12906) );
  AOI22_X1 U14811 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12842), .B1(
        n15170), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12904) );
  AOI22_X1 U14812 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n17377), .B1(
        n19406), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U14813 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19534), .B1(
        n19417), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12902) );
  OAI22_X1 U14814 ( .A1(n12899), .A2(n12898), .B1(n19443), .B2(n12897), .ZN(
        n12900) );
  INV_X1 U14815 ( .A(n12900), .ZN(n12901) );
  NAND4_X1 U14816 ( .A1(n12904), .A2(n12903), .A3(n12902), .A4(n12901), .ZN(
        n12905) );
  INV_X1 U14817 ( .A(n12907), .ZN(n13977) );
  NAND2_X1 U14818 ( .A1(n13977), .A2(n15667), .ZN(n12908) );
  OR2_X1 U14819 ( .A1(n12911), .A2(n12910), .ZN(n12912) );
  NAND2_X1 U14820 ( .A1(n12920), .A2(n12912), .ZN(n18507) );
  INV_X1 U14821 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15249) );
  XNOR2_X1 U14822 ( .A(n12913), .B(n15249), .ZN(n15235) );
  NAND2_X1 U14823 ( .A1(n12913), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12914) );
  AND2_X1 U14824 ( .A1(n13858), .A2(n12915), .ZN(n12916) );
  OR2_X1 U14825 ( .A1(n12916), .A2(n11080), .ZN(n18528) );
  INV_X1 U14826 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14208) );
  OR2_X1 U14827 ( .A1(n16730), .A2(n14208), .ZN(n12917) );
  NOR2_X1 U14828 ( .A1(n18528), .A2(n12917), .ZN(n17426) );
  INV_X1 U14829 ( .A(n12918), .ZN(n12919) );
  XNOR2_X1 U14830 ( .A(n12920), .B(n12919), .ZN(n18520) );
  OAI21_X1 U14831 ( .B1(n18528), .B2(n16730), .A(n14208), .ZN(n17425) );
  OR2_X1 U14832 ( .A1(n18520), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15300) );
  AND2_X1 U14833 ( .A1(n17425), .A2(n15300), .ZN(n12921) );
  XNOR2_X1 U14834 ( .A(n11080), .B(n11107), .ZN(n18542) );
  AOI21_X1 U14835 ( .B1(n18542), .B2(n13859), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17031) );
  INV_X1 U14836 ( .A(n12922), .ZN(n12923) );
  XNOR2_X1 U14837 ( .A(n12924), .B(n12923), .ZN(n18550) );
  NAND2_X1 U14838 ( .A1(n18550), .A2(n13859), .ZN(n12930) );
  INV_X1 U14839 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18814) );
  NAND2_X1 U14840 ( .A1(n12930), .A2(n18814), .ZN(n17445) );
  NAND2_X1 U14841 ( .A1(n12926), .A2(n12925), .ZN(n12927) );
  NAND2_X1 U14842 ( .A1(n12934), .A2(n12927), .ZN(n18564) );
  INV_X1 U14843 ( .A(n12928), .ZN(n12929) );
  NAND2_X1 U14844 ( .A1(n12929), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17010) );
  OR2_X1 U14845 ( .A1(n12930), .A2(n18814), .ZN(n17446) );
  INV_X1 U14846 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17020) );
  NOR2_X1 U14847 ( .A1(n16730), .A2(n17020), .ZN(n12931) );
  NAND2_X1 U14848 ( .A1(n18542), .A2(n12931), .ZN(n17029) );
  AND2_X1 U14849 ( .A1(n17446), .A2(n17029), .ZN(n17007) );
  XNOR2_X1 U14850 ( .A(n12934), .B(n11418), .ZN(n18576) );
  INV_X1 U14851 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17002) );
  NOR2_X1 U14852 ( .A1(n16995), .A2(n17002), .ZN(n12968) );
  XNOR2_X1 U14853 ( .A(n11073), .B(n11108), .ZN(n18665) );
  NAND2_X1 U14854 ( .A1(n18665), .A2(n13859), .ZN(n12969) );
  INV_X1 U14855 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16861) );
  NAND2_X1 U14856 ( .A1(n12969), .A2(n16861), .ZN(n16670) );
  XNOR2_X1 U14857 ( .A(n12938), .B(n11424), .ZN(n18645) );
  NAND2_X1 U14858 ( .A1(n18645), .A2(n13859), .ZN(n12970) );
  INV_X1 U14859 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16888) );
  NAND2_X1 U14860 ( .A1(n12970), .A2(n16888), .ZN(n16687) );
  OR2_X1 U14861 ( .A1(n12959), .A2(n12936), .ZN(n12937) );
  NAND2_X1 U14862 ( .A1(n12938), .A2(n12937), .ZN(n18633) );
  INV_X1 U14863 ( .A(n18633), .ZN(n12939) );
  NAND2_X1 U14864 ( .A1(n12939), .A2(n13859), .ZN(n16690) );
  INV_X1 U14865 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16907) );
  NAND2_X1 U14866 ( .A1(n16690), .A2(n16907), .ZN(n12940) );
  AND2_X1 U14867 ( .A1(n16687), .A2(n12940), .ZN(n16664) );
  INV_X1 U14868 ( .A(n12941), .ZN(n12942) );
  XNOR2_X1 U14869 ( .A(n11061), .B(n12942), .ZN(n18658) );
  NAND2_X1 U14870 ( .A1(n18658), .A2(n13859), .ZN(n16667) );
  INV_X1 U14871 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16883) );
  NAND2_X1 U14872 ( .A1(n11051), .A2(n12943), .ZN(n12944) );
  NAND2_X1 U14873 ( .A1(n12958), .A2(n12944), .ZN(n16353) );
  NOR2_X1 U14874 ( .A1(n16353), .A2(n16730), .ZN(n12945) );
  NAND2_X1 U14875 ( .A1(n12945), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16662) );
  INV_X1 U14876 ( .A(n12945), .ZN(n12946) );
  INV_X1 U14877 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16943) );
  NAND2_X1 U14878 ( .A1(n12946), .A2(n16943), .ZN(n12947) );
  OR2_X1 U14879 ( .A1(n12954), .A2(n12948), .ZN(n12949) );
  NAND2_X1 U14880 ( .A1(n11058), .A2(n12949), .ZN(n18598) );
  OR2_X1 U14881 ( .A1(n18598), .A2(n16730), .ZN(n12950) );
  INV_X1 U14882 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16957) );
  NAND2_X1 U14883 ( .A1(n12950), .A2(n16957), .ZN(n16728) );
  NOR2_X1 U14884 ( .A1(n12952), .A2(n12951), .ZN(n12953) );
  OR2_X1 U14885 ( .A1(n12954), .A2(n12953), .ZN(n18589) );
  INV_X1 U14886 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16990) );
  OAI21_X1 U14887 ( .B1(n18589), .B2(n16730), .A(n16990), .ZN(n16740) );
  OAI211_X1 U14888 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n12955), .A(
        n16728), .B(n16740), .ZN(n12956) );
  INV_X1 U14889 ( .A(n12956), .ZN(n12964) );
  AND2_X1 U14890 ( .A1(n12958), .A2(n12957), .ZN(n12960) );
  OR2_X1 U14891 ( .A1(n12960), .A2(n12959), .ZN(n12972) );
  INV_X1 U14892 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16922) );
  OAI21_X1 U14893 ( .B1(n12972), .B2(n16730), .A(n16922), .ZN(n16708) );
  NAND2_X1 U14894 ( .A1(n11058), .A2(n12961), .ZN(n12962) );
  NAND2_X1 U14895 ( .A1(n11051), .A2(n12962), .ZN(n18612) );
  OR2_X1 U14896 ( .A1(n18612), .A2(n16730), .ZN(n12963) );
  INV_X1 U14897 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16913) );
  NAND2_X1 U14898 ( .A1(n12963), .A2(n16913), .ZN(n16729) );
  NAND4_X1 U14899 ( .A1(n16715), .A2(n12964), .A3(n16708), .A4(n16729), .ZN(
        n12965) );
  AOI21_X1 U14900 ( .B1(n16667), .B2(n16883), .A(n12965), .ZN(n12966) );
  AND3_X1 U14901 ( .A1(n16670), .A2(n16664), .A3(n12966), .ZN(n12967) );
  OR2_X1 U14902 ( .A1(n12969), .A2(n16861), .ZN(n16671) );
  OR2_X1 U14903 ( .A1(n12970), .A2(n16888), .ZN(n16688) );
  INV_X1 U14904 ( .A(n16690), .ZN(n16700) );
  NAND2_X1 U14905 ( .A1(n16700), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12971) );
  AND2_X1 U14906 ( .A1(n16688), .A2(n12971), .ZN(n16666) );
  INV_X1 U14907 ( .A(n16667), .ZN(n16669) );
  INV_X1 U14908 ( .A(n12972), .ZN(n18626) );
  NOR2_X1 U14909 ( .A1(n16730), .A2(n16922), .ZN(n12973) );
  NAND2_X1 U14910 ( .A1(n18626), .A2(n12973), .ZN(n16707) );
  OR2_X1 U14911 ( .A1(n18612), .A2(n16913), .ZN(n16731) );
  INV_X1 U14912 ( .A(n18589), .ZN(n12974) );
  NAND2_X1 U14913 ( .A1(n12974), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16724) );
  OR2_X1 U14914 ( .A1(n18598), .A2(n16957), .ZN(n16726) );
  NAND3_X1 U14915 ( .A1(n16731), .A2(n16724), .A3(n16726), .ZN(n12975) );
  NAND2_X1 U14916 ( .A1(n12975), .A2(n13859), .ZN(n16660) );
  NAND3_X1 U14917 ( .A1(n16707), .A2(n16662), .A3(n16660), .ZN(n12976) );
  AOI21_X1 U14918 ( .B1(n16669), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12976), .ZN(n12977) );
  AND3_X1 U14919 ( .A1(n16671), .A2(n16666), .A3(n12977), .ZN(n12978) );
  NAND2_X1 U14920 ( .A1(n12980), .A2(n12979), .ZN(n12981) );
  AND2_X1 U14921 ( .A1(n12985), .A2(n12981), .ZN(n18682) );
  NAND2_X1 U14922 ( .A1(n18682), .A2(n13859), .ZN(n12982) );
  INV_X1 U14923 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16847) );
  XNOR2_X1 U14924 ( .A(n12982), .B(n16847), .ZN(n16651) );
  NAND2_X1 U14925 ( .A1(n12982), .A2(n16847), .ZN(n12983) );
  XNOR2_X1 U14926 ( .A(n12986), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16644) );
  INV_X1 U14927 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16833) );
  INV_X1 U14928 ( .A(n12987), .ZN(n12988) );
  XNOR2_X1 U14929 ( .A(n12989), .B(n12988), .ZN(n18708) );
  INV_X1 U14930 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16818) );
  NOR2_X1 U14931 ( .A1(n16730), .A2(n16818), .ZN(n12990) );
  NAND2_X1 U14932 ( .A1(n18708), .A2(n12990), .ZN(n16631) );
  NAND2_X1 U14933 ( .A1(n18708), .A2(n13859), .ZN(n12991) );
  NAND2_X1 U14934 ( .A1(n12991), .A2(n16818), .ZN(n16632) );
  INV_X1 U14935 ( .A(n12993), .ZN(n12994) );
  NAND2_X1 U14936 ( .A1(n18734), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16587) );
  OR2_X1 U14937 ( .A1(n16587), .A2(n16730), .ZN(n13011) );
  NAND2_X1 U14938 ( .A1(n18734), .A2(n13859), .ZN(n12996) );
  INV_X1 U14939 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16799) );
  NAND2_X1 U14940 ( .A1(n12996), .A2(n16799), .ZN(n12997) );
  NAND2_X1 U14941 ( .A1(n13011), .A2(n12997), .ZN(n16611) );
  INV_X1 U14942 ( .A(n12998), .ZN(n12999) );
  XNOR2_X1 U14943 ( .A(n13000), .B(n12999), .ZN(n18721) );
  NAND2_X1 U14944 ( .A1(n18721), .A2(n13859), .ZN(n13012) );
  INV_X1 U14945 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16798) );
  AND2_X1 U14946 ( .A1(n13002), .A2(n13001), .ZN(n13003) );
  OR2_X1 U14947 ( .A1(n13003), .A2(n13007), .ZN(n18751) );
  NOR2_X1 U14948 ( .A1(n18751), .A2(n16730), .ZN(n16589) );
  NOR2_X1 U14949 ( .A1(n13007), .A2(n13006), .ZN(n13008) );
  OR2_X1 U14950 ( .A1(n13853), .A2(n13008), .ZN(n18763) );
  NOR2_X1 U14951 ( .A1(n18763), .A2(n16730), .ZN(n16591) );
  OAI21_X1 U14952 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n16591), .ZN(n13009) );
  INV_X1 U14953 ( .A(n16591), .ZN(n13010) );
  INV_X1 U14954 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16595) );
  NAND2_X1 U14955 ( .A1(n13010), .A2(n16595), .ZN(n13014) );
  INV_X1 U14956 ( .A(n13011), .ZN(n13013) );
  NOR2_X1 U14957 ( .A1(n13012), .A2(n16798), .ZN(n16620) );
  AND2_X1 U14958 ( .A1(n15667), .A2(n16336), .ZN(n14663) );
  INV_X1 U14959 ( .A(n14663), .ZN(n13016) );
  NOR2_X1 U14960 ( .A1(n13015), .A2(n13016), .ZN(n14233) );
  NAND2_X1 U14961 ( .A1(n13018), .A2(n13017), .ZN(n13862) );
  INV_X1 U14962 ( .A(n13862), .ZN(n13026) );
  INV_X1 U14963 ( .A(n13028), .ZN(n13870) );
  OAI21_X1 U14964 ( .B1(n13020), .B2(n13870), .A(n13019), .ZN(n13025) );
  INV_X1 U14965 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17102) );
  AND2_X1 U14966 ( .A1(n17102), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13021) );
  AOI21_X1 U14967 ( .B1(n13026), .B2(n13025), .A(n13886), .ZN(n14645) );
  NAND2_X1 U14968 ( .A1(n14233), .A2(n14645), .ZN(n13908) );
  NOR2_X1 U14969 ( .A1(n13015), .A2(n13861), .ZN(n14637) );
  XNOR2_X1 U14970 ( .A(n13028), .B(n13027), .ZN(n13864) );
  NAND4_X1 U14971 ( .A1(n13880), .A2(n13863), .A3(n13876), .A4(n13864), .ZN(
        n13030) );
  NAND2_X1 U14972 ( .A1(n13030), .A2(n13029), .ZN(n14638) );
  NAND4_X1 U14973 ( .A1(n13880), .A2(n13863), .A3(n13865), .A4(n13876), .ZN(
        n13031) );
  NAND2_X1 U14974 ( .A1(n13031), .A2(n18890), .ZN(n13032) );
  OR2_X1 U14975 ( .A1(n14638), .A2(n13032), .ZN(n13036) );
  AND2_X1 U14976 ( .A1(n14656), .A2(n13033), .ZN(n14291) );
  NAND2_X1 U14977 ( .A1(n15484), .A2(n14291), .ZN(n13034) );
  INV_X1 U14978 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18912) );
  AOI21_X1 U14979 ( .B1(n13034), .B2(n18912), .A(n18890), .ZN(n17483) );
  INV_X1 U14980 ( .A(n17483), .ZN(n13035) );
  NAND2_X1 U14981 ( .A1(n13036), .A2(n13035), .ZN(n17101) );
  NAND2_X1 U14982 ( .A1(n14637), .A2(n17101), .ZN(n13037) );
  NAND2_X1 U14983 ( .A1(n13908), .A2(n13037), .ZN(n14659) );
  OR2_X2 U14984 ( .A1(n18911), .A2(n15667), .ZN(n17461) );
  INV_X1 U14985 ( .A(n13038), .ZN(n13040) );
  AND2_X1 U14986 ( .A1(n13040), .A2(n13039), .ZN(n13041) );
  INV_X1 U14987 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n18835) );
  NAND2_X1 U14988 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13044) );
  AOI22_X1 U14989 ( .A1(n13047), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13043) );
  OAI211_X1 U14990 ( .C1(n13124), .C2(n18835), .A(n13044), .B(n13043), .ZN(
        n15430) );
  INV_X1 U14991 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15219) );
  NAND2_X1 U14992 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13046) );
  AOI22_X1 U14993 ( .A1(n14180), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13045) );
  OAI211_X1 U14994 ( .C1(n13124), .C2(n15219), .A(n13046), .B(n13045), .ZN(
        n15216) );
  NAND2_X1 U14995 ( .A1(n15433), .A2(n15216), .ZN(n14475) );
  INV_X1 U14996 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U14997 ( .A1(n13047), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13048) );
  OAI21_X1 U14998 ( .B1(n13124), .B2(n13049), .A(n13048), .ZN(n13050) );
  INV_X1 U14999 ( .A(n13050), .ZN(n13052) );
  NAND2_X1 U15000 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13051) );
  INV_X1 U15001 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U15002 ( .A1(n14180), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13055) );
  OAI21_X1 U15003 ( .B1(n13124), .B2(n13056), .A(n13055), .ZN(n13057) );
  AOI21_X1 U15004 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n14179), .A(
        n13057), .ZN(n14507) );
  AOI22_X1 U15005 ( .A1(n14180), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13059) );
  NAND2_X1 U15006 ( .A1(n10999), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n13058) );
  OAI211_X1 U15007 ( .C1(n13042), .C2(n14208), .A(n13059), .B(n13058), .ZN(
        n14595) );
  INV_X1 U15008 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U15009 ( .A1(n14180), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13060) );
  OAI21_X1 U15010 ( .B1(n13124), .B2(n13061), .A(n13060), .ZN(n13062) );
  INV_X1 U15011 ( .A(n13062), .ZN(n13064) );
  NAND2_X1 U15012 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13063) );
  AOI22_X1 U15013 ( .A1(n14180), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n13066) );
  NAND2_X1 U15014 ( .A1(n10999), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n13065) );
  OAI211_X1 U15015 ( .C1(n13042), .C2(n18814), .A(n13066), .B(n13065), .ZN(
        n14873) );
  INV_X1 U15016 ( .A(n14872), .ZN(n14895) );
  INV_X1 U15017 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n13069) );
  NAND2_X1 U15018 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13068) );
  AOI22_X1 U15019 ( .A1(n14180), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n13067) );
  OAI211_X1 U15020 ( .C1(n13124), .C2(n13069), .A(n13068), .B(n13067), .ZN(
        n14896) );
  NAND2_X1 U15021 ( .A1(n14895), .A2(n14896), .ZN(n14926) );
  INV_X1 U15022 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U15023 ( .A1(n14180), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n13070) );
  OAI21_X1 U15024 ( .B1(n13124), .B2(n13071), .A(n13070), .ZN(n13072) );
  INV_X1 U15025 ( .A(n13072), .ZN(n13074) );
  NAND2_X1 U15026 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13073) );
  INV_X1 U15027 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U15028 ( .A1(n14180), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n13075) );
  OAI21_X1 U15029 ( .B1(n13124), .B2(n13076), .A(n13075), .ZN(n13077) );
  INV_X1 U15030 ( .A(n13077), .ZN(n13079) );
  NAND2_X1 U15031 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13078) );
  INV_X1 U15032 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n13083) );
  NAND2_X1 U15033 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13082) );
  AOI22_X1 U15034 ( .A1(n14180), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n13081) );
  OAI211_X1 U15035 ( .C1(n13124), .C2(n13083), .A(n13082), .B(n13081), .ZN(
        n15138) );
  INV_X1 U15036 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n17556) );
  NAND2_X1 U15037 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13085) );
  AOI22_X1 U15038 ( .A1(n14180), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n13084) );
  OAI211_X1 U15039 ( .C1(n13124), .C2(n17556), .A(n13085), .B(n13084), .ZN(
        n15228) );
  INV_X1 U15040 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n17557) );
  AOI22_X1 U15041 ( .A1(n14180), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n13086) );
  OAI21_X1 U15042 ( .B1(n13124), .B2(n17557), .A(n13086), .ZN(n13087) );
  INV_X1 U15043 ( .A(n13087), .ZN(n13089) );
  NAND2_X1 U15044 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13088) );
  INV_X1 U15045 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U15046 ( .A1(n14180), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n13090) );
  OAI21_X1 U15047 ( .B1(n13124), .B2(n13091), .A(n13090), .ZN(n13092) );
  INV_X1 U15048 ( .A(n13092), .ZN(n13094) );
  NAND2_X1 U15049 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13093) );
  INV_X1 U15050 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n17558) );
  AOI22_X1 U15051 ( .A1(n14180), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n13095) );
  OAI21_X1 U15052 ( .B1(n13124), .B2(n17558), .A(n13095), .ZN(n13096) );
  INV_X1 U15053 ( .A(n13096), .ZN(n13098) );
  NAND2_X1 U15054 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13097) );
  INV_X1 U15055 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n18647) );
  NAND2_X1 U15056 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13100) );
  AOI22_X1 U15057 ( .A1(n14180), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n13099) );
  OAI211_X1 U15058 ( .C1(n13124), .C2(n18647), .A(n13100), .B(n13099), .ZN(
        n16470) );
  NAND2_X1 U15059 ( .A1(n16471), .A2(n16470), .ZN(n16463) );
  INV_X1 U15060 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n14158) );
  AOI22_X1 U15061 ( .A1(n14180), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n13101) );
  OAI21_X1 U15062 ( .B1(n12743), .B2(n14158), .A(n13101), .ZN(n13102) );
  INV_X1 U15063 ( .A(n13102), .ZN(n13104) );
  NAND2_X1 U15064 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13103) );
  INV_X1 U15065 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U15066 ( .A1(n14180), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n13105) );
  OAI21_X1 U15067 ( .B1(n12743), .B2(n13106), .A(n13105), .ZN(n13107) );
  INV_X1 U15068 ( .A(n13107), .ZN(n13109) );
  NAND2_X1 U15069 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13108) );
  INV_X1 U15070 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16652) );
  NAND2_X1 U15071 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13111) );
  AOI22_X1 U15072 ( .A1(n14180), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n13110) );
  OAI211_X1 U15073 ( .C1(n13124), .C2(n16652), .A(n13111), .B(n13110), .ZN(
        n16444) );
  INV_X1 U15074 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n18687) );
  NAND2_X1 U15075 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13113) );
  AOI22_X1 U15076 ( .A1(n14180), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n13112) );
  OAI211_X1 U15077 ( .C1(n13124), .C2(n18687), .A(n13113), .B(n13112), .ZN(
        n16436) );
  INV_X1 U15078 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17565) );
  AOI22_X1 U15079 ( .A1(n14180), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n13114) );
  OAI21_X1 U15080 ( .B1(n12743), .B2(n17565), .A(n13114), .ZN(n13115) );
  INV_X1 U15081 ( .A(n13115), .ZN(n13117) );
  NAND2_X1 U15082 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13116) );
  INV_X1 U15083 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n18717) );
  AOI22_X1 U15084 ( .A1(n14180), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n13118) );
  OAI21_X1 U15085 ( .B1(n12743), .B2(n18717), .A(n13118), .ZN(n13119) );
  INV_X1 U15086 ( .A(n13119), .ZN(n13121) );
  NAND2_X1 U15087 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13120) );
  INV_X1 U15088 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17566) );
  NAND2_X1 U15089 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13123) );
  AOI22_X1 U15090 ( .A1(n14180), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n13122) );
  OAI211_X1 U15091 ( .C1(n13124), .C2(n17566), .A(n13123), .B(n13122), .ZN(
        n16410) );
  NAND2_X1 U15092 ( .A1(n16422), .A2(n16410), .ZN(n16412) );
  INV_X1 U15093 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n18739) );
  AOI22_X1 U15094 ( .A1(n14180), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n13125) );
  OAI21_X1 U15095 ( .B1(n12743), .B2(n18739), .A(n13125), .ZN(n13126) );
  INV_X1 U15096 ( .A(n13126), .ZN(n13128) );
  NAND2_X1 U15097 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13127) );
  AND2_X1 U15098 ( .A1(n13128), .A2(n13127), .ZN(n16407) );
  INV_X1 U15099 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U15100 ( .A1(n14180), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n13129) );
  OAI21_X1 U15101 ( .B1(n12743), .B2(n13130), .A(n13129), .ZN(n13131) );
  INV_X1 U15102 ( .A(n13131), .ZN(n13133) );
  NAND2_X1 U15103 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13132) );
  AND2_X1 U15104 ( .A1(n13133), .A2(n13132), .ZN(n16398) );
  INV_X1 U15105 ( .A(n16398), .ZN(n13134) );
  INV_X1 U15106 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n18764) );
  NAND2_X1 U15107 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13136) );
  AOI22_X1 U15108 ( .A1(n14180), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n13135) );
  OAI211_X1 U15109 ( .C1(n12743), .C2(n18764), .A(n13136), .B(n13135), .ZN(
        n13138) );
  OAI21_X1 U15110 ( .B1(n13137), .B2(n13138), .A(n15707), .ZN(n16390) );
  NAND2_X1 U15111 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n14840) );
  NAND2_X1 U15112 ( .A1(n19472), .A2(n14840), .ZN(n17480) );
  OR2_X1 U15113 ( .A1(n17480), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13139) );
  AND2_X1 U15114 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13140) );
  AND2_X2 U15115 ( .A1(n17459), .A2(n13140), .ZN(n17474) );
  INV_X1 U15116 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18766) );
  INV_X1 U15117 ( .A(n14438), .ZN(n14839) );
  INV_X1 U15118 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n14662) );
  NAND2_X1 U15119 ( .A1(n14662), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13141) );
  NAND2_X1 U15120 ( .A1(n14839), .A2(n13141), .ZN(n14301) );
  INV_X1 U15121 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16694) );
  INV_X1 U15122 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18622) );
  INV_X1 U15123 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17414) );
  INV_X1 U15124 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18688) );
  NAND2_X1 U15125 ( .A1(n16314), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16316) );
  INV_X1 U15126 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16625) );
  INV_X1 U15127 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16614) );
  INV_X1 U15128 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18740) );
  INV_X1 U15129 ( .A(n16323), .ZN(n13143) );
  AOI21_X1 U15130 ( .B1(n18766), .B2(n13143), .A(n16324), .ZN(n18770) );
  NAND2_X1 U15131 ( .A1(n17453), .A2(n18770), .ZN(n13145) );
  AND2_X1 U15132 ( .A1(n13144), .A2(n19508), .ZN(n16328) );
  INV_X1 U15133 ( .A(n18848), .ZN(n16675) );
  NAND2_X1 U15134 ( .A1(n16675), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16761) );
  OAI211_X1 U15135 ( .C1(n17459), .C2(n18766), .A(n13145), .B(n16761), .ZN(
        n13146) );
  OAI21_X1 U15136 ( .B1(n16771), .B2(n17461), .A(n13147), .ZN(n13188) );
  INV_X1 U15137 ( .A(n13952), .ZN(n13149) );
  NAND2_X1 U15138 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14307), .ZN(
        n14306) );
  NOR2_X1 U15139 ( .A1(n13952), .A2(n14306), .ZN(n13151) );
  INV_X1 U15140 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17065) );
  NOR2_X1 U15141 ( .A1(n13148), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13150) );
  XOR2_X1 U15142 ( .A(n13150), .B(n13149), .Z(n14272) );
  NOR2_X1 U15143 ( .A1(n17065), .A2(n14272), .ZN(n14271) );
  NOR2_X1 U15144 ( .A1(n13151), .A2(n14271), .ZN(n14333) );
  INV_X1 U15145 ( .A(n13962), .ZN(n13152) );
  XNOR2_X1 U15146 ( .A(n13153), .B(n13152), .ZN(n14334) );
  OAI21_X1 U15147 ( .B1(n14333), .B2(n14334), .A(n13154), .ZN(n13155) );
  NAND2_X1 U15148 ( .A1(n14333), .A2(n14334), .ZN(n14332) );
  NAND2_X1 U15149 ( .A1(n13155), .A2(n14332), .ZN(n17393) );
  OR2_X1 U15150 ( .A1(n17393), .A2(n18860), .ZN(n13156) );
  NAND2_X1 U15151 ( .A1(n17392), .A2(n13156), .ZN(n13158) );
  NAND2_X1 U15152 ( .A1(n17393), .A2(n18860), .ZN(n13157) );
  NAND2_X1 U15153 ( .A1(n13158), .A2(n13157), .ZN(n13163) );
  NAND2_X1 U15154 ( .A1(n13159), .A2(n13939), .ZN(n13160) );
  NAND2_X1 U15155 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  XNOR2_X1 U15156 ( .A(n13163), .B(n13162), .ZN(n17405) );
  NAND2_X1 U15157 ( .A1(n13163), .A2(n13162), .ZN(n13164) );
  NAND2_X1 U15158 ( .A1(n13165), .A2(n15215), .ZN(n15209) );
  INV_X1 U15159 ( .A(n13166), .ZN(n13167) );
  MUX2_X1 U15160 ( .A(n13173), .B(n15215), .S(n13165), .Z(n13169) );
  OAI21_X1 U15161 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n13166), .A(
        n13169), .ZN(n13170) );
  OR2_X1 U15162 ( .A1(n13165), .A2(n15215), .ZN(n15210) );
  NAND3_X1 U15163 ( .A1(n13171), .A2(n13166), .A3(n15209), .ZN(n13172) );
  NAND2_X1 U15164 ( .A1(n17415), .A2(n13172), .ZN(n15315) );
  XNOR2_X1 U15165 ( .A(n13178), .B(n16730), .ZN(n13175) );
  XNOR2_X1 U15166 ( .A(n13175), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15314) );
  INV_X1 U15167 ( .A(n13175), .ZN(n13176) );
  NAND2_X1 U15168 ( .A1(n13176), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13177) );
  INV_X1 U15169 ( .A(n13178), .ZN(n13179) );
  XNOR2_X1 U15170 ( .A(n13180), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17431) );
  INV_X1 U15171 ( .A(n13180), .ZN(n13181) );
  NAND3_X1 U15172 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16967) );
  NAND2_X1 U15173 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13182) );
  NOR2_X1 U15174 ( .A1(n16967), .A2(n13182), .ZN(n16968) );
  AND2_X1 U15175 ( .A1(n16968), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16921) );
  AND2_X1 U15176 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16923) );
  AND2_X1 U15177 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16875) );
  AND2_X1 U15178 ( .A1(n16875), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16873) );
  NAND2_X1 U15179 ( .A1(n16873), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14216) );
  AND2_X1 U15180 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14223) );
  AND2_X1 U15181 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16797) );
  AND2_X2 U15182 ( .A1(n16612), .A2(n16797), .ZN(n16613) );
  INV_X1 U15184 ( .A(n16605), .ZN(n13184) );
  AOI21_X1 U15185 ( .B1(n13184), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13186) );
  NAND2_X1 U15186 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13185) );
  NOR2_X1 U15187 ( .A1(n16769), .A2(n17463), .ZN(n13187) );
  OR2_X1 U15188 ( .A1(n13188), .A2(n13187), .ZN(P2_U2985) );
  NAND2_X1 U15189 ( .A1(n13190), .A2(n13189), .ZN(n18143) );
  OAI21_X1 U15190 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n13191), .A(
        n13192), .ZN(n18125) );
  INV_X1 U15191 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18139) );
  AOI21_X1 U15192 ( .B1(n13223), .B2(n13226), .A(n18139), .ZN(n13218) );
  OAI21_X1 U15193 ( .B1(n20982), .B2(n21137), .A(n11701), .ZN(n21071) );
  NAND4_X1 U15194 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A4(n21071), .ZN(n21091) );
  NOR2_X1 U15195 ( .A1(n21112), .A2(n21091), .ZN(n21113) );
  NAND3_X1 U15196 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21113), .ZN(n21131) );
  NOR2_X1 U15197 ( .A1(n21322), .A2(n21131), .ZN(n21313) );
  NAND2_X1 U15198 ( .A1(n21313), .A2(n13193), .ZN(n21267) );
  NAND3_X1 U15199 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n13194), .ZN(n13198) );
  OAI21_X1 U15200 ( .B1(n21267), .B2(n13198), .A(n21386), .ZN(n13840) );
  NAND2_X1 U15201 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n13840), .ZN(
        n21233) );
  INV_X1 U15202 ( .A(n21002), .ZN(n13196) );
  OAI21_X1 U15203 ( .B1(n13196), .B2(n13195), .A(n21010), .ZN(n21075) );
  NOR2_X1 U15204 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21363), .ZN(
        n21117) );
  INV_X1 U15205 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18004) );
  NOR2_X1 U15206 ( .A1(n11701), .A2(n20982), .ZN(n21072) );
  NAND4_X1 U15207 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A4(n21072), .ZN(n21093) );
  NOR2_X1 U15208 ( .A1(n21112), .A2(n21093), .ZN(n21114) );
  NAND2_X1 U15209 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21114), .ZN(
        n21366) );
  NOR2_X1 U15210 ( .A1(n21122), .A2(n21366), .ZN(n21136) );
  NAND2_X1 U15211 ( .A1(n21136), .A2(n21183), .ZN(n21180) );
  NOR2_X1 U15212 ( .A1(n18004), .A2(n21180), .ZN(n21035) );
  INV_X1 U15213 ( .A(n21035), .ZN(n21316) );
  NOR3_X1 U15214 ( .A1(n21117), .A2(n13197), .A3(n21316), .ZN(n21196) );
  NOR2_X1 U15215 ( .A1(n21362), .A2(n21196), .ZN(n21271) );
  AOI21_X1 U15216 ( .B1(n21321), .B2(n13198), .A(n21271), .ZN(n21231) );
  OAI21_X1 U15217 ( .B1(n21362), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n21231), .ZN(n13839) );
  AOI21_X1 U15218 ( .B1(n21386), .B2(n21233), .A(n13839), .ZN(n21253) );
  XNOR2_X1 U15219 ( .A(n20779), .B(n19177), .ZN(n13199) );
  OAI21_X1 U15220 ( .B1(n13199), .B2(n20312), .A(n21907), .ZN(n21404) );
  NOR3_X1 U15221 ( .A1(n13201), .A2(n13200), .A3(n21404), .ZN(n13217) );
  AOI211_X1 U15222 ( .C1(n20787), .C2(n17576), .A(n13203), .B(n13202), .ZN(
        n13205) );
  AOI21_X1 U15223 ( .B1(n13206), .B2(n13205), .A(n13204), .ZN(n13207) );
  AOI211_X1 U15224 ( .C1(n13210), .C2(n13209), .A(n13208), .B(n13207), .ZN(
        n15377) );
  NOR2_X1 U15225 ( .A1(n19220), .A2(n13211), .ZN(n13214) );
  OAI211_X1 U15226 ( .C1(n13214), .C2(n13213), .A(n13212), .B(n19177), .ZN(
        n13215) );
  OAI211_X1 U15227 ( .C1(n19095), .C2(n21385), .A(n15377), .B(n13215), .ZN(
        n13216) );
  OAI211_X1 U15228 ( .C1(n13818), .C2(n13218), .A(n21253), .B(n21275), .ZN(
        n13220) );
  NAND2_X1 U15229 ( .A1(n21084), .A2(n20812), .ZN(n21219) );
  OAI22_X1 U15230 ( .A1(n21244), .A2(n21219), .B1(n21245), .B2(n21268), .ZN(
        n13219) );
  INV_X1 U15231 ( .A(n17987), .ZN(n17986) );
  AOI22_X1 U15232 ( .A1(n21293), .A2(n21135), .B1(n21384), .B2(n21132), .ZN(
        n21141) );
  NAND2_X1 U15233 ( .A1(n21380), .A2(n11083), .ZN(n21367) );
  NOR2_X1 U15234 ( .A1(n21316), .A2(n21162), .ZN(n13835) );
  INV_X1 U15235 ( .A(n13835), .ZN(n13221) );
  OAI21_X1 U15236 ( .B1(n21141), .B2(n21322), .A(n13221), .ZN(n13222) );
  NOR2_X1 U15237 ( .A1(n21316), .A2(n21137), .ZN(n21178) );
  NAND2_X1 U15238 ( .A1(n17986), .A2(n21178), .ZN(n21041) );
  NAND2_X1 U15239 ( .A1(n17986), .A2(n21313), .ZN(n21037) );
  OAI22_X1 U15240 ( .A1(n21363), .A2(n21041), .B1(n21312), .B2(n21037), .ZN(
        n13834) );
  AOI21_X1 U15241 ( .B1(n17986), .B2(n13222), .A(n13834), .ZN(n21031) );
  NOR2_X1 U15242 ( .A1(n21031), .A2(n13833), .ZN(n21276) );
  NAND2_X1 U15243 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18112), .ZN(
        n21206) );
  NOR2_X1 U15244 ( .A1(n21206), .A2(n21205), .ZN(n18162) );
  NAND2_X1 U15245 ( .A1(n21276), .A2(n18162), .ZN(n21218) );
  NOR2_X1 U15246 ( .A1(n21218), .A2(n21229), .ZN(n21237) );
  AOI22_X1 U15247 ( .A1(n13191), .A2(n13223), .B1(n21237), .B2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13224) );
  NOR2_X1 U15248 ( .A1(n13224), .A2(n21263), .ZN(n13225) );
  NAND3_X1 U15249 ( .A1(n13227), .A2(n21373), .A3(n18125), .ZN(n13228) );
  INV_X2 U15250 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n13234) );
  INV_X1 U15251 ( .A(n13417), .ZN(n13373) );
  NAND2_X1 U15252 ( .A1(n13752), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13268) );
  INV_X1 U15253 ( .A(n13253), .ZN(n13231) );
  INV_X1 U15254 ( .A(n13242), .ZN(n13244) );
  INV_X1 U15255 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13232) );
  NAND2_X1 U15256 ( .A1(n13232), .A2(n13253), .ZN(n13233) );
  NAND2_X1 U15257 ( .A1(n13244), .A2(n13233), .ZN(n21667) );
  AOI22_X1 U15258 ( .A1(n21667), .A2(n13757), .B1(n13724), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13236) );
  NOR2_X2 U15259 ( .A1(n14683), .A2(n13234), .ZN(n13276) );
  NAND2_X1 U15260 ( .A1(n13276), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n13235) );
  OAI211_X1 U15261 ( .C1(n13268), .C2(n15008), .A(n13236), .B(n13235), .ZN(
        n13237) );
  INV_X1 U15262 ( .A(n13237), .ZN(n13238) );
  INV_X1 U15263 ( .A(n14727), .ZN(n13250) );
  NAND2_X1 U15264 ( .A1(n13234), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13240) );
  NAND2_X1 U15265 ( .A1(n13725), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n13239) );
  OAI211_X1 U15266 ( .C1(n13268), .C2(n17084), .A(n13240), .B(n13239), .ZN(
        n13241) );
  NAND2_X1 U15267 ( .A1(n13241), .A2(n11099), .ZN(n13247) );
  INV_X1 U15268 ( .A(n13277), .ZN(n13278) );
  INV_X1 U15269 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13243) );
  NAND2_X1 U15270 ( .A1(n13244), .A2(n13243), .ZN(n13245) );
  NAND2_X1 U15271 ( .A1(n13278), .A2(n13245), .ZN(n21676) );
  NAND2_X1 U15272 ( .A1(n21676), .A2(n13757), .ZN(n13246) );
  NAND2_X1 U15273 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  AOI21_X1 U15274 ( .B1(n13249), .B2(n13417), .A(n13248), .ZN(n14885) );
  NAND2_X1 U15275 ( .A1(n13251), .A2(n13417), .ZN(n13252) );
  NAND2_X1 U15276 ( .A1(n13252), .A2(n13344), .ZN(n13271) );
  INV_X2 U15277 ( .A(n11099), .ZN(n13757) );
  OAI21_X1 U15278 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13253), .ZN(n20150) );
  AOI22_X1 U15279 ( .A1(n13757), .A2(n20150), .B1(n13724), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13255) );
  NAND2_X1 U15280 ( .A1(n13725), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n13254) );
  OAI211_X1 U15281 ( .C1(n13268), .C2(n12023), .A(n13255), .B(n13254), .ZN(
        n13272) );
  XNOR2_X1 U15282 ( .A(n13271), .B(n13272), .ZN(n14704) );
  INV_X1 U15283 ( .A(n14704), .ZN(n13270) );
  INV_X1 U15284 ( .A(n13256), .ZN(n13258) );
  XNOR2_X2 U15285 ( .A(n13258), .B(n13257), .ZN(n14667) );
  NAND2_X1 U15286 ( .A1(n14667), .A2(n13417), .ZN(n13263) );
  AOI22_X1 U15287 ( .A1(n13725), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n13234), .ZN(n13261) );
  INV_X1 U15288 ( .A(n13268), .ZN(n13259) );
  NAND2_X1 U15289 ( .A1(n13259), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13260) );
  AND2_X1 U15290 ( .A1(n13261), .A2(n13260), .ZN(n13262) );
  NAND2_X1 U15291 ( .A1(n13263), .A2(n13262), .ZN(n14482) );
  AOI21_X1 U15292 ( .B1(n11025), .B2(n11859), .A(n13234), .ZN(n14523) );
  NAND2_X1 U15293 ( .A1(n13265), .A2(n13417), .ZN(n13267) );
  AOI22_X1 U15294 ( .A1(n13725), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13234), .ZN(n13266) );
  OAI211_X1 U15295 ( .C1(n13268), .C2(n15385), .A(n13267), .B(n13266), .ZN(
        n14524) );
  MUX2_X1 U15296 ( .A(n13757), .B(n14523), .S(n14524), .Z(n14481) );
  NAND2_X1 U15297 ( .A1(n14482), .A2(n14481), .ZN(n14480) );
  INV_X1 U15298 ( .A(n14480), .ZN(n13269) );
  NAND2_X1 U15299 ( .A1(n13270), .A2(n13269), .ZN(n13274) );
  NAND2_X1 U15300 ( .A1(n13271), .A2(n13272), .ZN(n13273) );
  NAND2_X1 U15301 ( .A1(n13275), .A2(n14726), .ZN(n14884) );
  INV_X1 U15302 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13283) );
  INV_X1 U15303 ( .A(n13287), .ZN(n13280) );
  INV_X1 U15304 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21688) );
  NAND2_X1 U15305 ( .A1(n13278), .A2(n21688), .ZN(n13279) );
  NAND2_X1 U15306 ( .A1(n13280), .A2(n13279), .ZN(n21689) );
  NOR2_X1 U15307 ( .A1(n13344), .A2(n21688), .ZN(n13281) );
  AOI21_X1 U15308 ( .B1(n21689), .B2(n13757), .A(n13281), .ZN(n13282) );
  OAI21_X1 U15309 ( .B1(n13583), .B2(n13283), .A(n13282), .ZN(n13284) );
  AOI21_X1 U15310 ( .B1(n13285), .B2(n13417), .A(n13284), .ZN(n14910) );
  INV_X1 U15311 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13290) );
  NAND2_X1 U15312 ( .A1(n13286), .A2(n13417), .ZN(n13289) );
  OAI21_X1 U15313 ( .B1(n13287), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13291), .ZN(n21702) );
  AOI22_X1 U15314 ( .A1(n21702), .A2(n13757), .B1(n13724), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13288) );
  OAI211_X1 U15315 ( .C1(n13583), .C2(n13290), .A(n13289), .B(n13288), .ZN(
        n14917) );
  INV_X1 U15316 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13294) );
  OAI21_X1 U15317 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13292), .A(
        n13313), .ZN(n21712) );
  AOI22_X1 U15318 ( .A1(n13757), .A2(n21712), .B1(n13724), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13293) );
  OAI21_X1 U15319 ( .B1(n13583), .B2(n13294), .A(n13293), .ZN(n13295) );
  AOI21_X1 U15320 ( .B1(n13296), .B2(n13417), .A(n13295), .ZN(n15114) );
  INV_X1 U15321 ( .A(n15114), .ZN(n13297) );
  XOR2_X1 U15322 ( .A(n13312), .B(n13313), .Z(n21725) );
  AOI22_X1 U15323 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U15324 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n13709), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U15325 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13701), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U15326 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13299) );
  NAND4_X1 U15327 ( .A1(n13302), .A2(n13301), .A3(n13300), .A4(n13299), .ZN(
        n13308) );
  AOI22_X1 U15328 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U15329 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U15330 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13702), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U15331 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11037), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13303) );
  NAND4_X1 U15332 ( .A1(n13306), .A2(n13305), .A3(n13304), .A4(n13303), .ZN(
        n13307) );
  OR2_X1 U15333 ( .A1(n13308), .A2(n13307), .ZN(n13309) );
  AOI22_X1 U15334 ( .A1(n13417), .A2(n13309), .B1(n13724), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13311) );
  NAND2_X1 U15335 ( .A1(n13276), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13310) );
  OAI211_X1 U15336 ( .C1(n21725), .C2(n11099), .A(n13311), .B(n13310), .ZN(
        n15122) );
  INV_X1 U15337 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21731) );
  XNOR2_X1 U15338 ( .A(n13329), .B(n21731), .ZN(n21740) );
  OR2_X1 U15339 ( .A1(n21740), .A2(n11099), .ZN(n13328) );
  AOI22_X1 U15340 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U15341 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U15342 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13315) );
  AOI22_X1 U15343 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13314) );
  NAND4_X1 U15344 ( .A1(n13317), .A2(n13316), .A3(n13315), .A4(n13314), .ZN(
        n13323) );
  AOI22_X1 U15345 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U15346 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13320) );
  AOI22_X1 U15347 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13319) );
  AOI22_X1 U15348 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13318) );
  NAND4_X1 U15349 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n13318), .ZN(
        n13322) );
  OAI21_X1 U15350 ( .B1(n13323), .B2(n13322), .A(n13417), .ZN(n13326) );
  NAND2_X1 U15351 ( .A1(n13276), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13325) );
  NAND2_X1 U15352 ( .A1(n13724), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13324) );
  NAND2_X1 U15353 ( .A1(n13328), .A2(n13327), .ZN(n15131) );
  XOR2_X1 U15354 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n13343), .Z(
        n20186) );
  AOI22_X1 U15355 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13333) );
  AOI22_X1 U15356 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U15357 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13331) );
  AOI22_X1 U15358 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13330) );
  NAND4_X1 U15359 ( .A1(n13333), .A2(n13332), .A3(n13331), .A4(n13330), .ZN(
        n13339) );
  AOI22_X1 U15360 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U15361 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13336) );
  AOI22_X1 U15362 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13335) );
  AOI22_X1 U15363 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13334) );
  NAND4_X1 U15364 ( .A1(n13337), .A2(n13336), .A3(n13335), .A4(n13334), .ZN(
        n13338) );
  OR2_X1 U15365 ( .A1(n13339), .A2(n13338), .ZN(n13340) );
  AOI22_X1 U15366 ( .A1(n13417), .A2(n13340), .B1(n13724), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13342) );
  NAND2_X1 U15367 ( .A1(n13276), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n13341) );
  OAI211_X1 U15368 ( .C1(n20186), .C2(n11099), .A(n13342), .B(n13341), .ZN(
        n15148) );
  XNOR2_X1 U15369 ( .A(n13369), .B(n15262), .ZN(n20193) );
  INV_X1 U15370 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20057) );
  OAI22_X1 U15371 ( .A1(n13583), .A2(n20057), .B1(n13344), .B2(n15262), .ZN(
        n13345) );
  AOI21_X1 U15372 ( .B1(n20193), .B2(n13757), .A(n13345), .ZN(n13357) );
  AOI22_X1 U15373 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13349) );
  AOI22_X1 U15374 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U15375 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13347) );
  AOI22_X1 U15376 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13346) );
  NAND4_X1 U15377 ( .A1(n13349), .A2(n13348), .A3(n13347), .A4(n13346), .ZN(
        n13355) );
  AOI22_X1 U15378 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13353) );
  AOI22_X1 U15379 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13352) );
  AOI22_X1 U15380 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13351) );
  AOI22_X1 U15381 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13350) );
  NAND4_X1 U15382 ( .A1(n13353), .A2(n13352), .A3(n13351), .A4(n13350), .ZN(
        n13354) );
  OR2_X1 U15383 ( .A1(n13355), .A2(n13354), .ZN(n13356) );
  NAND2_X1 U15384 ( .A1(n13417), .A2(n13356), .ZN(n15254) );
  AOI22_X1 U15385 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13362) );
  AOI22_X1 U15386 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13361) );
  AOI22_X1 U15387 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13360) );
  AOI22_X1 U15388 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13359) );
  NAND4_X1 U15389 ( .A1(n13362), .A2(n13361), .A3(n13360), .A4(n13359), .ZN(
        n13368) );
  AOI22_X1 U15390 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U15391 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U15392 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U15393 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13363) );
  NAND4_X1 U15394 ( .A1(n13366), .A2(n13365), .A3(n13364), .A4(n13363), .ZN(
        n13367) );
  NOR2_X1 U15395 ( .A1(n13368), .A2(n13367), .ZN(n13372) );
  XNOR2_X1 U15396 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n13374), .ZN(
        n20202) );
  AOI22_X1 U15397 ( .A1(n13757), .A2(n20202), .B1(n13724), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13371) );
  NAND2_X1 U15398 ( .A1(n13725), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n13370) );
  OAI211_X1 U15399 ( .C1(n13373), .C2(n13372), .A(n13371), .B(n13370), .ZN(
        n15328) );
  XOR2_X1 U15400 ( .A(n15863), .B(n13390), .Z(n15868) );
  INV_X1 U15401 ( .A(n15868), .ZN(n16151) );
  AOI22_X1 U15402 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13378) );
  AOI22_X1 U15403 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13377) );
  AOI22_X1 U15404 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U15405 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13375) );
  NAND4_X1 U15406 ( .A1(n13378), .A2(n13377), .A3(n13376), .A4(n13375), .ZN(
        n13384) );
  AOI22_X1 U15407 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13659), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13382) );
  AOI22_X1 U15408 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13381) );
  AOI22_X1 U15409 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13380) );
  AOI22_X1 U15410 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13379) );
  NAND4_X1 U15411 ( .A1(n13382), .A2(n13381), .A3(n13380), .A4(n13379), .ZN(
        n13383) );
  OAI21_X1 U15412 ( .B1(n13384), .B2(n13383), .A(n13417), .ZN(n13387) );
  NAND2_X1 U15413 ( .A1(n13725), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13386) );
  NAND2_X1 U15414 ( .A1(n13724), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13385) );
  NAND3_X1 U15415 ( .A1(n13387), .A2(n13386), .A3(n13385), .ZN(n13388) );
  AOI21_X1 U15416 ( .B1(n16151), .B2(n13757), .A(n13388), .ZN(n15855) );
  XNOR2_X1 U15417 ( .A(n13405), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16139) );
  AOI22_X1 U15418 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U15419 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13393) );
  AOI22_X1 U15420 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13392) );
  AOI22_X1 U15421 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13391) );
  NAND4_X1 U15422 ( .A1(n13394), .A2(n13393), .A3(n13392), .A4(n13391), .ZN(
        n13400) );
  AOI22_X1 U15423 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U15424 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13397) );
  AOI22_X1 U15425 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U15426 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13395) );
  NAND4_X1 U15427 ( .A1(n13398), .A2(n13397), .A3(n13396), .A4(n13395), .ZN(
        n13399) );
  OAI21_X1 U15428 ( .B1(n13400), .B2(n13399), .A(n13417), .ZN(n13403) );
  NAND2_X1 U15429 ( .A1(n13725), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13402) );
  NAND2_X1 U15430 ( .A1(n13724), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13401) );
  NAND3_X1 U15431 ( .A1(n13403), .A2(n13402), .A3(n13401), .ZN(n13404) );
  AOI21_X1 U15432 ( .B1(n16139), .B2(n13757), .A(n13404), .ZN(n15846) );
  XOR2_X1 U15433 ( .A(n15839), .B(n13420), .Z(n20210) );
  AOI22_X1 U15434 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13409) );
  AOI22_X1 U15435 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13408) );
  AOI22_X1 U15436 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U15437 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13406) );
  NAND4_X1 U15438 ( .A1(n13409), .A2(n13408), .A3(n13407), .A4(n13406), .ZN(
        n13415) );
  AOI22_X1 U15439 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U15440 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U15441 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U15442 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13410) );
  NAND4_X1 U15443 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n13410), .ZN(
        n13414) );
  OR2_X1 U15444 ( .A1(n13415), .A2(n13414), .ZN(n13416) );
  AOI22_X1 U15445 ( .A1(n13417), .A2(n13416), .B1(n13724), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13419) );
  NAND2_X1 U15446 ( .A1(n13725), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13418) );
  OAI211_X1 U15447 ( .C1(n20210), .C2(n11099), .A(n13419), .B(n13418), .ZN(
        n15832) );
  INV_X1 U15448 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n13421) );
  XNOR2_X1 U15449 ( .A(n13438), .B(n13421), .ZN(n21751) );
  OR2_X1 U15450 ( .A1(n21751), .A2(n11099), .ZN(n13437) );
  AOI22_X1 U15451 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13659), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U15452 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U15453 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U15454 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13423) );
  NAND4_X1 U15455 ( .A1(n13426), .A2(n13425), .A3(n13424), .A4(n13423), .ZN(
        n13432) );
  AOI22_X1 U15456 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U15457 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13701), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13429) );
  AOI22_X1 U15458 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U15459 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13427) );
  NAND4_X1 U15460 ( .A1(n13430), .A2(n13429), .A3(n13428), .A4(n13427), .ZN(
        n13431) );
  NOR2_X1 U15461 ( .A1(n13432), .A2(n13431), .ZN(n13434) );
  AOI22_X1 U15462 ( .A1(n13725), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13234), .ZN(n13433) );
  OAI21_X1 U15463 ( .B1(n13694), .B2(n13434), .A(n13433), .ZN(n13435) );
  NAND2_X1 U15464 ( .A1(n13435), .A2(n11099), .ZN(n13436) );
  XOR2_X1 U15465 ( .A(n15826), .B(n13453), .Z(n20221) );
  AOI22_X1 U15466 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13442) );
  AOI22_X1 U15467 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13441) );
  AOI22_X1 U15468 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U15469 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13439) );
  NAND4_X1 U15470 ( .A1(n13442), .A2(n13441), .A3(n13440), .A4(n13439), .ZN(
        n13448) );
  AOI22_X1 U15471 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U15472 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13445) );
  AOI22_X1 U15473 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13444) );
  AOI22_X1 U15474 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13443) );
  NAND4_X1 U15475 ( .A1(n13446), .A2(n13445), .A3(n13444), .A4(n13443), .ZN(
        n13447) );
  NOR2_X1 U15476 ( .A1(n13448), .A2(n13447), .ZN(n13450) );
  AOI22_X1 U15477 ( .A1(n13725), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13724), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13449) );
  OAI21_X1 U15478 ( .B1(n13694), .B2(n13450), .A(n13449), .ZN(n13451) );
  INV_X1 U15479 ( .A(n15817), .ZN(n13452) );
  AND2_X2 U15480 ( .A1(n15814), .A2(n13452), .ZN(n15815) );
  XNOR2_X1 U15481 ( .A(n13481), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21762) );
  AOI21_X1 U15482 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21756), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13454) );
  AOI21_X1 U15483 ( .B1(n13276), .B2(P1_EAX_REG_18__SCAN_IN), .A(n13454), .ZN(
        n13466) );
  AOI22_X1 U15484 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13458) );
  AOI22_X1 U15485 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13659), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U15486 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U15487 ( .A1(n13681), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13455) );
  NAND4_X1 U15488 ( .A1(n13458), .A2(n13457), .A3(n13456), .A4(n13455), .ZN(
        n13464) );
  AOI22_X1 U15489 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13462) );
  AOI22_X1 U15490 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13461) );
  AOI22_X1 U15491 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13460) );
  AOI22_X1 U15492 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13459) );
  NAND4_X1 U15493 ( .A1(n13462), .A2(n13461), .A3(n13460), .A4(n13459), .ZN(
        n13463) );
  OAI21_X1 U15494 ( .B1(n13464), .B2(n13463), .A(n13718), .ZN(n13465) );
  AOI22_X1 U15495 ( .A1(n21762), .A2(n13757), .B1(n13466), .B2(n13465), .ZN(
        n15933) );
  AOI22_X1 U15496 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13470) );
  AOI22_X1 U15497 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13469) );
  AOI22_X1 U15498 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U15499 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13467) );
  NAND4_X1 U15500 ( .A1(n13470), .A2(n13469), .A3(n13468), .A4(n13467), .ZN(
        n13476) );
  AOI22_X1 U15501 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13474) );
  AOI22_X1 U15502 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13473) );
  AOI22_X1 U15503 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13472) );
  AOI22_X1 U15504 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13471) );
  NAND4_X1 U15505 ( .A1(n13474), .A2(n13473), .A3(n13472), .A4(n13471), .ZN(
        n13475) );
  NOR2_X1 U15506 ( .A1(n13476), .A2(n13475), .ZN(n13480) );
  NAND2_X1 U15507 ( .A1(n13234), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13477) );
  NAND2_X1 U15508 ( .A1(n11099), .A2(n13477), .ZN(n13478) );
  AOI21_X1 U15509 ( .B1(n13276), .B2(P1_EAX_REG_19__SCAN_IN), .A(n13478), .ZN(
        n13479) );
  OAI21_X1 U15510 ( .B1(n13694), .B2(n13480), .A(n13479), .ZN(n13485) );
  OAI21_X1 U15511 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n13482), .A(
        n13518), .ZN(n21767) );
  INV_X1 U15512 ( .A(n21767), .ZN(n13483) );
  NAND2_X1 U15513 ( .A1(n13483), .A2(n13757), .ZN(n13484) );
  NAND2_X1 U15514 ( .A1(n13485), .A2(n13484), .ZN(n15929) );
  AOI22_X1 U15515 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13489) );
  AOI22_X1 U15516 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13488) );
  AOI22_X1 U15517 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U15518 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13486) );
  NAND4_X1 U15519 ( .A1(n13489), .A2(n13488), .A3(n13487), .A4(n13486), .ZN(
        n13495) );
  AOI22_X1 U15520 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13493) );
  AOI22_X1 U15521 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13492) );
  AOI22_X1 U15522 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13491) );
  AOI22_X1 U15523 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13490) );
  NAND4_X1 U15524 ( .A1(n13493), .A2(n13492), .A3(n13491), .A4(n13490), .ZN(
        n13494) );
  NOR2_X1 U15525 ( .A1(n13495), .A2(n13494), .ZN(n13499) );
  NOR2_X1 U15526 ( .A1(n13517), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13496) );
  OR2_X1 U15527 ( .A1(n13757), .A2(n13496), .ZN(n13497) );
  AOI21_X1 U15528 ( .B1(n13276), .B2(P1_EAX_REG_20__SCAN_IN), .A(n13497), .ZN(
        n13498) );
  OAI21_X1 U15529 ( .B1(n13694), .B2(n13499), .A(n13498), .ZN(n13501) );
  XNOR2_X1 U15530 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n13518), .ZN(
        n21786) );
  NAND2_X1 U15531 ( .A1(n13757), .A2(n21786), .ZN(n13500) );
  AOI22_X1 U15532 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13506) );
  AOI22_X1 U15533 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13505) );
  AOI22_X1 U15534 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13504) );
  AOI22_X1 U15535 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13503) );
  NAND4_X1 U15536 ( .A1(n13506), .A2(n13505), .A3(n13504), .A4(n13503), .ZN(
        n13512) );
  AOI22_X1 U15537 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13510) );
  AOI22_X1 U15538 ( .A1(n13681), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13509) );
  AOI22_X1 U15539 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13508) );
  AOI22_X1 U15540 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13642), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13507) );
  NAND4_X1 U15541 ( .A1(n13510), .A2(n13509), .A3(n13508), .A4(n13507), .ZN(
        n13511) );
  NOR2_X1 U15542 ( .A1(n13512), .A2(n13511), .ZN(n13516) );
  NAND2_X1 U15543 ( .A1(n13234), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13513) );
  NAND2_X1 U15544 ( .A1(n11099), .A2(n13513), .ZN(n13514) );
  AOI21_X1 U15545 ( .B1(n13276), .B2(P1_EAX_REG_21__SCAN_IN), .A(n13514), .ZN(
        n13515) );
  OAI21_X1 U15546 ( .B1(n13694), .B2(n13516), .A(n13515), .ZN(n13522) );
  OAI21_X1 U15547 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n13519), .A(
        n13563), .ZN(n21796) );
  INV_X1 U15548 ( .A(n21796), .ZN(n13520) );
  NAND2_X1 U15549 ( .A1(n13520), .A2(n13757), .ZN(n13521) );
  NAND2_X1 U15550 ( .A1(n13522), .A2(n13521), .ZN(n15916) );
  INV_X1 U15551 ( .A(n15916), .ZN(n13523) );
  AOI22_X1 U15552 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U15553 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13526) );
  AOI22_X1 U15554 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U15555 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13524) );
  NAND4_X1 U15556 ( .A1(n13527), .A2(n13526), .A3(n13525), .A4(n13524), .ZN(
        n13533) );
  AOI22_X1 U15557 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13531) );
  AOI22_X1 U15558 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13530) );
  AOI22_X1 U15559 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13529) );
  AOI22_X1 U15560 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13528) );
  NAND4_X1 U15561 ( .A1(n13531), .A2(n13530), .A3(n13529), .A4(n13528), .ZN(
        n13532) );
  NOR2_X1 U15562 ( .A1(n13533), .A2(n13532), .ZN(n13536) );
  INV_X1 U15563 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21821) );
  AOI21_X1 U15564 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21821), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13534) );
  AOI21_X1 U15565 ( .B1(n13276), .B2(P1_EAX_REG_22__SCAN_IN), .A(n13534), .ZN(
        n13535) );
  OAI21_X1 U15566 ( .B1(n13694), .B2(n13536), .A(n13535), .ZN(n13538) );
  XNOR2_X1 U15567 ( .A(n13563), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n21817) );
  NAND2_X1 U15568 ( .A1(n21817), .A2(n13757), .ZN(n13537) );
  AOI22_X1 U15569 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13542) );
  AOI22_X1 U15570 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U15571 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U15572 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13539) );
  NAND4_X1 U15573 ( .A1(n13542), .A2(n13541), .A3(n13540), .A4(n13539), .ZN(
        n13548) );
  AOI22_X1 U15574 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13546) );
  AOI22_X1 U15575 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13545) );
  AOI22_X1 U15576 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13544) );
  AOI22_X1 U15577 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13543) );
  NAND4_X1 U15578 ( .A1(n13546), .A2(n13545), .A3(n13544), .A4(n13543), .ZN(
        n13547) );
  NOR2_X1 U15579 ( .A1(n13548), .A2(n13547), .ZN(n13571) );
  AOI22_X1 U15580 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13552) );
  AOI22_X1 U15581 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n13701), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13551) );
  AOI22_X1 U15582 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13550) );
  AOI22_X1 U15583 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13549) );
  NAND4_X1 U15584 ( .A1(n13552), .A2(n13551), .A3(n13550), .A4(n13549), .ZN(
        n13558) );
  AOI22_X1 U15585 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13699), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13556) );
  AOI22_X1 U15586 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13681), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13555) );
  AOI22_X1 U15587 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13659), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13554) );
  AOI22_X1 U15588 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13553) );
  NAND4_X1 U15589 ( .A1(n13556), .A2(n13555), .A3(n13554), .A4(n13553), .ZN(
        n13557) );
  NOR2_X1 U15590 ( .A1(n13558), .A2(n13557), .ZN(n13572) );
  XNOR2_X1 U15591 ( .A(n13571), .B(n13572), .ZN(n13562) );
  NAND2_X1 U15592 ( .A1(n13234), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13559) );
  NAND2_X1 U15593 ( .A1(n11099), .A2(n13559), .ZN(n13560) );
  AOI21_X1 U15594 ( .B1(n13276), .B2(P1_EAX_REG_23__SCAN_IN), .A(n13560), .ZN(
        n13561) );
  OAI21_X1 U15595 ( .B1(n13694), .B2(n13562), .A(n13561), .ZN(n13570) );
  INV_X1 U15596 ( .A(n13565), .ZN(n13567) );
  INV_X1 U15597 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13566) );
  NAND2_X1 U15598 ( .A1(n13567), .A2(n13566), .ZN(n13568) );
  AND2_X1 U15599 ( .A1(n13606), .A2(n13568), .ZN(n15804) );
  NAND2_X1 U15600 ( .A1(n15804), .A2(n13757), .ZN(n13569) );
  NAND2_X1 U15601 ( .A1(n15799), .A2(n15800), .ZN(n15784) );
  NOR2_X1 U15602 ( .A1(n13572), .A2(n13571), .ZN(n13591) );
  AOI22_X1 U15603 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13576) );
  AOI22_X1 U15604 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13575) );
  AOI22_X1 U15605 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13574) );
  AOI22_X1 U15606 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13573) );
  NAND4_X1 U15607 ( .A1(n13576), .A2(n13575), .A3(n13574), .A4(n13573), .ZN(
        n13582) );
  AOI22_X1 U15608 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13580) );
  AOI22_X1 U15609 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U15610 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13578) );
  AOI22_X1 U15611 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13577) );
  NAND4_X1 U15612 ( .A1(n13580), .A2(n13579), .A3(n13578), .A4(n13577), .ZN(
        n13581) );
  OR2_X1 U15613 ( .A1(n13582), .A2(n13581), .ZN(n13590) );
  XNOR2_X1 U15614 ( .A(n13591), .B(n13590), .ZN(n13587) );
  INV_X1 U15615 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13584) );
  AOI21_X1 U15616 ( .B1(n13584), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13585) );
  AOI21_X1 U15617 ( .B1(n13276), .B2(P1_EAX_REG_24__SCAN_IN), .A(n13585), .ZN(
        n13586) );
  OAI21_X1 U15618 ( .B1(n13587), .B2(n13694), .A(n13586), .ZN(n13589) );
  XNOR2_X1 U15619 ( .A(n13606), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15790) );
  NAND2_X1 U15620 ( .A1(n15790), .A2(n13757), .ZN(n13588) );
  NAND2_X1 U15621 ( .A1(n13589), .A2(n13588), .ZN(n15786) );
  NAND2_X1 U15622 ( .A1(n13591), .A2(n13590), .ZN(n13624) );
  AOI22_X1 U15623 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13595) );
  AOI22_X1 U15624 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U15625 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13593) );
  AOI22_X1 U15626 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13592) );
  NAND4_X1 U15627 ( .A1(n13595), .A2(n13594), .A3(n13593), .A4(n13592), .ZN(
        n13601) );
  AOI22_X1 U15628 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13599) );
  AOI22_X1 U15629 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U15630 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13597) );
  AOI22_X1 U15631 ( .A1(n11037), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13596) );
  NAND4_X1 U15632 ( .A1(n13599), .A2(n13598), .A3(n13597), .A4(n13596), .ZN(
        n13600) );
  NOR2_X1 U15633 ( .A1(n13601), .A2(n13600), .ZN(n13625) );
  XNOR2_X1 U15634 ( .A(n13624), .B(n13625), .ZN(n13605) );
  NAND2_X1 U15635 ( .A1(n13234), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13602) );
  NAND2_X1 U15636 ( .A1(n11099), .A2(n13602), .ZN(n13603) );
  AOI21_X1 U15637 ( .B1(n13276), .B2(P1_EAX_REG_25__SCAN_IN), .A(n13603), .ZN(
        n13604) );
  OAI21_X1 U15638 ( .B1(n13605), .B2(n13694), .A(n13604), .ZN(n13612) );
  INV_X1 U15639 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U15640 ( .A1(n13609), .A2(n13608), .ZN(n13610) );
  NAND2_X1 U15641 ( .A1(n13631), .A2(n13610), .ZN(n16076) );
  AOI22_X1 U15642 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13617) );
  AOI22_X1 U15643 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13616) );
  AOI22_X1 U15644 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13615) );
  AOI22_X1 U15645 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13614) );
  NAND4_X1 U15646 ( .A1(n13617), .A2(n13616), .A3(n13615), .A4(n13614), .ZN(
        n13623) );
  AOI22_X1 U15647 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13621) );
  AOI22_X1 U15648 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13620) );
  AOI22_X1 U15649 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13619) );
  AOI22_X1 U15650 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13618) );
  NAND4_X1 U15651 ( .A1(n13621), .A2(n13620), .A3(n13619), .A4(n13618), .ZN(
        n13622) );
  OR2_X1 U15652 ( .A1(n13623), .A2(n13622), .ZN(n13649) );
  NOR2_X1 U15653 ( .A1(n13625), .A2(n13624), .ZN(n13650) );
  XOR2_X1 U15654 ( .A(n13649), .B(n13650), .Z(n13626) );
  NAND2_X1 U15655 ( .A1(n13626), .A2(n13718), .ZN(n13630) );
  INV_X1 U15656 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13627) );
  AOI21_X1 U15657 ( .B1(n13627), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13628) );
  AOI21_X1 U15658 ( .B1(n13276), .B2(P1_EAX_REG_26__SCAN_IN), .A(n13628), .ZN(
        n13629) );
  XNOR2_X1 U15659 ( .A(n13631), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15763) );
  INV_X1 U15660 ( .A(n13631), .ZN(n13632) );
  NAND2_X1 U15661 ( .A1(n13632), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13634) );
  INV_X1 U15662 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13633) );
  NAND2_X1 U15663 ( .A1(n13634), .A2(n13633), .ZN(n13635) );
  NAND2_X1 U15664 ( .A1(n13673), .A2(n13635), .ZN(n16060) );
  AOI22_X1 U15665 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13641) );
  AOI22_X1 U15666 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13680), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U15667 ( .A1(n13699), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13639) );
  AOI22_X1 U15668 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13638) );
  NAND4_X1 U15669 ( .A1(n13641), .A2(n13640), .A3(n13639), .A4(n13638), .ZN(
        n13648) );
  AOI22_X1 U15670 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13646) );
  AOI22_X1 U15671 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13645) );
  AOI22_X1 U15672 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13644) );
  AOI22_X1 U15673 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13643) );
  NAND4_X1 U15674 ( .A1(n13646), .A2(n13645), .A3(n13644), .A4(n13643), .ZN(
        n13647) );
  NOR2_X1 U15675 ( .A1(n13648), .A2(n13647), .ZN(n13667) );
  NAND2_X1 U15676 ( .A1(n13650), .A2(n13649), .ZN(n13666) );
  XNOR2_X1 U15677 ( .A(n13667), .B(n13666), .ZN(n13653) );
  AOI21_X1 U15678 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n13234), .A(
        n13757), .ZN(n13652) );
  NAND2_X1 U15679 ( .A1(n13725), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n13651) );
  OAI211_X1 U15680 ( .C1(n13653), .C2(n13694), .A(n13652), .B(n13651), .ZN(
        n13654) );
  OAI21_X1 U15681 ( .B1(n11099), .B2(n16060), .A(n13654), .ZN(n15751) );
  AOI22_X1 U15682 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U15683 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13657) );
  AOI22_X1 U15684 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13656) );
  AOI22_X1 U15685 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13655) );
  NAND4_X1 U15686 ( .A1(n13658), .A2(n13657), .A3(n13656), .A4(n13655), .ZN(
        n13665) );
  AOI22_X1 U15687 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U15688 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13662) );
  AOI22_X1 U15689 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U15690 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13660) );
  NAND4_X1 U15691 ( .A1(n13663), .A2(n13662), .A3(n13661), .A4(n13660), .ZN(
        n13664) );
  OR2_X1 U15692 ( .A1(n13665), .A2(n13664), .ZN(n13678) );
  NOR2_X1 U15693 ( .A1(n13667), .A2(n13666), .ZN(n13679) );
  XOR2_X1 U15694 ( .A(n13678), .B(n13679), .Z(n13668) );
  NAND2_X1 U15695 ( .A1(n13668), .A2(n13718), .ZN(n13672) );
  INV_X1 U15696 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13669) );
  AOI21_X1 U15697 ( .B1(n13669), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13670) );
  AOI21_X1 U15698 ( .B1(n13276), .B2(P1_EAX_REG_28__SCAN_IN), .A(n13670), .ZN(
        n13671) );
  XNOR2_X1 U15699 ( .A(n13673), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15739) );
  INV_X1 U15700 ( .A(n13673), .ZN(n13674) );
  NAND2_X1 U15701 ( .A1(n13674), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13676) );
  INV_X1 U15702 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U15703 ( .A1(n13676), .A2(n13675), .ZN(n13677) );
  NAND2_X1 U15704 ( .A1(n13760), .A2(n13677), .ZN(n16040) );
  NAND2_X1 U15705 ( .A1(n13679), .A2(n13678), .ZN(n13697) );
  AOI22_X1 U15706 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13685) );
  AOI22_X1 U15707 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12054), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13684) );
  AOI22_X1 U15708 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13683) );
  AOI22_X1 U15709 ( .A1(n13681), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13682) );
  NAND4_X1 U15710 ( .A1(n13685), .A2(n13684), .A3(n13683), .A4(n13682), .ZN(
        n13691) );
  AOI22_X1 U15711 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13689) );
  AOI22_X1 U15712 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U15713 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13687) );
  AOI22_X1 U15714 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13686) );
  NAND4_X1 U15715 ( .A1(n13689), .A2(n13688), .A3(n13687), .A4(n13686), .ZN(
        n13690) );
  NOR2_X1 U15716 ( .A1(n13691), .A2(n13690), .ZN(n13698) );
  XNOR2_X1 U15717 ( .A(n13697), .B(n13698), .ZN(n13695) );
  AOI21_X1 U15718 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n13234), .A(
        n13757), .ZN(n13693) );
  NAND2_X1 U15719 ( .A1(n13725), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n13692) );
  OAI211_X1 U15720 ( .C1(n13695), .C2(n13694), .A(n13693), .B(n13692), .ZN(
        n13696) );
  OAI21_X1 U15721 ( .B1(n11099), .B2(n16040), .A(n13696), .ZN(n15726) );
  NOR2_X1 U15722 ( .A1(n13698), .A2(n13697), .ZN(n13717) );
  AOI22_X1 U15723 ( .A1(n13700), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13699), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13706) );
  AOI22_X1 U15724 ( .A1(n13701), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13681), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U15725 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13702), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U15726 ( .A1(n13659), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13703) );
  NAND4_X1 U15727 ( .A1(n13706), .A2(n13705), .A3(n13704), .A4(n13703), .ZN(
        n13715) );
  AOI22_X1 U15728 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U15729 ( .A1(n12054), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11037), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13712) );
  AOI22_X1 U15730 ( .A1(n13680), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13711) );
  AOI22_X1 U15731 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13710) );
  NAND4_X1 U15732 ( .A1(n13713), .A2(n13712), .A3(n13711), .A4(n13710), .ZN(
        n13714) );
  NOR2_X1 U15733 ( .A1(n13715), .A2(n13714), .ZN(n13716) );
  XNOR2_X1 U15734 ( .A(n13717), .B(n13716), .ZN(n13719) );
  NAND2_X1 U15735 ( .A1(n13719), .A2(n13718), .ZN(n13723) );
  INV_X1 U15736 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15717) );
  AOI21_X1 U15737 ( .B1(n15717), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13720) );
  AOI21_X1 U15738 ( .B1(n13276), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13720), .ZN(
        n13722) );
  XNOR2_X1 U15739 ( .A(n13760), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16025) );
  AOI22_X1 U15740 ( .A1(n13725), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13724), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13726) );
  INV_X1 U15741 ( .A(n13726), .ZN(n13727) );
  INV_X1 U15742 ( .A(n21455), .ZN(n21866) );
  OAI21_X1 U15743 ( .B1(n13730), .B2(n21866), .A(n13729), .ZN(n13731) );
  NAND2_X1 U15744 ( .A1(n13731), .A2(n15389), .ZN(n13732) );
  INV_X1 U15745 ( .A(n14683), .ZN(n15956) );
  NAND4_X1 U15746 ( .A1(n11930), .A2(n13734), .A3(n15956), .A4(n14689), .ZN(
        n14513) );
  NOR2_X1 U15747 ( .A1(n14513), .A2(n13735), .ZN(n13736) );
  AND2_X1 U15748 ( .A1(n16015), .A2(n15956), .ZN(n13738) );
  NAND2_X1 U15749 ( .A1(n13790), .A2(n13738), .ZN(n13756) );
  NOR4_X1 U15750 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13742) );
  NOR4_X1 U15751 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13741) );
  NOR4_X1 U15752 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13740) );
  NOR4_X1 U15753 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13739) );
  AND4_X1 U15754 ( .A1(n13742), .A2(n13741), .A3(n13740), .A4(n13739), .ZN(
        n13747) );
  NOR4_X1 U15755 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13745) );
  NOR4_X1 U15756 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13744) );
  NOR4_X1 U15757 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13743) );
  INV_X1 U15758 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20068) );
  AND4_X1 U15759 ( .A1(n13745), .A2(n13744), .A3(n13743), .A4(n20068), .ZN(
        n13746) );
  NAND2_X1 U15760 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  NOR3_X1 U15761 ( .A1(n16019), .A2(n14789), .A3(n13749), .ZN(n13750) );
  AOI22_X1 U15762 ( .A1(n16008), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16019), .ZN(n13751) );
  INV_X1 U15763 ( .A(n13751), .ZN(n13754) );
  NAND3_X1 U15764 ( .A1(n16015), .A2(n13752), .A3(n14789), .ZN(n15955) );
  INV_X1 U15765 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20308) );
  NOR2_X1 U15766 ( .A1(n15955), .A2(n20308), .ZN(n13753) );
  NOR2_X1 U15767 ( .A1(n13754), .A2(n13753), .ZN(n13755) );
  NAND2_X1 U15768 ( .A1(n13756), .A2(n13755), .ZN(P1_U2873) );
  AND2_X1 U15769 ( .A1(n12208), .A2(n14396), .ZN(n14298) );
  NAND2_X1 U15770 ( .A1(n14298), .A2(n15390), .ZN(n14295) );
  NAND2_X1 U15771 ( .A1(n17154), .A2(n13234), .ZN(n21451) );
  INV_X1 U15772 ( .A(n21451), .ZN(n21838) );
  AOI21_X1 U15773 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21838), .A(n21832), 
        .ZN(n17150) );
  AOI21_X1 U15774 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n13757), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n13758) );
  NOR2_X1 U15775 ( .A1(n17150), .A2(n13758), .ZN(n13759) );
  INV_X2 U15776 ( .A(n21596), .ZN(n21639) );
  INV_X1 U15777 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13780) );
  INV_X1 U15778 ( .A(n15150), .ZN(n13762) );
  NAND2_X1 U15779 ( .A1(n13762), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13763) );
  NAND2_X1 U15780 ( .A1(n13790), .A2(n21771), .ZN(n13788) );
  MUX2_X1 U15781 ( .A(n13765), .B(n13764), .S(n15722), .Z(n13768) );
  AOI22_X1 U15782 ( .A1(n13766), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14512), .ZN(n13767) );
  XNOR2_X1 U15783 ( .A(n13768), .B(n13767), .ZN(n16161) );
  AND2_X1 U15784 ( .A1(n14749), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13776) );
  INV_X1 U15785 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n22050) );
  NAND2_X1 U15786 ( .A1(n21455), .A2(n22050), .ZN(n17143) );
  NAND4_X1 U15787 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_4__SCAN_IN), .ZN(n21684)
         );
  INV_X1 U15788 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21696) );
  NOR2_X1 U15789 ( .A1(n21684), .A2(n21696), .ZN(n21698) );
  NAND2_X1 U15790 ( .A1(n21698), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n21708) );
  INV_X1 U15791 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21717) );
  NOR2_X1 U15792 ( .A1(n21708), .A2(n21717), .ZN(n21719) );
  NAND2_X1 U15793 ( .A1(n21719), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n21733) );
  INV_X1 U15794 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21743) );
  NOR2_X1 U15795 ( .A1(n21733), .A2(n21743), .ZN(n15159) );
  NAND2_X1 U15796 ( .A1(n15159), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15255) );
  NOR2_X1 U15797 ( .A1(n21720), .A2(n15255), .ZN(n15335) );
  NAND2_X1 U15798 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n15823) );
  NAND2_X1 U15799 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15824) );
  INV_X1 U15800 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21775) );
  INV_X1 U15801 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21757) );
  NOR4_X1 U15802 ( .A1(n15823), .A2(n15824), .A3(n21775), .A4(n21757), .ZN(
        n21791) );
  NAND2_X1 U15803 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n15859) );
  INV_X1 U15804 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20082) );
  NOR2_X1 U15805 ( .A1(n15859), .A2(n20082), .ZN(n15822) );
  NAND4_X1 U15806 ( .A1(n15335), .A2(n21791), .A3(n15822), .A4(
        P1_REIP_REG_20__SCAN_IN), .ZN(n21782) );
  INV_X1 U15807 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21807) );
  NOR2_X1 U15808 ( .A1(n21782), .A2(n21807), .ZN(n21805) );
  AND4_X1 U15809 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_25__SCAN_IN), .A4(P1_REIP_REG_26__SCAN_IN), .ZN(n13770) );
  AND2_X1 U15810 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n13771) );
  NAND2_X1 U15811 ( .A1(n15752), .A2(n13771), .ZN(n15729) );
  NAND2_X1 U15812 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n13772) );
  NOR2_X1 U15813 ( .A1(n15729), .A2(n13772), .ZN(n13781) );
  OR2_X1 U15814 ( .A1(n13773), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13778) );
  INV_X1 U15815 ( .A(n13778), .ZN(n13774) );
  NOR2_X1 U15816 ( .A1(n13781), .A2(n21804), .ZN(n15721) );
  INV_X1 U15817 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n22021) );
  INV_X1 U15818 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15897) );
  INV_X1 U15819 ( .A(n13775), .ZN(n13777) );
  NOR2_X1 U15820 ( .A1(n13777), .A2(n13776), .ZN(n13779) );
  OAI22_X1 U15821 ( .A1(n21820), .A2(n13780), .B1(n15897), .B2(n21765), .ZN(
        n13784) );
  INV_X1 U15822 ( .A(n13781), .ZN(n13782) );
  NOR3_X1 U15823 ( .A1(n13782), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21732), 
        .ZN(n13783) );
  AOI211_X1 U15824 ( .C1(n15721), .C2(P1_REIP_REG_31__SCAN_IN), .A(n13784), 
        .B(n13783), .ZN(n13785) );
  OAI21_X1 U15825 ( .B1(n16161), .B2(n21812), .A(n13785), .ZN(n13786) );
  INV_X1 U15826 ( .A(n13786), .ZN(n13787) );
  NAND2_X1 U15827 ( .A1(n13788), .A2(n13787), .ZN(P1_U2809) );
  NOR2_X2 U15828 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22077) );
  NAND2_X1 U15829 ( .A1(n13790), .A2(n20236), .ZN(n13817) );
  NAND2_X1 U15830 ( .A1(n20231), .A2(n16174), .ZN(n13791) );
  AND2_X1 U15831 ( .A1(n20231), .A2(n13792), .ZN(n16035) );
  INV_X1 U15832 ( .A(n13800), .ZN(n13797) );
  NOR2_X1 U15833 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13794) );
  XNOR2_X1 U15834 ( .A(n12179), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13799) );
  INV_X1 U15835 ( .A(n13799), .ZN(n13793) );
  INV_X1 U15836 ( .A(n13795), .ZN(n13796) );
  NAND2_X1 U15837 ( .A1(n13797), .A2(n13796), .ZN(n13806) );
  NAND2_X1 U15838 ( .A1(n20231), .A2(n13798), .ZN(n13801) );
  NAND3_X1 U15839 ( .A1(n13800), .A2(n13799), .A3(n13801), .ZN(n13805) );
  INV_X1 U15840 ( .A(n13801), .ZN(n13802) );
  AOI211_X1 U15841 ( .C1(n11209), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16034), .B(n13802), .ZN(n13803) );
  NAND3_X1 U15842 ( .A1(n13806), .A2(n13805), .A3(n13804), .ZN(n16172) );
  INV_X1 U15843 ( .A(n16172), .ZN(n13809) );
  NAND2_X1 U15844 ( .A1(n13809), .A2(n20237), .ZN(n13816) );
  NAND2_X1 U15845 ( .A1(n22043), .A2(n13810), .ZN(n21454) );
  NAND2_X1 U15846 ( .A1(n21454), .A2(n21832), .ZN(n13811) );
  NAND2_X1 U15847 ( .A1(n21832), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17149) );
  NAND2_X1 U15848 ( .A1(n22050), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13812) );
  NAND2_X1 U15849 ( .A1(n17149), .A2(n13812), .ZN(n14528) );
  INV_X1 U15850 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n17264) );
  NOR2_X1 U15851 ( .A1(n21596), .A2(n17264), .ZN(n16163) );
  AOI21_X1 U15852 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16163), .ZN(n13813) );
  OAI21_X1 U15853 ( .B1(n20240), .B2(n15150), .A(n13813), .ZN(n13814) );
  INV_X1 U15854 ( .A(n13814), .ZN(n13815) );
  NAND3_X1 U15855 ( .A1(n13817), .A2(n13816), .A3(n13815), .ZN(P1_U2968) );
  INV_X1 U15856 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20983) );
  NAND2_X1 U15857 ( .A1(n13818), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n18168) );
  NAND2_X1 U15858 ( .A1(n13819), .A2(n21250), .ZN(n18169) );
  INV_X1 U15859 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n18178) );
  XNOR2_X1 U15860 ( .A(n20983), .B(n13820), .ZN(n13831) );
  NAND2_X1 U15861 ( .A1(n13831), .A2(n18261), .ZN(n13830) );
  NAND3_X1 U15862 ( .A1(n21244), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13821) );
  XOR2_X1 U15863 ( .A(n13821), .B(n20983), .Z(n13838) );
  NAND3_X1 U15864 ( .A1(n21245), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13822) );
  NAND2_X1 U15865 ( .A1(n10995), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n13845) );
  INV_X1 U15866 ( .A(n13845), .ZN(n13828) );
  OR2_X1 U15867 ( .A1(n13823), .A2(n18132), .ZN(n18174) );
  XNOR2_X1 U15868 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13826) );
  NOR2_X1 U15869 ( .A1(n13825), .A2(n13824), .ZN(n18173) );
  OAI22_X1 U15870 ( .A1(n18174), .A2(n13826), .B1(n18173), .B2(n20763), .ZN(
        n13827) );
  AOI211_X1 U15871 ( .C1(n20580), .C2(n18171), .A(n13828), .B(n13827), .ZN(
        n13829) );
  NAND2_X1 U15872 ( .A1(n13831), .A2(n21373), .ZN(n13849) );
  NAND2_X1 U15873 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13832) );
  NOR2_X1 U15874 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13832), .ZN(
        n13837) );
  INV_X1 U15875 ( .A(n13833), .ZN(n18113) );
  AOI22_X1 U15876 ( .A1(n13835), .A2(n18048), .B1(n18113), .B2(n13834), .ZN(
        n21207) );
  NOR4_X1 U15877 ( .A1(n21207), .A2(n18138), .A3(n21206), .A4(n13836), .ZN(
        n21243) );
  AOI22_X1 U15878 ( .A1(n21293), .A2(n13838), .B1(n13837), .B2(n21243), .ZN(
        n13843) );
  NOR2_X1 U15879 ( .A1(n13839), .A2(n18178), .ZN(n13841) );
  OAI211_X1 U15880 ( .C1(n21285), .C2(n18167), .A(n13841), .B(n13840), .ZN(
        n21259) );
  NAND3_X1 U15881 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21336), .A3(
        n21259), .ZN(n13842) );
  OAI211_X1 U15882 ( .C1(n13844), .C2(n21268), .A(n13843), .B(n13842), .ZN(
        n13847) );
  OAI21_X1 U15883 ( .B1(n21275), .B2(n20983), .A(n13845), .ZN(n13846) );
  NAND2_X1 U15884 ( .A1(n13849), .A2(n13848), .ZN(P3_U2831) );
  NAND2_X1 U15885 ( .A1(n13853), .A2(n13852), .ZN(n13856) );
  INV_X1 U15886 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n18789) );
  NOR2_X1 U15887 ( .A1(n14857), .A2(n18789), .ZN(n13854) );
  XNOR2_X1 U15888 ( .A(n13856), .B(n13854), .ZN(n18801) );
  OR2_X1 U15889 ( .A1(n18801), .A2(n16730), .ZN(n13855) );
  NAND2_X1 U15890 ( .A1(n13855), .A2(n11275), .ZN(n16578) );
  NOR3_X1 U15891 ( .A1(n18801), .A2(n16730), .A3(n11275), .ZN(n16577) );
  NOR2_X1 U15892 ( .A1(n13856), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13857) );
  MUX2_X1 U15893 ( .A(n13858), .B(n13857), .S(n11028), .Z(n16286) );
  NAND2_X1 U15894 ( .A1(n16286), .A2(n13859), .ZN(n13860) );
  NAND2_X1 U15895 ( .A1(n13862), .A2(n13861), .ZN(n13879) );
  AOI21_X1 U15896 ( .B1(n13885), .B2(n16334), .A(n13863), .ZN(n13874) );
  INV_X1 U15897 ( .A(n13863), .ZN(n13867) );
  OAI21_X1 U15898 ( .B1(n16334), .B2(n13865), .A(n13864), .ZN(n13866) );
  OAI21_X1 U15899 ( .B1(n16334), .B2(n13867), .A(n13866), .ZN(n13868) );
  NAND2_X1 U15900 ( .A1(n13868), .A2(n19872), .ZN(n13872) );
  OAI21_X1 U15901 ( .B1(n13870), .B2(n13869), .A(n16287), .ZN(n13871) );
  NAND2_X1 U15902 ( .A1(n13872), .A2(n13871), .ZN(n13873) );
  OAI21_X1 U15903 ( .B1(n13875), .B2(n13874), .A(n13873), .ZN(n13877) );
  NAND2_X1 U15904 ( .A1(n13877), .A2(n13876), .ZN(n13878) );
  NAND2_X1 U15905 ( .A1(n13879), .A2(n13878), .ZN(n13883) );
  INV_X1 U15906 ( .A(n13880), .ZN(n13881) );
  AOI21_X1 U15907 ( .B1(n16287), .B2(n13881), .A(n13886), .ZN(n13882) );
  NAND2_X1 U15908 ( .A1(n13883), .A2(n13882), .ZN(n13884) );
  MUX2_X1 U15909 ( .A(n13884), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n14841), .Z(n13890) );
  NAND2_X1 U15910 ( .A1(n14647), .A2(n16334), .ZN(n14421) );
  NOR2_X1 U15911 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n17541) );
  NAND2_X2 U15912 ( .A1(n13888), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n17572) );
  NOR2_X2 U15913 ( .A1(n17572), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n17563) );
  AOI21_X1 U15914 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n17541), .A(n17563), 
        .ZN(n21893) );
  OAI22_X1 U15915 ( .A1(n14421), .A2(n21893), .B1(n16334), .B2(n14638), .ZN(
        n13889) );
  NAND2_X1 U15916 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n18899) );
  NAND3_X1 U15917 ( .A1(n13889), .A2(n18899), .A3(n15031), .ZN(n13911) );
  AOI21_X1 U15918 ( .B1(n13890), .B2(n19872), .A(n19671), .ZN(n13891) );
  NAND2_X1 U15919 ( .A1(n14421), .A2(n13891), .ZN(n13909) );
  NOR2_X1 U15920 ( .A1(n13892), .A2(n14638), .ZN(n13904) );
  INV_X1 U15921 ( .A(n18899), .ZN(n21883) );
  NOR2_X1 U15922 ( .A1(n21883), .A2(n21893), .ZN(n14661) );
  NAND2_X1 U15923 ( .A1(n11013), .A2(n14197), .ZN(n13894) );
  NAND2_X1 U15924 ( .A1(n14292), .A2(n13894), .ZN(n13898) );
  INV_X1 U15925 ( .A(n12687), .ZN(n14575) );
  OR2_X1 U15926 ( .A1(n13895), .A2(n14575), .ZN(n13896) );
  NAND2_X1 U15927 ( .A1(n13896), .A2(n14663), .ZN(n14192) );
  NAND3_X1 U15928 ( .A1(n13898), .A2(n13897), .A3(n14192), .ZN(n14190) );
  INV_X1 U15929 ( .A(n14190), .ZN(n13902) );
  OAI211_X1 U15930 ( .C1(n19872), .C2(n14575), .A(n13900), .B(n14197), .ZN(
        n13901) );
  NAND3_X1 U15931 ( .A1(n13902), .A2(n11007), .A3(n13901), .ZN(n13903) );
  AOI21_X1 U15932 ( .B1(n13904), .B2(n14661), .A(n13903), .ZN(n14286) );
  INV_X1 U15933 ( .A(n13904), .ZN(n13905) );
  INV_X1 U15934 ( .A(n17101), .ZN(n18894) );
  OAI22_X1 U15935 ( .A1(n13905), .A2(n21883), .B1(n18894), .B2(n13015), .ZN(
        n13906) );
  NAND2_X1 U15936 ( .A1(n13906), .A2(n16334), .ZN(n13907) );
  NAND2_X1 U15937 ( .A1(n13911), .A2(n13910), .ZN(n13912) );
  INV_X1 U15938 ( .A(n14637), .ZN(n13913) );
  NAND2_X1 U15939 ( .A1(n14170), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n13936) );
  NOR2_X1 U15940 ( .A1(n13931), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13915) );
  AOI22_X1 U15941 ( .A1(n15509), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15508), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13919) );
  AOI22_X1 U15942 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U15943 ( .A1(n15512), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13917) );
  NAND2_X1 U15944 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13916) );
  AND4_X1 U15945 ( .A1(n13919), .A2(n13918), .A3(n13917), .A4(n13916), .ZN(
        n13930) );
  INV_X1 U15946 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13922) );
  NAND2_X1 U15947 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13921) );
  NAND2_X1 U15948 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13920) );
  OAI211_X1 U15949 ( .C1(n13922), .C2(n15484), .A(n13921), .B(n13920), .ZN(
        n13928) );
  NAND2_X1 U15950 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n13926) );
  AOI22_X1 U15951 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U15952 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13924) );
  NAND2_X1 U15953 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13923) );
  NAND4_X1 U15954 ( .A1(n13926), .A2(n13925), .A3(n13924), .A4(n13923), .ZN(
        n13927) );
  NOR2_X1 U15955 ( .A1(n13928), .A2(n13927), .ZN(n13929) );
  NAND2_X1 U15956 ( .A1(n14171), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n13933) );
  NAND2_X1 U15957 ( .A1(n14155), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13932) );
  OAI211_X1 U15958 ( .C1(n14145), .C2(n15083), .A(n13933), .B(n13932), .ZN(
        n13934) );
  INV_X1 U15959 ( .A(n13934), .ZN(n13935) );
  NAND2_X1 U15960 ( .A1(n13936), .A2(n13935), .ZN(n16982) );
  NAND2_X1 U15961 ( .A1(n14170), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n13942) );
  NAND2_X1 U15962 ( .A1(n14171), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n13938) );
  NAND2_X1 U15963 ( .A1(n14155), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13937) );
  OAI211_X1 U15964 ( .C1(n14145), .C2(n13939), .A(n13938), .B(n13937), .ZN(
        n13940) );
  INV_X1 U15965 ( .A(n13940), .ZN(n13941) );
  NAND2_X1 U15966 ( .A1(n16334), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13946) );
  INV_X1 U15967 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n17501) );
  NAND2_X1 U15968 ( .A1(n13948), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13945) );
  INV_X1 U15969 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n17514) );
  INV_X1 U15970 ( .A(n13943), .ZN(n13944) );
  NAND3_X1 U15971 ( .A1(n13946), .A2(n13945), .A3(n13944), .ZN(n14561) );
  INV_X1 U15972 ( .A(n12688), .ZN(n14572) );
  NAND2_X1 U15973 ( .A1(n14572), .A2(n14155), .ZN(n13961) );
  MUX2_X1 U15974 ( .A(n12687), .B(n17485), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13947) );
  INV_X1 U15975 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n18464) );
  NAND2_X1 U15976 ( .A1(n13948), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U15977 ( .A1(n13949), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n14155), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U15978 ( .A1(n13951), .A2(n13950), .ZN(n13956) );
  OR2_X1 U15979 ( .A1(n13952), .A2(n14145), .ZN(n13955) );
  NAND2_X1 U15980 ( .A1(n12688), .A2(n12687), .ZN(n13953) );
  MUX2_X1 U15981 ( .A(n13953), .B(n19488), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13954) );
  NAND2_X1 U15982 ( .A1(n13955), .A2(n13954), .ZN(n14558) );
  NOR2_X1 U15983 ( .A1(n14559), .A2(n14558), .ZN(n13959) );
  NOR2_X1 U15984 ( .A1(n13957), .A2(n13956), .ZN(n13958) );
  NOR2_X2 U15985 ( .A1(n13959), .A2(n13958), .ZN(n13966) );
  NAND2_X1 U15986 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13960) );
  OAI211_X1 U15987 ( .C1(n14145), .C2(n13962), .A(n13961), .B(n13960), .ZN(
        n13965) );
  XNOR2_X1 U15988 ( .A(n13966), .B(n13965), .ZN(n14562) );
  NAND2_X1 U15989 ( .A1(n14170), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13964) );
  AOI22_X1 U15990 ( .A1(n14171), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n14155), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13963) );
  NAND2_X1 U15991 ( .A1(n13964), .A2(n13963), .ZN(n14563) );
  NOR2_X1 U15992 ( .A1(n14562), .A2(n14563), .ZN(n13968) );
  NOR2_X1 U15993 ( .A1(n13966), .A2(n13965), .ZN(n13967) );
  INV_X1 U15994 ( .A(n14145), .ZN(n13970) );
  AOI22_X1 U15995 ( .A1(n13970), .A2(n13969), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14155), .ZN(n13973) );
  NAND2_X1 U15996 ( .A1(n14170), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13972) );
  AOI22_X1 U15997 ( .A1(n14171), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13971) );
  NAND2_X1 U15998 ( .A1(n14170), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n13975) );
  AOI22_X1 U15999 ( .A1(n14171), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n14155), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13974) );
  OAI211_X1 U16000 ( .C1(n13976), .C2(n14145), .A(n13975), .B(n13974), .ZN(
        n15218) );
  OR2_X1 U16001 ( .A1(n14145), .A2(n13977), .ZN(n13978) );
  NAND2_X1 U16002 ( .A1(n14170), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n13981) );
  AOI22_X1 U16003 ( .A1(n14171), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n14155), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13980) );
  NAND2_X1 U16004 ( .A1(n13981), .A2(n13980), .ZN(n15241) );
  NAND2_X1 U16005 ( .A1(n15242), .A2(n15241), .ZN(n13983) );
  OR2_X1 U16006 ( .A1(n14145), .A2(n16730), .ZN(n13982) );
  NAND2_X1 U16007 ( .A1(n14170), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n13985) );
  AOI22_X1 U16008 ( .A1(n14171), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n14155), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13984) );
  NAND2_X1 U16009 ( .A1(n13985), .A2(n13984), .ZN(n15304) );
  NAND2_X1 U16010 ( .A1(n15305), .A2(n15304), .ZN(n15306) );
  INV_X1 U16011 ( .A(n15499), .ZN(n14079) );
  INV_X1 U16012 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13987) );
  INV_X1 U16013 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13986) );
  OAI22_X1 U16014 ( .A1(n14079), .A2(n13987), .B1(n14078), .B2(n13986), .ZN(
        n13990) );
  OAI22_X1 U16015 ( .A1(n14057), .A2(n13988), .B1(n14462), .B2(n15531), .ZN(
        n13989) );
  NOR2_X1 U16016 ( .A1(n13990), .A2(n13989), .ZN(n14005) );
  INV_X1 U16017 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13993) );
  NAND2_X1 U16018 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13992) );
  NAND2_X1 U16019 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13991) );
  OAI211_X1 U16020 ( .C1(n13993), .C2(n15484), .A(n13992), .B(n13991), .ZN(
        n13994) );
  INV_X1 U16021 ( .A(n13994), .ZN(n14004) );
  NAND2_X1 U16022 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13998) );
  AOI22_X1 U16023 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13997) );
  AOI22_X1 U16024 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13996) );
  NAND2_X1 U16025 ( .A1(n15509), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13995) );
  AND4_X1 U16026 ( .A1(n13998), .A2(n13997), .A3(n13996), .A4(n13995), .ZN(
        n14003) );
  INV_X1 U16027 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15524) );
  NAND2_X1 U16028 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14000) );
  NAND2_X1 U16029 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13999) );
  OAI211_X1 U16030 ( .C1(n15524), .C2(n14081), .A(n14000), .B(n13999), .ZN(
        n14001) );
  INV_X1 U16031 ( .A(n14001), .ZN(n14002) );
  NAND4_X1 U16032 ( .A1(n14005), .A2(n14004), .A3(n14003), .A4(n14002), .ZN(
        n14599) );
  INV_X1 U16033 ( .A(n14599), .ZN(n14008) );
  NAND2_X1 U16034 ( .A1(n14170), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n14007) );
  AOI22_X1 U16035 ( .A1(n14171), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n14155), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14006) );
  OAI211_X1 U16036 ( .C1(n14008), .C2(n14145), .A(n14007), .B(n14006), .ZN(
        n14009) );
  INV_X1 U16037 ( .A(n14009), .ZN(n18531) );
  NOR2_X2 U16038 ( .A1(n15306), .A2(n18531), .ZN(n18530) );
  AOI22_X1 U16039 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n15508), .B1(
        n15509), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14013) );
  AOI22_X1 U16040 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14012) );
  AOI22_X1 U16041 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12802), .B1(
        n15512), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14011) );
  NAND2_X1 U16042 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14010) );
  AND4_X1 U16043 ( .A1(n14013), .A2(n14012), .A3(n14011), .A4(n14010), .ZN(
        n14025) );
  INV_X1 U16044 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14016) );
  NAND2_X1 U16045 ( .A1(n15504), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14015) );
  NAND2_X1 U16046 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n14014) );
  OAI211_X1 U16047 ( .C1(n14017), .C2(n14016), .A(n14015), .B(n14014), .ZN(
        n14023) );
  NAND2_X1 U16048 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n14021) );
  AOI22_X1 U16049 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12479), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14020) );
  AOI22_X1 U16050 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n15498), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14019) );
  NAND2_X1 U16051 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14018) );
  NAND4_X1 U16052 ( .A1(n14021), .A2(n14020), .A3(n14019), .A4(n14018), .ZN(
        n14022) );
  NOR2_X1 U16053 ( .A1(n14023), .A2(n14022), .ZN(n14024) );
  NAND2_X1 U16054 ( .A1(n14170), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n14027) );
  AOI22_X1 U16055 ( .A1(n14171), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n14155), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14026) );
  OAI211_X1 U16056 ( .C1(n14862), .C2(n14145), .A(n14027), .B(n14026), .ZN(
        n17035) );
  NAND2_X1 U16057 ( .A1(n18530), .A2(n17035), .ZN(n18555) );
  NAND2_X1 U16058 ( .A1(n14170), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n14053) );
  INV_X1 U16059 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14028) );
  OAI22_X1 U16060 ( .A1(n14082), .A2(n14029), .B1(n14078), .B2(n14028), .ZN(
        n14033) );
  INV_X1 U16061 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14030) );
  OAI22_X1 U16062 ( .A1(n14057), .A2(n14031), .B1(n14081), .B2(n14030), .ZN(
        n14032) );
  NOR2_X1 U16063 ( .A1(n14033), .A2(n14032), .ZN(n14048) );
  INV_X1 U16064 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14036) );
  NAND2_X1 U16065 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14035) );
  NAND2_X1 U16066 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n14034) );
  OAI211_X1 U16067 ( .C1(n14036), .C2(n15484), .A(n14035), .B(n14034), .ZN(
        n14037) );
  INV_X1 U16068 ( .A(n14037), .ZN(n14047) );
  NAND2_X1 U16069 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n14041) );
  AOI22_X1 U16070 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U16071 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14039) );
  NAND2_X1 U16072 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n14038) );
  AND4_X1 U16073 ( .A1(n14041), .A2(n14040), .A3(n14039), .A4(n14038), .ZN(
        n14046) );
  NAND2_X1 U16074 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14043) );
  NAND2_X1 U16075 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14042) );
  OAI211_X1 U16076 ( .C1(n15574), .C2(n14462), .A(n14043), .B(n14042), .ZN(
        n14044) );
  INV_X1 U16077 ( .A(n14044), .ZN(n14045) );
  NAND4_X1 U16078 ( .A1(n14048), .A2(n14047), .A3(n14046), .A4(n14045), .ZN(
        n14899) );
  INV_X1 U16079 ( .A(n14899), .ZN(n14902) );
  NAND2_X1 U16080 ( .A1(n14171), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n14050) );
  NAND2_X1 U16081 ( .A1(n14155), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14049) );
  OAI211_X1 U16082 ( .C1(n14145), .C2(n14902), .A(n14050), .B(n14049), .ZN(
        n14051) );
  INV_X1 U16083 ( .A(n14051), .ZN(n14052) );
  INV_X1 U16084 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14054) );
  OAI22_X1 U16085 ( .A1(n14082), .A2(n14055), .B1(n14078), .B2(n14054), .ZN(
        n14059) );
  INV_X1 U16086 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15590) );
  OAI22_X1 U16087 ( .A1(n14057), .A2(n14056), .B1(n14081), .B2(n15590), .ZN(
        n14058) );
  NOR2_X1 U16088 ( .A1(n14059), .A2(n14058), .ZN(n14074) );
  INV_X1 U16089 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14062) );
  NAND2_X1 U16090 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14061) );
  NAND2_X1 U16091 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14060) );
  OAI211_X1 U16092 ( .C1(n14062), .C2(n15484), .A(n14061), .B(n14060), .ZN(
        n14063) );
  INV_X1 U16093 ( .A(n14063), .ZN(n14073) );
  NAND2_X1 U16094 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n14067) );
  AOI22_X1 U16095 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14066) );
  AOI22_X1 U16096 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14065) );
  NAND2_X1 U16097 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14064) );
  AND4_X1 U16098 ( .A1(n14067), .A2(n14066), .A3(n14065), .A4(n14064), .ZN(
        n14072) );
  NAND2_X1 U16099 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n14069) );
  NAND2_X1 U16100 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14068) );
  OAI211_X1 U16101 ( .C1(n15597), .C2(n14462), .A(n14069), .B(n14068), .ZN(
        n14070) );
  INV_X1 U16102 ( .A(n14070), .ZN(n14071) );
  NAND4_X1 U16103 ( .A1(n14074), .A2(n14073), .A3(n14072), .A4(n14071), .ZN(
        n14898) );
  INV_X1 U16104 ( .A(n14898), .ZN(n14901) );
  NAND2_X1 U16105 ( .A1(n14170), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n14076) );
  AOI22_X1 U16106 ( .A1(n14171), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n14155), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14075) );
  OAI211_X1 U16107 ( .C1(n14901), .C2(n14145), .A(n14076), .B(n14075), .ZN(
        n17018) );
  NAND2_X1 U16108 ( .A1(n17017), .A2(n17018), .ZN(n16998) );
  NAND2_X1 U16109 ( .A1(n14170), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n14106) );
  INV_X1 U16110 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14077) );
  OAI22_X1 U16111 ( .A1(n14080), .A2(n14079), .B1(n14078), .B2(n14077), .ZN(
        n14085) );
  INV_X1 U16112 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14083) );
  INV_X1 U16113 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15611) );
  OAI22_X1 U16114 ( .A1(n14083), .A2(n14082), .B1(n14081), .B2(n15611), .ZN(
        n14084) );
  NOR2_X1 U16115 ( .A1(n14085), .A2(n14084), .ZN(n14101) );
  INV_X1 U16116 ( .A(n14086), .ZN(n14114) );
  INV_X1 U16117 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14089) );
  NAND2_X1 U16118 ( .A1(n15504), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14088) );
  NAND2_X1 U16119 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14087) );
  OAI211_X1 U16120 ( .C1(n14114), .C2(n14089), .A(n14088), .B(n14087), .ZN(
        n14090) );
  INV_X1 U16121 ( .A(n14090), .ZN(n14100) );
  NAND2_X1 U16122 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14094) );
  AOI22_X1 U16123 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n15498), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14093) );
  AOI22_X1 U16124 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12479), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14092) );
  NAND2_X1 U16125 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14091) );
  AND4_X1 U16126 ( .A1(n14094), .A2(n14093), .A3(n14092), .A4(n14091), .ZN(
        n14099) );
  NAND2_X1 U16127 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n14096) );
  NAND2_X1 U16128 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14095) );
  OAI211_X1 U16129 ( .C1(n14462), .C2(n15618), .A(n14096), .B(n14095), .ZN(
        n14097) );
  INV_X1 U16130 ( .A(n14097), .ZN(n14098) );
  NAND4_X1 U16131 ( .A1(n14101), .A2(n14100), .A3(n14099), .A4(n14098), .ZN(
        n14930) );
  NAND2_X1 U16132 ( .A1(n14171), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n14103) );
  NAND2_X1 U16133 ( .A1(n14155), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14102) );
  OAI211_X1 U16134 ( .C1(n14145), .C2(n11435), .A(n14103), .B(n14102), .ZN(
        n14104) );
  INV_X1 U16135 ( .A(n14104), .ZN(n14105) );
  NAND2_X1 U16136 ( .A1(n16982), .A2(n16981), .ZN(n16984) );
  NAND2_X1 U16137 ( .A1(n14170), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n14127) );
  AOI22_X1 U16138 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n15499), .B1(
        n15508), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14110) );
  AOI22_X1 U16139 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14109) );
  AOI22_X1 U16140 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12802), .B1(
        n15512), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14108) );
  NAND2_X1 U16141 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14107) );
  AND4_X1 U16142 ( .A1(n14110), .A2(n14109), .A3(n14108), .A4(n14107), .ZN(
        n14122) );
  INV_X1 U16143 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14113) );
  NAND2_X1 U16144 ( .A1(n15504), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14112) );
  NAND2_X1 U16145 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n14111) );
  OAI211_X1 U16146 ( .C1(n14114), .C2(n14113), .A(n14112), .B(n14111), .ZN(
        n14120) );
  NAND2_X1 U16147 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14118) );
  AOI22_X1 U16148 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12479), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U16149 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n15498), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14116) );
  NAND2_X1 U16150 ( .A1(n15509), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14115) );
  NAND4_X1 U16151 ( .A1(n14118), .A2(n14117), .A3(n14116), .A4(n14115), .ZN(
        n14119) );
  NOR2_X1 U16152 ( .A1(n14120), .A2(n14119), .ZN(n14121) );
  NAND2_X1 U16153 ( .A1(n14171), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n14124) );
  NAND2_X1 U16154 ( .A1(n14155), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14123) );
  OAI211_X1 U16155 ( .C1(n14145), .C2(n15141), .A(n14124), .B(n14123), .ZN(
        n14125) );
  INV_X1 U16156 ( .A(n14125), .ZN(n14126) );
  NAND2_X1 U16157 ( .A1(n14170), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U16158 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n15509), .B1(
        n15508), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14131) );
  AOI22_X1 U16159 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14130) );
  AOI22_X1 U16160 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12802), .B1(
        n15512), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14129) );
  NAND2_X1 U16161 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14128) );
  AND4_X1 U16162 ( .A1(n14131), .A2(n14130), .A3(n14129), .A4(n14128), .ZN(
        n14142) );
  INV_X1 U16163 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14134) );
  NAND2_X1 U16164 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14133) );
  NAND2_X1 U16165 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n14132) );
  OAI211_X1 U16166 ( .C1(n14134), .C2(n15484), .A(n14133), .B(n14132), .ZN(
        n14140) );
  NAND2_X1 U16167 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n14138) );
  AOI22_X1 U16168 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U16169 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n15498), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14136) );
  NAND2_X1 U16170 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14135) );
  NAND4_X1 U16171 ( .A1(n14138), .A2(n14137), .A3(n14136), .A4(n14135), .ZN(
        n14139) );
  NOR2_X1 U16172 ( .A1(n14140), .A2(n14139), .ZN(n14141) );
  NAND2_X1 U16173 ( .A1(n14171), .A2(P2_EAX_REG_15__SCAN_IN), .ZN(n14144) );
  NAND2_X1 U16174 ( .A1(n14155), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14143) );
  OAI211_X1 U16175 ( .C1(n14145), .C2(n15230), .A(n14144), .B(n14143), .ZN(
        n14146) );
  INV_X1 U16176 ( .A(n14146), .ZN(n14147) );
  AOI22_X1 U16177 ( .A1(n14171), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n14155), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14149) );
  OAI21_X1 U16178 ( .B1(n14150), .B2(n17557), .A(n14149), .ZN(n16348) );
  AOI22_X1 U16179 ( .A1(n14171), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n14155), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14151) );
  OAI21_X1 U16180 ( .B1(n14150), .B2(n13091), .A(n14151), .ZN(n16554) );
  INV_X1 U16181 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14153) );
  OAI22_X1 U16182 ( .A1(n14167), .A2(n14153), .B1(n16907), .B2(n14152), .ZN(
        n14154) );
  AOI21_X1 U16183 ( .B1(n14170), .B2(P2_REIP_REG_18__SCAN_IN), .A(n14154), 
        .ZN(n16902) );
  INV_X1 U16184 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16548) );
  OAI22_X1 U16185 ( .A1(n14167), .A2(n16548), .B1(n16888), .B2(n14152), .ZN(
        n14156) );
  AOI21_X1 U16186 ( .B1(n14170), .B2(P2_REIP_REG_19__SCAN_IN), .A(n14156), 
        .ZN(n16546) );
  NOR2_X4 U16187 ( .A1(n16901), .A2(n16546), .ZN(n16877) );
  AOI22_X1 U16188 ( .A1(n14171), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n14155), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14157) );
  OAI21_X1 U16189 ( .B1(n14150), .B2(n14158), .A(n14157), .ZN(n16876) );
  INV_X1 U16190 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n16541) );
  OAI22_X1 U16191 ( .A1(n14167), .A2(n16541), .B1(n16861), .B2(n14152), .ZN(
        n14159) );
  AOI21_X1 U16192 ( .B1(n14170), .B2(P2_REIP_REG_21__SCAN_IN), .A(n14159), 
        .ZN(n16540) );
  INV_X1 U16193 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14160) );
  OAI22_X1 U16194 ( .A1(n14167), .A2(n14160), .B1(n16847), .B2(n14152), .ZN(
        n14161) );
  AOI21_X1 U16195 ( .B1(n14170), .B2(P2_REIP_REG_22__SCAN_IN), .A(n14161), 
        .ZN(n16841) );
  INV_X1 U16196 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16530) );
  OAI22_X1 U16197 ( .A1(n14167), .A2(n16530), .B1(n16833), .B2(n14152), .ZN(
        n14162) );
  AOI21_X1 U16198 ( .B1(n14170), .B2(P2_REIP_REG_23__SCAN_IN), .A(n14162), 
        .ZN(n16527) );
  AOI22_X1 U16199 ( .A1(n14171), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n14155), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14163) );
  OAI21_X1 U16200 ( .B1(n14150), .B2(n17565), .A(n14163), .ZN(n16521) );
  AND2_X2 U16201 ( .A1(n16529), .A2(n16521), .ZN(n16512) );
  AOI22_X1 U16202 ( .A1(n14171), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n14155), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14164) );
  OAI21_X1 U16203 ( .B1(n14150), .B2(n18717), .A(n14164), .ZN(n16511) );
  AOI22_X1 U16204 ( .A1(n14171), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n14155), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14165) );
  OAI21_X1 U16205 ( .B1(n14150), .B2(n17566), .A(n14165), .ZN(n16505) );
  INV_X1 U16206 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n16495) );
  INV_X1 U16207 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16764) );
  OAI22_X1 U16208 ( .A1(n14167), .A2(n16495), .B1(n16764), .B2(n14152), .ZN(
        n14166) );
  AOI21_X1 U16209 ( .B1(n14170), .B2(P2_REIP_REG_27__SCAN_IN), .A(n14166), 
        .ZN(n16500) );
  INV_X1 U16210 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n16485) );
  OAI22_X1 U16211 ( .A1(n14167), .A2(n16485), .B1(n16595), .B2(n14152), .ZN(
        n14168) );
  AOI21_X1 U16212 ( .B1(n14170), .B2(P2_REIP_REG_28__SCAN_IN), .A(n14168), 
        .ZN(n16491) );
  AOI22_X1 U16213 ( .A1(n14171), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n14155), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14169) );
  OAI21_X1 U16214 ( .B1(n14150), .B2(n18764), .A(n14169), .ZN(n16475) );
  AOI222_X1 U16215 ( .A1(n14170), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14155), .C1(n14171), .C2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n15703) );
  AOI222_X1 U16216 ( .A1(n14170), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n14171), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n14155), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14172) );
  AND2_X1 U16217 ( .A1(n14639), .A2(n16334), .ZN(n14175) );
  NOR2_X1 U16218 ( .A1(n14648), .A2(n14175), .ZN(n14176) );
  INV_X1 U16219 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n18790) );
  NAND2_X1 U16220 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14178) );
  AOI22_X1 U16221 ( .A1(n14180), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n14177) );
  OAI211_X1 U16222 ( .C1(n12743), .C2(n18790), .A(n14178), .B(n14177), .ZN(
        n15706) );
  INV_X1 U16223 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n17568) );
  NAND2_X1 U16224 ( .A1(n14179), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14182) );
  AOI22_X1 U16225 ( .A1(n14180), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14181) );
  OAI211_X1 U16226 ( .C1(n12743), .C2(n17568), .A(n14182), .B(n14181), .ZN(
        n14183) );
  INV_X1 U16227 ( .A(n14185), .ZN(n14186) );
  NAND2_X1 U16228 ( .A1(n14260), .A2(n14186), .ZN(n14621) );
  AOI21_X1 U16229 ( .B1(n14621), .B2(n15667), .A(n14187), .ZN(n14188) );
  INV_X1 U16230 ( .A(n18849), .ZN(n14189) );
  INV_X1 U16231 ( .A(n14640), .ZN(n14191) );
  NAND2_X1 U16232 ( .A1(n14614), .A2(n14192), .ZN(n14194) );
  NAND2_X1 U16233 ( .A1(n14194), .A2(n14193), .ZN(n14205) );
  INV_X1 U16234 ( .A(n14195), .ZN(n14204) );
  OR2_X1 U16235 ( .A1(n16279), .A2(n19671), .ZN(n14203) );
  INV_X1 U16236 ( .A(n16279), .ZN(n14268) );
  OAI21_X1 U16237 ( .B1(n14196), .B2(n14268), .A(n19720), .ZN(n14198) );
  NAND2_X1 U16238 ( .A1(n14198), .A2(n14197), .ZN(n14201) );
  INV_X1 U16239 ( .A(n14199), .ZN(n14200) );
  NAND2_X1 U16240 ( .A1(n14201), .A2(n14200), .ZN(n14202) );
  NAND4_X1 U16241 ( .A1(n14205), .A2(n14204), .A3(n14203), .A4(n14202), .ZN(
        n14623) );
  NOR2_X1 U16242 ( .A1(n14623), .A2(n14453), .ZN(n14206) );
  NAND2_X1 U16243 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16762) );
  NAND2_X1 U16244 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14207) );
  NOR2_X1 U16245 ( .A1(n16762), .A2(n14207), .ZN(n14232) );
  INV_X1 U16246 ( .A(n16797), .ZN(n14225) );
  NOR2_X1 U16247 ( .A1(n17065), .A2(n17048), .ZN(n18864) );
  NAND2_X1 U16248 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18864), .ZN(
        n14213) );
  NOR2_X1 U16249 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18864), .ZN(
        n18876) );
  NOR4_X1 U16250 ( .A1(n18876), .A2(n18860), .A3(n18844), .A4(n15215), .ZN(
        n15239) );
  NAND2_X1 U16251 ( .A1(n18847), .A2(n15239), .ZN(n15237) );
  INV_X1 U16252 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15310) );
  NOR2_X1 U16253 ( .A1(n15310), .A2(n14208), .ZN(n14211) );
  NAND2_X1 U16254 ( .A1(n16921), .A2(n11476), .ZN(n14217) );
  INV_X1 U16255 ( .A(n14216), .ZN(n14209) );
  NAND2_X1 U16256 ( .A1(n16908), .A2(n14209), .ZN(n16848) );
  NAND2_X1 U16257 ( .A1(n14223), .A2(n16818), .ZN(n14210) );
  OR2_X1 U16258 ( .A1(n16848), .A2(n14210), .ZN(n16824) );
  NAND2_X1 U16259 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15239), .ZN(
        n14214) );
  INV_X1 U16260 ( .A(n14211), .ZN(n18828) );
  NOR2_X1 U16261 ( .A1(n14214), .A2(n18828), .ZN(n14212) );
  NAND2_X1 U16262 ( .A1(n14234), .A2(n18848), .ZN(n18804) );
  OAI21_X1 U16263 ( .B1(n16912), .B2(n14212), .A(n18804), .ZN(n16870) );
  INV_X1 U16264 ( .A(n14213), .ZN(n18877) );
  INV_X1 U16265 ( .A(n14214), .ZN(n15309) );
  NAND2_X1 U16266 ( .A1(n18877), .A2(n15309), .ZN(n15238) );
  NOR2_X1 U16267 ( .A1(n18828), .A2(n15238), .ZN(n16868) );
  NOR2_X1 U16268 ( .A1(n16917), .A2(n16868), .ZN(n14215) );
  OR2_X1 U16269 ( .A1(n16870), .A2(n14215), .ZN(n17043) );
  OR2_X1 U16270 ( .A1(n14217), .A2(n14216), .ZN(n14218) );
  AND2_X1 U16271 ( .A1(n18808), .A2(n14218), .ZN(n14219) );
  NOR2_X1 U16272 ( .A1(n17043), .A2(n14219), .ZN(n16862) );
  INV_X1 U16273 ( .A(n14223), .ZN(n16830) );
  NAND2_X1 U16274 ( .A1(n18808), .A2(n16830), .ZN(n14220) );
  AND2_X1 U16275 ( .A1(n16862), .A2(n14220), .ZN(n16819) );
  NAND2_X1 U16276 ( .A1(n16824), .A2(n16819), .ZN(n16814) );
  AOI21_X1 U16277 ( .B1(n18808), .B2(n14225), .A(n16814), .ZN(n16782) );
  OAI21_X1 U16278 ( .B1(n17047), .B2(n14232), .A(n16782), .ZN(n16753) );
  INV_X1 U16279 ( .A(n16753), .ZN(n14222) );
  INV_X1 U16280 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14221) );
  NOR2_X1 U16281 ( .A1(n14222), .A2(n14221), .ZN(n14228) );
  NAND2_X1 U16282 ( .A1(n14223), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14224) );
  NOR2_X1 U16283 ( .A1(n16809), .A2(n14225), .ZN(n16766) );
  NAND3_X1 U16284 ( .A1(n16766), .A2(n14232), .A3(n14221), .ZN(n14226) );
  NAND2_X1 U16285 ( .A1(n16675), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n16569) );
  NAND2_X1 U16286 ( .A1(n14226), .A2(n16569), .ZN(n14227) );
  NOR2_X1 U16287 ( .A1(n14228), .A2(n14227), .ZN(n14229) );
  OAI211_X1 U16288 ( .C1(n16341), .C2(n18870), .A(n14230), .B(n14229), .ZN(
        n14231) );
  INV_X1 U16289 ( .A(n14231), .ZN(n14235) );
  INV_X1 U16290 ( .A(n14233), .ZN(n14644) );
  INV_X1 U16291 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22396) );
  NOR3_X1 U16292 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n22396), .ZN(n14237) );
  NOR4_X1 U16293 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14236) );
  NAND4_X1 U16294 ( .A1(n14789), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n14237), .A4(
        n14236), .ZN(U214) );
  NOR4_X1 U16295 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n14241) );
  NOR4_X1 U16296 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n14240) );
  NOR4_X1 U16297 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n14239) );
  NOR4_X1 U16298 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n14238) );
  NAND4_X1 U16299 ( .A1(n14241), .A2(n14240), .A3(n14239), .A4(n14238), .ZN(
        n14246) );
  NOR4_X1 U16300 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n14244) );
  NOR4_X1 U16301 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n14243) );
  NOR4_X1 U16302 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n14242) );
  INV_X1 U16303 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n17544) );
  NAND4_X1 U16304 ( .A1(n14244), .A2(n14243), .A3(n14242), .A4(n17544), .ZN(
        n14245) );
  NOR2_X1 U16305 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14248) );
  NOR4_X1 U16306 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14247) );
  NAND4_X1 U16307 ( .A1(n14248), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14247), .ZN(n14249) );
  OR2_X1 U16308 ( .A1(n14361), .A2(n14249), .ZN(n20243) );
  INV_X2 U16309 ( .A(U214), .ZN(n20296) );
  AOI211_X1 U16310 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n20591), .A(n20597), .B(
        n20764), .ZN(n14259) );
  AOI22_X1 U16311 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n14250) );
  INV_X1 U16312 ( .A(n14250), .ZN(n14258) );
  NAND2_X1 U16313 ( .A1(n14251), .A2(n20576), .ZN(n14256) );
  INV_X1 U16314 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18433) );
  NOR2_X1 U16315 ( .A1(n20719), .A2(n14252), .ZN(n20614) );
  INV_X1 U16316 ( .A(n20614), .ZN(n20606) );
  OAI211_X1 U16317 ( .C1(n18195), .C2(n14254), .A(n20741), .B(n14253), .ZN(
        n14255) );
  OAI221_X1 U16318 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n14256), .C1(n18433), 
        .C2(n20606), .A(n14255), .ZN(n14257) );
  OR4_X1 U16319 ( .A1(n10995), .A2(n14259), .A3(n14258), .A4(n14257), .ZN(
        P3_U2654) );
  INV_X1 U16320 ( .A(n18907), .ZN(n18904) );
  NOR2_X1 U16321 ( .A1(n14292), .A2(n18904), .ZN(n14423) );
  INV_X1 U16322 ( .A(n14638), .ZN(n14636) );
  NAND2_X1 U16323 ( .A1(n14423), .A2(n14636), .ZN(n18485) );
  INV_X1 U16324 ( .A(n18485), .ZN(n18472) );
  INV_X1 U16325 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14263) );
  INV_X1 U16326 ( .A(n14260), .ZN(n14261) );
  NOR2_X1 U16327 ( .A1(n19532), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14265) );
  INV_X1 U16328 ( .A(n14265), .ZN(n14262) );
  OAI211_X1 U16329 ( .C1(n18472), .C2(n14263), .A(n14278), .B(n14262), .ZN(
        P2_U2814) );
  INV_X1 U16330 ( .A(n17388), .ZN(n14267) );
  OAI21_X1 U16331 ( .B1(n14265), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n14267), 
        .ZN(n14266) );
  OAI21_X1 U16332 ( .B1(n14268), .B2(n14267), .A(n14266), .ZN(P2_U3612) );
  OAI21_X1 U16333 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14270), .A(
        n14269), .ZN(n17046) );
  INV_X1 U16334 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18473) );
  AOI21_X1 U16335 ( .B1(n17065), .B2(n14272), .A(n14271), .ZN(n17051) );
  INV_X1 U16336 ( .A(n17051), .ZN(n14274) );
  OR2_X1 U16337 ( .A1(n17459), .A2(n18473), .ZN(n14273) );
  NAND2_X1 U16338 ( .A1(n16328), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n17054) );
  OAI211_X1 U16339 ( .C1(n17463), .C2(n14274), .A(n14273), .B(n17054), .ZN(
        n14275) );
  AOI21_X1 U16340 ( .B1(n17453), .B2(n18473), .A(n14275), .ZN(n14277) );
  NAND2_X1 U16341 ( .A1(n18470), .A2(n17474), .ZN(n14276) );
  OAI211_X1 U16342 ( .C1(n17046), .C2(n17461), .A(n14277), .B(n14276), .ZN(
        P2_U3013) );
  INV_X1 U16343 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14283) );
  NOR2_X1 U16344 ( .A1(n14278), .A2(n21883), .ZN(n14279) );
  OR2_X1 U16345 ( .A1(n14382), .A2(n14279), .ZN(n14341) );
  INV_X1 U16346 ( .A(n14279), .ZN(n14280) );
  NOR2_X2 U16347 ( .A1(n14280), .A2(n15667), .ZN(n14367) );
  INV_X1 U16348 ( .A(n14367), .ZN(n14282) );
  AOI22_X1 U16349 ( .A1(n15695), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14361), .ZN(n19368) );
  INV_X1 U16350 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n14281) );
  OAI222_X1 U16351 ( .A1(n14283), .A2(n14341), .B1(n14282), .B2(n19368), .C1(
        n14281), .C2(n14319), .ZN(P2_U2982) );
  INV_X1 U16352 ( .A(n14292), .ZN(n14284) );
  NAND2_X1 U16353 ( .A1(n14284), .A2(n14661), .ZN(n14288) );
  NAND2_X1 U16354 ( .A1(n14647), .A2(n14640), .ZN(n14568) );
  AND2_X1 U16355 ( .A1(n16279), .A2(n18899), .ZN(n14634) );
  NAND3_X1 U16356 ( .A1(n14639), .A2(n14634), .A3(n14636), .ZN(n14285) );
  AND3_X1 U16357 ( .A1(n14286), .A2(n14568), .A3(n14285), .ZN(n14287) );
  INV_X1 U16358 ( .A(n14647), .ZN(n14641) );
  NAND2_X1 U16359 ( .A1(n14641), .A2(n14648), .ZN(n14409) );
  OAI211_X1 U16360 ( .C1(n14421), .C2(n14288), .A(n14287), .B(n14409), .ZN(
        n14655) );
  NAND2_X1 U16361 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18912), .ZN(n14290) );
  NOR2_X1 U16362 ( .A1(n14841), .A2(n14840), .ZN(n17099) );
  INV_X1 U16363 ( .A(n17099), .ZN(n18893) );
  OAI21_X1 U16364 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n19472), .A(n18893), 
        .ZN(n14289) );
  AOI22_X1 U16365 ( .A1(n14655), .A2(n18907), .B1(n14290), .B2(n14289), .ZN(
        n17073) );
  INV_X1 U16366 ( .A(n17073), .ZN(n14294) );
  NOR2_X1 U16367 ( .A1(n14292), .A2(n14291), .ZN(n14649) );
  NOR2_X1 U16368 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17387) );
  NAND4_X1 U16369 ( .A1(n14294), .A2(n15667), .A3(n14649), .A4(n17387), .ZN(
        n14293) );
  OAI21_X1 U16370 ( .B1(n14656), .B2(n14294), .A(n14293), .ZN(P2_U3595) );
  INV_X1 U16371 ( .A(n14295), .ZN(n14297) );
  INV_X1 U16372 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22397) );
  NOR2_X1 U16373 ( .A1(n22043), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14386) );
  INV_X1 U16374 ( .A(n14386), .ZN(n14296) );
  OAI211_X1 U16375 ( .C1(n14297), .C2(n22397), .A(n14740), .B(n14296), .ZN(
        P1_U2801) );
  OAI22_X1 U16376 ( .A1(n14298), .A2(n11103), .B1(n15876), .B2(n15389), .ZN(
        n14391) );
  NOR2_X1 U16377 ( .A1(n14391), .A2(n21844), .ZN(n14300) );
  INV_X1 U16378 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n17172) );
  NAND3_X1 U16379 ( .A1(n17081), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13234), 
        .ZN(n14299) );
  OAI21_X1 U16380 ( .B1(n14300), .B2(n17172), .A(n14299), .ZN(P1_U2803) );
  INV_X1 U16381 ( .A(n17474), .ZN(n17449) );
  OAI21_X1 U16382 ( .B1(n17470), .B2(n14301), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14302) );
  OAI21_X1 U16383 ( .B1(n18805), .B2(n17449), .A(n14302), .ZN(n14310) );
  INV_X1 U16384 ( .A(n14303), .ZN(n14305) );
  NAND2_X1 U16385 ( .A1(n18453), .A2(n17048), .ZN(n14304) );
  NAND2_X1 U16386 ( .A1(n14305), .A2(n14304), .ZN(n18803) );
  NOR2_X1 U16387 ( .A1(n17461), .A2(n18803), .ZN(n14309) );
  OAI21_X1 U16388 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14307), .A(
        n14306), .ZN(n18811) );
  NAND2_X1 U16389 ( .A1(n16675), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18809) );
  OAI21_X1 U16390 ( .B1(n17463), .B2(n18811), .A(n18809), .ZN(n14308) );
  OR3_X1 U16391 ( .A1(n14310), .A2(n14309), .A3(n14308), .ZN(P2_U3014) );
  INV_X1 U16392 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17532) );
  NAND2_X1 U16393 ( .A1(n14383), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14313) );
  NAND2_X1 U16394 ( .A1(n15697), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14312) );
  INV_X1 U16395 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20265) );
  OR2_X1 U16396 ( .A1(n14361), .A2(n20265), .ZN(n14311) );
  NAND2_X1 U16397 ( .A1(n14312), .A2(n14311), .ZN(n19384) );
  NAND2_X1 U16398 ( .A1(n14367), .A2(n19384), .ZN(n14314) );
  OAI211_X1 U16399 ( .C1(n17532), .C2(n14319), .A(n14313), .B(n14314), .ZN(
        P2_U2977) );
  INV_X1 U16400 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14498) );
  NAND2_X1 U16401 ( .A1(n14383), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14315) );
  OAI211_X1 U16402 ( .C1(n14498), .C2(n14319), .A(n14315), .B(n14314), .ZN(
        P2_U2962) );
  AOI22_X1 U16403 ( .A1(n14383), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n14382), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U16404 ( .A1(n15695), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15697), .ZN(n14855) );
  INV_X1 U16405 ( .A(n14855), .ZN(n19607) );
  NAND2_X1 U16406 ( .A1(n14367), .A2(n19607), .ZN(n14344) );
  NAND2_X1 U16407 ( .A1(n14316), .A2(n14344), .ZN(P2_U2957) );
  AOI22_X1 U16408 ( .A1(n14383), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n14369), .ZN(n14318) );
  AOI22_X1 U16409 ( .A1(n15695), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n15697), .ZN(n19380) );
  INV_X1 U16410 ( .A(n19380), .ZN(n14317) );
  NAND2_X1 U16411 ( .A1(n14367), .A2(n14317), .ZN(n14376) );
  NAND2_X1 U16412 ( .A1(n14318), .A2(n14376), .ZN(P2_U2978) );
  AOI22_X1 U16413 ( .A1(n14383), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n14382), .ZN(n14320) );
  INV_X1 U16414 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20253) );
  INV_X1 U16415 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20829) );
  AOI22_X1 U16416 ( .A1(n15695), .A2(n20253), .B1(n20829), .B2(n15697), .ZN(
        n19662) );
  NAND2_X1 U16417 ( .A1(n14367), .A2(n19662), .ZN(n14321) );
  NAND2_X1 U16418 ( .A1(n14320), .A2(n14321), .ZN(P2_U2971) );
  AOI22_X1 U16419 ( .A1(n14383), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n14382), .ZN(n14322) );
  NAND2_X1 U16420 ( .A1(n14322), .A2(n14321), .ZN(P2_U2956) );
  AOI22_X1 U16421 ( .A1(n14383), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n14382), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n14324) );
  AOI22_X1 U16422 ( .A1(n15695), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15697), .ZN(n19816) );
  INV_X1 U16423 ( .A(n19816), .ZN(n14323) );
  NAND2_X1 U16424 ( .A1(n14367), .A2(n14323), .ZN(n14350) );
  NAND2_X1 U16425 ( .A1(n14324), .A2(n14350), .ZN(P2_U2953) );
  AOI22_X1 U16426 ( .A1(n14383), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n14382), .ZN(n14325) );
  OAI22_X1 U16427 ( .A1(n15697), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15695), .ZN(n15029) );
  INV_X1 U16428 ( .A(n15029), .ZN(n19762) );
  NAND2_X1 U16429 ( .A1(n14367), .A2(n19762), .ZN(n14342) );
  NAND2_X1 U16430 ( .A1(n14325), .A2(n14342), .ZN(P2_U2954) );
  AOI22_X1 U16431 ( .A1(n14383), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n14382), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n14326) );
  AOI22_X1 U16432 ( .A1(n15695), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15697), .ZN(n19394) );
  INV_X1 U16433 ( .A(n19394), .ZN(n16533) );
  NAND2_X1 U16434 ( .A1(n14367), .A2(n16533), .ZN(n14355) );
  NAND2_X1 U16435 ( .A1(n14326), .A2(n14355), .ZN(P2_U2974) );
  AOI22_X1 U16436 ( .A1(n14383), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n14382), .ZN(n14328) );
  AOI22_X1 U16437 ( .A1(n15695), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15697), .ZN(n19870) );
  INV_X1 U16438 ( .A(n19870), .ZN(n14327) );
  NAND2_X1 U16439 ( .A1(n14367), .A2(n14327), .ZN(n14374) );
  NAND2_X1 U16440 ( .A1(n14328), .A2(n14374), .ZN(P2_U2952) );
  XNOR2_X1 U16441 ( .A(n14330), .B(n14329), .ZN(n18868) );
  INV_X1 U16442 ( .A(n14331), .ZN(n18863) );
  OAI21_X1 U16443 ( .B1(n14334), .B2(n14333), .A(n14332), .ZN(n14335) );
  XOR2_X1 U16444 ( .A(n14335), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(
        n18880) );
  NOR2_X1 U16445 ( .A1(n18848), .A2(n14336), .ZN(n18862) );
  OAI21_X1 U16446 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16293), .ZN(n16373) );
  NOR2_X1 U16447 ( .A1(n17479), .A2(n16373), .ZN(n14337) );
  AOI211_X1 U16448 ( .C1(n17470), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n18862), .B(n14337), .ZN(n14338) );
  OAI21_X1 U16449 ( .B1(n18880), .B2(n17463), .A(n14338), .ZN(n14339) );
  AOI21_X1 U16450 ( .B1(n18863), .B2(n17474), .A(n14339), .ZN(n14340) );
  OAI21_X1 U16451 ( .B1(n17461), .B2(n18868), .A(n14340), .ZN(P2_U3012) );
  INV_X2 U16452 ( .A(n14341), .ZN(n14383) );
  AOI22_X1 U16453 ( .A1(n14383), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n14382), .ZN(n14343) );
  NAND2_X1 U16454 ( .A1(n14343), .A2(n14342), .ZN(P2_U2969) );
  AOI22_X1 U16455 ( .A1(n14383), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n14382), .ZN(n14345) );
  NAND2_X1 U16456 ( .A1(n14345), .A2(n14344), .ZN(P2_U2972) );
  AOI22_X1 U16457 ( .A1(n14383), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n14382), .ZN(n14347) );
  AOI22_X1 U16458 ( .A1(n15695), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n14361), .ZN(n19391) );
  INV_X1 U16459 ( .A(n19391), .ZN(n14346) );
  NAND2_X1 U16460 ( .A1(n14367), .A2(n14346), .ZN(n14359) );
  NAND2_X1 U16461 ( .A1(n14347), .A2(n14359), .ZN(P2_U2960) );
  AOI22_X1 U16462 ( .A1(n14383), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n14382), .ZN(n14349) );
  AOI22_X1 U16463 ( .A1(n15695), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n15697), .ZN(n19371) );
  INV_X1 U16464 ( .A(n19371), .ZN(n14348) );
  NAND2_X1 U16465 ( .A1(n14367), .A2(n14348), .ZN(n14380) );
  NAND2_X1 U16466 ( .A1(n14349), .A2(n14380), .ZN(P2_U2981) );
  AOI22_X1 U16467 ( .A1(n14383), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n14382), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n14351) );
  NAND2_X1 U16468 ( .A1(n14351), .A2(n14350), .ZN(P2_U2968) );
  AOI22_X1 U16469 ( .A1(n14383), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n14382), .ZN(n14353) );
  AOI22_X1 U16470 ( .A1(n15695), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15697), .ZN(n19719) );
  INV_X1 U16471 ( .A(n19719), .ZN(n14352) );
  NAND2_X1 U16472 ( .A1(n14367), .A2(n14352), .ZN(n14364) );
  NAND2_X1 U16473 ( .A1(n14353), .A2(n14364), .ZN(P2_U2970) );
  AOI22_X1 U16474 ( .A1(n14383), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n14369), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n14354) );
  INV_X1 U16475 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20257) );
  INV_X1 U16476 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20865) );
  AOI22_X1 U16477 ( .A1(n15695), .A2(n20257), .B1(n20865), .B2(n15697), .ZN(
        n19555) );
  NAND2_X1 U16478 ( .A1(n14367), .A2(n19555), .ZN(n14384) );
  NAND2_X1 U16479 ( .A1(n14354), .A2(n14384), .ZN(P2_U2973) );
  AOI22_X1 U16480 ( .A1(n14383), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n14382), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n14356) );
  NAND2_X1 U16481 ( .A1(n14356), .A2(n14355), .ZN(P2_U2959) );
  AOI22_X1 U16482 ( .A1(n14383), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n14382), .ZN(n14358) );
  INV_X1 U16483 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20263) );
  NOR2_X1 U16484 ( .A1(n14361), .A2(n20263), .ZN(n14357) );
  AOI21_X1 U16485 ( .B1(n14361), .B2(BUF2_REG_9__SCAN_IN), .A(n14357), .ZN(
        n19387) );
  INV_X1 U16486 ( .A(n19387), .ZN(n16517) );
  NAND2_X1 U16487 ( .A1(n14367), .A2(n16517), .ZN(n14372) );
  NAND2_X1 U16488 ( .A1(n14358), .A2(n14372), .ZN(P2_U2976) );
  AOI22_X1 U16489 ( .A1(n14383), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n14382), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n14360) );
  NAND2_X1 U16490 ( .A1(n14360), .A2(n14359), .ZN(P2_U2975) );
  AOI22_X1 U16491 ( .A1(n14383), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n14382), .ZN(n14363) );
  AOI22_X1 U16492 ( .A1(n15695), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n14361), .ZN(n19377) );
  INV_X1 U16493 ( .A(n19377), .ZN(n14362) );
  NAND2_X1 U16494 ( .A1(n14367), .A2(n14362), .ZN(n14370) );
  NAND2_X1 U16495 ( .A1(n14363), .A2(n14370), .ZN(P2_U2964) );
  AOI22_X1 U16496 ( .A1(n14383), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n14382), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n14365) );
  NAND2_X1 U16497 ( .A1(n14365), .A2(n14364), .ZN(P2_U2955) );
  AOI22_X1 U16498 ( .A1(n14383), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n14369), .ZN(n14368) );
  AOI22_X1 U16499 ( .A1(n15695), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n15697), .ZN(n19374) );
  INV_X1 U16500 ( .A(n19374), .ZN(n14366) );
  NAND2_X1 U16501 ( .A1(n14367), .A2(n14366), .ZN(n14378) );
  NAND2_X1 U16502 ( .A1(n14368), .A2(n14378), .ZN(P2_U2980) );
  AOI22_X1 U16503 ( .A1(n14383), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n14369), .ZN(n14371) );
  NAND2_X1 U16504 ( .A1(n14371), .A2(n14370), .ZN(P2_U2979) );
  AOI22_X1 U16505 ( .A1(n14383), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n14382), .ZN(n14373) );
  NAND2_X1 U16506 ( .A1(n14373), .A2(n14372), .ZN(P2_U2961) );
  AOI22_X1 U16507 ( .A1(n14383), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n14382), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U16508 ( .A1(n14375), .A2(n14374), .ZN(P2_U2967) );
  AOI22_X1 U16509 ( .A1(n14383), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n14382), .ZN(n14377) );
  NAND2_X1 U16510 ( .A1(n14377), .A2(n14376), .ZN(P2_U2963) );
  AOI22_X1 U16511 ( .A1(n14383), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n14382), .ZN(n14379) );
  NAND2_X1 U16512 ( .A1(n14379), .A2(n14378), .ZN(P2_U2965) );
  AOI22_X1 U16513 ( .A1(n14383), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n14382), .ZN(n14381) );
  NAND2_X1 U16514 ( .A1(n14381), .A2(n14380), .ZN(P2_U2966) );
  AOI22_X1 U16515 ( .A1(n14383), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n14382), .ZN(n14385) );
  NAND2_X1 U16516 ( .A1(n14385), .A2(n14384), .ZN(P2_U2958) );
  INV_X1 U16517 ( .A(n21453), .ZN(n14388) );
  OAI21_X1 U16518 ( .B1(n14386), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n14388), 
        .ZN(n14387) );
  OAI21_X1 U16519 ( .B1(n14389), .B2(n14388), .A(n14387), .ZN(P1_U3487) );
  NAND2_X1 U16520 ( .A1(n21446), .A2(n21448), .ZN(n14534) );
  AOI21_X1 U16521 ( .B1(n14534), .B2(n21875), .A(n21866), .ZN(n14390) );
  OR2_X1 U16522 ( .A1(n14391), .A2(n14390), .ZN(n17134) );
  AND2_X1 U16523 ( .A1(n17134), .A2(n15390), .ZN(n21824) );
  INV_X1 U16524 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17135) );
  NAND3_X1 U16525 ( .A1(n14392), .A2(n12110), .A3(n11027), .ZN(n14393) );
  NAND2_X1 U16526 ( .A1(n14394), .A2(n14393), .ZN(n14395) );
  NAND2_X1 U16527 ( .A1(n14395), .A2(n14548), .ZN(n14400) );
  INV_X1 U16528 ( .A(n14396), .ZN(n14398) );
  AOI22_X1 U16529 ( .A1(n12208), .A2(n14398), .B1(n14397), .B2(n15389), .ZN(
        n14399) );
  AOI21_X1 U16530 ( .B1(n14400), .B2(n14399), .A(n15956), .ZN(n17136) );
  NAND2_X1 U16531 ( .A1(n21824), .A2(n17136), .ZN(n14401) );
  OAI21_X1 U16532 ( .B1(n21824), .B2(n17135), .A(n14401), .ZN(P1_U3484) );
  NAND2_X1 U16533 ( .A1(n14468), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14402) );
  NOR2_X1 U16534 ( .A1(n19532), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n14403) );
  AOI21_X1 U16535 ( .B1(n14440), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n14403), .ZN(n14404) );
  NAND2_X1 U16536 ( .A1(n16334), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14406) );
  AND4_X1 U16537 ( .A1(n14406), .A2(n19562), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19472), .ZN(n14407) );
  INV_X1 U16538 ( .A(n14453), .ZN(n14408) );
  NAND2_X1 U16539 ( .A1(n14409), .A2(n14408), .ZN(n14410) );
  MUX2_X1 U16540 ( .A(n18805), .B(n14411), .S(n16433), .Z(n14412) );
  OAI21_X1 U16541 ( .B1(n17481), .B2(n16474), .A(n14412), .ZN(P2_U2887) );
  NAND2_X1 U16542 ( .A1(n14440), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14413) );
  NAND2_X1 U16543 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17485), .ZN(
        n19495) );
  NAND2_X1 U16544 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19488), .ZN(
        n19529) );
  NAND2_X1 U16545 ( .A1(n19495), .A2(n19529), .ZN(n19442) );
  NAND2_X1 U16546 ( .A1(n19508), .A2(n19442), .ZN(n19497) );
  NAND2_X1 U16547 ( .A1(n14413), .A2(n19497), .ZN(n14414) );
  NAND2_X1 U16548 ( .A1(n15627), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14430) );
  XNOR2_X1 U16549 ( .A(n14429), .B(n14430), .ZN(n14417) );
  NAND2_X1 U16550 ( .A1(n18470), .A2(n16448), .ZN(n14420) );
  NAND2_X1 U16551 ( .A1(n16433), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n14419) );
  OAI211_X1 U16552 ( .C1(n19420), .C2(n16474), .A(n14420), .B(n14419), .ZN(
        P2_U2886) );
  INV_X1 U16553 ( .A(n14421), .ZN(n14422) );
  NAND2_X1 U16554 ( .A1(n17512), .A2(n16277), .ZN(n14504) );
  NOR2_X1 U16555 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14840), .ZN(n17530) );
  AOI22_X1 U16556 ( .A1(n17530), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14425) );
  OAI21_X1 U16557 ( .B1(n14153), .B2(n14504), .A(n14425), .ZN(P2_U2933) );
  NAND2_X1 U16558 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n14980) );
  XNOR2_X1 U16559 ( .A(n14980), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15090) );
  AOI22_X1 U16560 ( .A1(n14440), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19508), .B2(n15090), .ZN(n14427) );
  NAND2_X1 U16561 ( .A1(n15627), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14445) );
  INV_X1 U16562 ( .A(n14429), .ZN(n17058) );
  NAND2_X1 U16563 ( .A1(n17058), .A2(n14430), .ZN(n14431) );
  NAND2_X1 U16564 ( .A1(n14434), .A2(n14433), .ZN(n14449) );
  INV_X1 U16565 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14436) );
  MUX2_X1 U16566 ( .A(n14436), .B(n14331), .S(n16448), .Z(n14437) );
  OAI21_X1 U16567 ( .B1(n19611), .B2(n16474), .A(n14437), .ZN(P2_U2885) );
  OAI21_X1 U16568 ( .B1(n14980), .B2(n17490), .A(n19432), .ZN(n14439) );
  INV_X1 U16569 ( .A(n14980), .ZN(n19471) );
  NAND2_X1 U16570 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19408) );
  INV_X1 U16571 ( .A(n19408), .ZN(n19415) );
  NAND2_X1 U16572 ( .A1(n19471), .A2(n19415), .ZN(n19400) );
  AND3_X1 U16573 ( .A1(n14439), .A2(n19400), .A3(n19508), .ZN(n19427) );
  AOI21_X1 U16574 ( .B1(n14440), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19427), .ZN(n14441) );
  NAND2_X1 U16575 ( .A1(n14443), .A2(n14442), .ZN(n14470) );
  INV_X1 U16576 ( .A(n14445), .ZN(n14446) );
  NAND2_X1 U16577 ( .A1(n14447), .A2(n14446), .ZN(n14448) );
  INV_X1 U16578 ( .A(n19613), .ZN(n19614) );
  MUX2_X1 U16579 ( .A(n17397), .B(P2_EBX_REG_3__SCAN_IN), .S(n16433), .Z(
        n14451) );
  AOI21_X1 U16580 ( .B1(n19614), .B2(n16457), .A(n14451), .ZN(n14452) );
  INV_X1 U16581 ( .A(n14452), .ZN(P2_U2884) );
  INV_X1 U16582 ( .A(n17397), .ZN(n18850) );
  INV_X1 U16583 ( .A(n14623), .ZN(n14463) );
  NOR2_X1 U16584 ( .A1(n14187), .A2(n14453), .ZN(n14607) );
  INV_X1 U16585 ( .A(n14603), .ZN(n14455) );
  NAND2_X1 U16586 ( .A1(n14621), .A2(n14455), .ZN(n14457) );
  INV_X1 U16587 ( .A(n12448), .ZN(n14456) );
  NAND2_X1 U16588 ( .A1(n14456), .A2(n11409), .ZN(n14602) );
  OAI211_X1 U16589 ( .C1(n14607), .C2(n11001), .A(n14457), .B(n14602), .ZN(
        n14458) );
  INV_X1 U16590 ( .A(n14458), .ZN(n14460) );
  OR2_X1 U16591 ( .A1(n14648), .A2(n14640), .ZN(n14610) );
  AOI22_X1 U16592 ( .A1(n14610), .A2(n14602), .B1(n14603), .B2(n14621), .ZN(
        n14459) );
  MUX2_X1 U16593 ( .A(n14460), .B(n14459), .S(n12648), .Z(n14461) );
  OAI211_X1 U16594 ( .C1(n18850), .C2(n14463), .A(n14462), .B(n14461), .ZN(
        n14631) );
  AOI22_X1 U16595 ( .A1(n19614), .A2(n18897), .B1(n17387), .B2(n14631), .ZN(
        n14465) );
  NAND2_X1 U16596 ( .A1(n17073), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14464) );
  OAI21_X1 U16597 ( .B1(n14465), .B2(n17073), .A(n14464), .ZN(P2_U3596) );
  NAND2_X1 U16598 ( .A1(n14466), .A2(n14467), .ZN(n14472) );
  NAND2_X1 U16599 ( .A1(n14468), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14469) );
  AND2_X1 U16600 ( .A1(n14470), .A2(n14469), .ZN(n14471) );
  NOR2_X1 U16601 ( .A1(n14473), .A2(n15469), .ZN(n14474) );
  OAI211_X1 U16602 ( .C1(n14474), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n16457), .B(n14596), .ZN(n14479) );
  NAND2_X1 U16603 ( .A1(n14475), .A2(n14476), .ZN(n14477) );
  AND2_X1 U16604 ( .A1(n14506), .A2(n14477), .ZN(n18514) );
  NAND2_X1 U16605 ( .A1(n18514), .A2(n16448), .ZN(n14478) );
  OAI211_X1 U16606 ( .C1(n16448), .C2(n18506), .A(n14479), .B(n14478), .ZN(
        P2_U2881) );
  NAND2_X1 U16607 ( .A1(n11920), .A2(n14683), .ZN(n14483) );
  OAI21_X1 U16608 ( .B1(n14482), .B2(n14481), .A(n14480), .ZN(n20137) );
  INV_X1 U16609 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20039) );
  INV_X1 U16610 ( .A(n14789), .ZN(n14732) );
  NAND2_X1 U16611 ( .A1(n14732), .A2(DATAI_1_), .ZN(n14485) );
  NAND2_X1 U16612 ( .A1(n14789), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14484) );
  AND2_X1 U16613 ( .A1(n14485), .A2(n14484), .ZN(n14769) );
  OAI222_X1 U16614 ( .A1(n16023), .A2(n20137), .B1(n16015), .B2(n20039), .C1(
        n16014), .C2(n14769), .ZN(P1_U2903) );
  INV_X1 U16615 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14487) );
  AOI22_X1 U16616 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n17538), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17537), .ZN(n14486) );
  OAI21_X1 U16617 ( .B1(n14487), .B2(n14504), .A(n14486), .ZN(P2_U2935) );
  AOI22_X1 U16618 ( .A1(n17538), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14488) );
  OAI21_X1 U16619 ( .B1(n14160), .B2(n14504), .A(n14488), .ZN(P2_U2929) );
  AOI22_X1 U16620 ( .A1(n17538), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14489) );
  OAI21_X1 U16621 ( .B1(n16485), .B2(n14504), .A(n14489), .ZN(P2_U2923) );
  AOI22_X1 U16622 ( .A1(n17538), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14490) );
  OAI21_X1 U16623 ( .B1(n16541), .B2(n14504), .A(n14490), .ZN(P2_U2930) );
  INV_X1 U16624 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U16625 ( .A1(n17538), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14491) );
  OAI21_X1 U16626 ( .B1(n14492), .B2(n14504), .A(n14491), .ZN(P2_U2931) );
  AOI22_X1 U16627 ( .A1(n17538), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14493) );
  OAI21_X1 U16628 ( .B1(n16495), .B2(n14504), .A(n14493), .ZN(P2_U2924) );
  INV_X1 U16629 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n16478) );
  AOI22_X1 U16630 ( .A1(n17538), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14494) );
  OAI21_X1 U16631 ( .B1(n16478), .B2(n14504), .A(n14494), .ZN(P2_U2922) );
  INV_X1 U16632 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n16515) );
  AOI22_X1 U16633 ( .A1(n17538), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14495) );
  OAI21_X1 U16634 ( .B1(n16515), .B2(n14504), .A(n14495), .ZN(P2_U2926) );
  INV_X1 U16635 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n16522) );
  AOI22_X1 U16636 ( .A1(n17538), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14496) );
  OAI21_X1 U16637 ( .B1(n16522), .B2(n14504), .A(n14496), .ZN(P2_U2927) );
  AOI22_X1 U16638 ( .A1(n17538), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14497) );
  OAI21_X1 U16639 ( .B1(n14498), .B2(n14504), .A(n14497), .ZN(P2_U2925) );
  AOI22_X1 U16640 ( .A1(n17538), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14499) );
  OAI21_X1 U16641 ( .B1(n16530), .B2(n14504), .A(n14499), .ZN(P2_U2928) );
  INV_X1 U16642 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14501) );
  AOI22_X1 U16643 ( .A1(n17530), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14500) );
  OAI21_X1 U16644 ( .B1(n14501), .B2(n14504), .A(n14500), .ZN(P2_U2934) );
  AOI22_X1 U16645 ( .A1(n17530), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14502) );
  OAI21_X1 U16646 ( .B1(n16548), .B2(n14504), .A(n14502), .ZN(P2_U2932) );
  INV_X1 U16647 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n15696) );
  AOI22_X1 U16648 ( .A1(n17530), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14503) );
  OAI21_X1 U16649 ( .B1(n15696), .B2(n14504), .A(n14503), .ZN(P2_U2921) );
  XOR2_X1 U16650 ( .A(n14596), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n14510)
         );
  INV_X1 U16651 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14508) );
  AOI21_X1 U16652 ( .B1(n14507), .B2(n14506), .A(n14505), .ZN(n18524) );
  INV_X1 U16653 ( .A(n18524), .ZN(n15321) );
  MUX2_X1 U16654 ( .A(n14508), .B(n15321), .S(n16448), .Z(n14509) );
  OAI21_X1 U16655 ( .B1(n14510), .B2(n16474), .A(n14509), .ZN(P2_U2880) );
  OR2_X1 U16656 ( .A1(n14513), .A2(n14512), .ZN(n14514) );
  OR2_X1 U16657 ( .A1(n21648), .A2(n12380), .ZN(n14516) );
  AND2_X1 U16658 ( .A1(n14517), .A2(n14516), .ZN(n21643) );
  INV_X1 U16659 ( .A(n21643), .ZN(n14518) );
  AOI22_X1 U16660 ( .A1(n20131), .A2(n14518), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n15949), .ZN(n14519) );
  OAI21_X1 U16661 ( .B1(n20137), .B2(n15954), .A(n14519), .ZN(P1_U2871) );
  NAND2_X1 U16662 ( .A1(n14520), .A2(n21472), .ZN(n14522) );
  NAND2_X1 U16663 ( .A1(n14522), .A2(n14521), .ZN(n15890) );
  INV_X1 U16664 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14525) );
  XOR2_X1 U16665 ( .A(n14524), .B(n14523), .Z(n15888) );
  INV_X1 U16666 ( .A(n15888), .ZN(n14581) );
  OAI222_X1 U16667 ( .A1(n15890), .A2(n15952), .B1(n14525), .B2(n20136), .C1(
        n15954), .C2(n14581), .ZN(P1_U2872) );
  OAI21_X1 U16668 ( .B1(n14527), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14526), .ZN(n14883) );
  NAND2_X1 U16669 ( .A1(n21639), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14876) );
  OAI21_X1 U16670 ( .B1(n20230), .B2(n14528), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14529) );
  OAI211_X1 U16671 ( .C1(n14883), .C2(n21822), .A(n14876), .B(n14529), .ZN(
        n14530) );
  AOI21_X1 U16672 ( .B1(n15888), .B2(n20236), .A(n14530), .ZN(n14531) );
  INV_X1 U16673 ( .A(n14531), .ZN(P1_U2999) );
  XNOR2_X1 U16674 ( .A(n12023), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14543) );
  NOR2_X1 U16675 ( .A1(n14532), .A2(n15380), .ZN(n15002) );
  INV_X1 U16676 ( .A(n14533), .ZN(n14535) );
  NOR2_X1 U16677 ( .A1(n14535), .A2(n14534), .ZN(n14998) );
  INV_X1 U16678 ( .A(n14584), .ZN(n14587) );
  NAND2_X1 U16679 ( .A1(n14587), .A2(n12023), .ZN(n14999) );
  NAND2_X1 U16680 ( .A1(n14584), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15001) );
  NAND2_X1 U16681 ( .A1(n14999), .A2(n15001), .ZN(n14544) );
  MUX2_X1 U16682 ( .A(n15002), .B(n14998), .S(n14544), .Z(n14542) );
  NOR2_X1 U16683 ( .A1(n14537), .A2(n17146), .ZN(n14538) );
  AND2_X1 U16684 ( .A1(n12287), .A2(n14538), .ZN(n14540) );
  AND2_X1 U16685 ( .A1(n14540), .A2(n14539), .ZN(n14583) );
  NOR2_X1 U16686 ( .A1(n14536), .A2(n14583), .ZN(n14541) );
  AOI211_X1 U16687 ( .C1(n17118), .C2(n14543), .A(n14542), .B(n14541), .ZN(
        n14993) );
  INV_X1 U16688 ( .A(n14993), .ZN(n14547) );
  NAND2_X1 U16689 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15383) );
  INV_X1 U16690 ( .A(n15383), .ZN(n14546) );
  INV_X1 U16691 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16164) );
  AOI22_X1 U16692 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n16164), .B2(n21632), .ZN(
        n14590) );
  INV_X1 U16693 ( .A(n21825), .ZN(n21839) );
  INV_X1 U16694 ( .A(n14544), .ZN(n14545) );
  AOI222_X1 U16695 ( .A1(n14547), .A2(n17081), .B1(n14546), .B2(n14590), .C1(
        n21839), .C2(n14545), .ZN(n14557) );
  NOR2_X1 U16696 ( .A1(n14548), .A2(n21875), .ZN(n14549) );
  OAI211_X1 U16697 ( .C1(n17118), .C2(n17146), .A(n14549), .B(n21455), .ZN(
        n14553) );
  OR2_X1 U16698 ( .A1(n21448), .A2(n11023), .ZN(n14550) );
  NAND4_X1 U16699 ( .A1(n14553), .A2(n14552), .A3(n14551), .A4(n14550), .ZN(
        n14555) );
  OR2_X1 U16700 ( .A1(n14555), .A2(n14554), .ZN(n15014) );
  INV_X1 U16701 ( .A(n15014), .ZN(n17121) );
  NAND2_X1 U16702 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21834), .ZN(n21835) );
  INV_X1 U16703 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21823) );
  OAI22_X1 U16704 ( .A1(n17121), .A2(n21844), .B1(n21835), .B2(n21823), .ZN(
        n17079) );
  AOI21_X1 U16705 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21832), .A(n17079), 
        .ZN(n15387) );
  NAND2_X1 U16706 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15387), .ZN(
        n14556) );
  OAI21_X1 U16707 ( .B1(n14557), .B2(n15387), .A(n14556), .ZN(P1_U3472) );
  XNOR2_X1 U16708 ( .A(n14559), .B(n14558), .ZN(n19809) );
  INV_X1 U16709 ( .A(n19809), .ZN(n18468) );
  XNOR2_X1 U16710 ( .A(n18471), .B(n19809), .ZN(n19811) );
  XNOR2_X1 U16711 ( .A(n14561), .B(n14560), .ZN(n18802) );
  NOR2_X1 U16712 ( .A1(n17481), .A2(n18802), .ZN(n19861) );
  NOR2_X1 U16713 ( .A1(n19811), .A2(n19861), .ZN(n19810) );
  AOI21_X1 U16714 ( .B1(n19420), .B2(n18468), .A(n19810), .ZN(n19609) );
  XNOR2_X1 U16715 ( .A(n14562), .B(n14563), .ZN(n19608) );
  XNOR2_X1 U16716 ( .A(n19609), .B(n19608), .ZN(n19612) );
  XNOR2_X1 U16717 ( .A(n19612), .B(n19611), .ZN(n14578) );
  NAND3_X1 U16718 ( .A1(n14566), .A2(n14565), .A3(n14564), .ZN(n14567) );
  NAND2_X1 U16719 ( .A1(n14568), .A2(n14567), .ZN(n14569) );
  NAND2_X1 U16720 ( .A1(n17388), .A2(n14634), .ZN(n14570) );
  AND2_X1 U16721 ( .A1(n11028), .A2(n12687), .ZN(n14573) );
  NOR2_X1 U16722 ( .A1(n14575), .A2(n19562), .ZN(n14574) );
  OR2_X1 U16723 ( .A1(n19763), .A2(n15698), .ZN(n19606) );
  AOI22_X1 U16724 ( .A1(n19606), .A2(n19762), .B1(n19859), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n14577) );
  NAND2_X1 U16725 ( .A1(n19608), .A2(n19860), .ZN(n14576) );
  OAI211_X1 U16726 ( .C1(n14578), .C2(n19812), .A(n14577), .B(n14576), .ZN(
        P2_U2917) );
  NAND2_X1 U16727 ( .A1(n14732), .A2(DATAI_0_), .ZN(n14580) );
  NAND2_X1 U16728 ( .A1(n14789), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14579) );
  AND2_X1 U16729 ( .A1(n14580), .A2(n14579), .ZN(n14771) );
  INV_X1 U16730 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20037) );
  OAI222_X1 U16731 ( .A1(n16014), .A2(n14771), .B1(n16023), .B2(n14581), .C1(
        n20037), .C2(n16015), .ZN(P1_U2904) );
  INV_X1 U16732 ( .A(n15387), .ZN(n21829) );
  INV_X1 U16733 ( .A(n14582), .ZN(n22053) );
  INV_X1 U16734 ( .A(n14583), .ZN(n15382) );
  INV_X1 U16735 ( .A(n17118), .ZN(n14997) );
  NOR2_X1 U16736 ( .A1(n14997), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14586) );
  NOR3_X1 U16737 ( .A1(n15380), .A2(n11823), .A3(n14584), .ZN(n14585) );
  AOI211_X1 U16738 ( .C1(n22053), .C2(n15382), .A(n14586), .B(n14585), .ZN(
        n17122) );
  INV_X1 U16739 ( .A(n17081), .ZN(n21827) );
  NOR2_X1 U16740 ( .A1(n17122), .A2(n21827), .ZN(n14592) );
  INV_X1 U16741 ( .A(n11823), .ZN(n14588) );
  NAND3_X1 U16742 ( .A1(n14588), .A2(n14587), .A3(n21839), .ZN(n14589) );
  OAI21_X1 U16743 ( .B1(n14590), .B2(n15383), .A(n14589), .ZN(n14591) );
  OAI21_X1 U16744 ( .B1(n14592), .B2(n14591), .A(n21829), .ZN(n14593) );
  OAI21_X1 U16745 ( .B1(n21829), .B2(n14594), .A(n14593), .ZN(P1_U3473) );
  OAI21_X1 U16746 ( .B1(n14505), .B2(n14595), .A(n14864), .ZN(n18538) );
  NAND2_X1 U16747 ( .A1(n14597), .A2(n14599), .ZN(n14861) );
  OAI211_X1 U16748 ( .C1(n14597), .C2(n14599), .A(n14598), .B(n16457), .ZN(
        n14601) );
  NAND2_X1 U16749 ( .A1(n16433), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14600) );
  OAI211_X1 U16750 ( .C1(n18538), .C2(n16433), .A(n14601), .B(n14600), .ZN(
        P2_U2879) );
  NAND2_X1 U16751 ( .A1(n18863), .A2(n14623), .ZN(n14612) );
  INV_X1 U16752 ( .A(n11001), .ZN(n15675) );
  NAND2_X1 U16753 ( .A1(n15675), .A2(n14602), .ZN(n14609) );
  NOR2_X1 U16754 ( .A1(n14604), .A2(n14603), .ZN(n14605) );
  NAND2_X1 U16755 ( .A1(n14621), .A2(n14605), .ZN(n14606) );
  OAI21_X1 U16756 ( .B1(n14607), .B2(n14609), .A(n14606), .ZN(n14608) );
  AOI21_X1 U16757 ( .B1(n14610), .B2(n14609), .A(n14608), .ZN(n14611) );
  NAND2_X1 U16758 ( .A1(n14612), .A2(n14611), .ZN(n17072) );
  INV_X1 U16759 ( .A(n17072), .ZN(n14627) );
  NAND2_X1 U16760 ( .A1(n18470), .A2(n14623), .ZN(n14618) );
  NOR2_X1 U16761 ( .A1(n14613), .A2(n12448), .ZN(n14615) );
  NAND2_X1 U16762 ( .A1(n14614), .A2(n14174), .ZN(n14620) );
  AOI22_X1 U16763 ( .A1(n14621), .A2(n14616), .B1(n14615), .B2(n14620), .ZN(
        n14617) );
  NAND2_X1 U16764 ( .A1(n14618), .A2(n14617), .ZN(n17067) );
  INV_X1 U16765 ( .A(n17067), .ZN(n14624) );
  MUX2_X1 U16766 ( .A(n14621), .B(n14620), .S(n14619), .Z(n14622) );
  AOI21_X1 U16767 ( .B1(n18452), .B2(n14623), .A(n14622), .ZN(n17057) );
  OAI211_X1 U16768 ( .C1(n14624), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n17057), .ZN(n14625) );
  OAI21_X1 U16769 ( .B1(n17067), .B2(n19488), .A(n14625), .ZN(n14626) );
  AOI21_X1 U16770 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14627), .A(
        n14626), .ZN(n14628) );
  MUX2_X1 U16771 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17072), .S(
        n14655), .Z(n14652) );
  AOI22_X1 U16772 ( .A1(n14628), .A2(n14655), .B1(n14652), .B2(n17490), .ZN(
        n14633) );
  INV_X1 U16773 ( .A(n14655), .ZN(n14630) );
  NAND2_X1 U16774 ( .A1(n14630), .A2(n12648), .ZN(n14629) );
  OAI21_X1 U16775 ( .B1(n14631), .B2(n14630), .A(n14629), .ZN(n14654) );
  OR2_X1 U16776 ( .A1(n14654), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14632) );
  AOI221_X1 U16777 ( .B1(n14633), .B2(n14632), .C1(n14654), .C2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n14660) );
  NOR2_X1 U16778 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n14651) );
  INV_X1 U16779 ( .A(n14661), .ZN(n16331) );
  INV_X1 U16780 ( .A(n14634), .ZN(n14635) );
  NAND4_X1 U16781 ( .A1(n14639), .A2(n14636), .A3(n16331), .A4(n14635), .ZN(
        n18906) );
  AOI22_X1 U16782 ( .A1(n14639), .A2(n14638), .B1(n14637), .B2(n18894), .ZN(
        n14643) );
  NAND2_X1 U16783 ( .A1(n14641), .A2(n14640), .ZN(n14642) );
  OAI211_X1 U16784 ( .C1(n14645), .C2(n14644), .A(n14643), .B(n14642), .ZN(
        n14646) );
  AOI21_X1 U16785 ( .B1(n14648), .B2(n14647), .A(n14646), .ZN(n18909) );
  NAND2_X1 U16786 ( .A1(n14649), .A2(n15667), .ZN(n14650) );
  OAI211_X1 U16787 ( .C1(n14651), .C2(n18906), .A(n18909), .B(n14650), .ZN(
        n14658) );
  INV_X1 U16788 ( .A(n14652), .ZN(n14653) );
  OAI22_X1 U16789 ( .A1(n14656), .A2(n14655), .B1(n14654), .B2(n14653), .ZN(
        n14657) );
  NOR4_X1 U16790 ( .A1(n14660), .A2(n14659), .A3(n14658), .A4(n14657), .ZN(
        n18905) );
  NAND3_X1 U16791 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18905), .A3(n18890), 
        .ZN(n14665) );
  NAND3_X1 U16792 ( .A1(n14663), .A2(n14662), .A3(n14661), .ZN(n16326) );
  NOR2_X1 U16793 ( .A1(n13892), .A2(n16326), .ZN(n14664) );
  AOI21_X1 U16794 ( .B1(n14665), .B2(n14839), .A(n14664), .ZN(n18896) );
  OAI21_X1 U16795 ( .B1(n18896), .B2(n14841), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14666) );
  NAND2_X1 U16796 ( .A1(n14666), .A2(n18893), .ZN(P2_U3593) );
  NAND2_X1 U16797 ( .A1(n15105), .A2(n15104), .ZN(n14939) );
  INV_X1 U16798 ( .A(n22041), .ZN(n21941) );
  INV_X1 U16799 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20304) );
  INV_X1 U16800 ( .A(DATAI_29_), .ZN(n17194) );
  OAI22_X1 U16801 ( .A1(n20304), .A2(n14748), .B1(n17194), .B2(n14747), .ZN(
        n22257) );
  INV_X1 U16802 ( .A(n22257), .ZN(n22267) );
  INV_X1 U16803 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20287) );
  INV_X1 U16804 ( .A(DATAI_21_), .ZN(n17309) );
  OAI22_X1 U16805 ( .A1(n20287), .A2(n14748), .B1(n17309), .B2(n14747), .ZN(
        n22264) );
  OR2_X1 U16806 ( .A1(n14939), .A2(n15043), .ZN(n14725) );
  NOR2_X1 U16807 ( .A1(n14536), .A2(n15010), .ZN(n21966) );
  INV_X1 U16808 ( .A(n21966), .ZN(n14935) );
  NAND2_X1 U16809 ( .A1(n14668), .A2(n10986), .ZN(n22064) );
  OAI21_X1 U16810 ( .B1(n14935), .B2(n22064), .A(n14751), .ZN(n14675) );
  NOR2_X1 U16811 ( .A1(n22067), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14678) );
  INV_X1 U16812 ( .A(n14678), .ZN(n14669) );
  NOR2_X1 U16813 ( .A1(n13234), .A2(n14669), .ZN(n14670) );
  AOI21_X1 U16814 ( .B1(n14675), .B2(n22077), .A(n14670), .ZN(n14752) );
  NAND2_X1 U16815 ( .A1(n14732), .A2(DATAI_5_), .ZN(n14672) );
  NAND2_X1 U16816 ( .A1(n14789), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14671) );
  AND2_X1 U16817 ( .A1(n14672), .A2(n14671), .ZN(n14915) );
  NAND2_X1 U16818 ( .A1(n14750), .A2(n11858), .ZN(n22262) );
  OAI22_X1 U16819 ( .A1(n14752), .A2(n22261), .B1(n14751), .B2(n22262), .ZN(
        n14674) );
  AOI21_X1 U16820 ( .B1(n22264), .B2(n22343), .A(n14674), .ZN(n14680) );
  NAND2_X1 U16821 ( .A1(n14667), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21952) );
  INV_X1 U16822 ( .A(n14675), .ZN(n14676) );
  OAI211_X1 U16823 ( .C1(n14939), .C2(n21952), .A(n22077), .B(n14676), .ZN(
        n14677) );
  OAI211_X1 U16824 ( .C1(n22077), .C2(n14678), .A(n14677), .B(n22035), .ZN(
        n14754) );
  NAND2_X1 U16825 ( .A1(n14754), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14679) );
  OAI211_X1 U16826 ( .C1(n14757), .C2(n22267), .A(n14680), .B(n14679), .ZN(
        P1_U3094) );
  INV_X1 U16827 ( .A(DATAI_31_), .ZN(n17290) );
  OAI22_X1 U16828 ( .A1(n20308), .A2(n14748), .B1(n17290), .B2(n14747), .ZN(
        n22377) );
  INV_X1 U16829 ( .A(n22377), .ZN(n22394) );
  INV_X1 U16830 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20291) );
  INV_X1 U16831 ( .A(DATAI_23_), .ZN(n17299) );
  OAI22_X1 U16832 ( .A1(n20291), .A2(n14748), .B1(n17299), .B2(n14747), .ZN(
        n22388) );
  NAND2_X1 U16833 ( .A1(n14732), .A2(DATAI_7_), .ZN(n14682) );
  NAND2_X1 U16834 ( .A1(n14789), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14681) );
  AND2_X1 U16835 ( .A1(n14682), .A2(n14681), .ZN(n15130) );
  NAND2_X1 U16836 ( .A1(n14750), .A2(n14683), .ZN(n22386) );
  OAI22_X1 U16837 ( .A1(n14752), .A2(n22383), .B1(n14751), .B2(n22386), .ZN(
        n14684) );
  AOI21_X1 U16838 ( .B1(n22388), .B2(n22343), .A(n14684), .ZN(n14686) );
  NAND2_X1 U16839 ( .A1(n14754), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14685) );
  OAI211_X1 U16840 ( .C1(n14757), .C2(n22394), .A(n14686), .B(n14685), .ZN(
        P1_U3096) );
  INV_X1 U16841 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20306) );
  INV_X1 U16842 ( .A(DATAI_30_), .ZN(n17188) );
  OAI22_X1 U16843 ( .A1(n20306), .A2(n14748), .B1(n17188), .B2(n14747), .ZN(
        n22294) );
  INV_X1 U16844 ( .A(n22294), .ZN(n22304) );
  INV_X1 U16845 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20289) );
  INV_X1 U16846 ( .A(DATAI_22_), .ZN(n17307) );
  OAI22_X1 U16847 ( .A1(n20289), .A2(n14748), .B1(n17307), .B2(n14747), .ZN(
        n22301) );
  NAND2_X1 U16848 ( .A1(n14732), .A2(DATAI_6_), .ZN(n14688) );
  NAND2_X1 U16849 ( .A1(n14789), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14687) );
  AND2_X1 U16850 ( .A1(n14688), .A2(n14687), .ZN(n14978) );
  NAND2_X1 U16851 ( .A1(n14750), .A2(n14689), .ZN(n22299) );
  OAI22_X1 U16852 ( .A1(n14752), .A2(n22298), .B1(n14751), .B2(n22299), .ZN(
        n14690) );
  AOI21_X1 U16853 ( .B1(n22301), .B2(n22343), .A(n14690), .ZN(n14692) );
  NAND2_X1 U16854 ( .A1(n14754), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14691) );
  OAI211_X1 U16855 ( .C1(n14757), .C2(n22304), .A(n14692), .B(n14691), .ZN(
        P1_U3095) );
  INV_X1 U16856 ( .A(n15107), .ZN(n14693) );
  INV_X1 U16857 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20277) );
  INV_X1 U16858 ( .A(DATAI_16_), .ZN(n17181) );
  OAI22_X1 U16859 ( .A1(n20277), .A2(n14748), .B1(n17181), .B2(n14747), .ZN(
        n22078) );
  INV_X1 U16860 ( .A(n22078), .ZN(n22062) );
  NOR3_X1 U16861 ( .A1(n12225), .A2(n21944), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22001) );
  NAND2_X1 U16862 ( .A1(n14694), .A2(n14536), .ZN(n21997) );
  OR2_X1 U16863 ( .A1(n21997), .A2(n22064), .ZN(n14696) );
  INV_X1 U16864 ( .A(n22001), .ZN(n14695) );
  OR2_X1 U16865 ( .A1(n22029), .A2(n14695), .ZN(n14832) );
  AND2_X1 U16866 ( .A1(n14696), .A2(n14832), .ZN(n14699) );
  OAI211_X1 U16867 ( .C1(n21993), .C2(n21952), .A(n22077), .B(n14699), .ZN(
        n14697) );
  OAI211_X1 U16868 ( .C1(n22077), .C2(n22001), .A(n14697), .B(n22035), .ZN(
        n14831) );
  NAND2_X1 U16869 ( .A1(n14831), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14703) );
  INV_X1 U16870 ( .A(DATAI_24_), .ZN(n14698) );
  INV_X1 U16871 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20293) );
  OAI22_X2 U16872 ( .A1(n14698), .A2(n14747), .B1(n20293), .B2(n14748), .ZN(
        n22059) );
  INV_X1 U16873 ( .A(n14699), .ZN(n14700) );
  AOI22_X1 U16874 ( .A1(n14700), .A2(n22077), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n22001), .ZN(n14833) );
  NAND2_X1 U16875 ( .A1(n14750), .A2(n11027), .ZN(n22070) );
  OAI22_X1 U16876 ( .A1(n14833), .A2(n22069), .B1(n22070), .B2(n14832), .ZN(
        n14701) );
  AOI21_X1 U16877 ( .B1(n22354), .B2(n22059), .A(n14701), .ZN(n14702) );
  OAI211_X1 U16878 ( .C1(n14812), .C2(n22062), .A(n14703), .B(n14702), .ZN(
        P1_U3121) );
  XOR2_X1 U16879 ( .A(n14480), .B(n14704), .Z(n20147) );
  INV_X1 U16880 ( .A(n20147), .ZN(n15887) );
  NAND2_X1 U16881 ( .A1(n14706), .A2(n14705), .ZN(n14707) );
  NAND2_X1 U16882 ( .A1(n14730), .A2(n14707), .ZN(n21474) );
  INV_X1 U16883 ( .A(n21474), .ZN(n14708) );
  AOI22_X1 U16884 ( .A1(n14708), .A2(n20131), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n15949), .ZN(n14709) );
  OAI21_X1 U16885 ( .B1(n15887), .B2(n15954), .A(n14709), .ZN(P1_U2870) );
  INV_X1 U16886 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20302) );
  INV_X1 U16887 ( .A(DATAI_28_), .ZN(n17192) );
  OAI22_X1 U16888 ( .A1(n20302), .A2(n14748), .B1(n17192), .B2(n14747), .ZN(
        n22220) );
  INV_X1 U16889 ( .A(n22220), .ZN(n22230) );
  INV_X1 U16890 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20285) );
  INV_X1 U16891 ( .A(DATAI_20_), .ZN(n17289) );
  OAI22_X1 U16892 ( .A1(n20285), .A2(n14748), .B1(n17289), .B2(n14747), .ZN(
        n22227) );
  NAND2_X1 U16893 ( .A1(n14732), .A2(DATAI_4_), .ZN(n14711) );
  NAND2_X1 U16894 ( .A1(n14789), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14710) );
  AND2_X1 U16895 ( .A1(n14711), .A2(n14710), .ZN(n14893) );
  NAND2_X1 U16896 ( .A1(n14750), .A2(n14712), .ZN(n22225) );
  OAI22_X1 U16897 ( .A1(n14752), .A2(n22224), .B1(n14751), .B2(n22225), .ZN(
        n14713) );
  AOI21_X1 U16898 ( .B1(n22227), .B2(n22343), .A(n14713), .ZN(n14715) );
  NAND2_X1 U16899 ( .A1(n14754), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14714) );
  OAI211_X1 U16900 ( .C1(n14757), .C2(n22230), .A(n14715), .B(n14714), .ZN(
        P1_U3093) );
  INV_X1 U16901 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20298) );
  INV_X1 U16902 ( .A(DATAI_26_), .ZN(n14716) );
  OAI22_X1 U16903 ( .A1(n20298), .A2(n14748), .B1(n14716), .B2(n14747), .ZN(
        n22145) );
  INV_X1 U16904 ( .A(n22145), .ZN(n22155) );
  INV_X1 U16905 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20281) );
  INV_X1 U16906 ( .A(DATAI_18_), .ZN(n17208) );
  OAI22_X1 U16907 ( .A1(n20281), .A2(n14748), .B1(n17208), .B2(n14747), .ZN(
        n22152) );
  NAND2_X1 U16908 ( .A1(n14732), .A2(DATAI_2_), .ZN(n14718) );
  NAND2_X1 U16909 ( .A1(n14789), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14717) );
  AND2_X1 U16910 ( .A1(n14718), .A2(n14717), .ZN(n14811) );
  NAND2_X1 U16911 ( .A1(n14750), .A2(n11023), .ZN(n22150) );
  OAI22_X1 U16912 ( .A1(n14752), .A2(n22149), .B1(n14751), .B2(n22150), .ZN(
        n14719) );
  AOI21_X1 U16913 ( .B1(n22152), .B2(n22343), .A(n14719), .ZN(n14721) );
  NAND2_X1 U16914 ( .A1(n14754), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14720) );
  OAI211_X1 U16915 ( .C1(n14757), .C2(n22155), .A(n14721), .B(n14720), .ZN(
        P1_U3091) );
  OAI22_X1 U16916 ( .A1(n14752), .A2(n22069), .B1(n14751), .B2(n22070), .ZN(
        n14722) );
  AOI21_X1 U16917 ( .B1(n22059), .B2(n22336), .A(n14722), .ZN(n14724) );
  NAND2_X1 U16918 ( .A1(n14754), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14723) );
  OAI211_X1 U16919 ( .C1(n14725), .C2(n22062), .A(n14724), .B(n14723), .ZN(
        P1_U3089) );
  NAND2_X1 U16920 ( .A1(n14726), .A2(n14727), .ZN(n14886) );
  OAI21_X1 U16921 ( .B1(n14726), .B2(n14727), .A(n14886), .ZN(n20155) );
  INV_X1 U16922 ( .A(n14728), .ZN(n14729) );
  XNOR2_X1 U16923 ( .A(n14730), .B(n14729), .ZN(n21661) );
  AOI22_X1 U16924 ( .A1(n21661), .A2(n20131), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n15949), .ZN(n14731) );
  OAI21_X1 U16925 ( .B1(n20155), .B2(n15954), .A(n14731), .ZN(P1_U2869) );
  INV_X1 U16926 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20300) );
  INV_X1 U16927 ( .A(DATAI_27_), .ZN(n17295) );
  OAI22_X1 U16928 ( .A1(n20300), .A2(n14748), .B1(n17295), .B2(n14747), .ZN(
        n22182) );
  INV_X1 U16929 ( .A(n22182), .ZN(n22192) );
  INV_X1 U16930 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20283) );
  INV_X1 U16931 ( .A(DATAI_19_), .ZN(n17186) );
  OAI22_X1 U16932 ( .A1(n20283), .A2(n14748), .B1(n17186), .B2(n14747), .ZN(
        n22189) );
  NAND2_X1 U16933 ( .A1(n14732), .A2(DATAI_3_), .ZN(n14734) );
  NAND2_X1 U16934 ( .A1(n14789), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14733) );
  AND2_X1 U16935 ( .A1(n14734), .A2(n14733), .ZN(n14838) );
  NAND2_X1 U16936 ( .A1(n14750), .A2(n14735), .ZN(n22187) );
  OAI22_X1 U16937 ( .A1(n14752), .A2(n22186), .B1(n14751), .B2(n22187), .ZN(
        n14736) );
  AOI21_X1 U16938 ( .B1(n22189), .B2(n22343), .A(n14736), .ZN(n14738) );
  NAND2_X1 U16939 ( .A1(n14754), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14737) );
  OAI211_X1 U16940 ( .C1(n14757), .C2(n22192), .A(n14738), .B(n14737), .ZN(
        P1_U3092) );
  INV_X1 U16941 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20067) );
  NOR2_X1 U16942 ( .A1(n17144), .A2(n21455), .ZN(n14739) );
  NOR2_X2 U16943 ( .A1(n14808), .A2(n14741), .ZN(n14790) );
  INV_X1 U16944 ( .A(n14790), .ZN(n14746) );
  INV_X1 U16945 ( .A(DATAI_15_), .ZN(n14742) );
  NOR2_X1 U16946 ( .A1(n14789), .A2(n14742), .ZN(n14743) );
  AOI21_X1 U16947 ( .B1(n14789), .B2(BUF1_REG_15__SCAN_IN), .A(n14743), .ZN(
        n16013) );
  INV_X1 U16948 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14744) );
  OAI222_X1 U16949 ( .A1(n14807), .A2(n20067), .B1(n14746), .B2(n16013), .C1(
        n14745), .C2(n14744), .ZN(P1_U2967) );
  INV_X1 U16950 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20295) );
  INV_X1 U16951 ( .A(DATAI_25_), .ZN(n17298) );
  OAI22_X1 U16952 ( .A1(n20295), .A2(n14748), .B1(n17298), .B2(n14747), .ZN(
        n22108) );
  INV_X1 U16953 ( .A(n22108), .ZN(n22118) );
  INV_X1 U16954 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20279) );
  INV_X1 U16955 ( .A(DATAI_17_), .ZN(n17315) );
  OAI22_X1 U16956 ( .A1(n20279), .A2(n14748), .B1(n17315), .B2(n14747), .ZN(
        n22115) );
  NAND2_X1 U16957 ( .A1(n14750), .A2(n14749), .ZN(n22113) );
  OAI22_X1 U16958 ( .A1(n14752), .A2(n22112), .B1(n14751), .B2(n22113), .ZN(
        n14753) );
  AOI21_X1 U16959 ( .B1(n22115), .B2(n22343), .A(n14753), .ZN(n14756) );
  NAND2_X1 U16960 ( .A1(n14754), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14755) );
  OAI211_X1 U16961 ( .C1(n14757), .C2(n22118), .A(n14756), .B(n14755), .ZN(
        P1_U3090) );
  INV_X1 U16962 ( .A(n14915), .ZN(n15990) );
  NAND2_X1 U16963 ( .A1(n14790), .A2(n15990), .ZN(n14793) );
  NAND2_X1 U16964 ( .A1(n14804), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n14758) );
  OAI211_X1 U16965 ( .C1(n13283), .C2(n14807), .A(n14793), .B(n14758), .ZN(
        P1_U2957) );
  INV_X1 U16966 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15400) );
  INV_X1 U16967 ( .A(n14838), .ZN(n15996) );
  NAND2_X1 U16968 ( .A1(n14790), .A2(n15996), .ZN(n14795) );
  NAND2_X1 U16969 ( .A1(n14808), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14759) );
  OAI211_X1 U16970 ( .C1(n15400), .C2(n14807), .A(n14795), .B(n14759), .ZN(
        P1_U2940) );
  INV_X1 U16971 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20050) );
  INV_X1 U16972 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20261) );
  NOR2_X1 U16973 ( .A1(n14789), .A2(DATAI_8_), .ZN(n14760) );
  AOI21_X1 U16974 ( .B1(n14789), .B2(n20261), .A(n14760), .ZN(n15980) );
  NAND2_X1 U16975 ( .A1(n14790), .A2(n15980), .ZN(n14803) );
  NAND2_X1 U16976 ( .A1(n14804), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14761) );
  OAI211_X1 U16977 ( .C1(n20050), .C2(n14807), .A(n14803), .B(n14761), .ZN(
        P1_U2960) );
  INV_X1 U16978 ( .A(n15130), .ZN(n15984) );
  NAND2_X1 U16979 ( .A1(n14790), .A2(n15984), .ZN(n14765) );
  NAND2_X1 U16980 ( .A1(n14808), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n14762) );
  OAI211_X1 U16981 ( .C1(n13294), .C2(n14807), .A(n14765), .B(n14762), .ZN(
        P1_U2959) );
  INV_X1 U16982 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20052) );
  MUX2_X1 U16983 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n14789), .Z(
        n15976) );
  NAND2_X1 U16984 ( .A1(n14790), .A2(n15976), .ZN(n14810) );
  NAND2_X1 U16985 ( .A1(n14804), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n14763) );
  OAI211_X1 U16986 ( .C1(n20052), .C2(n14807), .A(n14810), .B(n14763), .ZN(
        P1_U2961) );
  INV_X1 U16987 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n15408) );
  NAND2_X1 U16988 ( .A1(n14808), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14764) );
  OAI211_X1 U16989 ( .C1(n15408), .C2(n14807), .A(n14765), .B(n14764), .ZN(
        P1_U2944) );
  INV_X1 U16990 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15402) );
  INV_X1 U16991 ( .A(n14893), .ZN(n15993) );
  NAND2_X1 U16992 ( .A1(n14790), .A2(n15993), .ZN(n14777) );
  NAND2_X1 U16993 ( .A1(n14808), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14766) );
  OAI211_X1 U16994 ( .C1(n15402), .C2(n14807), .A(n14777), .B(n14766), .ZN(
        P1_U2941) );
  INV_X1 U16995 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15423) );
  MUX2_X1 U16996 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n14789), .Z(
        n16016) );
  NAND2_X1 U16997 ( .A1(n14790), .A2(n16016), .ZN(n14781) );
  NAND2_X1 U16998 ( .A1(n14804), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n14767) );
  OAI211_X1 U16999 ( .C1(n15423), .C2(n14807), .A(n14781), .B(n14767), .ZN(
        P1_U2951) );
  INV_X1 U17000 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20041) );
  INV_X1 U17001 ( .A(n14811), .ZN(n16000) );
  NAND2_X1 U17002 ( .A1(n14790), .A2(n16000), .ZN(n14786) );
  NAND2_X1 U17003 ( .A1(n14804), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n14768) );
  OAI211_X1 U17004 ( .C1(n20041), .C2(n14807), .A(n14786), .B(n14768), .ZN(
        P1_U2954) );
  INV_X1 U17005 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15396) );
  INV_X1 U17006 ( .A(n14769), .ZN(n16003) );
  NAND2_X1 U17007 ( .A1(n14790), .A2(n16003), .ZN(n14788) );
  NAND2_X1 U17008 ( .A1(n14808), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14770) );
  OAI211_X1 U17009 ( .C1(n15396), .C2(n14807), .A(n14788), .B(n14770), .ZN(
        P1_U2938) );
  INV_X1 U17010 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15394) );
  INV_X1 U17011 ( .A(n14771), .ZN(n16009) );
  NAND2_X1 U17012 ( .A1(n14790), .A2(n16009), .ZN(n14806) );
  NAND2_X1 U17013 ( .A1(n14808), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14772) );
  OAI211_X1 U17014 ( .C1(n15394), .C2(n14807), .A(n14806), .B(n14772), .ZN(
        P1_U2937) );
  INV_X1 U17015 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20055) );
  MUX2_X1 U17016 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n14789), .Z(
        n15972) );
  NAND2_X1 U17017 ( .A1(n14790), .A2(n15972), .ZN(n14801) );
  NAND2_X1 U17018 ( .A1(n14804), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n14773) );
  OAI211_X1 U17019 ( .C1(n20055), .C2(n14807), .A(n14801), .B(n14773), .ZN(
        P1_U2962) );
  INV_X1 U17020 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15420) );
  MUX2_X1 U17021 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n14789), .Z(
        n16020) );
  NAND2_X1 U17022 ( .A1(n14790), .A2(n16020), .ZN(n14783) );
  NAND2_X1 U17023 ( .A1(n14804), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n14774) );
  OAI211_X1 U17024 ( .C1(n15420), .C2(n14807), .A(n14783), .B(n14774), .ZN(
        P1_U2950) );
  INV_X1 U17025 ( .A(n14978), .ZN(n15987) );
  NAND2_X1 U17026 ( .A1(n14790), .A2(n15987), .ZN(n14779) );
  NAND2_X1 U17027 ( .A1(n14808), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n14775) );
  OAI211_X1 U17028 ( .C1(n13290), .C2(n14807), .A(n14779), .B(n14775), .ZN(
        P1_U2958) );
  INV_X1 U17029 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20045) );
  NAND2_X1 U17030 ( .A1(n14804), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n14776) );
  OAI211_X1 U17031 ( .C1(n20045), .C2(n14807), .A(n14777), .B(n14776), .ZN(
        P1_U2956) );
  INV_X1 U17032 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15406) );
  NAND2_X1 U17033 ( .A1(n14808), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14778) );
  OAI211_X1 U17034 ( .C1(n15406), .C2(n14807), .A(n14779), .B(n14778), .ZN(
        P1_U2943) );
  INV_X1 U17035 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20064) );
  NAND2_X1 U17036 ( .A1(n14804), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n14780) );
  OAI211_X1 U17037 ( .C1(n20064), .C2(n14807), .A(n14781), .B(n14780), .ZN(
        P1_U2966) );
  INV_X1 U17038 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20062) );
  NAND2_X1 U17039 ( .A1(n14804), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n14782) );
  OAI211_X1 U17040 ( .C1(n20062), .C2(n14807), .A(n14783), .B(n14782), .ZN(
        P1_U2965) );
  INV_X1 U17041 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20059) );
  MUX2_X1 U17042 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n14789), .Z(
        n15964) );
  NAND2_X1 U17043 ( .A1(n14790), .A2(n15964), .ZN(n14797) );
  NAND2_X1 U17044 ( .A1(n14804), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n14784) );
  OAI211_X1 U17045 ( .C1(n20059), .C2(n14807), .A(n14797), .B(n14784), .ZN(
        P1_U2964) );
  INV_X1 U17046 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15398) );
  NAND2_X1 U17047 ( .A1(n14808), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14785) );
  OAI211_X1 U17048 ( .C1(n15398), .C2(n14807), .A(n14786), .B(n14785), .ZN(
        P1_U2939) );
  NAND2_X1 U17049 ( .A1(n14804), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n14787) );
  OAI211_X1 U17050 ( .C1(n20039), .C2(n14807), .A(n14788), .B(n14787), .ZN(
        P1_U2953) );
  MUX2_X1 U17051 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n14789), .Z(
        n15968) );
  NAND2_X1 U17052 ( .A1(n14790), .A2(n15968), .ZN(n14799) );
  NAND2_X1 U17053 ( .A1(n14804), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n14791) );
  OAI211_X1 U17054 ( .C1(n14807), .C2(n20057), .A(n14799), .B(n14791), .ZN(
        P1_U2963) );
  INV_X1 U17055 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15404) );
  NAND2_X1 U17056 ( .A1(n14808), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14792) );
  OAI211_X1 U17057 ( .C1(n15404), .C2(n14807), .A(n14793), .B(n14792), .ZN(
        P1_U2942) );
  INV_X1 U17058 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20043) );
  NAND2_X1 U17059 ( .A1(n14804), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n14794) );
  OAI211_X1 U17060 ( .C1(n20043), .C2(n14807), .A(n14795), .B(n14794), .ZN(
        P1_U2955) );
  INV_X1 U17061 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15418) );
  NAND2_X1 U17062 ( .A1(n14804), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14796) );
  OAI211_X1 U17063 ( .C1(n15418), .C2(n14807), .A(n14797), .B(n14796), .ZN(
        P1_U2949) );
  INV_X1 U17064 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n15416) );
  NAND2_X1 U17065 ( .A1(n14804), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14798) );
  OAI211_X1 U17066 ( .C1(n15416), .C2(n14807), .A(n14799), .B(n14798), .ZN(
        P1_U2948) );
  INV_X1 U17067 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15414) );
  NAND2_X1 U17068 ( .A1(n14808), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14800) );
  OAI211_X1 U17069 ( .C1(n15414), .C2(n14807), .A(n14801), .B(n14800), .ZN(
        P1_U2947) );
  INV_X1 U17070 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15410) );
  NAND2_X1 U17071 ( .A1(n14808), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14802) );
  OAI211_X1 U17072 ( .C1(n15410), .C2(n14807), .A(n14803), .B(n14802), .ZN(
        P1_U2945) );
  NAND2_X1 U17073 ( .A1(n14804), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n14805) );
  OAI211_X1 U17074 ( .C1(n20037), .C2(n14807), .A(n14806), .B(n14805), .ZN(
        P1_U2952) );
  INV_X1 U17075 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15412) );
  NAND2_X1 U17076 ( .A1(n14808), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14809) );
  OAI211_X1 U17077 ( .C1(n15412), .C2(n14807), .A(n14810), .B(n14809), .ZN(
        P1_U2946) );
  OAI222_X1 U17078 ( .A1(n16023), .A2(n15887), .B1(n16015), .B2(n20041), .C1(
        n16014), .C2(n14811), .ZN(P1_U2902) );
  NAND2_X1 U17079 ( .A1(n14831), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14815) );
  OAI22_X1 U17080 ( .A1(n14833), .A2(n22261), .B1(n22262), .B2(n14832), .ZN(
        n14813) );
  AOI21_X1 U17081 ( .B1(n22362), .B2(n22264), .A(n14813), .ZN(n14814) );
  OAI211_X1 U17082 ( .C1(n14837), .C2(n22267), .A(n14815), .B(n14814), .ZN(
        P1_U3126) );
  NAND2_X1 U17083 ( .A1(n14831), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14818) );
  OAI22_X1 U17084 ( .A1(n14833), .A2(n22186), .B1(n22187), .B2(n14832), .ZN(
        n14816) );
  AOI21_X1 U17085 ( .B1(n22362), .B2(n22189), .A(n14816), .ZN(n14817) );
  OAI211_X1 U17086 ( .C1(n14837), .C2(n22192), .A(n14818), .B(n14817), .ZN(
        P1_U3124) );
  NAND2_X1 U17087 ( .A1(n14831), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n14821) );
  OAI22_X1 U17088 ( .A1(n14833), .A2(n22383), .B1(n22386), .B2(n14832), .ZN(
        n14819) );
  AOI21_X1 U17089 ( .B1(n22362), .B2(n22388), .A(n14819), .ZN(n14820) );
  OAI211_X1 U17090 ( .C1(n14837), .C2(n22394), .A(n14821), .B(n14820), .ZN(
        P1_U3128) );
  NAND2_X1 U17091 ( .A1(n14831), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14824) );
  OAI22_X1 U17092 ( .A1(n14833), .A2(n22224), .B1(n22225), .B2(n14832), .ZN(
        n14822) );
  AOI21_X1 U17093 ( .B1(n22362), .B2(n22227), .A(n14822), .ZN(n14823) );
  OAI211_X1 U17094 ( .C1(n14837), .C2(n22230), .A(n14824), .B(n14823), .ZN(
        P1_U3125) );
  NAND2_X1 U17095 ( .A1(n14831), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14827) );
  OAI22_X1 U17096 ( .A1(n14833), .A2(n22149), .B1(n22150), .B2(n14832), .ZN(
        n14825) );
  AOI21_X1 U17097 ( .B1(n22362), .B2(n22152), .A(n14825), .ZN(n14826) );
  OAI211_X1 U17098 ( .C1(n14837), .C2(n22155), .A(n14827), .B(n14826), .ZN(
        P1_U3123) );
  NAND2_X1 U17099 ( .A1(n14831), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14830) );
  OAI22_X1 U17100 ( .A1(n14833), .A2(n22298), .B1(n22299), .B2(n14832), .ZN(
        n14828) );
  AOI21_X1 U17101 ( .B1(n22362), .B2(n22301), .A(n14828), .ZN(n14829) );
  OAI211_X1 U17102 ( .C1(n14837), .C2(n22304), .A(n14830), .B(n14829), .ZN(
        P1_U3127) );
  NAND2_X1 U17103 ( .A1(n14831), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14836) );
  OAI22_X1 U17104 ( .A1(n14833), .A2(n22112), .B1(n22113), .B2(n14832), .ZN(
        n14834) );
  AOI21_X1 U17105 ( .B1(n22362), .B2(n22115), .A(n14834), .ZN(n14835) );
  OAI211_X1 U17106 ( .C1(n14837), .C2(n22118), .A(n14836), .B(n14835), .ZN(
        P1_U3122) );
  OAI222_X1 U17107 ( .A1(n16023), .A2(n20155), .B1(n16015), .B2(n20043), .C1(
        n16014), .C2(n14838), .ZN(P1_U2901) );
  NAND2_X1 U17108 ( .A1(n18471), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19489) );
  NOR2_X1 U17109 ( .A1(n17488), .A2(n19489), .ZN(n17487) );
  NAND2_X1 U17110 ( .A1(n17487), .A2(n19613), .ZN(n14851) );
  NAND2_X1 U17111 ( .A1(n19432), .A2(n17490), .ZN(n19528) );
  INV_X1 U17112 ( .A(n19528), .ZN(n15165) );
  NAND2_X1 U17113 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15165), .ZN(
        n14849) );
  NAND2_X1 U17114 ( .A1(n14851), .A2(n14849), .ZN(n14848) );
  NAND2_X1 U17115 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n14841), .ZN(n16281) );
  NAND2_X1 U17116 ( .A1(n14839), .A2(n16281), .ZN(n18900) );
  NAND2_X1 U17117 ( .A1(n19472), .A2(n14842), .ZN(n19535) );
  INV_X1 U17118 ( .A(n19535), .ZN(n15169) );
  NAND2_X1 U17119 ( .A1(n14852), .A2(n15169), .ZN(n14846) );
  NOR2_X1 U17120 ( .A1(n14980), .A2(n19528), .ZN(n19952) );
  OAI21_X1 U17121 ( .B1(n19508), .B2(n19952), .A(n19475), .ZN(n14845) );
  NAND2_X1 U17122 ( .A1(n14846), .A2(n14845), .ZN(n14847) );
  NAND2_X1 U17123 ( .A1(n14848), .A2(n14847), .ZN(n19955) );
  INV_X1 U17124 ( .A(n19955), .ZN(n19525) );
  INV_X1 U17125 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14860) );
  INV_X1 U17126 ( .A(n19655), .ZN(n19644) );
  INV_X1 U17127 ( .A(n14849), .ZN(n14850) );
  NAND3_X1 U17128 ( .A1(n14851), .A2(n19508), .A3(n14850), .ZN(n14854) );
  OAI21_X1 U17129 ( .B1(n14852), .B2(n19952), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14853) );
  NAND2_X1 U17130 ( .A1(n14854), .A2(n14853), .ZN(n19954) );
  NOR2_X2 U17131 ( .A1(n14855), .A2(n19869), .ZN(n19651) );
  AOI22_X1 U17132 ( .A1(n19644), .A2(n19953), .B1(n19954), .B2(n19651), .ZN(
        n14859) );
  INV_X1 U17133 ( .A(n19492), .ZN(n14856) );
  AOI22_X1 U17134 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19875), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19876), .ZN(n19635) );
  INV_X1 U17135 ( .A(n19871), .ZN(n15030) );
  AOI22_X1 U17136 ( .A1(n19846), .A2(n19652), .B1(n19650), .B2(n19952), .ZN(
        n14858) );
  OAI211_X1 U17137 ( .C1(n19525), .C2(n14860), .A(n14859), .B(n14858), .ZN(
        P2_U3077) );
  INV_X1 U17138 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n14871) );
  INV_X1 U17139 ( .A(n14862), .ZN(n14863) );
  OAI211_X1 U17140 ( .C1(n11436), .C2(n14863), .A(n16457), .B(n14900), .ZN(
        n14870) );
  NAND2_X1 U17141 ( .A1(n14865), .A2(n14864), .ZN(n14868) );
  INV_X1 U17142 ( .A(n14866), .ZN(n14867) );
  AND2_X1 U17143 ( .A1(n14868), .A2(n14867), .ZN(n18544) );
  NAND2_X1 U17144 ( .A1(n18544), .A2(n16448), .ZN(n14869) );
  OAI211_X1 U17145 ( .C1(n16448), .C2(n14871), .A(n14870), .B(n14869), .ZN(
        P2_U2878) );
  XNOR2_X1 U17146 ( .A(n14900), .B(n14902), .ZN(n14875) );
  INV_X1 U17147 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n18553) );
  OAI21_X1 U17148 ( .B1(n14873), .B2(n14866), .A(n14872), .ZN(n18817) );
  MUX2_X1 U17149 ( .A(n18553), .B(n18817), .S(n16448), .Z(n14874) );
  OAI21_X1 U17150 ( .B1(n14875), .B2(n16474), .A(n14874), .ZN(P2_U2877) );
  INV_X1 U17151 ( .A(n15890), .ZN(n14881) );
  INV_X1 U17152 ( .A(n14876), .ZN(n14880) );
  INV_X1 U17153 ( .A(n21554), .ZN(n21481) );
  AOI21_X1 U17154 ( .B1(n21575), .B2(n21472), .A(n21481), .ZN(n21630) );
  INV_X1 U17155 ( .A(n16268), .ZN(n14877) );
  NOR3_X1 U17156 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14877), .A3(
        n21575), .ZN(n14878) );
  AOI21_X1 U17157 ( .B1(n21630), .B2(n21608), .A(n14878), .ZN(n14879) );
  AOI211_X1 U17158 ( .C1(n21625), .C2(n14881), .A(n14880), .B(n14879), .ZN(
        n14882) );
  OAI21_X1 U17159 ( .B1(n14883), .B2(n21635), .A(n14882), .ZN(P1_U3031) );
  NAND2_X1 U17160 ( .A1(n14886), .A2(n14885), .ZN(n14887) );
  AND2_X1 U17161 ( .A1(n14909), .A2(n14887), .ZN(n21680) );
  OR2_X1 U17162 ( .A1(n14889), .A2(n14888), .ZN(n14890) );
  NAND2_X1 U17163 ( .A1(n14912), .A2(n14890), .ZN(n21668) );
  OAI22_X1 U17164 ( .A1(n21668), .A2(n15952), .B1(n21683), .B2(n20136), .ZN(
        n14891) );
  AOI21_X1 U17165 ( .B1(n21680), .B2(n20132), .A(n14891), .ZN(n14892) );
  INV_X1 U17166 ( .A(n14892), .ZN(P1_U2868) );
  INV_X1 U17167 ( .A(n21680), .ZN(n14894) );
  OAI222_X1 U17168 ( .A1(n16023), .A2(n14894), .B1(n16015), .B2(n20045), .C1(
        n16014), .C2(n14893), .ZN(P1_U2900) );
  OR2_X1 U17169 ( .A1(n14896), .A2(n14895), .ZN(n14897) );
  AND2_X1 U17170 ( .A1(n14926), .A2(n14897), .ZN(n18570) );
  INV_X1 U17171 ( .A(n18570), .ZN(n14907) );
  INV_X1 U17172 ( .A(n14928), .ZN(n14904) );
  OAI21_X1 U17173 ( .B1(n14900), .B2(n14902), .A(n14901), .ZN(n14903) );
  NAND3_X1 U17174 ( .A1(n14904), .A2(n16457), .A3(n14903), .ZN(n14906) );
  NAND2_X1 U17175 ( .A1(n16433), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14905) );
  OAI211_X1 U17176 ( .C1(n14907), .C2(n16433), .A(n14906), .B(n14905), .ZN(
        P2_U2876) );
  AOI21_X1 U17177 ( .B1(n14910), .B2(n14909), .A(n14908), .ZN(n20168) );
  INV_X1 U17178 ( .A(n20168), .ZN(n21691) );
  INV_X1 U17179 ( .A(n14920), .ZN(n14911) );
  AOI21_X1 U17180 ( .B1(n14913), .B2(n14912), .A(n14911), .ZN(n21685) );
  AOI22_X1 U17181 ( .A1(n21685), .A2(n20131), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n15949), .ZN(n14914) );
  OAI21_X1 U17182 ( .B1(n21691), .B2(n15954), .A(n14914), .ZN(P1_U2867) );
  OAI222_X1 U17183 ( .A1(n16023), .A2(n21691), .B1(n16015), .B2(n13283), .C1(
        n16014), .C2(n14915), .ZN(P1_U2899) );
  OR2_X1 U17184 ( .A1(n14908), .A2(n14917), .ZN(n14918) );
  AND2_X1 U17185 ( .A1(n14916), .A2(n14918), .ZN(n21704) );
  NAND2_X1 U17186 ( .A1(n14920), .A2(n14919), .ZN(n14921) );
  NAND2_X1 U17187 ( .A1(n15116), .A2(n14921), .ZN(n21699) );
  OAI22_X1 U17188 ( .A1(n21699), .A2(n15952), .B1(n21700), .B2(n20136), .ZN(
        n14922) );
  AOI21_X1 U17189 ( .B1(n21704), .B2(n20132), .A(n14922), .ZN(n14923) );
  INV_X1 U17190 ( .A(n14923), .ZN(P1_U2866) );
  NAND2_X1 U17191 ( .A1(n14926), .A2(n14925), .ZN(n14927) );
  AND2_X1 U17192 ( .A1(n15080), .A2(n14927), .ZN(n18580) );
  INV_X1 U17193 ( .A(n18580), .ZN(n14933) );
  OAI211_X1 U17194 ( .C1(n14928), .C2(n14930), .A(n14929), .B(n16457), .ZN(
        n14932) );
  NAND2_X1 U17195 ( .A1(n16433), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14931) );
  OAI211_X1 U17196 ( .C1(n14933), .C2(n16433), .A(n14932), .B(n14931), .ZN(
        P2_U2875) );
  OR3_X1 U17197 ( .A1(n22018), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15046) );
  INV_X1 U17198 ( .A(n22035), .ZN(n22072) );
  NOR2_X1 U17199 ( .A1(n14939), .A2(n22050), .ZN(n14936) );
  NOR2_X1 U17200 ( .A1(n22029), .A2(n15046), .ZN(n14971) );
  INV_X1 U17201 ( .A(n14971), .ZN(n14934) );
  OAI21_X1 U17202 ( .B1(n14935), .B2(n21933), .A(n14934), .ZN(n14940) );
  NOR3_X1 U17203 ( .A1(n14936), .A2(n22043), .A3(n14940), .ZN(n14937) );
  AOI211_X2 U17204 ( .C1(n22043), .C2(n15046), .A(n22072), .B(n14937), .ZN(
        n14977) );
  INV_X1 U17205 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14945) );
  OR2_X1 U17206 ( .A1(n14667), .A2(n11025), .ZN(n22037) );
  INV_X1 U17207 ( .A(n22115), .ZN(n22111) );
  INV_X1 U17208 ( .A(n14940), .ZN(n14941) );
  OAI22_X1 U17209 ( .A1(n14941), .A2(n22043), .B1(n15046), .B2(n13234), .ZN(
        n14970) );
  AOI22_X1 U17210 ( .A1(n22107), .A2(n14971), .B1(n14970), .B2(n22106), .ZN(
        n14942) );
  OAI21_X1 U17211 ( .B1(n22334), .B2(n22111), .A(n14942), .ZN(n14943) );
  AOI21_X1 U17212 ( .B1(n14974), .B2(n22108), .A(n14943), .ZN(n14944) );
  OAI21_X1 U17213 ( .B1(n14977), .B2(n14945), .A(n14944), .ZN(P1_U3074) );
  INV_X1 U17214 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14949) );
  INV_X1 U17215 ( .A(n22301), .ZN(n22297) );
  AOI22_X1 U17216 ( .A1(n22293), .A2(n14971), .B1(n14970), .B2(n22292), .ZN(
        n14946) );
  OAI21_X1 U17217 ( .B1(n22334), .B2(n22297), .A(n14946), .ZN(n14947) );
  AOI21_X1 U17218 ( .B1(n14974), .B2(n22294), .A(n14947), .ZN(n14948) );
  OAI21_X1 U17219 ( .B1(n14977), .B2(n14949), .A(n14948), .ZN(P1_U3079) );
  INV_X1 U17220 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14953) );
  INV_X1 U17221 ( .A(n22264), .ZN(n22260) );
  AOI22_X1 U17222 ( .A1(n22256), .A2(n14971), .B1(n14970), .B2(n22255), .ZN(
        n14950) );
  OAI21_X1 U17223 ( .B1(n22334), .B2(n22260), .A(n14950), .ZN(n14951) );
  AOI21_X1 U17224 ( .B1(n14974), .B2(n22257), .A(n14951), .ZN(n14952) );
  OAI21_X1 U17225 ( .B1(n14977), .B2(n14953), .A(n14952), .ZN(P1_U3078) );
  INV_X1 U17226 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14957) );
  INV_X1 U17227 ( .A(n22152), .ZN(n22148) );
  AOI22_X1 U17228 ( .A1(n22144), .A2(n14971), .B1(n14970), .B2(n22143), .ZN(
        n14954) );
  OAI21_X1 U17229 ( .B1(n22334), .B2(n22148), .A(n14954), .ZN(n14955) );
  AOI21_X1 U17230 ( .B1(n14974), .B2(n22145), .A(n14955), .ZN(n14956) );
  OAI21_X1 U17231 ( .B1(n14977), .B2(n14957), .A(n14956), .ZN(P1_U3075) );
  INV_X1 U17232 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14961) );
  INV_X1 U17233 ( .A(n22227), .ZN(n22223) );
  AOI22_X1 U17234 ( .A1(n22219), .A2(n14971), .B1(n14970), .B2(n22218), .ZN(
        n14958) );
  OAI21_X1 U17235 ( .B1(n22334), .B2(n22223), .A(n14958), .ZN(n14959) );
  AOI21_X1 U17236 ( .B1(n14974), .B2(n22220), .A(n14959), .ZN(n14960) );
  OAI21_X1 U17237 ( .B1(n14977), .B2(n14961), .A(n14960), .ZN(P1_U3077) );
  INV_X1 U17238 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14965) );
  INV_X1 U17239 ( .A(n22189), .ZN(n22185) );
  AOI22_X1 U17240 ( .A1(n22181), .A2(n14971), .B1(n14970), .B2(n22180), .ZN(
        n14962) );
  OAI21_X1 U17241 ( .B1(n22334), .B2(n22185), .A(n14962), .ZN(n14963) );
  AOI21_X1 U17242 ( .B1(n14974), .B2(n22182), .A(n14963), .ZN(n14964) );
  OAI21_X1 U17243 ( .B1(n14977), .B2(n14965), .A(n14964), .ZN(P1_U3076) );
  INV_X1 U17244 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14969) );
  AOI22_X1 U17245 ( .A1(n22049), .A2(n14971), .B1(n14970), .B2(n22048), .ZN(
        n14966) );
  OAI21_X1 U17246 ( .B1(n22334), .B2(n22062), .A(n14966), .ZN(n14967) );
  AOI21_X1 U17247 ( .B1(n14974), .B2(n22059), .A(n14967), .ZN(n14968) );
  OAI21_X1 U17248 ( .B1(n14977), .B2(n14969), .A(n14968), .ZN(P1_U3073) );
  INV_X1 U17249 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14976) );
  INV_X1 U17250 ( .A(n22388), .ZN(n22382) );
  AOI22_X1 U17251 ( .A1(n22376), .A2(n14971), .B1(n14970), .B2(n22374), .ZN(
        n14972) );
  OAI21_X1 U17252 ( .B1(n22334), .B2(n22382), .A(n14972), .ZN(n14973) );
  AOI21_X1 U17253 ( .B1(n14974), .B2(n22377), .A(n14973), .ZN(n14975) );
  OAI21_X1 U17254 ( .B1(n14977), .B2(n14976), .A(n14975), .ZN(P1_U3080) );
  INV_X1 U17255 ( .A(n21704), .ZN(n14979) );
  OAI222_X1 U17256 ( .A1(n16023), .A2(n14979), .B1(n16015), .B2(n13290), .C1(
        n16014), .C2(n14978), .ZN(P1_U2898) );
  NAND2_X1 U17257 ( .A1(n17490), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19454) );
  INV_X1 U17258 ( .A(n19454), .ZN(n19456) );
  AOI22_X1 U17259 ( .A1(n19614), .A2(n17487), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19456), .ZN(n14984) );
  NOR2_X1 U17260 ( .A1(n14980), .A2(n19454), .ZN(n19900) );
  NOR2_X1 U17261 ( .A1(n14981), .A2(n19535), .ZN(n14982) );
  AOI211_X1 U17262 ( .C1(n19900), .C2(n19475), .A(n19511), .B(n14982), .ZN(
        n14983) );
  INV_X1 U17263 ( .A(n19903), .ZN(n15037) );
  INV_X1 U17264 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14992) );
  NAND2_X1 U17265 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19456), .ZN(
        n14987) );
  OAI21_X1 U17266 ( .B1(n14985), .B2(n19900), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14986) );
  OAI21_X1 U17267 ( .B1(n14987), .B2(n19532), .A(n14986), .ZN(n19901) );
  INV_X1 U17268 ( .A(n19531), .ZN(n15094) );
  INV_X1 U17269 ( .A(n19900), .ZN(n15033) );
  AOI22_X1 U17270 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19875), .ZN(n19426) );
  NOR2_X2 U17271 ( .A1(n19455), .A2(n19467), .ZN(n19902) );
  INV_X1 U17272 ( .A(n19546), .ZN(n19521) );
  AOI22_X1 U17273 ( .A1(n19908), .A2(n19543), .B1(n19902), .B2(n19521), .ZN(
        n14989) );
  OAI21_X1 U17274 ( .B1(n15094), .B2(n15033), .A(n14989), .ZN(n14990) );
  AOI21_X1 U17275 ( .B1(n19901), .B2(n14988), .A(n14990), .ZN(n14991) );
  OAI21_X1 U17276 ( .B1(n15037), .B2(n14992), .A(n14991), .ZN(P2_U3143) );
  MUX2_X1 U17277 ( .A(n12023), .B(n14993), .S(n15014), .Z(n17128) );
  NAND2_X1 U17278 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14995) );
  INV_X1 U17279 ( .A(n14995), .ZN(n14994) );
  MUX2_X1 U17280 ( .A(n14995), .B(n14994), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14996) );
  NOR2_X1 U17281 ( .A1(n14997), .A2(n14996), .ZN(n15007) );
  INV_X1 U17282 ( .A(n14998), .ZN(n15005) );
  INV_X1 U17283 ( .A(n14999), .ZN(n15000) );
  XNOR2_X1 U17284 ( .A(n15000), .B(n15008), .ZN(n15004) );
  AOI21_X1 U17285 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n15001), .A(
        n12054), .ZN(n21826) );
  INV_X1 U17286 ( .A(n15002), .ZN(n15003) );
  OAI22_X1 U17287 ( .A1(n15005), .A2(n15004), .B1(n21826), .B2(n15003), .ZN(
        n15006) );
  MUX2_X1 U17288 ( .A(n15008), .B(n21828), .S(n15014), .Z(n17129) );
  NOR3_X1 U17289 ( .A1(n17128), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n17129), 
        .ZN(n15020) );
  NOR2_X1 U17290 ( .A1(n17154), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n15015) );
  INV_X1 U17291 ( .A(n15015), .ZN(n15018) );
  INV_X1 U17292 ( .A(n15009), .ZN(n15017) );
  INV_X1 U17293 ( .A(n15010), .ZN(n22015) );
  NOR2_X1 U17294 ( .A1(n15011), .A2(n22015), .ZN(n15012) );
  XNOR2_X1 U17295 ( .A(n15012), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21670) );
  OAI21_X1 U17296 ( .B1(n21670), .B2(n12287), .A(n15014), .ZN(n15013) );
  OAI211_X1 U17297 ( .C1(n15014), .C2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n15013), .B(n17154), .ZN(n15016) );
  NAND2_X1 U17298 ( .A1(n15015), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n15021) );
  OAI211_X1 U17299 ( .C1(n15018), .C2(n15017), .A(n15016), .B(n15021), .ZN(
        n15019) );
  OR2_X1 U17300 ( .A1(n15020), .A2(n15019), .ZN(n17139) );
  NAND2_X1 U17301 ( .A1(n15021), .A2(n11823), .ZN(n15022) );
  NAND2_X1 U17302 ( .A1(n17139), .A2(n15022), .ZN(n15024) );
  AND2_X1 U17303 ( .A1(n15024), .A2(n21823), .ZN(n15023) );
  AND2_X1 U17304 ( .A1(n15024), .A2(n21834), .ZN(n21842) );
  INV_X1 U17305 ( .A(n13265), .ZN(n15026) );
  NAND2_X1 U17306 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22021), .ZN(n15038) );
  INV_X1 U17307 ( .A(n15038), .ZN(n15025) );
  OAI22_X1 U17308 ( .A1(n11025), .A2(n22043), .B1(n15026), .B2(n15025), .ZN(
        n15027) );
  OAI21_X1 U17309 ( .B1(n21842), .B2(n15027), .A(n17155), .ZN(n15028) );
  OAI21_X1 U17310 ( .B1(n17155), .B2(n22029), .A(n15028), .ZN(P1_U3478) );
  NOR2_X2 U17311 ( .A1(n15029), .A2(n19869), .ZN(n19805) );
  INV_X1 U17312 ( .A(n19802), .ZN(n15034) );
  AOI22_X1 U17313 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19875), .ZN(n19801) );
  INV_X1 U17314 ( .A(n19801), .ZN(n19804) );
  AOI22_X1 U17315 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19875), .ZN(n19791) );
  AOI22_X1 U17316 ( .A1(n19902), .A2(n19804), .B1(n19908), .B2(n19803), .ZN(
        n15032) );
  OAI21_X1 U17317 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15035) );
  AOI21_X1 U17318 ( .B1(n19901), .B2(n19805), .A(n15035), .ZN(n15036) );
  OAI21_X1 U17319 ( .B1(n15037), .B2(n14028), .A(n15036), .ZN(P2_U3138) );
  NAND2_X1 U17320 ( .A1(n17155), .A2(n15038), .ZN(n15713) );
  INV_X1 U17321 ( .A(n17155), .ZN(n15039) );
  NAND2_X1 U17322 ( .A1(n15039), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15042) );
  XNOR2_X1 U17323 ( .A(n15105), .B(n21952), .ZN(n15040) );
  NAND3_X1 U17324 ( .A1(n17155), .A2(n22077), .A3(n15040), .ZN(n15041) );
  OAI211_X1 U17325 ( .C1(n15713), .C2(n14536), .A(n15042), .B(n15041), .ZN(
        P1_U3476) );
  AOI21_X1 U17326 ( .B1(n22326), .B2(n15078), .A(n22050), .ZN(n15044) );
  AOI21_X1 U17327 ( .B1(n21966), .B2(n14582), .A(n15044), .ZN(n15045) );
  NOR2_X1 U17328 ( .A1(n15045), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15047) );
  NOR2_X1 U17329 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15046), .ZN(
        n15048) );
  NOR2_X1 U17330 ( .A1(n15049), .A2(n13234), .ZN(n21999) );
  NAND2_X1 U17331 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n15053) );
  INV_X1 U17332 ( .A(n15048), .ZN(n15074) );
  NOR2_X1 U17333 ( .A1(n22053), .A2(n22043), .ZN(n15050) );
  INV_X1 U17334 ( .A(n21979), .ZN(n21998) );
  AND2_X1 U17335 ( .A1(n15049), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22044) );
  AOI22_X1 U17336 ( .A1(n21966), .A2(n15050), .B1(n11469), .B2(n22044), .ZN(
        n15073) );
  OAI22_X1 U17337 ( .A1(n22299), .A2(n15074), .B1(n15073), .B2(n22298), .ZN(
        n15051) );
  AOI21_X1 U17338 ( .B1(n22201), .B2(n22294), .A(n15051), .ZN(n15052) );
  OAI211_X1 U17339 ( .C1(n15078), .C2(n22297), .A(n15053), .B(n15052), .ZN(
        P1_U3071) );
  NAND2_X1 U17340 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n15056) );
  OAI22_X1 U17341 ( .A1(n22225), .A2(n15074), .B1(n15073), .B2(n22224), .ZN(
        n15054) );
  AOI21_X1 U17342 ( .B1(n22201), .B2(n22220), .A(n15054), .ZN(n15055) );
  OAI211_X1 U17343 ( .C1(n15078), .C2(n22223), .A(n15056), .B(n15055), .ZN(
        P1_U3069) );
  NAND2_X1 U17344 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n15059) );
  OAI22_X1 U17345 ( .A1(n22187), .A2(n15074), .B1(n15073), .B2(n22186), .ZN(
        n15057) );
  AOI21_X1 U17346 ( .B1(n22201), .B2(n22182), .A(n15057), .ZN(n15058) );
  OAI211_X1 U17347 ( .C1(n15078), .C2(n22185), .A(n15059), .B(n15058), .ZN(
        P1_U3068) );
  NAND2_X1 U17348 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n15062) );
  OAI22_X1 U17349 ( .A1(n22262), .A2(n15074), .B1(n15073), .B2(n22261), .ZN(
        n15060) );
  AOI21_X1 U17350 ( .B1(n22201), .B2(n22257), .A(n15060), .ZN(n15061) );
  OAI211_X1 U17351 ( .C1(n15078), .C2(n22260), .A(n15062), .B(n15061), .ZN(
        P1_U3070) );
  NAND2_X1 U17352 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n15065) );
  OAI22_X1 U17353 ( .A1(n22070), .A2(n15074), .B1(n15073), .B2(n22069), .ZN(
        n15063) );
  AOI21_X1 U17354 ( .B1(n22201), .B2(n22059), .A(n15063), .ZN(n15064) );
  OAI211_X1 U17355 ( .C1(n15078), .C2(n22062), .A(n15065), .B(n15064), .ZN(
        P1_U3065) );
  NAND2_X1 U17356 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n15068) );
  OAI22_X1 U17357 ( .A1(n22386), .A2(n15074), .B1(n15073), .B2(n22383), .ZN(
        n15066) );
  AOI21_X1 U17358 ( .B1(n22201), .B2(n22377), .A(n15066), .ZN(n15067) );
  OAI211_X1 U17359 ( .C1(n15078), .C2(n22382), .A(n15068), .B(n15067), .ZN(
        P1_U3072) );
  NAND2_X1 U17360 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n15071) );
  OAI22_X1 U17361 ( .A1(n22150), .A2(n15074), .B1(n15073), .B2(n22149), .ZN(
        n15069) );
  AOI21_X1 U17362 ( .B1(n22201), .B2(n22145), .A(n15069), .ZN(n15070) );
  OAI211_X1 U17363 ( .C1(n15078), .C2(n22148), .A(n15071), .B(n15070), .ZN(
        P1_U3067) );
  NAND2_X1 U17364 ( .A1(n15072), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n15077) );
  OAI22_X1 U17365 ( .A1(n22113), .A2(n15074), .B1(n15073), .B2(n22112), .ZN(
        n15075) );
  AOI21_X1 U17366 ( .B1(n22201), .B2(n22108), .A(n15075), .ZN(n15076) );
  OAI211_X1 U17367 ( .C1(n15078), .C2(n22111), .A(n15077), .B(n15076), .ZN(
        P1_U3066) );
  AND2_X1 U17368 ( .A1(n15080), .A2(n15079), .ZN(n15082) );
  OR2_X1 U17369 ( .A1(n15082), .A2(n15081), .ZN(n16980) );
  INV_X1 U17370 ( .A(n14929), .ZN(n15086) );
  INV_X1 U17371 ( .A(n15083), .ZN(n15085) );
  OAI211_X1 U17372 ( .C1(n15086), .C2(n15085), .A(n16457), .B(n15140), .ZN(
        n15088) );
  NAND2_X1 U17373 ( .A1(n16433), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n15087) );
  OAI211_X1 U17374 ( .C1(n16980), .C2(n16433), .A(n15088), .B(n15087), .ZN(
        P2_U2874) );
  NOR2_X1 U17375 ( .A1(n19946), .A2(n19953), .ZN(n15089) );
  OAI21_X1 U17376 ( .B1(n15089), .B2(n14662), .A(n19508), .ZN(n15099) );
  INV_X1 U17377 ( .A(n15099), .ZN(n15093) );
  INV_X1 U17378 ( .A(n19442), .ZN(n19500) );
  NAND2_X1 U17379 ( .A1(n15090), .A2(n19500), .ZN(n19433) );
  OR2_X1 U17380 ( .A1(n19433), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15098) );
  NAND2_X1 U17381 ( .A1(n19432), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19510) );
  INV_X1 U17382 ( .A(n19510), .ZN(n19483) );
  NAND3_X1 U17383 ( .A1(n19483), .A2(n19488), .A3(n17485), .ZN(n15096) );
  AOI21_X1 U17384 ( .B1(n15096), .B2(n19532), .A(n19869), .ZN(n15091) );
  AOI21_X1 U17385 ( .B1(n12842), .B2(n15169), .A(n15091), .ZN(n15092) );
  INV_X1 U17386 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15102) );
  OAI22_X1 U17387 ( .A1(n19426), .A2(n19849), .B1(n15094), .B2(n15096), .ZN(
        n15095) );
  AOI21_X1 U17388 ( .B1(n19946), .B2(n19521), .A(n15095), .ZN(n15101) );
  INV_X1 U17389 ( .A(n15096), .ZN(n19945) );
  OAI21_X1 U17390 ( .B1(n12842), .B2(n19945), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15097) );
  OAI21_X1 U17391 ( .B1(n15099), .B2(n15098), .A(n15097), .ZN(n19947) );
  NAND2_X1 U17392 ( .A1(n19947), .A2(n14988), .ZN(n15100) );
  OAI211_X1 U17393 ( .C1(n19951), .C2(n15102), .A(n15101), .B(n15100), .ZN(
        P2_U3087) );
  INV_X1 U17394 ( .A(n15713), .ZN(n15103) );
  NAND2_X1 U17395 ( .A1(n15103), .A2(n14694), .ZN(n15111) );
  INV_X1 U17396 ( .A(n21952), .ZN(n15106) );
  AOI21_X1 U17397 ( .B1(n22042), .B2(n15106), .A(n22043), .ZN(n22074) );
  OAI21_X1 U17398 ( .B1(n15108), .B2(n21952), .A(n15107), .ZN(n15109) );
  NAND3_X1 U17399 ( .A1(n17155), .A2(n22074), .A3(n15109), .ZN(n15110) );
  OAI211_X1 U17400 ( .C1(n12225), .C2(n17155), .A(n15111), .B(n15110), .ZN(
        P1_U3475) );
  INV_X1 U17401 ( .A(n15112), .ZN(n15113) );
  AOI21_X1 U17402 ( .B1(n15114), .B2(n14916), .A(n15113), .ZN(n20180) );
  INV_X1 U17403 ( .A(n15126), .ZN(n15118) );
  NAND2_X1 U17404 ( .A1(n15116), .A2(n15115), .ZN(n15117) );
  NAND2_X1 U17405 ( .A1(n15118), .A2(n15117), .ZN(n21711) );
  OAI22_X1 U17406 ( .A1(n21711), .A2(n15952), .B1(n15119), .B2(n20136), .ZN(
        n15120) );
  AOI21_X1 U17407 ( .B1(n20180), .B2(n20132), .A(n15120), .ZN(n15121) );
  INV_X1 U17408 ( .A(n15121), .ZN(P1_U2865) );
  XNOR2_X1 U17409 ( .A(n15112), .B(n15122), .ZN(n21726) );
  INV_X1 U17410 ( .A(n21726), .ZN(n15124) );
  AOI22_X1 U17411 ( .A1(n16021), .A2(n15980), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16019), .ZN(n15123) );
  OAI21_X1 U17412 ( .B1(n15124), .B2(n16023), .A(n15123), .ZN(P1_U2896) );
  OR2_X1 U17413 ( .A1(n15126), .A2(n15125), .ZN(n15127) );
  NAND2_X1 U17414 ( .A1(n15135), .A2(n15127), .ZN(n21722) );
  OAI22_X1 U17415 ( .A1(n21722), .A2(n15952), .B1(n21723), .B2(n20136), .ZN(
        n15128) );
  AOI21_X1 U17416 ( .B1(n21726), .B2(n20132), .A(n15128), .ZN(n15129) );
  INV_X1 U17417 ( .A(n15129), .ZN(P1_U2864) );
  INV_X1 U17418 ( .A(n20180), .ZN(n21713) );
  OAI222_X1 U17419 ( .A1(n16023), .A2(n21713), .B1(n16015), .B2(n13294), .C1(
        n16014), .C2(n15130), .ZN(P1_U2897) );
  NOR2_X1 U17420 ( .A1(n11085), .A2(n15131), .ZN(n15132) );
  OR2_X1 U17421 ( .A1(n11043), .A2(n15132), .ZN(n21738) );
  INV_X1 U17422 ( .A(n15156), .ZN(n15133) );
  AOI21_X1 U17423 ( .B1(n15135), .B2(n15134), .A(n15133), .ZN(n21736) );
  AOI22_X1 U17424 ( .A1(n21736), .A2(n20131), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n15949), .ZN(n15136) );
  OAI21_X1 U17425 ( .B1(n21738), .B2(n15954), .A(n15136), .ZN(P1_U2863) );
  AOI22_X1 U17426 ( .A1(n16021), .A2(n15976), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n16019), .ZN(n15137) );
  OAI21_X1 U17427 ( .B1(n21738), .B2(n16023), .A(n15137), .ZN(P1_U2895) );
  NOR2_X1 U17428 ( .A1(n15081), .A2(n15138), .ZN(n15139) );
  OR2_X1 U17429 ( .A1(n15229), .A2(n15139), .ZN(n17471) );
  NAND2_X1 U17430 ( .A1(n15143), .A2(n15142), .ZN(n15188) );
  OAI211_X1 U17431 ( .C1(n15143), .C2(n15142), .A(n16457), .B(n15144), .ZN(
        n15146) );
  NAND2_X1 U17432 ( .A1(n16433), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15145) );
  OAI211_X1 U17433 ( .C1(n17471), .C2(n16433), .A(n15146), .B(n15145), .ZN(
        P2_U2873) );
  OAI21_X1 U17434 ( .B1(n11043), .B2(n15148), .A(n15147), .ZN(n15184) );
  AOI22_X1 U17435 ( .A1(n16021), .A2(n15972), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n16019), .ZN(n15149) );
  OAI21_X1 U17436 ( .B1(n15184), .B2(n16023), .A(n15149), .ZN(P1_U2894) );
  NOR2_X1 U17437 ( .A1(n15335), .A2(n21804), .ZN(n15260) );
  INV_X1 U17438 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15153) );
  NAND2_X1 U17439 ( .A1(n15150), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15151) );
  NOR3_X2 U17440 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21720), .A3(n22043), 
        .ZN(n21769) );
  AOI21_X1 U17441 ( .B1(n21816), .B2(n20186), .A(n21769), .ZN(n15152) );
  OAI21_X1 U17442 ( .B1(n15153), .B2(n21820), .A(n15152), .ZN(n15162) );
  INV_X1 U17443 ( .A(n15154), .ZN(n15258) );
  NAND2_X1 U17444 ( .A1(n15156), .A2(n15155), .ZN(n15157) );
  NAND2_X1 U17445 ( .A1(n15258), .A2(n15157), .ZN(n21548) );
  NOR2_X1 U17446 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n21732), .ZN(n15158) );
  AOI22_X1 U17447 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n21810), .B1(n15159), 
        .B2(n15158), .ZN(n15160) );
  OAI21_X1 U17448 ( .B1(n21812), .B2(n21548), .A(n15160), .ZN(n15161) );
  AOI211_X1 U17449 ( .C1(n15260), .C2(P1_REIP_REG_10__SCAN_IN), .A(n15162), 
        .B(n15161), .ZN(n15163) );
  OAI21_X1 U17450 ( .B1(n15184), .B2(n21813), .A(n15163), .ZN(P1_U2830) );
  NOR2_X2 U17451 ( .A1(n19539), .A2(n19414), .ZN(n19978) );
  OAI21_X1 U17452 ( .B1(n19975), .B2(n19978), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15164) );
  NAND2_X1 U17453 ( .A1(n15164), .A2(n19508), .ZN(n15168) );
  NAND2_X1 U17454 ( .A1(n15165), .A2(n19488), .ZN(n19537) );
  NOR2_X1 U17455 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19537), .ZN(
        n19974) );
  OAI21_X1 U17456 ( .B1(n15170), .B2(n19974), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15167) );
  INV_X1 U17457 ( .A(n19974), .ZN(n15166) );
  AND2_X1 U17458 ( .A1(n19400), .A2(n15166), .ZN(n15173) );
  INV_X1 U17459 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19473) );
  AOI22_X1 U17460 ( .A1(n15168), .A2(n15167), .B1(n15173), .B2(n19473), .ZN(
        n19979) );
  INV_X1 U17461 ( .A(n15168), .ZN(n15174) );
  AOI21_X1 U17462 ( .B1(n19974), .B2(n19475), .A(n19511), .ZN(n15172) );
  NAND2_X1 U17463 ( .A1(n15170), .A2(n15169), .ZN(n15171) );
  AOI22_X1 U17464 ( .A1(n19644), .A2(n19978), .B1(n19974), .B2(n19650), .ZN(
        n15176) );
  NAND2_X1 U17465 ( .A1(n19975), .A2(n19652), .ZN(n15175) );
  OAI211_X1 U17466 ( .C1(n19984), .C2(n15469), .A(n15176), .B(n15175), .ZN(
        n15177) );
  AOI21_X1 U17467 ( .B1(n19979), .B2(n19651), .A(n15177), .ZN(n15178) );
  INV_X1 U17468 ( .A(n15178), .ZN(P2_U3053) );
  AOI22_X1 U17469 ( .A1(n19521), .A2(n19978), .B1(n19531), .B2(n19974), .ZN(
        n15180) );
  NAND2_X1 U17470 ( .A1(n19975), .A2(n19543), .ZN(n15179) );
  OAI211_X1 U17471 ( .C1(n19984), .C2(n15181), .A(n15180), .B(n15179), .ZN(
        n15182) );
  AOI21_X1 U17472 ( .B1(n14988), .B2(n19979), .A(n15182), .ZN(n15183) );
  INV_X1 U17473 ( .A(n15183), .ZN(P2_U3055) );
  INV_X1 U17474 ( .A(n15184), .ZN(n20187) );
  OAI22_X1 U17475 ( .A1(n21548), .A2(n15952), .B1(n15185), .B2(n20136), .ZN(
        n15186) );
  AOI21_X1 U17476 ( .B1(n20187), .B2(n20132), .A(n15186), .ZN(n15187) );
  INV_X1 U17477 ( .A(n15187), .ZN(P1_U2862) );
  NAND2_X1 U17478 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n15192) );
  AOI22_X1 U17479 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U17480 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15190) );
  NAND2_X1 U17481 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n15189) );
  AND4_X1 U17482 ( .A1(n15192), .A2(n15191), .A3(n15190), .A4(n15189), .ZN(
        n15195) );
  AOI22_X1 U17483 ( .A1(n15504), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12793), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U17484 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n15193) );
  NAND3_X1 U17485 ( .A1(n15195), .A2(n15194), .A3(n15193), .ZN(n15201) );
  AOI22_X1 U17486 ( .A1(n15509), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15508), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15199) );
  AOI22_X1 U17487 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15198) );
  AOI22_X1 U17488 ( .A1(n15512), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U17489 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n15196) );
  NAND4_X1 U17490 ( .A1(n15199), .A2(n15198), .A3(n15197), .A4(n15196), .ZN(
        n15200) );
  NAND2_X1 U17491 ( .A1(n15202), .A2(n15204), .ZN(n15283) );
  OAI21_X1 U17492 ( .B1(n15202), .B2(n15204), .A(n15203), .ZN(n16567) );
  NAND2_X1 U17493 ( .A1(n15227), .A2(n15205), .ZN(n15206) );
  NAND2_X1 U17494 ( .A1(n15267), .A2(n15206), .ZN(n16717) );
  NOR2_X1 U17495 ( .A1(n16717), .A2(n16433), .ZN(n15207) );
  AOI21_X1 U17496 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n16433), .A(n15207), .ZN(
        n15208) );
  OAI21_X1 U17497 ( .B1(n16567), .B2(n16474), .A(n15208), .ZN(P2_U2871) );
  NAND2_X1 U17498 ( .A1(n15210), .A2(n15209), .ZN(n15211) );
  XNOR2_X1 U17499 ( .A(n15212), .B(n15211), .ZN(n17410) );
  XNOR2_X1 U17500 ( .A(n15214), .B(n15213), .ZN(n17409) );
  INV_X1 U17501 ( .A(n17409), .ZN(n15225) );
  INV_X1 U17502 ( .A(n18876), .ZN(n18846) );
  NAND3_X1 U17503 ( .A1(n18847), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18846), .ZN(n18845) );
  AOI221_X1 U17504 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n18844), .C2(n15215), .A(
        n18845), .ZN(n15224) );
  INV_X1 U17505 ( .A(n16912), .ZN(n18875) );
  NOR2_X1 U17506 ( .A1(n16917), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18865) );
  OAI21_X1 U17507 ( .B1(n16917), .B2(n18864), .A(n18804), .ZN(n18874) );
  AOI211_X1 U17508 ( .C1(n18876), .C2(n18875), .A(n18865), .B(n18874), .ZN(
        n18859) );
  OAI21_X1 U17509 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17047), .A(
        n18859), .ZN(n18834) );
  NAND2_X1 U17510 ( .A1(n18834), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15222) );
  OR2_X1 U17511 ( .A1(n15433), .A2(n15216), .ZN(n15217) );
  AND2_X1 U17512 ( .A1(n14475), .A2(n15217), .ZN(n18503) );
  XNOR2_X1 U17513 ( .A(n15218), .B(n18479), .ZN(n19619) );
  OAI22_X1 U17514 ( .A1(n18870), .A2(n19619), .B1(n18848), .B2(n15219), .ZN(
        n15220) );
  AOI21_X1 U17515 ( .B1(n18503), .B2(n14189), .A(n15220), .ZN(n15221) );
  NAND2_X1 U17516 ( .A1(n15222), .A2(n15221), .ZN(n15223) );
  AOI211_X1 U17517 ( .C1(n15225), .C2(n18856), .A(n15224), .B(n15223), .ZN(
        n15226) );
  OAI21_X1 U17518 ( .B1(n18881), .B2(n17410), .A(n15226), .ZN(P2_U3041) );
  OAI21_X1 U17519 ( .B1(n15229), .B2(n15228), .A(n15227), .ZN(n16946) );
  NOR2_X1 U17520 ( .A1(n16946), .A2(n16433), .ZN(n15232) );
  AOI211_X1 U17521 ( .C1(n15230), .C2(n15144), .A(n16474), .B(n15202), .ZN(
        n15231) );
  AOI211_X1 U17522 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n16433), .A(n15232), .B(
        n15231), .ZN(n15233) );
  INV_X1 U17523 ( .A(n15233), .ZN(P2_U2872) );
  XNOR2_X1 U17524 ( .A(n15235), .B(n15234), .ZN(n17419) );
  NAND2_X1 U17525 ( .A1(n15236), .A2(n15249), .ZN(n17416) );
  NAND3_X1 U17526 ( .A1(n17416), .A2(n18825), .A3(n17415), .ZN(n15252) );
  INV_X1 U17527 ( .A(n15237), .ZN(n15250) );
  INV_X1 U17528 ( .A(n18514), .ZN(n15247) );
  INV_X1 U17529 ( .A(n16917), .ZN(n16872) );
  INV_X1 U17530 ( .A(n18804), .ZN(n17052) );
  AOI21_X1 U17531 ( .B1(n16872), .B2(n15238), .A(n17052), .ZN(n15308) );
  OAI21_X1 U17532 ( .B1(n15239), .B2(n16912), .A(n15308), .ZN(n15240) );
  NAND2_X1 U17533 ( .A1(n15240), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15246) );
  XNOR2_X1 U17534 ( .A(n15242), .B(n15241), .ZN(n19558) );
  INV_X1 U17535 ( .A(n19558), .ZN(n15244) );
  NOR2_X1 U17536 ( .A1(n13049), .A2(n18848), .ZN(n15243) );
  AOI21_X1 U17537 ( .B1(n18852), .B2(n15244), .A(n15243), .ZN(n15245) );
  OAI211_X1 U17538 ( .C1(n15247), .C2(n18849), .A(n15246), .B(n15245), .ZN(
        n15248) );
  AOI21_X1 U17539 ( .B1(n15250), .B2(n15249), .A(n15248), .ZN(n15251) );
  OAI211_X1 U17540 ( .C1(n17419), .C2(n18869), .A(n15252), .B(n15251), .ZN(
        P2_U3040) );
  XOR2_X1 U17541 ( .A(n15254), .B(n15253), .Z(n20195) );
  INV_X1 U17542 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20078) );
  INV_X1 U17543 ( .A(n15256), .ZN(n15259) );
  AOI21_X1 U17544 ( .B1(n15259), .B2(n15258), .A(n15257), .ZN(n21565) );
  INV_X1 U17545 ( .A(n21565), .ZN(n15296) );
  OAI22_X1 U17546 ( .A1(n15296), .A2(n21812), .B1(n20193), .B2(n21795), .ZN(
        n15264) );
  AOI22_X1 U17547 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n21810), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n15260), .ZN(n15261) );
  INV_X1 U17548 ( .A(n21769), .ZN(n21686) );
  OAI211_X1 U17549 ( .C1(n21820), .C2(n15262), .A(n15261), .B(n21686), .ZN(
        n15263) );
  AOI211_X1 U17550 ( .C1(n15857), .C2(n20078), .A(n15264), .B(n15263), .ZN(
        n15265) );
  OAI21_X1 U17551 ( .B1(n15297), .B2(n21813), .A(n15265), .ZN(P1_U2829) );
  NAND2_X1 U17552 ( .A1(n15267), .A2(n15266), .ZN(n15268) );
  AND2_X1 U17553 ( .A1(n15347), .A2(n15268), .ZN(n18628) );
  INV_X1 U17554 ( .A(n18628), .ZN(n16926) );
  AOI22_X1 U17555 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n15509), .B1(
        n15508), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15272) );
  AOI22_X1 U17556 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15271) );
  AOI22_X1 U17557 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n15512), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15270) );
  NAND2_X1 U17558 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n15269) );
  AND4_X1 U17559 ( .A1(n15272), .A2(n15271), .A3(n15270), .A4(n15269), .ZN(
        n15282) );
  INV_X1 U17560 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19858) );
  NAND2_X1 U17561 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n15274) );
  NAND2_X1 U17562 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n15273) );
  OAI211_X1 U17563 ( .C1(n15484), .C2(n19858), .A(n15274), .B(n15273), .ZN(
        n15280) );
  NAND2_X1 U17564 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n15278) );
  AOI22_X1 U17565 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12479), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15277) );
  AOI22_X1 U17566 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n15498), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15276) );
  NAND2_X1 U17567 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n15275) );
  NAND4_X1 U17568 ( .A1(n15278), .A2(n15277), .A3(n15276), .A4(n15275), .ZN(
        n15279) );
  NOR2_X1 U17569 ( .A1(n15280), .A2(n15279), .ZN(n15281) );
  AND2_X1 U17570 ( .A1(n15282), .A2(n15281), .ZN(n15285) );
  INV_X1 U17571 ( .A(n15285), .ZN(n15284) );
  AOI21_X1 U17572 ( .B1(n15285), .B2(n15203), .A(n11448), .ZN(n16559) );
  NAND2_X1 U17573 ( .A1(n16559), .A2(n16457), .ZN(n15287) );
  NAND2_X1 U17574 ( .A1(n16433), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15286) );
  OAI211_X1 U17575 ( .C1(n16926), .C2(n16433), .A(n15287), .B(n15286), .ZN(
        P2_U2870) );
  OAI21_X1 U17576 ( .B1(n15290), .B2(n15289), .A(n15288), .ZN(n21520) );
  INV_X1 U17577 ( .A(n21725), .ZN(n15292) );
  AOI22_X1 U17578 ( .A1(n20230), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n21639), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15291) );
  OAI21_X1 U17579 ( .B1(n20240), .B2(n15292), .A(n15291), .ZN(n15293) );
  AOI21_X1 U17580 ( .B1(n21726), .B2(n20236), .A(n15293), .ZN(n15294) );
  OAI21_X1 U17581 ( .B1(n21520), .B2(n21822), .A(n15294), .ZN(P1_U2991) );
  INV_X1 U17582 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15295) );
  OAI222_X1 U17583 ( .A1(n15296), .A2(n15952), .B1(n15954), .B2(n15297), .C1(
        n15295), .C2(n20136), .ZN(P1_U2861) );
  INV_X1 U17584 ( .A(n15968), .ZN(n15298) );
  OAI222_X1 U17585 ( .A1(n16014), .A2(n15298), .B1(n16023), .B2(n15297), .C1(
        n20057), .C2(n16015), .ZN(P1_U2893) );
  AND2_X1 U17586 ( .A1(n15299), .A2(n15300), .ZN(n17424) );
  INV_X1 U17587 ( .A(n17424), .ZN(n15303) );
  INV_X1 U17588 ( .A(n15300), .ZN(n15301) );
  NOR2_X1 U17589 ( .A1(n15301), .A2(n17423), .ZN(n15302) );
  OAI22_X1 U17590 ( .A1(n15303), .A2(n17423), .B1(n15302), .B2(n15299), .ZN(
        n15326) );
  OR2_X1 U17591 ( .A1(n15305), .A2(n15304), .ZN(n15307) );
  NAND2_X1 U17592 ( .A1(n15307), .A2(n15306), .ZN(n19396) );
  OAI21_X1 U17593 ( .B1(n15309), .B2(n16912), .A(n15308), .ZN(n18823) );
  NAND2_X1 U17594 ( .A1(n18823), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15312) );
  AOI22_X1 U17595 ( .A1(n16675), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n18829), 
        .B2(n15310), .ZN(n15311) );
  OAI211_X1 U17596 ( .C1(n18870), .C2(n19396), .A(n15312), .B(n15311), .ZN(
        n15313) );
  AOI21_X1 U17597 ( .B1(n18524), .B2(n14189), .A(n15313), .ZN(n15318) );
  OR2_X1 U17598 ( .A1(n15315), .A2(n15314), .ZN(n15319) );
  NAND3_X1 U17599 ( .A1(n15319), .A2(n18825), .A3(n15316), .ZN(n15317) );
  OAI211_X1 U17600 ( .C1(n15326), .C2(n18869), .A(n15318), .B(n15317), .ZN(
        P2_U3039) );
  NAND3_X1 U17601 ( .A1(n15319), .A2(n17473), .A3(n15316), .ZN(n15325) );
  AOI21_X1 U17602 ( .B1(n15320), .B2(n16296), .A(n16299), .ZN(n18518) );
  OAI22_X1 U17603 ( .A1(n15320), .A2(n17459), .B1(n13056), .B2(n18848), .ZN(
        n15323) );
  NOR2_X1 U17604 ( .A1(n15321), .A2(n17449), .ZN(n15322) );
  AOI211_X1 U17605 ( .C1(n17453), .C2(n18518), .A(n15323), .B(n15322), .ZN(
        n15324) );
  OAI211_X1 U17606 ( .C1(n15326), .C2(n17461), .A(n15325), .B(n15324), .ZN(
        P2_U3007) );
  OR2_X1 U17607 ( .A1(n15329), .A2(n15328), .ZN(n15330) );
  AND2_X1 U17608 ( .A1(n15327), .A2(n15330), .ZN(n20204) );
  OR2_X1 U17609 ( .A1(n15257), .A2(n15331), .ZN(n15332) );
  NAND2_X1 U17610 ( .A1(n15865), .A2(n15332), .ZN(n21564) );
  OAI22_X1 U17611 ( .A1(n21564), .A2(n15952), .B1(n15337), .B2(n20136), .ZN(
        n15333) );
  AOI21_X1 U17612 ( .B1(n20204), .B2(n20132), .A(n15333), .ZN(n15334) );
  INV_X1 U17613 ( .A(n15334), .ZN(P1_U2860) );
  INV_X1 U17614 ( .A(n20204), .ZN(n15346) );
  INV_X1 U17615 ( .A(n20202), .ZN(n15343) );
  NAND2_X1 U17616 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15857), .ZN(n15341) );
  INV_X1 U17617 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15340) );
  INV_X1 U17618 ( .A(n15335), .ZN(n15336) );
  OAI21_X1 U17619 ( .B1(n15336), .B2(n15859), .A(n21781), .ZN(n15860) );
  OAI22_X1 U17620 ( .A1(n15337), .A2(n21765), .B1(n21812), .B2(n21564), .ZN(
        n15338) );
  AOI211_X1 U17621 ( .C1(n21792), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21769), .B(n15338), .ZN(n15339) );
  OAI221_X1 U17622 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n15341), .C1(n15340), 
        .C2(n15860), .A(n15339), .ZN(n15342) );
  AOI21_X1 U17623 ( .B1(n21816), .B2(n15343), .A(n15342), .ZN(n15344) );
  OAI21_X1 U17624 ( .B1(n15346), .B2(n21813), .A(n15344), .ZN(P1_U2828) );
  AOI22_X1 U17625 ( .A1(n16021), .A2(n15964), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n16019), .ZN(n15345) );
  OAI21_X1 U17626 ( .B1(n15346), .B2(n16023), .A(n15345), .ZN(P1_U2892) );
  AOI21_X1 U17627 ( .B1(n15348), .B2(n15347), .A(n16471), .ZN(n16704) );
  INV_X1 U17628 ( .A(n16704), .ZN(n18641) );
  AOI22_X1 U17629 ( .A1(n15509), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15508), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15352) );
  AOI22_X1 U17630 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15351) );
  AOI22_X1 U17631 ( .A1(n15512), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15350) );
  NAND2_X1 U17632 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n15349) );
  AND4_X1 U17633 ( .A1(n15352), .A2(n15351), .A3(n15350), .A4(n15349), .ZN(
        n15362) );
  NAND2_X1 U17634 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n15354) );
  NAND2_X1 U17635 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n15353) );
  OAI211_X1 U17636 ( .C1(n15484), .C2(n19808), .A(n15354), .B(n15353), .ZN(
        n15360) );
  NAND2_X1 U17637 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n15358) );
  AOI22_X1 U17638 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15357) );
  AOI22_X1 U17639 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15356) );
  NAND2_X1 U17640 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n15355) );
  NAND4_X1 U17641 ( .A1(n15358), .A2(n15357), .A3(n15356), .A4(n15355), .ZN(
        n15359) );
  NOR2_X1 U17642 ( .A1(n15360), .A2(n15359), .ZN(n15361) );
  AOI21_X1 U17643 ( .B1(n15364), .B2(n15363), .A(n15449), .ZN(n19767) );
  NAND2_X1 U17644 ( .A1(n19767), .A2(n16457), .ZN(n15366) );
  NAND2_X1 U17645 ( .A1(n16433), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15365) );
  OAI211_X1 U17646 ( .C1(n18641), .C2(n16433), .A(n15366), .B(n15365), .ZN(
        P2_U2869) );
  NOR2_X1 U17647 ( .A1(n21438), .A2(n15367), .ZN(n21424) );
  AOI211_X1 U17648 ( .C1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n21013), .A(
        n17771), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17973) );
  INV_X1 U17649 ( .A(n17973), .ZN(n15368) );
  NAND2_X1 U17650 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18306) );
  NAND2_X1 U17651 ( .A1(n20319), .A2(n18306), .ZN(n15369) );
  OAI21_X1 U17652 ( .B1(n18980), .B2(n21426), .A(n15369), .ZN(n18353) );
  INV_X1 U17653 ( .A(n18353), .ZN(n15370) );
  NOR2_X1 U17654 ( .A1(n18356), .A2(n15370), .ZN(n15372) );
  INV_X1 U17655 ( .A(n18976), .ZN(n17076) );
  NAND2_X1 U17656 ( .A1(n18980), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17975) );
  INV_X1 U17657 ( .A(n17975), .ZN(n18942) );
  OR3_X1 U17658 ( .A1(n17076), .A2(n18942), .A3(n18356), .ZN(n15371) );
  MUX2_X1 U17659 ( .A(n15372), .B(n15371), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AOI21_X1 U17660 ( .B1(n21013), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15374) );
  OR2_X1 U17661 ( .A1(n15374), .A2(n15373), .ZN(n21406) );
  NAND2_X1 U17662 ( .A1(n18347), .A2(n21426), .ZN(n20996) );
  NOR2_X1 U17663 ( .A1(n21406), .A2(n20996), .ZN(n15379) );
  OAI211_X1 U17664 ( .C1(n17091), .C2(n20781), .A(n21405), .B(n21907), .ZN(
        n15376) );
  OAI211_X1 U17665 ( .C1(n21385), .C2(n17574), .A(n15377), .B(n15376), .ZN(
        n21412) );
  INV_X1 U17666 ( .A(n21412), .ZN(n21393) );
  NAND2_X1 U17667 ( .A1(n21438), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18940) );
  NAND2_X1 U17668 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n21424), .ZN(n15378) );
  OAI211_X1 U17669 ( .C1(n21414), .C2(n21393), .A(n18940), .B(n15378), .ZN(
        n21027) );
  INV_X1 U17670 ( .A(n21027), .ZN(n21030) );
  MUX2_X1 U17671 ( .A(n15379), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n21030), .Z(P3_U3284) );
  NOR2_X1 U17672 ( .A1(n15380), .A2(n11008), .ZN(n15381) );
  AOI21_X1 U17673 ( .B1(n10986), .B2(n15382), .A(n15381), .ZN(n17120) );
  OAI21_X1 U17674 ( .B1(n17120), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n17154), 
        .ZN(n15384) );
  AOI22_X1 U17675 ( .A1(n15384), .A2(n15383), .B1(n15385), .B2(n21839), .ZN(
        n15388) );
  AOI21_X1 U17676 ( .B1(n17118), .B2(n17081), .A(n15387), .ZN(n15386) );
  OAI22_X1 U17677 ( .A1(n15388), .A2(n15387), .B1(n15386), .B2(n15385), .ZN(
        P1_U3474) );
  NAND3_X1 U17678 ( .A1(n17118), .A2(n15390), .A3(n15389), .ZN(n15391) );
  NAND2_X1 U17679 ( .A1(n20035), .A2(n11027), .ZN(n15422) );
  INV_X1 U17680 ( .A(n21834), .ZN(n17152) );
  NOR2_X4 U17681 ( .A1(n20035), .A2(n21456), .ZN(n20060) );
  AOI22_X1 U17682 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20053), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20060), .ZN(n15393) );
  OAI21_X1 U17683 ( .B1(n15394), .B2(n15422), .A(n15393), .ZN(P1_U2920) );
  AOI22_X1 U17684 ( .A1(n21456), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n15395) );
  OAI21_X1 U17685 ( .B1(n15396), .B2(n15422), .A(n15395), .ZN(P1_U2919) );
  AOI22_X1 U17686 ( .A1(n21456), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n15397) );
  OAI21_X1 U17687 ( .B1(n15398), .B2(n15422), .A(n15397), .ZN(P1_U2918) );
  AOI22_X1 U17688 ( .A1(n21456), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15399) );
  OAI21_X1 U17689 ( .B1(n15400), .B2(n15422), .A(n15399), .ZN(P1_U2917) );
  AOI22_X1 U17690 ( .A1(n21456), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15401) );
  OAI21_X1 U17691 ( .B1(n15402), .B2(n15422), .A(n15401), .ZN(P1_U2916) );
  AOI22_X1 U17692 ( .A1(n21456), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15403) );
  OAI21_X1 U17693 ( .B1(n15404), .B2(n15422), .A(n15403), .ZN(P1_U2915) );
  AOI22_X1 U17694 ( .A1(n21456), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n15405) );
  OAI21_X1 U17695 ( .B1(n15406), .B2(n15422), .A(n15405), .ZN(P1_U2914) );
  AOI22_X1 U17696 ( .A1(n21456), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n15407) );
  OAI21_X1 U17697 ( .B1(n15408), .B2(n15422), .A(n15407), .ZN(P1_U2913) );
  AOI22_X1 U17698 ( .A1(n21456), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n15409) );
  OAI21_X1 U17699 ( .B1(n15410), .B2(n15422), .A(n15409), .ZN(P1_U2912) );
  AOI22_X1 U17700 ( .A1(n21456), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n15411) );
  OAI21_X1 U17701 ( .B1(n15412), .B2(n15422), .A(n15411), .ZN(P1_U2911) );
  AOI22_X1 U17702 ( .A1(n21456), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n15413) );
  OAI21_X1 U17703 ( .B1(n15414), .B2(n15422), .A(n15413), .ZN(P1_U2910) );
  AOI22_X1 U17704 ( .A1(n21456), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15415) );
  OAI21_X1 U17705 ( .B1(n15416), .B2(n15422), .A(n15415), .ZN(P1_U2909) );
  AOI22_X1 U17706 ( .A1(n21456), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15417) );
  OAI21_X1 U17707 ( .B1(n15418), .B2(n15422), .A(n15417), .ZN(P1_U2908) );
  AOI22_X1 U17708 ( .A1(n21456), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15419) );
  OAI21_X1 U17709 ( .B1(n15420), .B2(n15422), .A(n15419), .ZN(P1_U2907) );
  AOI22_X1 U17710 ( .A1(n21456), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15421) );
  OAI21_X1 U17711 ( .B1(n15423), .B2(n15422), .A(n15421), .ZN(P1_U2906) );
  XOR2_X1 U17712 ( .A(n14473), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n15426)
         );
  NAND2_X1 U17713 ( .A1(n16433), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n15425) );
  NAND2_X1 U17714 ( .A1(n18503), .A2(n16448), .ZN(n15424) );
  OAI211_X1 U17715 ( .C1(n15426), .C2(n16474), .A(n15425), .B(n15424), .ZN(
        P2_U2882) );
  OR2_X1 U17716 ( .A1(n15428), .A2(n15427), .ZN(n15429) );
  NAND2_X1 U17717 ( .A1(n14473), .A2(n15429), .ZN(n19665) );
  NOR2_X1 U17718 ( .A1(n15431), .A2(n15430), .ZN(n15432) );
  OR2_X1 U17719 ( .A1(n15433), .A2(n15432), .ZN(n18484) );
  MUX2_X1 U17720 ( .A(n18484), .B(n15434), .S(n16433), .Z(n15435) );
  OAI21_X1 U17721 ( .B1(n19665), .B2(n16474), .A(n15435), .ZN(P2_U2883) );
  NAND2_X1 U17722 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n15439) );
  AOI22_X1 U17723 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15438) );
  AOI22_X1 U17724 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15437) );
  NAND2_X1 U17725 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n15436) );
  AND4_X1 U17726 ( .A1(n15439), .A2(n15438), .A3(n15437), .A4(n15436), .ZN(
        n15442) );
  AOI22_X1 U17727 ( .A1(n15504), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12793), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15441) );
  NAND2_X1 U17728 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n15440) );
  NAND3_X1 U17729 ( .A1(n15442), .A2(n15441), .A3(n15440), .ZN(n15448) );
  AOI22_X1 U17730 ( .A1(n15509), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15508), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15446) );
  AOI22_X1 U17731 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15445) );
  AOI22_X1 U17732 ( .A1(n15512), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15444) );
  NAND2_X1 U17733 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n15443) );
  NAND4_X1 U17734 ( .A1(n15446), .A2(n15445), .A3(n15444), .A4(n15443), .ZN(
        n15447) );
  OR2_X1 U17735 ( .A1(n15448), .A2(n15447), .ZN(n16469) );
  NAND2_X1 U17736 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n15453) );
  AOI22_X1 U17737 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12479), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15452) );
  AOI22_X1 U17738 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n15498), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U17739 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n15450) );
  AND4_X1 U17740 ( .A1(n15453), .A2(n15452), .A3(n15451), .A4(n15450), .ZN(
        n15456) );
  AOI22_X1 U17741 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n15504), .B1(
        n12793), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15455) );
  NAND2_X1 U17742 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n15454) );
  NAND3_X1 U17743 ( .A1(n15456), .A2(n15455), .A3(n15454), .ZN(n15462) );
  AOI22_X1 U17744 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n15508), .B1(
        n15509), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15460) );
  AOI22_X1 U17745 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U17746 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n15512), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15458) );
  NAND2_X1 U17747 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n15457) );
  NAND4_X1 U17748 ( .A1(n15460), .A2(n15459), .A3(n15458), .A4(n15457), .ZN(
        n15461) );
  OR2_X1 U17749 ( .A1(n15462), .A2(n15461), .ZN(n16462) );
  AOI22_X1 U17750 ( .A1(n15509), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15508), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U17751 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15465) );
  AOI22_X1 U17752 ( .A1(n15512), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15464) );
  NAND2_X1 U17753 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n15463) );
  AND4_X1 U17754 ( .A1(n15466), .A2(n15465), .A3(n15464), .A4(n15463), .ZN(
        n15477) );
  NAND2_X1 U17755 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n15468) );
  NAND2_X1 U17756 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n15467) );
  OAI211_X1 U17757 ( .C1(n15484), .C2(n15469), .A(n15468), .B(n15467), .ZN(
        n15475) );
  NAND2_X1 U17758 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n15473) );
  AOI22_X1 U17759 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U17760 ( .A1(n15498), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15471) );
  NAND2_X1 U17761 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n15470) );
  NAND4_X1 U17762 ( .A1(n15473), .A2(n15472), .A3(n15471), .A4(n15470), .ZN(
        n15474) );
  NOR2_X1 U17763 ( .A1(n15475), .A2(n15474), .ZN(n15476) );
  AND2_X1 U17764 ( .A1(n15477), .A2(n15476), .ZN(n16456) );
  AOI22_X1 U17765 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n15508), .B1(
        n15509), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15481) );
  AOI22_X1 U17766 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15480) );
  AOI22_X1 U17767 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n15512), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15479) );
  NAND2_X1 U17768 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n15478) );
  AND4_X1 U17769 ( .A1(n15481), .A2(n15480), .A3(n15479), .A4(n15478), .ZN(
        n15494) );
  NAND2_X1 U17770 ( .A1(n12793), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n15483) );
  NAND2_X1 U17771 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n15482) );
  OAI211_X1 U17772 ( .C1(n15484), .C2(n19605), .A(n15483), .B(n15482), .ZN(
        n15492) );
  NAND2_X1 U17773 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n15490) );
  AOI22_X1 U17774 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12479), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15489) );
  AOI22_X1 U17775 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n15498), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15488) );
  NAND2_X1 U17776 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n15487) );
  NAND4_X1 U17777 ( .A1(n15490), .A2(n15489), .A3(n15488), .A4(n15487), .ZN(
        n15491) );
  NOR2_X1 U17778 ( .A1(n15492), .A2(n15491), .ZN(n15493) );
  AND2_X1 U17779 ( .A1(n15494), .A2(n15493), .ZN(n16442) );
  NAND2_X1 U17780 ( .A1(n14086), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n15503) );
  AOI22_X1 U17781 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12479), .B1(
        n15485), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15502) );
  AOI22_X1 U17782 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n15498), .B1(
        n15486), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15501) );
  NAND2_X1 U17783 ( .A1(n15499), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n15500) );
  AND4_X1 U17784 ( .A1(n15503), .A2(n15502), .A3(n15501), .A4(n15500), .ZN(
        n15507) );
  AOI22_X1 U17785 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n15504), .B1(
        n12793), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15506) );
  NAND2_X1 U17786 ( .A1(n12500), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n15505) );
  NAND3_X1 U17787 ( .A1(n15507), .A2(n15506), .A3(n15505), .ZN(n15519) );
  AOI22_X1 U17788 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n15509), .B1(
        n15508), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15517) );
  AOI22_X1 U17789 ( .A1(n15511), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15510), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15516) );
  AOI22_X1 U17790 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n15512), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15515) );
  NAND2_X1 U17791 ( .A1(n15513), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n15514) );
  NAND4_X1 U17792 ( .A1(n15517), .A2(n15516), .A3(n15515), .A4(n15514), .ZN(
        n15518) );
  OR2_X1 U17793 ( .A1(n15519), .A2(n15518), .ZN(n15540) );
  AOI22_X1 U17794 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15529) );
  INV_X1 U17795 ( .A(n15649), .ZN(n15654) );
  AOI22_X1 U17796 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15528) );
  INV_X1 U17797 ( .A(n15683), .ZN(n15619) );
  NAND2_X1 U17798 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n15523) );
  INV_X1 U17799 ( .A(n15520), .ZN(n15522) );
  NAND2_X1 U17800 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15521) );
  NAND2_X1 U17801 ( .A1(n15522), .A2(n15521), .ZN(n15682) );
  OAI211_X1 U17802 ( .C1(n15619), .C2(n15524), .A(n15523), .B(n15682), .ZN(
        n15525) );
  INV_X1 U17803 ( .A(n15525), .ZN(n15527) );
  AOI22_X1 U17804 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15526) );
  NAND4_X1 U17805 ( .A1(n15529), .A2(n15528), .A3(n15527), .A4(n15526), .ZN(
        n15538) );
  AOI22_X1 U17806 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15536) );
  AOI22_X1 U17807 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15535) );
  INV_X1 U17808 ( .A(n15682), .ZN(n15672) );
  NAND2_X1 U17809 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n15530) );
  OAI211_X1 U17810 ( .C1(n15619), .C2(n15531), .A(n15672), .B(n15530), .ZN(
        n15532) );
  INV_X1 U17811 ( .A(n15532), .ZN(n15534) );
  AOI22_X1 U17812 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15533) );
  NAND4_X1 U17813 ( .A1(n15536), .A2(n15535), .A3(n15534), .A4(n15533), .ZN(
        n15537) );
  AND2_X1 U17814 ( .A1(n15538), .A2(n15537), .ZN(n15539) );
  XNOR2_X1 U17815 ( .A(n15540), .B(n15539), .ZN(n16435) );
  NAND2_X1 U17816 ( .A1(n15540), .A2(n15539), .ZN(n15562) );
  AOI22_X1 U17817 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15550) );
  AOI22_X1 U17818 ( .A1(n15566), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n15676), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15549) );
  INV_X1 U17819 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15545) );
  NAND2_X1 U17820 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n15544) );
  OAI211_X1 U17821 ( .C1(n15619), .C2(n15545), .A(n15682), .B(n15544), .ZN(
        n15546) );
  INV_X1 U17822 ( .A(n15546), .ZN(n15548) );
  AOI22_X1 U17823 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15547) );
  NAND4_X1 U17824 ( .A1(n15550), .A2(n15549), .A3(n15548), .A4(n15547), .ZN(
        n15559) );
  AOI22_X1 U17825 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15557) );
  AOI22_X1 U17826 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15556) );
  INV_X1 U17827 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15552) );
  NAND2_X1 U17828 ( .A1(n15681), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n15551) );
  OAI211_X1 U17829 ( .C1(n15619), .C2(n15552), .A(n15672), .B(n15551), .ZN(
        n15553) );
  INV_X1 U17830 ( .A(n15553), .ZN(n15555) );
  AOI22_X1 U17831 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15554) );
  NAND4_X1 U17832 ( .A1(n15557), .A2(n15556), .A3(n15555), .A4(n15554), .ZN(
        n15558) );
  NAND2_X1 U17833 ( .A1(n15559), .A2(n15558), .ZN(n15561) );
  INV_X1 U17834 ( .A(n15561), .ZN(n15560) );
  AND2_X1 U17835 ( .A1(n15541), .A2(n15560), .ZN(n15565) );
  NAND2_X1 U17836 ( .A1(n15565), .A2(n16334), .ZN(n15564) );
  OAI21_X1 U17837 ( .B1(n15582), .B2(n15562), .A(n15561), .ZN(n15563) );
  AND2_X1 U17838 ( .A1(n15564), .A2(n15563), .ZN(n16427) );
  INV_X1 U17839 ( .A(n15565), .ZN(n15583) );
  AOI22_X1 U17840 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U17841 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15571) );
  NAND2_X1 U17842 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n15567) );
  OAI211_X1 U17843 ( .C1(n15619), .C2(n14030), .A(n15682), .B(n15567), .ZN(
        n15568) );
  INV_X1 U17844 ( .A(n15568), .ZN(n15570) );
  AOI22_X1 U17845 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15569) );
  NAND4_X1 U17846 ( .A1(n15572), .A2(n15571), .A3(n15570), .A4(n15569), .ZN(
        n15581) );
  AOI22_X1 U17847 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15579) );
  AOI22_X1 U17848 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15578) );
  NAND2_X1 U17849 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n15573) );
  OAI211_X1 U17850 ( .C1(n15619), .C2(n15574), .A(n15672), .B(n15573), .ZN(
        n15575) );
  INV_X1 U17851 ( .A(n15575), .ZN(n15577) );
  AOI22_X1 U17852 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15576) );
  NAND4_X1 U17853 ( .A1(n15579), .A2(n15578), .A3(n15577), .A4(n15576), .ZN(
        n15580) );
  NAND2_X1 U17854 ( .A1(n15581), .A2(n15580), .ZN(n15584) );
  NOR2_X1 U17855 ( .A1(n15583), .A2(n15584), .ZN(n15587) );
  AOI211_X1 U17856 ( .C1(n15583), .C2(n15584), .A(n15582), .B(n15587), .ZN(
        n15585) );
  NOR2_X1 U17857 ( .A1(n16334), .A2(n15584), .ZN(n16420) );
  INV_X1 U17858 ( .A(n15585), .ZN(n15586) );
  INV_X1 U17859 ( .A(n15587), .ZN(n15609) );
  AOI22_X1 U17860 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15678), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15595) );
  AOI22_X1 U17861 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15588), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15594) );
  NAND2_X1 U17862 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n15589) );
  OAI211_X1 U17863 ( .C1(n15619), .C2(n15590), .A(n15682), .B(n15589), .ZN(
        n15591) );
  INV_X1 U17864 ( .A(n15591), .ZN(n15593) );
  AOI22_X1 U17865 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15592) );
  NAND4_X1 U17866 ( .A1(n15595), .A2(n15594), .A3(n15593), .A4(n15592), .ZN(
        n15604) );
  AOI22_X1 U17867 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15602) );
  AOI22_X1 U17868 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15601) );
  NAND2_X1 U17869 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n15596) );
  OAI211_X1 U17870 ( .C1(n15619), .C2(n15597), .A(n15672), .B(n15596), .ZN(
        n15598) );
  INV_X1 U17871 ( .A(n15598), .ZN(n15600) );
  AOI22_X1 U17872 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15599) );
  NAND4_X1 U17873 ( .A1(n15602), .A2(n15601), .A3(n15600), .A4(n15599), .ZN(
        n15603) );
  AND2_X1 U17874 ( .A1(n15604), .A2(n15603), .ZN(n15607) );
  XNOR2_X1 U17875 ( .A(n15609), .B(n15607), .ZN(n15605) );
  NAND2_X1 U17876 ( .A1(n15667), .A2(n15607), .ZN(n16415) );
  INV_X1 U17877 ( .A(n15607), .ZN(n15608) );
  NOR2_X1 U17878 ( .A1(n15609), .A2(n15608), .ZN(n15628) );
  AOI22_X1 U17879 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15616) );
  AOI22_X1 U17880 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15615) );
  NAND2_X1 U17881 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n15610) );
  OAI211_X1 U17882 ( .C1(n15619), .C2(n15611), .A(n15610), .B(n15682), .ZN(
        n15612) );
  INV_X1 U17883 ( .A(n15612), .ZN(n15614) );
  AOI22_X1 U17884 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15613) );
  NAND4_X1 U17885 ( .A1(n15616), .A2(n15615), .A3(n15614), .A4(n15613), .ZN(
        n15626) );
  AOI22_X1 U17886 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15624) );
  AOI22_X1 U17887 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15623) );
  NAND2_X1 U17888 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n15617) );
  OAI211_X1 U17889 ( .C1(n15619), .C2(n15618), .A(n15672), .B(n15617), .ZN(
        n15620) );
  INV_X1 U17890 ( .A(n15620), .ZN(n15622) );
  AOI22_X1 U17891 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15621) );
  NAND4_X1 U17892 ( .A1(n15624), .A2(n15623), .A3(n15622), .A4(n15621), .ZN(
        n15625) );
  AND2_X1 U17893 ( .A1(n15626), .A2(n15625), .ZN(n15629) );
  NAND2_X1 U17894 ( .A1(n15628), .A2(n15629), .ZN(n16394) );
  OAI211_X1 U17895 ( .C1(n15628), .C2(n15629), .A(n15627), .B(n16394), .ZN(
        n15645) );
  INV_X1 U17896 ( .A(n15629), .ZN(n15630) );
  NOR2_X1 U17897 ( .A1(n16334), .A2(n15630), .ZN(n16405) );
  AOI22_X1 U17898 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15632) );
  AOI22_X1 U17899 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15631) );
  NAND2_X1 U17900 ( .A1(n15632), .A2(n15631), .ZN(n15644) );
  INV_X1 U17901 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15635) );
  AOI21_X1 U17902 ( .B1(n15683), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n15672), .ZN(n15634) );
  AOI22_X1 U17903 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15633) );
  OAI211_X1 U17904 ( .C1(n15687), .C2(n15635), .A(n15634), .B(n15633), .ZN(
        n15643) );
  AOI22_X1 U17905 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15637) );
  AOI22_X1 U17906 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15636) );
  NAND2_X1 U17907 ( .A1(n15637), .A2(n15636), .ZN(n15642) );
  AOI22_X1 U17908 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15639) );
  AOI21_X1 U17909 ( .B1(n15683), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n15682), .ZN(n15638) );
  OAI211_X1 U17910 ( .C1(n15687), .C2(n15640), .A(n15639), .B(n15638), .ZN(
        n15641) );
  OAI22_X1 U17911 ( .A1(n15644), .A2(n15643), .B1(n15642), .B2(n15641), .ZN(
        n15666) );
  INV_X1 U17912 ( .A(n15666), .ZN(n16395) );
  NAND2_X1 U17913 ( .A1(n15646), .A2(n15645), .ZN(n16402) );
  AOI22_X1 U17914 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15566), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15648) );
  NAND2_X1 U17915 ( .A1(n15677), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n15647) );
  OAI211_X1 U17916 ( .C1(n15649), .C2(n19605), .A(n15648), .B(n15647), .ZN(
        n15663) );
  INV_X1 U17917 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15653) );
  AOI21_X1 U17918 ( .B1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n15683), .A(
        n15672), .ZN(n15652) );
  AOI22_X1 U17919 ( .A1(n12657), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15651) );
  OAI211_X1 U17920 ( .C1(n15653), .C2(n15650), .A(n15652), .B(n15651), .ZN(
        n15662) );
  AOI22_X1 U17921 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15678), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U17922 ( .A1(n15654), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U17923 ( .A1(n15656), .A2(n15655), .ZN(n15661) );
  INV_X1 U17924 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15659) );
  AOI22_X1 U17925 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15658) );
  AOI21_X1 U17926 ( .B1(n15683), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n15682), .ZN(n15657) );
  OAI211_X1 U17927 ( .C1(n15650), .C2(n15659), .A(n15658), .B(n15657), .ZN(
        n15660) );
  OAI22_X1 U17928 ( .A1(n15663), .A2(n15662), .B1(n15661), .B2(n15660), .ZN(
        n15664) );
  NOR2_X1 U17929 ( .A1(n15665), .A2(n15664), .ZN(n16387) );
  INV_X1 U17930 ( .A(n16387), .ZN(n15669) );
  NAND2_X1 U17931 ( .A1(n15665), .A2(n15664), .ZN(n16385) );
  NOR3_X1 U17932 ( .A1(n16394), .A2(n15667), .A3(n15666), .ZN(n16388) );
  NAND2_X1 U17933 ( .A1(n16385), .A2(n16388), .ZN(n15668) );
  NAND2_X1 U17934 ( .A1(n15669), .A2(n15668), .ZN(n15694) );
  AOI22_X1 U17935 ( .A1(n15683), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15671) );
  AOI22_X1 U17936 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15676), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15670) );
  NAND2_X1 U17937 ( .A1(n15671), .A2(n15670), .ZN(n15691) );
  INV_X1 U17938 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n19524) );
  AOI21_X1 U17939 ( .B1(n12667), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n15672), .ZN(n15674) );
  AOI22_X1 U17940 ( .A1(n12618), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15673) );
  OAI211_X1 U17941 ( .C1(n15675), .C2(n19524), .A(n15674), .B(n15673), .ZN(
        n15690) );
  AOI22_X1 U17942 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15676), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U17943 ( .A1(n15678), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15677), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15679) );
  NAND2_X1 U17944 ( .A1(n15680), .A2(n15679), .ZN(n15689) );
  AOI22_X1 U17945 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15681), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15685) );
  AOI21_X1 U17946 ( .B1(n15683), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n15682), .ZN(n15684) );
  OAI211_X1 U17947 ( .C1(n15687), .C2(n15686), .A(n15685), .B(n15684), .ZN(
        n15688) );
  OAI22_X1 U17948 ( .A1(n15691), .A2(n15690), .B1(n15689), .B2(n15688), .ZN(
        n15692) );
  INV_X1 U17949 ( .A(n15692), .ZN(n15693) );
  XNOR2_X1 U17950 ( .A(n15694), .B(n15693), .ZN(n15710) );
  OAI22_X1 U17951 ( .A1(n16564), .A2(n19371), .B1(n19556), .B2(n15696), .ZN(
        n15701) );
  INV_X1 U17952 ( .A(n19764), .ZN(n16487) );
  INV_X1 U17953 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n15699) );
  NOR2_X1 U17954 ( .A1(n16487), .A2(n15699), .ZN(n15700) );
  AOI211_X1 U17955 ( .C1(BUF1_REG_30__SCAN_IN), .C2(n19765), .A(n15701), .B(
        n15700), .ZN(n15705) );
  AOI21_X1 U17956 ( .B1(n15703), .B2(n16477), .A(n15702), .ZN(n16751) );
  NAND2_X1 U17957 ( .A1(n16751), .A2(n19860), .ZN(n15704) );
  OAI211_X1 U17958 ( .C1(n15710), .C2(n19812), .A(n15705), .B(n15704), .ZN(
        P2_U2889) );
  XNOR2_X1 U17959 ( .A(n15707), .B(n15706), .ZN(n18797) );
  NAND2_X1 U17960 ( .A1(n18797), .A2(n16448), .ZN(n15709) );
  NAND2_X1 U17961 ( .A1(n16433), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15708) );
  OAI211_X1 U17962 ( .C1(n15710), .C2(n16474), .A(n15709), .B(n15708), .ZN(
        P2_U2857) );
  OAI211_X1 U17963 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n14667), .A(n21952), 
        .B(n22077), .ZN(n15711) );
  MUX2_X1 U17964 ( .A(n21944), .B(n15711), .S(n17155), .Z(n15712) );
  OAI21_X1 U17965 ( .B1(n14582), .B2(n15713), .A(n15712), .ZN(P1_U3477) );
  INV_X1 U17966 ( .A(n15714), .ZN(n15715) );
  XNOR2_X1 U17967 ( .A(n15725), .B(n15715), .ZN(n16030) );
  INV_X1 U17968 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n17359) );
  OAI21_X1 U17969 ( .B1(n15729), .B2(n17359), .A(n17357), .ZN(n15720) );
  AOI22_X1 U17970 ( .A1(n21816), .A2(n16025), .B1(n21810), .B2(
        P1_EBX_REG_30__SCAN_IN), .ZN(n15716) );
  OAI21_X1 U17971 ( .B1(n15717), .B2(n21820), .A(n15716), .ZN(n15719) );
  OAI21_X1 U17972 ( .B1(n15734), .B2(n15723), .A(n15722), .ZN(n16178) );
  AOI21_X2 U17973 ( .B1(n15726), .B2(n15724), .A(n15725), .ZN(n16042) );
  NAND2_X1 U17974 ( .A1(n16042), .A2(n21771), .ZN(n15733) );
  INV_X1 U17975 ( .A(n15729), .ZN(n15727) );
  NOR2_X1 U17976 ( .A1(n15727), .A2(n21804), .ZN(n15740) );
  AOI22_X1 U17977 ( .A1(n21792), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n21810), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n15728) );
  OAI21_X1 U17978 ( .B1(n16040), .B2(n21795), .A(n15728), .ZN(n15731) );
  NOR3_X1 U17979 ( .A1(n15729), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n21732), 
        .ZN(n15730) );
  AOI211_X1 U17980 ( .C1(n15740), .C2(P1_REIP_REG_29__SCAN_IN), .A(n15731), 
        .B(n15730), .ZN(n15732) );
  OAI211_X1 U17981 ( .C1(n21812), .C2(n16178), .A(n15733), .B(n15732), .ZN(
        P1_U2811) );
  INV_X1 U17982 ( .A(n15734), .ZN(n15735) );
  OAI21_X1 U17983 ( .B1(n15748), .B2(n15736), .A(n15735), .ZN(n16188) );
  OAI21_X2 U17984 ( .B1(n15737), .B2(n15738), .A(n15724), .ZN(n15967) );
  INV_X1 U17985 ( .A(n15967), .ZN(n16054) );
  NAND2_X1 U17986 ( .A1(n16054), .A2(n21771), .ZN(n15746) );
  INV_X1 U17987 ( .A(n15739), .ZN(n16052) );
  INV_X1 U17988 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15900) );
  OAI22_X1 U17989 ( .A1(n21795), .A2(n16052), .B1(n21765), .B2(n15900), .ZN(
        n15744) );
  INV_X1 U17990 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n17362) );
  NAND2_X1 U17991 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n15752), .ZN(n15742) );
  INV_X1 U17992 ( .A(n15740), .ZN(n15741) );
  AOI21_X1 U17993 ( .B1(n17362), .B2(n15742), .A(n15741), .ZN(n15743) );
  AOI211_X1 U17994 ( .C1(n21792), .C2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15744), .B(n15743), .ZN(n15745) );
  OAI211_X1 U17995 ( .C1(n16188), .C2(n21812), .A(n15746), .B(n15745), .ZN(
        P1_U2812) );
  AND2_X1 U17996 ( .A1(n15760), .A2(n15747), .ZN(n15749) );
  OR2_X1 U17997 ( .A1(n15749), .A2(n15748), .ZN(n16193) );
  AOI21_X1 U17998 ( .B1(n15751), .B2(n15750), .A(n15737), .ZN(n16062) );
  NAND2_X1 U17999 ( .A1(n16062), .A2(n21771), .ZN(n15757) );
  NOR2_X1 U18000 ( .A1(n15752), .A2(n21804), .ZN(n15768) );
  INV_X1 U18001 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n16058) );
  NAND3_X1 U18002 ( .A1(n15752), .A2(n21721), .A3(n16058), .ZN(n15754) );
  AOI22_X1 U18003 ( .A1(n21792), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n21810), .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n15753) );
  OAI211_X1 U18004 ( .C1(n21795), .C2(n16060), .A(n15754), .B(n15753), .ZN(
        n15755) );
  AOI21_X1 U18005 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n15768), .A(n15755), 
        .ZN(n15756) );
  OAI211_X1 U18006 ( .C1(n16193), .C2(n21812), .A(n15757), .B(n15756), .ZN(
        P1_U2813) );
  NAND2_X1 U18007 ( .A1(n15772), .A2(n15758), .ZN(n15759) );
  NAND2_X1 U18008 ( .A1(n15760), .A2(n15759), .ZN(n16208) );
  OAI21_X1 U18009 ( .B1(n15761), .B2(n15762), .A(n15750), .ZN(n15975) );
  INV_X1 U18010 ( .A(n15975), .ZN(n16069) );
  NAND2_X1 U18011 ( .A1(n16069), .A2(n21771), .ZN(n15770) );
  INV_X1 U18012 ( .A(n15763), .ZN(n16067) );
  AOI22_X1 U18013 ( .A1(n21792), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n21810), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n15764) );
  OAI21_X1 U18014 ( .B1(n16067), .B2(n21795), .A(n15764), .ZN(n15767) );
  NAND2_X1 U18015 ( .A1(n15778), .A2(n21721), .ZN(n15809) );
  NAND3_X1 U18016 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_25__SCAN_IN), .ZN(n15765) );
  NOR3_X1 U18017 ( .A1(n15809), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n15765), 
        .ZN(n15766) );
  AOI211_X1 U18018 ( .C1(n15768), .C2(P1_REIP_REG_26__SCAN_IN), .A(n15767), 
        .B(n15766), .ZN(n15769) );
  OAI211_X1 U18019 ( .C1(n16208), .C2(n21812), .A(n15770), .B(n15769), .ZN(
        P1_U2814) );
  INV_X1 U18020 ( .A(n15788), .ZN(n15774) );
  INV_X1 U18021 ( .A(n15771), .ZN(n15773) );
  OAI21_X1 U18022 ( .B1(n15774), .B2(n15773), .A(n15772), .ZN(n16213) );
  INV_X1 U18023 ( .A(n15775), .ZN(n15776) );
  AOI21_X1 U18024 ( .B1(n15777), .B2(n15776), .A(n15761), .ZN(n16078) );
  NAND2_X1 U18025 ( .A1(n16078), .A2(n21771), .ZN(n15783) );
  NAND2_X1 U18026 ( .A1(n15778), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15787) );
  NAND2_X1 U18027 ( .A1(n15787), .A2(n21781), .ZN(n15808) );
  OAI21_X1 U18028 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n21732), .A(n15808), 
        .ZN(n15796) );
  AOI22_X1 U18029 ( .A1(n21792), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n21810), .B2(P1_EBX_REG_25__SCAN_IN), .ZN(n15779) );
  OAI21_X1 U18030 ( .B1(n16076), .B2(n21795), .A(n15779), .ZN(n15781) );
  INV_X1 U18031 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n17161) );
  INV_X1 U18032 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n17260) );
  NOR4_X1 U18033 ( .A1(n15809), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n17161), 
        .A4(n17260), .ZN(n15780) );
  AOI211_X1 U18034 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n15796), .A(n15781), 
        .B(n15780), .ZN(n15782) );
  OAI211_X1 U18035 ( .C1(n16213), .C2(n21812), .A(n15783), .B(n15782), .ZN(
        P1_U2815) );
  AOI21_X1 U18037 ( .B1(n15786), .B2(n15785), .A(n15775), .ZN(n16086) );
  INV_X1 U18038 ( .A(n16086), .ZN(n15983) );
  INV_X1 U18039 ( .A(n15787), .ZN(n15797) );
  OAI21_X1 U18040 ( .B1(n15803), .B2(n15789), .A(n15788), .ZN(n16222) );
  INV_X1 U18041 ( .A(n15790), .ZN(n16084) );
  OAI22_X1 U18042 ( .A1(n21795), .A2(n16084), .B1(n15791), .B2(n21765), .ZN(
        n15793) );
  NOR2_X1 U18043 ( .A1(n15808), .A2(n17161), .ZN(n15792) );
  AOI211_X1 U18044 ( .C1(n21792), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15793), .B(n15792), .ZN(n15794) );
  OAI21_X1 U18045 ( .B1(n16222), .B2(n21812), .A(n15794), .ZN(n15795) );
  AOI21_X1 U18046 ( .B1(n15797), .B2(n15796), .A(n15795), .ZN(n15798) );
  OAI21_X1 U18047 ( .B1(n15983), .B2(n21813), .A(n15798), .ZN(P1_U2816) );
  OAI21_X1 U18048 ( .B1(n15799), .B2(n15800), .A(n15785), .ZN(n16090) );
  AND2_X1 U18049 ( .A1(n15912), .A2(n15801), .ZN(n15802) );
  OR2_X1 U18050 ( .A1(n15803), .A2(n15802), .ZN(n15904) );
  INV_X1 U18051 ( .A(n15904), .ZN(n16239) );
  INV_X1 U18052 ( .A(n15804), .ZN(n16092) );
  NAND2_X1 U18053 ( .A1(n21792), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15806) );
  NAND2_X1 U18054 ( .A1(n21810), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n15805) );
  OAI211_X1 U18055 ( .C1(n21795), .C2(n16092), .A(n15806), .B(n15805), .ZN(
        n15807) );
  AOI21_X1 U18056 ( .B1(n16239), .B2(n21801), .A(n15807), .ZN(n15813) );
  INV_X1 U18057 ( .A(n15808), .ZN(n15811) );
  NAND2_X1 U18058 ( .A1(n15809), .A2(n17260), .ZN(n15810) );
  NAND2_X1 U18059 ( .A1(n15811), .A2(n15810), .ZN(n15812) );
  OAI211_X1 U18060 ( .C1(n16090), .C2(n21813), .A(n15813), .B(n15812), .ZN(
        P1_U2817) );
  AOI21_X1 U18062 ( .B1(n15817), .B2(n11125), .A(n15816), .ZN(n20223) );
  INV_X1 U18063 ( .A(n20223), .ZN(n16006) );
  OR2_X1 U18064 ( .A1(n15946), .A2(n15818), .ZN(n15819) );
  AND2_X1 U18065 ( .A1(n15935), .A2(n15819), .ZN(n21592) );
  AOI21_X1 U18066 ( .B1(n21810), .B2(P1_EBX_REG_17__SCAN_IN), .A(n21769), .ZN(
        n15820) );
  OAI21_X1 U18067 ( .B1(n21795), .B2(n15821), .A(n15820), .ZN(n15828) );
  INV_X1 U18068 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21745) );
  NAND2_X1 U18069 ( .A1(n15822), .A2(n15857), .ZN(n15838) );
  NOR2_X1 U18070 ( .A1(n15823), .A2(n15838), .ZN(n15841) );
  INV_X1 U18071 ( .A(n15841), .ZN(n21746) );
  NOR2_X1 U18072 ( .A1(n21745), .A2(n21746), .ZN(n21744) );
  NOR2_X1 U18073 ( .A1(n15824), .A2(n21746), .ZN(n21776) );
  NOR2_X1 U18074 ( .A1(n21804), .A2(n21776), .ZN(n21774) );
  OAI21_X1 U18075 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n21744), .A(n21774), 
        .ZN(n15825) );
  OAI21_X1 U18076 ( .B1(n21820), .B2(n15826), .A(n15825), .ZN(n15827) );
  AOI211_X1 U18077 ( .C1(n21592), .C2(n21801), .A(n15828), .B(n15827), .ZN(
        n15829) );
  OAI21_X1 U18078 ( .B1(n16006), .B2(n21813), .A(n15829), .ZN(P1_U2823) );
  OAI21_X1 U18079 ( .B1(n15830), .B2(n15832), .A(n15831), .ZN(n20209) );
  INV_X1 U18080 ( .A(n15867), .ZN(n15834) );
  AOI21_X1 U18081 ( .B1(n15834), .B2(n15847), .A(n15833), .ZN(n15835) );
  NOR2_X1 U18082 ( .A1(n15835), .A2(n15944), .ZN(n21577) );
  INV_X1 U18083 ( .A(n20210), .ZN(n15837) );
  AOI21_X1 U18084 ( .B1(n21810), .B2(P1_EBX_REG_15__SCAN_IN), .A(n21769), .ZN(
        n15836) );
  OAI21_X1 U18085 ( .B1(n21795), .B2(n15837), .A(n15836), .ZN(n15843) );
  INV_X1 U18086 ( .A(n15838), .ZN(n21790) );
  AOI22_X1 U18087 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n21781), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21790), .ZN(n15840) );
  OAI22_X1 U18088 ( .A1(n15841), .A2(n15840), .B1(n15839), .B2(n21820), .ZN(
        n15842) );
  AOI211_X1 U18089 ( .C1(n21577), .C2(n21801), .A(n15843), .B(n15842), .ZN(
        n15844) );
  OAI21_X1 U18090 ( .B1(n20209), .B2(n21813), .A(n15844), .ZN(P1_U2825) );
  AOI21_X1 U18091 ( .B1(n15846), .B2(n15845), .A(n15830), .ZN(n16141) );
  INV_X1 U18092 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15849) );
  XNOR2_X1 U18093 ( .A(n15867), .B(n15847), .ZN(n21460) );
  AOI22_X1 U18094 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(n21810), .B1(n21801), 
        .B2(n21460), .ZN(n15848) );
  OAI21_X1 U18095 ( .B1(n15849), .B2(n21820), .A(n15848), .ZN(n15853) );
  NAND2_X1 U18096 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n21790), .ZN(n15850) );
  OAI211_X1 U18097 ( .C1(n21790), .C2(P1_REIP_REG_14__SCAN_IN), .A(n15850), 
        .B(n21781), .ZN(n15851) );
  OAI211_X1 U18098 ( .C1(n21795), .C2(n16139), .A(n15851), .B(n21686), .ZN(
        n15852) );
  AOI211_X1 U18099 ( .C1(n16141), .C2(n21771), .A(n15853), .B(n15852), .ZN(
        n15854) );
  INV_X1 U18100 ( .A(n15854), .ZN(P1_U2826) );
  NAND2_X1 U18101 ( .A1(n15327), .A2(n15855), .ZN(n15856) );
  AND2_X1 U18102 ( .A1(n15845), .A2(n15856), .ZN(n20133) );
  INV_X1 U18103 ( .A(n20133), .ZN(n16024) );
  INV_X1 U18104 ( .A(n15857), .ZN(n15858) );
  NOR2_X1 U18105 ( .A1(n15859), .A2(n15858), .ZN(n15862) );
  INV_X1 U18106 ( .A(n15860), .ZN(n15861) );
  MUX2_X1 U18107 ( .A(n15862), .B(n15861), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n15873) );
  OAI21_X1 U18108 ( .B1(n21820), .B2(n15863), .A(n21686), .ZN(n15872) );
  NAND2_X1 U18109 ( .A1(n15865), .A2(n15864), .ZN(n15866) );
  AND2_X1 U18110 ( .A1(n15867), .A2(n15866), .ZN(n20130) );
  INV_X1 U18111 ( .A(n20130), .ZN(n15870) );
  AOI22_X1 U18112 ( .A1(n21816), .A2(n15868), .B1(n21810), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15869) );
  OAI21_X1 U18113 ( .B1(n15870), .B2(n21812), .A(n15869), .ZN(n15871) );
  NOR3_X1 U18114 ( .A1(n15873), .A2(n15872), .A3(n15871), .ZN(n15874) );
  OAI21_X1 U18115 ( .B1(n16024), .B2(n21813), .A(n15874), .ZN(P1_U2827) );
  NAND2_X1 U18116 ( .A1(n15876), .A2(n15875), .ZN(n15877) );
  NOR2_X1 U18117 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n21732), .ZN(n15885) );
  OR2_X1 U18118 ( .A1(n21448), .A2(n15878), .ZN(n21669) );
  INV_X1 U18119 ( .A(n20150), .ZN(n15879) );
  AOI22_X1 U18120 ( .A1(n21816), .A2(n15879), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n21810), .ZN(n15881) );
  NAND2_X1 U18121 ( .A1(n21792), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15880) );
  OAI211_X1 U18122 ( .C1(n14536), .C2(n21669), .A(n15881), .B(n15880), .ZN(
        n15884) );
  INV_X1 U18123 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21674) );
  AOI21_X1 U18124 ( .B1(n21721), .B2(n21674), .A(n21720), .ZN(n15882) );
  INV_X1 U18125 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21673) );
  OAI22_X1 U18126 ( .A1(n15882), .A2(n21673), .B1(n21812), .B2(n21474), .ZN(
        n15883) );
  AOI211_X1 U18127 ( .C1(P1_REIP_REG_1__SCAN_IN), .C2(n15885), .A(n15884), .B(
        n15883), .ZN(n15886) );
  OAI21_X1 U18128 ( .B1(n15887), .B2(n21690), .A(n15886), .ZN(P1_U2838) );
  NAND2_X1 U18129 ( .A1(n15888), .A2(n21679), .ZN(n15896) );
  NAND2_X1 U18130 ( .A1(n21810), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n15889) );
  OAI21_X1 U18131 ( .B1(n15890), .B2(n21812), .A(n15889), .ZN(n15891) );
  AOI21_X1 U18132 ( .B1(n21781), .B2(P1_REIP_REG_0__SCAN_IN), .A(n15891), .ZN(
        n15895) );
  INV_X1 U18133 ( .A(n21669), .ZN(n21647) );
  NAND2_X1 U18134 ( .A1(n10986), .A2(n21647), .ZN(n15894) );
  NAND2_X1 U18135 ( .A1(n21820), .A2(n21795), .ZN(n15892) );
  NAND2_X1 U18136 ( .A1(n15892), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15893) );
  NAND4_X1 U18137 ( .A1(n15896), .A2(n15895), .A3(n15894), .A4(n15893), .ZN(
        P1_U2840) );
  OAI22_X1 U18138 ( .A1(n16161), .A2(n15952), .B1(n20136), .B2(n15897), .ZN(
        P1_U2841) );
  INV_X1 U18139 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15898) );
  OAI222_X1 U18140 ( .A1(n15960), .A2(n15954), .B1(n15898), .B2(n20136), .C1(
        n15952), .C2(n15718), .ZN(P1_U2842) );
  INV_X1 U18141 ( .A(n16042), .ZN(n15963) );
  INV_X1 U18142 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15899) );
  OAI222_X1 U18143 ( .A1(n15954), .A2(n15963), .B1(n15899), .B2(n20136), .C1(
        n16178), .C2(n15952), .ZN(P1_U2843) );
  OAI222_X1 U18144 ( .A1(n15967), .A2(n15954), .B1(n15900), .B2(n20136), .C1(
        n16188), .C2(n15952), .ZN(P1_U2844) );
  INV_X1 U18145 ( .A(n16062), .ZN(n15971) );
  INV_X1 U18146 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15901) );
  OAI222_X1 U18147 ( .A1(n15954), .A2(n15971), .B1(n15901), .B2(n20136), .C1(
        n16193), .C2(n15952), .ZN(P1_U2845) );
  OAI222_X1 U18148 ( .A1(n15975), .A2(n15954), .B1(n15902), .B2(n20136), .C1(
        n16208), .C2(n15952), .ZN(P1_U2846) );
  INV_X1 U18149 ( .A(n16078), .ZN(n15979) );
  INV_X1 U18150 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15903) );
  OAI222_X1 U18151 ( .A1(n15979), .A2(n15954), .B1(n15903), .B2(n20136), .C1(
        n16213), .C2(n15952), .ZN(P1_U2847) );
  OAI222_X1 U18152 ( .A1(n15983), .A2(n15954), .B1(n20136), .B2(n15791), .C1(
        n16222), .C2(n15952), .ZN(P1_U2848) );
  INV_X1 U18153 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15905) );
  OAI222_X1 U18154 ( .A1(n16090), .A2(n15954), .B1(n15905), .B2(n20136), .C1(
        n15904), .C2(n15952), .ZN(P1_U2849) );
  BUF_X1 U18155 ( .A(n15906), .Z(n15907) );
  INV_X1 U18156 ( .A(n15799), .ZN(n15908) );
  OAI21_X1 U18157 ( .B1(n15909), .B2(n15907), .A(n15908), .ZN(n21814) );
  NAND2_X1 U18158 ( .A1(n15920), .A2(n15910), .ZN(n15911) );
  NAND2_X1 U18159 ( .A1(n15912), .A2(n15911), .ZN(n21811) );
  OAI22_X1 U18160 ( .A1(n21811), .A2(n15952), .B1(n15913), .B2(n20136), .ZN(
        n15914) );
  INV_X1 U18161 ( .A(n15914), .ZN(n15915) );
  OAI21_X1 U18162 ( .B1(n21814), .B2(n15954), .A(n15915), .ZN(P1_U2850) );
  AND2_X1 U18163 ( .A1(n11056), .A2(n15916), .ZN(n15917) );
  NOR2_X1 U18164 ( .A1(n15907), .A2(n15917), .ZN(n20235) );
  INV_X1 U18165 ( .A(n20235), .ZN(n21797) );
  OR2_X1 U18166 ( .A1(n15924), .A2(n15918), .ZN(n15919) );
  AND2_X1 U18167 ( .A1(n15920), .A2(n15919), .ZN(n21800) );
  AOI22_X1 U18168 ( .A1(n21800), .A2(n20131), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n15949), .ZN(n15921) );
  OAI21_X1 U18169 ( .B1(n21797), .B2(n15954), .A(n15921), .ZN(P1_U2851) );
  OAI21_X1 U18170 ( .B1(n11042), .B2(n11113), .A(n11056), .ZN(n21784) );
  NOR2_X1 U18171 ( .A1(n15930), .A2(n15922), .ZN(n15923) );
  OR2_X1 U18172 ( .A1(n15924), .A2(n15923), .ZN(n21783) );
  OAI22_X1 U18173 ( .A1(n21783), .A2(n15952), .B1(n15925), .B2(n20136), .ZN(
        n15926) );
  INV_X1 U18174 ( .A(n15926), .ZN(n15927) );
  OAI21_X1 U18175 ( .B1(n21784), .B2(n15954), .A(n15927), .ZN(P1_U2852) );
  AOI21_X1 U18176 ( .B1(n15929), .B2(n15928), .A(n11042), .ZN(n21772) );
  INV_X1 U18177 ( .A(n21772), .ZN(n15999) );
  AOI21_X1 U18178 ( .B1(n15931), .B2(n15937), .A(n15930), .ZN(n21770) );
  AOI22_X1 U18179 ( .A1(n21770), .A2(n20131), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n15949), .ZN(n15932) );
  OAI21_X1 U18180 ( .B1(n15999), .B2(n15954), .A(n15932), .ZN(P1_U2853) );
  OAI21_X1 U18181 ( .B1(n15816), .B2(n15933), .A(n15928), .ZN(n21760) );
  NAND2_X1 U18182 ( .A1(n15935), .A2(n15934), .ZN(n15936) );
  NAND2_X1 U18183 ( .A1(n15937), .A2(n15936), .ZN(n21764) );
  OAI22_X1 U18184 ( .A1(n21764), .A2(n15952), .B1(n15938), .B2(n20136), .ZN(
        n15939) );
  INV_X1 U18185 ( .A(n15939), .ZN(n15940) );
  OAI21_X1 U18186 ( .B1(n21760), .B2(n15954), .A(n15940), .ZN(P1_U2854) );
  AOI22_X1 U18187 ( .A1(n21592), .A2(n20131), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n15949), .ZN(n15941) );
  OAI21_X1 U18188 ( .B1(n16006), .B2(n15954), .A(n15941), .ZN(P1_U2855) );
  AOI21_X1 U18189 ( .B1(n15942), .B2(n15831), .A(n15814), .ZN(n16129) );
  INV_X1 U18190 ( .A(n16129), .ZN(n21749) );
  NOR2_X1 U18191 ( .A1(n15944), .A2(n15943), .ZN(n15945) );
  OR2_X1 U18192 ( .A1(n15946), .A2(n15945), .ZN(n21748) );
  OAI22_X1 U18193 ( .A1(n21748), .A2(n15952), .B1(n21754), .B2(n20136), .ZN(
        n15947) );
  INV_X1 U18194 ( .A(n15947), .ZN(n15948) );
  OAI21_X1 U18195 ( .B1(n21749), .B2(n15954), .A(n15948), .ZN(P1_U2856) );
  AOI22_X1 U18196 ( .A1(n21577), .A2(n20131), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n15949), .ZN(n15950) );
  OAI21_X1 U18197 ( .B1(n20209), .B2(n15954), .A(n15950), .ZN(P1_U2857) );
  INV_X1 U18198 ( .A(n16141), .ZN(n16018) );
  INV_X1 U18199 ( .A(n21460), .ZN(n15951) );
  OAI222_X1 U18200 ( .A1(n16018), .A2(n15954), .B1(n15953), .B2(n20136), .C1(
        n15952), .C2(n15951), .ZN(P1_U2858) );
  AOI22_X1 U18201 ( .A1(n16007), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n16019), .ZN(n15959) );
  NOR3_X1 U18202 ( .A1(n16019), .A2(n15956), .A3(n11858), .ZN(n15957) );
  AOI22_X1 U18203 ( .A1(n16010), .A2(n16016), .B1(n16008), .B2(DATAI_30_), 
        .ZN(n15958) );
  OAI211_X1 U18204 ( .C1(n15960), .C2(n16023), .A(n15959), .B(n15958), .ZN(
        P1_U2874) );
  AOI22_X1 U18205 ( .A1(n16007), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n16019), .ZN(n15962) );
  AOI22_X1 U18206 ( .A1(n16010), .A2(n16020), .B1(n16008), .B2(DATAI_29_), 
        .ZN(n15961) );
  OAI211_X1 U18207 ( .C1(n15963), .C2(n16023), .A(n15962), .B(n15961), .ZN(
        P1_U2875) );
  AOI22_X1 U18208 ( .A1(n16007), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n16019), .ZN(n15966) );
  AOI22_X1 U18209 ( .A1(n16010), .A2(n15964), .B1(n16008), .B2(DATAI_28_), 
        .ZN(n15965) );
  OAI211_X1 U18210 ( .C1(n15967), .C2(n16023), .A(n15966), .B(n15965), .ZN(
        P1_U2876) );
  AOI22_X1 U18211 ( .A1(n16007), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n16019), .ZN(n15970) );
  AOI22_X1 U18212 ( .A1(n16010), .A2(n15968), .B1(n16008), .B2(DATAI_27_), 
        .ZN(n15969) );
  OAI211_X1 U18213 ( .C1(n15971), .C2(n16023), .A(n15970), .B(n15969), .ZN(
        P1_U2877) );
  AOI22_X1 U18214 ( .A1(n16007), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n16019), .ZN(n15974) );
  AOI22_X1 U18215 ( .A1(n16010), .A2(n15972), .B1(n16008), .B2(DATAI_26_), 
        .ZN(n15973) );
  OAI211_X1 U18216 ( .C1(n15975), .C2(n16023), .A(n15974), .B(n15973), .ZN(
        P1_U2878) );
  AOI22_X1 U18217 ( .A1(n16007), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n16019), .ZN(n15978) );
  AOI22_X1 U18218 ( .A1(n16010), .A2(n15976), .B1(n16008), .B2(DATAI_25_), 
        .ZN(n15977) );
  OAI211_X1 U18219 ( .C1(n15979), .C2(n16023), .A(n15978), .B(n15977), .ZN(
        P1_U2879) );
  AOI22_X1 U18220 ( .A1(n16007), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n16019), .ZN(n15982) );
  AOI22_X1 U18221 ( .A1(n16010), .A2(n15980), .B1(n16008), .B2(DATAI_24_), 
        .ZN(n15981) );
  OAI211_X1 U18222 ( .C1(n15983), .C2(n16023), .A(n15982), .B(n15981), .ZN(
        P1_U2880) );
  AOI22_X1 U18223 ( .A1(n16007), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n16019), .ZN(n15986) );
  AOI22_X1 U18224 ( .A1(n16010), .A2(n15984), .B1(n16008), .B2(DATAI_23_), 
        .ZN(n15985) );
  OAI211_X1 U18225 ( .C1(n16090), .C2(n16023), .A(n15986), .B(n15985), .ZN(
        P1_U2881) );
  AOI22_X1 U18226 ( .A1(n16007), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n16019), .ZN(n15989) );
  AOI22_X1 U18227 ( .A1(n16010), .A2(n15987), .B1(n16008), .B2(DATAI_22_), 
        .ZN(n15988) );
  OAI211_X1 U18228 ( .C1(n21814), .C2(n16023), .A(n15989), .B(n15988), .ZN(
        P1_U2882) );
  AOI22_X1 U18229 ( .A1(n16007), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n16019), .ZN(n15992) );
  AOI22_X1 U18230 ( .A1(n16010), .A2(n15990), .B1(n16008), .B2(DATAI_21_), 
        .ZN(n15991) );
  OAI211_X1 U18231 ( .C1(n21797), .C2(n16023), .A(n15992), .B(n15991), .ZN(
        P1_U2883) );
  AOI22_X1 U18232 ( .A1(n16007), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n16019), .ZN(n15995) );
  AOI22_X1 U18233 ( .A1(n16010), .A2(n15993), .B1(n16008), .B2(DATAI_20_), 
        .ZN(n15994) );
  OAI211_X1 U18234 ( .C1(n21784), .C2(n16023), .A(n15995), .B(n15994), .ZN(
        P1_U2884) );
  AOI22_X1 U18235 ( .A1(n16007), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n16019), .ZN(n15998) );
  AOI22_X1 U18236 ( .A1(n16010), .A2(n15996), .B1(n16008), .B2(DATAI_19_), 
        .ZN(n15997) );
  OAI211_X1 U18237 ( .C1(n15999), .C2(n16023), .A(n15998), .B(n15997), .ZN(
        P1_U2885) );
  AOI22_X1 U18238 ( .A1(n16007), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n16019), .ZN(n16002) );
  AOI22_X1 U18239 ( .A1(n16010), .A2(n16000), .B1(n16008), .B2(DATAI_18_), 
        .ZN(n16001) );
  OAI211_X1 U18240 ( .C1(n21760), .C2(n16023), .A(n16002), .B(n16001), .ZN(
        P1_U2886) );
  AOI22_X1 U18241 ( .A1(n16007), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n16019), .ZN(n16005) );
  AOI22_X1 U18242 ( .A1(n16010), .A2(n16003), .B1(n16008), .B2(DATAI_17_), 
        .ZN(n16004) );
  OAI211_X1 U18243 ( .C1(n16006), .C2(n16023), .A(n16005), .B(n16004), .ZN(
        P1_U2887) );
  AOI22_X1 U18244 ( .A1(n16007), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n16019), .ZN(n16012) );
  AOI22_X1 U18245 ( .A1(n16010), .A2(n16009), .B1(n16008), .B2(DATAI_16_), 
        .ZN(n16011) );
  OAI211_X1 U18246 ( .C1(n21749), .C2(n16023), .A(n16012), .B(n16011), .ZN(
        P1_U2888) );
  OAI222_X1 U18247 ( .A1(n16023), .A2(n20209), .B1(n16015), .B2(n20067), .C1(
        n16014), .C2(n16013), .ZN(P1_U2889) );
  AOI22_X1 U18248 ( .A1(n16021), .A2(n16016), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n16019), .ZN(n16017) );
  OAI21_X1 U18249 ( .B1(n16018), .B2(n16023), .A(n16017), .ZN(P1_U2890) );
  AOI22_X1 U18250 ( .A1(n16021), .A2(n16020), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n16019), .ZN(n16022) );
  OAI21_X1 U18251 ( .B1(n16024), .B2(n16023), .A(n16022), .ZN(P1_U2891) );
  INV_X1 U18252 ( .A(n16025), .ZN(n16028) );
  AOI21_X1 U18253 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16026), .ZN(n16027) );
  OAI21_X1 U18254 ( .B1(n20240), .B2(n16028), .A(n16027), .ZN(n16029) );
  AOI21_X1 U18255 ( .B1(n16030), .B2(n20236), .A(n16029), .ZN(n16031) );
  OAI21_X1 U18256 ( .B1(n16032), .B2(n21822), .A(n16031), .ZN(P1_U2969) );
  INV_X1 U18257 ( .A(n16034), .ZN(n16037) );
  INV_X1 U18258 ( .A(n16035), .ZN(n16036) );
  NAND2_X1 U18259 ( .A1(n16037), .A2(n16036), .ZN(n16038) );
  XNOR2_X1 U18260 ( .A(n16033), .B(n16038), .ZN(n16182) );
  NOR2_X1 U18261 ( .A1(n21596), .A2(n17359), .ZN(n16176) );
  AOI21_X1 U18262 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16176), .ZN(n16039) );
  OAI21_X1 U18263 ( .B1(n20240), .B2(n16040), .A(n16039), .ZN(n16041) );
  AOI21_X1 U18264 ( .B1(n16042), .B2(n20236), .A(n16041), .ZN(n16043) );
  OAI21_X1 U18265 ( .B1(n21822), .B2(n16182), .A(n16043), .ZN(P1_U2970) );
  NAND2_X1 U18266 ( .A1(n16044), .A2(n16045), .ZN(n16049) );
  OAI21_X1 U18267 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n16046), .A(
        n16049), .ZN(n16048) );
  INV_X1 U18268 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16198) );
  MUX2_X1 U18269 ( .A(n16198), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n20231), .Z(n16047) );
  OAI211_X1 U18270 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16049), .A(
        n16048), .B(n16047), .ZN(n16050) );
  XOR2_X1 U18271 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n16050), .Z(
        n16192) );
  NOR2_X1 U18272 ( .A1(n21596), .A2(n17362), .ZN(n16186) );
  AOI21_X1 U18273 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16186), .ZN(n16051) );
  OAI21_X1 U18274 ( .B1(n20240), .B2(n16052), .A(n16051), .ZN(n16053) );
  AOI21_X1 U18275 ( .B1(n16054), .B2(n20236), .A(n16053), .ZN(n16055) );
  OAI21_X1 U18276 ( .B1(n21822), .B2(n16192), .A(n16055), .ZN(P1_U2971) );
  XNOR2_X1 U18277 ( .A(n12179), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16056) );
  XNOR2_X1 U18278 ( .A(n16057), .B(n16056), .ZN(n16203) );
  NOR2_X1 U18279 ( .A1(n21596), .A2(n16058), .ZN(n16195) );
  AOI21_X1 U18280 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16195), .ZN(n16059) );
  OAI21_X1 U18281 ( .B1(n20240), .B2(n16060), .A(n16059), .ZN(n16061) );
  AOI21_X1 U18282 ( .B1(n16062), .B2(n20236), .A(n16061), .ZN(n16063) );
  OAI21_X1 U18283 ( .B1(n16203), .B2(n21822), .A(n16063), .ZN(P1_U2972) );
  OAI21_X1 U18284 ( .B1(n11075), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16064), .ZN(n16212) );
  INV_X1 U18285 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n16065) );
  NOR2_X1 U18286 ( .A1(n21596), .A2(n16065), .ZN(n16206) );
  AOI21_X1 U18287 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16206), .ZN(n16066) );
  OAI21_X1 U18288 ( .B1(n20240), .B2(n16067), .A(n16066), .ZN(n16068) );
  AOI21_X1 U18289 ( .B1(n16069), .B2(n20236), .A(n16068), .ZN(n16070) );
  OAI21_X1 U18290 ( .B1(n21822), .B2(n16212), .A(n16070), .ZN(P1_U2973) );
  NOR2_X1 U18291 ( .A1(n16044), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16072) );
  NAND2_X1 U18292 ( .A1(n11209), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16088) );
  OAI211_X1 U18293 ( .C1(n16072), .C2(n16214), .A(n16071), .B(n16088), .ZN(
        n16074) );
  XNOR2_X1 U18294 ( .A(n16074), .B(n16073), .ZN(n16221) );
  INV_X1 U18295 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n17367) );
  NOR2_X1 U18296 ( .A1(n21596), .A2(n17367), .ZN(n16218) );
  AOI21_X1 U18297 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16218), .ZN(n16075) );
  OAI21_X1 U18298 ( .B1(n20240), .B2(n16076), .A(n16075), .ZN(n16077) );
  AOI21_X1 U18299 ( .B1(n16078), .B2(n20236), .A(n16077), .ZN(n16079) );
  OAI21_X1 U18300 ( .B1(n21822), .B2(n16221), .A(n16079), .ZN(P1_U2974) );
  NAND2_X1 U18301 ( .A1(n11209), .A2(n16223), .ZN(n16081) );
  NAND3_X1 U18302 ( .A1(n16044), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n20231), .ZN(n16080) );
  OAI21_X1 U18303 ( .B1(n16044), .B2(n16081), .A(n16080), .ZN(n16082) );
  XNOR2_X1 U18304 ( .A(n16082), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16233) );
  NOR2_X1 U18305 ( .A1(n21596), .A2(n17161), .ZN(n16224) );
  AOI21_X1 U18306 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16224), .ZN(n16083) );
  OAI21_X1 U18307 ( .B1(n20240), .B2(n16084), .A(n16083), .ZN(n16085) );
  AOI21_X1 U18308 ( .B1(n16086), .B2(n20236), .A(n16085), .ZN(n16087) );
  OAI21_X1 U18309 ( .B1(n16233), .B2(n21822), .A(n16087), .ZN(P1_U2975) );
  OAI21_X1 U18310 ( .B1(n11209), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16088), .ZN(n16089) );
  XOR2_X1 U18311 ( .A(n16089), .B(n16044), .Z(n16241) );
  INV_X1 U18312 ( .A(n16090), .ZN(n16094) );
  NOR2_X1 U18313 ( .A1(n21596), .A2(n17260), .ZN(n16234) );
  AOI21_X1 U18314 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16234), .ZN(n16091) );
  OAI21_X1 U18315 ( .B1(n20240), .B2(n16092), .A(n16091), .ZN(n16093) );
  AOI21_X1 U18316 ( .B1(n16094), .B2(n20236), .A(n16093), .ZN(n16095) );
  OAI21_X1 U18317 ( .B1(n16241), .B2(n21822), .A(n16095), .ZN(P1_U2976) );
  NAND2_X1 U18318 ( .A1(n16096), .A2(n16097), .ZN(n16099) );
  XNOR2_X1 U18319 ( .A(n16099), .B(n16098), .ZN(n16260) );
  INV_X1 U18320 ( .A(n21814), .ZN(n16103) );
  INV_X1 U18321 ( .A(n21817), .ZN(n16101) );
  INV_X1 U18322 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21803) );
  NOR2_X1 U18323 ( .A1(n21596), .A2(n21803), .ZN(n16250) );
  AOI21_X1 U18324 ( .B1(n20230), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16250), .ZN(n16100) );
  OAI21_X1 U18325 ( .B1(n20240), .B2(n16101), .A(n16100), .ZN(n16102) );
  AOI21_X1 U18326 ( .B1(n16103), .B2(n20236), .A(n16102), .ZN(n16104) );
  OAI21_X1 U18327 ( .B1(n21822), .B2(n16260), .A(n16104), .ZN(P1_U2977) );
  INV_X1 U18328 ( .A(n10984), .ZN(n16112) );
  MUX2_X1 U18329 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n12349), .S(
        n20231), .Z(n16113) );
  AOI21_X1 U18330 ( .B1(n11209), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16111), .ZN(n20227) );
  OAI22_X1 U18331 ( .A1(n20227), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n11209), .B2(n16111), .ZN(n20233) );
  AOI21_X1 U18332 ( .B1(n11209), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n20233), .ZN(n16106) );
  XNOR2_X1 U18333 ( .A(n16106), .B(n12355), .ZN(n21611) );
  AOI22_X1 U18334 ( .A1(n20230), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n21639), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n16108) );
  NAND2_X1 U18335 ( .A1(n20222), .A2(n21786), .ZN(n16107) );
  OAI211_X1 U18336 ( .C1(n21784), .C2(n16118), .A(n16108), .B(n16107), .ZN(
        n16109) );
  AOI21_X1 U18337 ( .B1(n21611), .B2(n20237), .A(n16109), .ZN(n16110) );
  INV_X1 U18338 ( .A(n16110), .ZN(P1_U2979) );
  AOI21_X1 U18339 ( .B1(n16113), .B2(n16112), .A(n16111), .ZN(n21581) );
  NAND2_X1 U18340 ( .A1(n21581), .A2(n20237), .ZN(n16117) );
  OAI22_X1 U18341 ( .A1(n16114), .A2(n21756), .B1(n21596), .B2(n21757), .ZN(
        n16115) );
  AOI21_X1 U18342 ( .B1(n21762), .B2(n20222), .A(n16115), .ZN(n16116) );
  OAI211_X1 U18343 ( .C1(n16118), .C2(n21760), .A(n16117), .B(n16116), .ZN(
        P1_U2981) );
  NAND2_X1 U18344 ( .A1(n11209), .A2(n21597), .ZN(n16124) );
  NAND2_X1 U18345 ( .A1(n20231), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16123) );
  INV_X1 U18346 ( .A(n16120), .ZN(n16134) );
  AOI211_X1 U18347 ( .C1(n11209), .C2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16134), .B(n16132), .ZN(n16121) );
  OAI21_X1 U18348 ( .B1(n11024), .B2(n16122), .A(n16121), .ZN(n20208) );
  MUX2_X1 U18349 ( .A(n16124), .B(n16123), .S(n20208), .Z(n16125) );
  XNOR2_X1 U18350 ( .A(n16125), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n21601) );
  INV_X1 U18351 ( .A(n21601), .ZN(n16131) );
  INV_X1 U18352 ( .A(n21751), .ZN(n16127) );
  AOI22_X1 U18353 ( .A1(n20230), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n21639), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16126) );
  OAI21_X1 U18354 ( .B1(n16127), .B2(n20240), .A(n16126), .ZN(n16128) );
  AOI21_X1 U18355 ( .B1(n16129), .B2(n20236), .A(n16128), .ZN(n16130) );
  OAI21_X1 U18356 ( .B1(n16131), .B2(n21822), .A(n16130), .ZN(P1_U2983) );
  INV_X1 U18357 ( .A(n16132), .ZN(n16133) );
  NAND2_X1 U18358 ( .A1(n11024), .A2(n16133), .ZN(n20216) );
  AOI21_X1 U18359 ( .B1(n20216), .B2(n16135), .A(n16134), .ZN(n16137) );
  XNOR2_X1 U18360 ( .A(n12179), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16136) );
  XNOR2_X1 U18361 ( .A(n16137), .B(n16136), .ZN(n21459) );
  INV_X1 U18362 ( .A(n21459), .ZN(n16143) );
  AOI22_X1 U18363 ( .A1(n20230), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n21639), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16138) );
  OAI21_X1 U18364 ( .B1(n20240), .B2(n16139), .A(n16138), .ZN(n16140) );
  AOI21_X1 U18365 ( .B1(n16141), .B2(n20236), .A(n16140), .ZN(n16142) );
  OAI21_X1 U18366 ( .B1(n16143), .B2(n21822), .A(n16142), .ZN(P1_U2985) );
  INV_X1 U18367 ( .A(n11024), .ZN(n20183) );
  INV_X1 U18368 ( .A(n16144), .ZN(n16145) );
  AOI21_X1 U18369 ( .B1(n20183), .B2(n16146), .A(n16145), .ZN(n20200) );
  NAND2_X1 U18370 ( .A1(n20200), .A2(n20199), .ZN(n20198) );
  XNOR2_X1 U18371 ( .A(n16149), .B(n16148), .ZN(n16276) );
  AOI22_X1 U18372 ( .A1(n20230), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n21639), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n16150) );
  OAI21_X1 U18373 ( .B1(n20240), .B2(n16151), .A(n16150), .ZN(n16152) );
  AOI21_X1 U18374 ( .B1(n20133), .B2(n20236), .A(n16152), .ZN(n16153) );
  OAI21_X1 U18375 ( .B1(n16276), .B2(n21822), .A(n16153), .ZN(P1_U2986) );
  INV_X1 U18376 ( .A(n11483), .ZN(n20184) );
  AOI21_X1 U18377 ( .B1(n16155), .B2(n16154), .A(n20184), .ZN(n21531) );
  INV_X1 U18378 ( .A(n21738), .ZN(n16159) );
  INV_X1 U18379 ( .A(n21740), .ZN(n16157) );
  AOI22_X1 U18380 ( .A1(n20230), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n21639), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n16156) );
  OAI21_X1 U18381 ( .B1(n20240), .B2(n16157), .A(n16156), .ZN(n16158) );
  AOI21_X1 U18382 ( .B1(n16159), .B2(n20236), .A(n16158), .ZN(n16160) );
  OAI21_X1 U18383 ( .B1(n21531), .B2(n21822), .A(n16160), .ZN(P1_U2990) );
  INV_X1 U18384 ( .A(n16161), .ZN(n16170) );
  OAI211_X1 U18385 ( .C1(n16162), .C2(n16174), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n21515), .ZN(n16168) );
  INV_X1 U18386 ( .A(n16163), .ZN(n16167) );
  NAND3_X1 U18387 ( .A1(n16165), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16164), .ZN(n16166) );
  NAND3_X1 U18388 ( .A1(n16168), .A2(n16167), .A3(n16166), .ZN(n16169) );
  AOI21_X1 U18389 ( .B1(n16170), .B2(n21625), .A(n16169), .ZN(n16171) );
  OAI21_X1 U18390 ( .B1(n16172), .B2(n21635), .A(n16171), .ZN(P1_U3000) );
  INV_X1 U18391 ( .A(n16173), .ZN(n16177) );
  NOR3_X1 U18392 ( .A1(n16194), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16174), .ZN(n16175) );
  AOI211_X1 U18393 ( .C1(n16177), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16176), .B(n16175), .ZN(n16181) );
  INV_X1 U18394 ( .A(n16178), .ZN(n16179) );
  NAND2_X1 U18395 ( .A1(n16179), .A2(n21625), .ZN(n16180) );
  OAI211_X1 U18396 ( .C1(n16182), .C2(n21635), .A(n16181), .B(n16180), .ZN(
        P1_U3002) );
  INV_X1 U18397 ( .A(n16199), .ZN(n16187) );
  NOR3_X1 U18398 ( .A1(n16194), .A2(n16184), .A3(n16183), .ZN(n16185) );
  AOI211_X1 U18399 ( .C1(n16187), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16186), .B(n16185), .ZN(n16191) );
  INV_X1 U18400 ( .A(n16188), .ZN(n16189) );
  NAND2_X1 U18401 ( .A1(n16189), .A2(n21625), .ZN(n16190) );
  OAI211_X1 U18402 ( .C1(n16192), .C2(n21635), .A(n16191), .B(n16190), .ZN(
        P1_U3003) );
  INV_X1 U18403 ( .A(n16193), .ZN(n16201) );
  INV_X1 U18404 ( .A(n16194), .ZN(n16196) );
  AOI21_X1 U18405 ( .B1(n16196), .B2(n16198), .A(n16195), .ZN(n16197) );
  OAI21_X1 U18406 ( .B1(n16199), .B2(n16198), .A(n16197), .ZN(n16200) );
  AOI21_X1 U18407 ( .B1(n16201), .B2(n21625), .A(n16200), .ZN(n16202) );
  OAI21_X1 U18408 ( .B1(n16203), .B2(n21635), .A(n16202), .ZN(P1_U3004) );
  INV_X1 U18409 ( .A(n16216), .ZN(n16207) );
  INV_X1 U18410 ( .A(n16225), .ZN(n16237) );
  NOR3_X1 U18411 ( .A1(n16237), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n16204), .ZN(n16205) );
  AOI211_X1 U18412 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n16207), .A(
        n16206), .B(n16205), .ZN(n16211) );
  INV_X1 U18413 ( .A(n16208), .ZN(n16209) );
  NAND2_X1 U18414 ( .A1(n16209), .A2(n21625), .ZN(n16210) );
  OAI211_X1 U18415 ( .C1(n16212), .C2(n21635), .A(n16211), .B(n16210), .ZN(
        P1_U3005) );
  INV_X1 U18416 ( .A(n16213), .ZN(n16219) );
  AOI21_X1 U18417 ( .B1(n16225), .B2(n16214), .A(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16215) );
  NOR2_X1 U18418 ( .A1(n16216), .A2(n16215), .ZN(n16217) );
  AOI211_X1 U18419 ( .C1(n16219), .C2(n21625), .A(n16218), .B(n16217), .ZN(
        n16220) );
  OAI21_X1 U18420 ( .B1(n16221), .B2(n21635), .A(n16220), .ZN(P1_U3006) );
  INV_X1 U18421 ( .A(n16222), .ZN(n16231) );
  AOI21_X1 U18422 ( .B1(n21573), .B2(n16223), .A(n16235), .ZN(n16229) );
  INV_X1 U18423 ( .A(n16224), .ZN(n16227) );
  NAND3_X1 U18424 ( .A1(n16225), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n16228), .ZN(n16226) );
  OAI211_X1 U18425 ( .C1(n16229), .C2(n16228), .A(n16227), .B(n16226), .ZN(
        n16230) );
  AOI21_X1 U18426 ( .B1(n16231), .B2(n21625), .A(n16230), .ZN(n16232) );
  OAI21_X1 U18427 ( .B1(n16233), .B2(n21635), .A(n16232), .ZN(P1_U3007) );
  AOI21_X1 U18428 ( .B1(n16235), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16234), .ZN(n16236) );
  OAI21_X1 U18429 ( .B1(n16237), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16236), .ZN(n16238) );
  AOI21_X1 U18430 ( .B1(n16239), .B2(n21625), .A(n16238), .ZN(n16240) );
  OAI21_X1 U18431 ( .B1(n16241), .B2(n21635), .A(n16240), .ZN(P1_U3008) );
  INV_X1 U18432 ( .A(n21811), .ZN(n16251) );
  INV_X1 U18433 ( .A(n16273), .ZN(n16242) );
  OR2_X1 U18434 ( .A1(n21501), .A2(n16242), .ZN(n16244) );
  NAND2_X1 U18435 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16264), .ZN(
        n16265) );
  OR2_X1 U18436 ( .A1(n16268), .A2(n16265), .ZN(n16243) );
  NAND2_X1 U18437 ( .A1(n16244), .A2(n16243), .ZN(n16262) );
  NAND2_X1 U18438 ( .A1(n16262), .A2(n16245), .ZN(n21615) );
  OR2_X1 U18439 ( .A1(n21608), .A2(n21616), .ZN(n16246) );
  NAND2_X1 U18440 ( .A1(n21615), .A2(n16246), .ZN(n21606) );
  INV_X1 U18441 ( .A(n21606), .ZN(n16248) );
  NOR3_X1 U18442 ( .A1(n16248), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n16247), .ZN(n16249) );
  AOI211_X1 U18443 ( .C1(n16251), .C2(n21625), .A(n16250), .B(n16249), .ZN(
        n16259) );
  NAND2_X1 U18444 ( .A1(n16264), .A2(n16252), .ZN(n21571) );
  AND2_X1 U18445 ( .A1(n16252), .A2(n16273), .ZN(n21574) );
  OAI21_X1 U18446 ( .B1(n21574), .B2(n21501), .A(n21554), .ZN(n16253) );
  AOI21_X1 U18447 ( .B1(n21551), .B2(n21571), .A(n16253), .ZN(n21576) );
  OAI21_X1 U18448 ( .B1(n21585), .B2(n21534), .A(n21576), .ZN(n21591) );
  AOI21_X1 U18449 ( .B1(n12349), .B2(n21633), .A(n21591), .ZN(n21621) );
  INV_X1 U18450 ( .A(n21621), .ZN(n16254) );
  NAND2_X1 U18451 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16255) );
  OAI21_X1 U18452 ( .B1(n16254), .B2(n16255), .A(n21515), .ZN(n21628) );
  INV_X1 U18453 ( .A(n21628), .ZN(n16257) );
  NOR2_X1 U18454 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n16255), .ZN(
        n16256) );
  AND2_X1 U18455 ( .A1(n21606), .A2(n16256), .ZN(n21622) );
  OAI21_X1 U18456 ( .B1(n16257), .B2(n21622), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16258) );
  OAI211_X1 U18457 ( .C1(n16260), .C2(n21635), .A(n16259), .B(n16258), .ZN(
        P1_U3009) );
  NOR3_X1 U18458 ( .A1(n12189), .A2(n12191), .A3(n21556), .ZN(n21465) );
  AOI21_X1 U18459 ( .B1(n16261), .B2(n21465), .A(n21608), .ZN(n16270) );
  NOR2_X1 U18460 ( .A1(n21596), .A2(n20082), .ZN(n16263) );
  AND2_X1 U18461 ( .A1(n12189), .A2(n16262), .ZN(n21467) );
  AOI211_X1 U18462 ( .C1(n16264), .C2(n16270), .A(n16263), .B(n21467), .ZN(
        n16275) );
  INV_X1 U18463 ( .A(n16265), .ZN(n16267) );
  OAI21_X1 U18464 ( .B1(n16268), .B2(n16267), .A(n16266), .ZN(n16269) );
  INV_X1 U18465 ( .A(n16269), .ZN(n16272) );
  INV_X1 U18466 ( .A(n16270), .ZN(n16271) );
  OAI211_X1 U18467 ( .C1(n16273), .C2(n21501), .A(n16272), .B(n16271), .ZN(
        n21466) );
  AOI22_X1 U18468 ( .A1(n21466), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n21625), .B2(n20130), .ZN(n16274) );
  OAI211_X1 U18469 ( .C1(n16276), .C2(n21635), .A(n16275), .B(n16274), .ZN(
        P1_U3018) );
  AOI22_X1 U18470 ( .A1(n21893), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16277), 
        .B2(n14662), .ZN(n16280) );
  NAND2_X1 U18471 ( .A1(n18899), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16282) );
  INV_X1 U18472 ( .A(n16282), .ZN(n16278) );
  OAI22_X1 U18473 ( .A1(n16280), .A2(n16279), .B1(n16278), .B2(n18900), .ZN(
        n16285) );
  OAI22_X1 U18474 ( .A1(n18907), .A2(n17480), .B1(n16282), .B2(n16281), .ZN(
        n16283) );
  NOR2_X1 U18475 ( .A1(n17388), .A2(n16283), .ZN(n16284) );
  MUX2_X1 U18476 ( .A(n16285), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n16284), 
        .Z(P2_U3610) );
  INV_X1 U18477 ( .A(n16286), .ZN(n16345) );
  AND2_X1 U18478 ( .A1(n17388), .A2(n16287), .ZN(n16290) );
  AND2_X1 U18479 ( .A1(n14662), .A2(n18899), .ZN(n16332) );
  INV_X1 U18480 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16384) );
  NOR2_X1 U18481 ( .A1(n16332), .A2(n16384), .ZN(n16288) );
  NAND4_X1 U18482 ( .A1(n14662), .A2(n14841), .A3(n19473), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n18888) );
  INV_X1 U18483 ( .A(n18888), .ZN(n18784) );
  AOI21_X1 U18484 ( .B1(n18740), .B2(n16319), .A(n16321), .ZN(n18743) );
  INV_X1 U18485 ( .A(n16317), .ZN(n16291) );
  AOI21_X1 U18486 ( .B1(n16625), .B2(n16316), .A(n16291), .ZN(n18715) );
  AOI21_X1 U18487 ( .B1(n18688), .B2(n16312), .A(n16314), .ZN(n18691) );
  INV_X1 U18488 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16292) );
  AOI21_X1 U18489 ( .B1(n16310), .B2(n16292), .A(n16313), .ZN(n18671) );
  AOI21_X1 U18490 ( .B1(n16694), .B2(n16308), .A(n16311), .ZN(n18644) );
  AOI21_X1 U18491 ( .B1(n18622), .B2(n16306), .A(n16309), .ZN(n18621) );
  AOI21_X1 U18492 ( .B1(n18604), .B2(n16304), .A(n16307), .ZN(n18615) );
  AOI21_X1 U18493 ( .B1(n16302), .B2(n16745), .A(n16305), .ZN(n18591) );
  AOI21_X1 U18494 ( .B1(n17460), .B2(n16300), .A(n16303), .ZN(n18568) );
  AOI21_X1 U18495 ( .B1(n17441), .B2(n16298), .A(n16301), .ZN(n18540) );
  AOI21_X1 U18496 ( .B1(n17414), .B2(n16294), .A(n16297), .ZN(n18501) );
  AOI21_X1 U18497 ( .B1(n17400), .B2(n16293), .A(n16295), .ZN(n17389) );
  OAI22_X1 U18498 ( .A1(n14841), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n18462) );
  OAI22_X1 U18499 ( .A1(n14841), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n18473), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17064) );
  AND2_X1 U18500 ( .A1(n18462), .A2(n17064), .ZN(n16371) );
  NAND2_X1 U18501 ( .A1(n16371), .A2(n16373), .ZN(n16359) );
  NOR2_X1 U18502 ( .A1(n17389), .A2(n16359), .ZN(n18488) );
  OAI21_X1 U18503 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16295), .A(
        n16294), .ZN(n18487) );
  NAND2_X1 U18504 ( .A1(n18488), .A2(n18487), .ZN(n18499) );
  NOR2_X1 U18505 ( .A1(n18501), .A2(n18499), .ZN(n18510) );
  OAI21_X1 U18506 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16297), .A(
        n16296), .ZN(n18511) );
  NAND2_X1 U18507 ( .A1(n18510), .A2(n18511), .ZN(n18517) );
  NOR2_X1 U18508 ( .A1(n18518), .A2(n18517), .ZN(n18532) );
  OAI21_X1 U18509 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16299), .A(
        n16298), .ZN(n18533) );
  NAND2_X1 U18510 ( .A1(n18532), .A2(n18533), .ZN(n18539) );
  NOR2_X1 U18511 ( .A1(n18540), .A2(n18539), .ZN(n18557) );
  OAI21_X1 U18512 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16301), .A(
        n16300), .ZN(n18558) );
  NAND2_X1 U18513 ( .A1(n18557), .A2(n18558), .ZN(n18566) );
  NOR2_X1 U18514 ( .A1(n18568), .A2(n18566), .ZN(n18573) );
  OAI21_X1 U18515 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16303), .A(
        n16302), .ZN(n18574) );
  NAND2_X1 U18516 ( .A1(n18573), .A2(n18574), .ZN(n18585) );
  NOR2_X1 U18517 ( .A1(n18591), .A2(n18585), .ZN(n18584) );
  OAI21_X1 U18518 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16305), .A(
        n16304), .ZN(n18595) );
  NAND2_X1 U18519 ( .A1(n18584), .A2(n18595), .ZN(n18608) );
  NOR2_X1 U18520 ( .A1(n18615), .A2(n18608), .ZN(n16346) );
  OAI21_X1 U18521 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16307), .A(
        n16306), .ZN(n16719) );
  NAND2_X1 U18522 ( .A1(n16346), .A2(n16719), .ZN(n18619) );
  NOR2_X1 U18523 ( .A1(n18621), .A2(n18619), .ZN(n18635) );
  OAI21_X1 U18524 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16309), .A(
        n16308), .ZN(n18636) );
  NAND2_X1 U18525 ( .A1(n18635), .A2(n18636), .ZN(n18642) );
  NOR2_X1 U18526 ( .A1(n18644), .A2(n18642), .ZN(n18654) );
  OAI21_X1 U18527 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n16311), .A(
        n16310), .ZN(n18656) );
  NAND2_X1 U18528 ( .A1(n18654), .A2(n18656), .ZN(n18668) );
  NOR2_X1 U18529 ( .A1(n18671), .A2(n18668), .ZN(n18676) );
  OAI21_X1 U18530 ( .B1(n16313), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16312), .ZN(n18677) );
  NAND2_X1 U18531 ( .A1(n18676), .A2(n18677), .ZN(n18689) );
  NOR2_X1 U18532 ( .A1(n18691), .A2(n18689), .ZN(n18701) );
  OR2_X1 U18533 ( .A1(n16314), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16315) );
  AND2_X1 U18534 ( .A1(n16316), .A2(n16315), .ZN(n18703) );
  INV_X1 U18535 ( .A(n18703), .ZN(n16635) );
  NAND2_X1 U18536 ( .A1(n18701), .A2(n16635), .ZN(n18712) );
  NOR2_X1 U18537 ( .A1(n18715), .A2(n18712), .ZN(n18725) );
  NAND2_X1 U18538 ( .A1(n16317), .A2(n16614), .ZN(n16318) );
  AND2_X1 U18539 ( .A1(n16319), .A2(n16318), .ZN(n18727) );
  INV_X1 U18540 ( .A(n18727), .ZN(n16320) );
  NAND2_X1 U18541 ( .A1(n18725), .A2(n16320), .ZN(n18741) );
  NOR2_X1 U18542 ( .A1(n18743), .A2(n18741), .ZN(n18752) );
  NOR2_X1 U18543 ( .A1(n16321), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16322) );
  OR2_X1 U18544 ( .A1(n16323), .A2(n16322), .ZN(n18754) );
  NAND2_X1 U18545 ( .A1(n18752), .A2(n18754), .ZN(n18767) );
  NOR2_X1 U18546 ( .A1(n18770), .A2(n18767), .ZN(n18782) );
  XNOR2_X1 U18547 ( .A(n16324), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18787) );
  INV_X1 U18548 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16338) );
  AND4_X1 U18549 ( .A1(n18784), .A2(n18782), .A3(n18787), .A4(n11029), .ZN(
        n16343) );
  INV_X1 U18550 ( .A(n16326), .ZN(n16327) );
  NAND2_X1 U18551 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19473), .ZN(n18891) );
  OR3_X1 U18552 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19472), .A3(n18891), 
        .ZN(n16329) );
  NAND3_X1 U18553 ( .A1(n18888), .A2(n18848), .A3(n16329), .ZN(n16330) );
  NOR2_X1 U18554 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n16331), .ZN(n16333) );
  OAI22_X1 U18555 ( .A1(n16334), .A2(n16333), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n16332), .ZN(n16335) );
  AND2_X1 U18556 ( .A1(n16336), .A2(n16335), .ZN(n16337) );
  NAND2_X1 U18557 ( .A1(n17388), .A2(n16337), .ZN(n18788) );
  OAI22_X1 U18558 ( .A1(n18788), .A2(n16384), .B1(n18765), .B2(n16338), .ZN(
        n16339) );
  AOI21_X1 U18559 ( .B1(P2_REIP_REG_31__SCAN_IN), .B2(n18755), .A(n16339), 
        .ZN(n16340) );
  OAI21_X1 U18560 ( .B1(n16341), .B2(n18780), .A(n16340), .ZN(n16342) );
  OAI21_X1 U18561 ( .B1(n16345), .B2(n18800), .A(n16344), .ZN(P2_U2824) );
  OR2_X1 U18562 ( .A1(n18783), .A2(n16346), .ZN(n18607) );
  XOR2_X1 U18563 ( .A(n16719), .B(n18607), .Z(n16352) );
  NOR2_X1 U18564 ( .A1(n16349), .A2(n16348), .ZN(n16350) );
  OR2_X1 U18565 ( .A1(n16347), .A2(n16350), .ZN(n16934) );
  OAI22_X1 U18566 ( .A1(n16717), .A2(n18737), .B1(n16934), .B2(n18780), .ZN(
        n16351) );
  AOI21_X1 U18567 ( .B1(n16352), .B2(n18784), .A(n16351), .ZN(n16358) );
  NOR2_X1 U18568 ( .A1(n18788), .A2(n12606), .ZN(n16356) );
  INV_X1 U18569 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16354) );
  OAI22_X1 U18570 ( .A1(n16354), .A2(n18765), .B1(n16353), .B2(n18800), .ZN(
        n16355) );
  NOR3_X1 U18571 ( .A1(n16356), .A2(n16675), .A3(n16355), .ZN(n16357) );
  OAI211_X1 U18572 ( .C1(n17557), .C2(n18791), .A(n16358), .B(n16357), .ZN(
        P2_U2839) );
  NAND2_X1 U18573 ( .A1(n11029), .A2(n16359), .ZN(n16360) );
  XNOR2_X1 U18574 ( .A(n17389), .B(n16360), .ZN(n16361) );
  NAND2_X1 U18575 ( .A1(n16361), .A2(n18784), .ZN(n16370) );
  XNOR2_X1 U18576 ( .A(n16362), .B(n11118), .ZN(n19712) );
  INV_X1 U18577 ( .A(n16363), .ZN(n16364) );
  AOI22_X1 U18578 ( .A1(n18776), .A2(n16364), .B1(P2_EBX_REG_3__SCAN_IN), .B2(
        n18774), .ZN(n16365) );
  OAI21_X1 U18579 ( .B1(n18850), .B2(n18737), .A(n16365), .ZN(n16368) );
  INV_X1 U18580 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n16366) );
  OAI22_X1 U18581 ( .A1(n17400), .A2(n18765), .B1(n16366), .B2(n18791), .ZN(
        n16367) );
  AOI211_X1 U18582 ( .C1(n18795), .C2(n19712), .A(n16368), .B(n16367), .ZN(
        n16369) );
  OAI211_X1 U18583 ( .C1(n19613), .C2(n18485), .A(n16370), .B(n16369), .ZN(
        P2_U2852) );
  INV_X1 U18584 ( .A(n16373), .ZN(n16374) );
  INV_X1 U18585 ( .A(n17063), .ZN(n16372) );
  AOI221_X1 U18586 ( .B1(n16374), .B2(n17063), .C1(n16373), .C2(n16372), .A(
        n18888), .ZN(n16375) );
  INV_X1 U18587 ( .A(n16375), .ZN(n16382) );
  AOI22_X1 U18588 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18794), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n18755), .ZN(n16377) );
  NAND2_X1 U18589 ( .A1(n18774), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n16376) );
  OAI211_X1 U18590 ( .C1(n18800), .C2(n16378), .A(n16377), .B(n16376), .ZN(
        n16380) );
  NOR2_X1 U18591 ( .A1(n14331), .A2(n18737), .ZN(n16379) );
  AOI211_X1 U18592 ( .C1(n19608), .C2(n18795), .A(n16380), .B(n16379), .ZN(
        n16381) );
  OAI211_X1 U18593 ( .C1(n19611), .C2(n18485), .A(n16382), .B(n16381), .ZN(
        P2_U2853) );
  NAND2_X1 U18594 ( .A1(n16289), .A2(n16448), .ZN(n16383) );
  OAI21_X1 U18595 ( .B1(n16448), .B2(n16384), .A(n16383), .ZN(P2_U2856) );
  INV_X1 U18596 ( .A(n16385), .ZN(n16386) );
  NOR2_X1 U18597 ( .A1(n16387), .A2(n16386), .ZN(n16389) );
  XNOR2_X1 U18598 ( .A(n16389), .B(n16388), .ZN(n16484) );
  NOR2_X1 U18599 ( .A1(n16390), .A2(n16433), .ZN(n16391) );
  AOI21_X1 U18600 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n16433), .A(n16391), .ZN(
        n16392) );
  OAI21_X1 U18601 ( .B1(n16484), .B2(n16474), .A(n16392), .ZN(P2_U2858) );
  INV_X1 U18602 ( .A(n16393), .ZN(n16403) );
  NAND2_X1 U18603 ( .A1(n16403), .A2(n16394), .ZN(n16396) );
  XNOR2_X1 U18604 ( .A(n16396), .B(n16395), .ZN(n16494) );
  INV_X1 U18605 ( .A(n16397), .ZN(n16406) );
  AND2_X1 U18606 ( .A1(n16406), .A2(n16398), .ZN(n16399) );
  OR2_X1 U18607 ( .A1(n13137), .A2(n16399), .ZN(n16775) );
  NOR2_X1 U18608 ( .A1(n16775), .A2(n16433), .ZN(n16400) );
  AOI21_X1 U18609 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16433), .A(n16400), .ZN(
        n16401) );
  OAI21_X1 U18610 ( .B1(n16494), .B2(n16474), .A(n16401), .ZN(P2_U2859) );
  NAND2_X1 U18611 ( .A1(n16403), .A2(n16402), .ZN(n16404) );
  XOR2_X1 U18612 ( .A(n16405), .B(n16404), .Z(n16503) );
  NAND2_X1 U18613 ( .A1(n16433), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16409) );
  AOI21_X1 U18614 ( .B1(n16407), .B2(n16412), .A(n16397), .ZN(n18748) );
  NAND2_X1 U18615 ( .A1(n18748), .A2(n16448), .ZN(n16408) );
  OAI211_X1 U18616 ( .C1(n16503), .C2(n16474), .A(n16409), .B(n16408), .ZN(
        P2_U2860) );
  OR2_X1 U18617 ( .A1(n16422), .A2(n16410), .ZN(n16411) );
  NAND2_X1 U18618 ( .A1(n16412), .A2(n16411), .ZN(n18738) );
  AOI21_X1 U18619 ( .B1(n16413), .B2(n16415), .A(n16414), .ZN(n16504) );
  NAND2_X1 U18620 ( .A1(n16504), .A2(n16457), .ZN(n16417) );
  NAND2_X1 U18621 ( .A1(n16433), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16416) );
  OAI211_X1 U18622 ( .C1(n18738), .C2(n16433), .A(n16417), .B(n16416), .ZN(
        P2_U2861) );
  OAI21_X1 U18623 ( .B1(n16418), .B2(n16420), .A(n16419), .ZN(n16520) );
  AND2_X1 U18624 ( .A1(n16431), .A2(n16421), .ZN(n16423) );
  OR2_X1 U18625 ( .A1(n16423), .A2(n16422), .ZN(n16623) );
  NOR2_X1 U18626 ( .A1(n16623), .A2(n16433), .ZN(n16424) );
  AOI21_X1 U18627 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n16433), .A(n16424), .ZN(
        n16425) );
  OAI21_X1 U18628 ( .B1(n16520), .B2(n16474), .A(n16425), .ZN(P2_U2862) );
  OAI21_X1 U18629 ( .B1(n16428), .B2(n16427), .A(n16426), .ZN(n16526) );
  NAND2_X1 U18630 ( .A1(n16438), .A2(n16429), .ZN(n16430) );
  AND2_X1 U18631 ( .A1(n16431), .A2(n16430), .ZN(n18707) );
  INV_X1 U18632 ( .A(n18707), .ZN(n16825) );
  NOR2_X1 U18633 ( .A1(n16825), .A2(n16433), .ZN(n16432) );
  AOI21_X1 U18634 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16433), .A(n16432), .ZN(
        n16434) );
  OAI21_X1 U18635 ( .B1(n16526), .B2(n16474), .A(n16434), .ZN(P2_U2863) );
  XNOR2_X1 U18636 ( .A(n11079), .B(n16435), .ZN(n16536) );
  NAND2_X1 U18637 ( .A1(n16433), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16440) );
  OR2_X1 U18638 ( .A1(n16445), .A2(n16436), .ZN(n16437) );
  AND2_X1 U18639 ( .A1(n16438), .A2(n16437), .ZN(n18696) );
  NAND2_X1 U18640 ( .A1(n18696), .A2(n16448), .ZN(n16439) );
  OAI211_X1 U18641 ( .C1(n16536), .C2(n16474), .A(n16440), .B(n16439), .ZN(
        P2_U2864) );
  INV_X1 U18642 ( .A(n16441), .ZN(n16455) );
  NAND2_X1 U18643 ( .A1(n16455), .A2(n16442), .ZN(n16443) );
  NAND2_X1 U18644 ( .A1(n11079), .A2(n16443), .ZN(n19550) );
  NAND2_X1 U18645 ( .A1(n16433), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16450) );
  INV_X1 U18646 ( .A(n16444), .ZN(n16447) );
  INV_X1 U18647 ( .A(n16452), .ZN(n16446) );
  AOI21_X1 U18648 ( .B1(n16447), .B2(n16446), .A(n16445), .ZN(n18683) );
  NAND2_X1 U18649 ( .A1(n18683), .A2(n16448), .ZN(n16449) );
  OAI211_X1 U18650 ( .C1(n19550), .C2(n16474), .A(n16450), .B(n16449), .ZN(
        P2_U2865) );
  AND2_X1 U18651 ( .A1(n11050), .A2(n16451), .ZN(n16453) );
  OR2_X1 U18652 ( .A1(n16453), .A2(n16452), .ZN(n16674) );
  AOI21_X1 U18653 ( .B1(n16456), .B2(n16461), .A(n16441), .ZN(n16537) );
  NAND2_X1 U18654 ( .A1(n16537), .A2(n16457), .ZN(n16459) );
  NAND2_X1 U18655 ( .A1(n16433), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16458) );
  OAI211_X1 U18656 ( .C1(n16674), .C2(n16433), .A(n16459), .B(n16458), .ZN(
        P2_U2866) );
  OAI21_X1 U18657 ( .B1(n16460), .B2(n16462), .A(n16461), .ZN(n19656) );
  NAND2_X1 U18658 ( .A1(n16463), .A2(n16464), .ZN(n16465) );
  NAND2_X1 U18659 ( .A1(n11050), .A2(n16465), .ZN(n18661) );
  NOR2_X1 U18660 ( .A1(n18661), .A2(n16433), .ZN(n16466) );
  AOI21_X1 U18661 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n16433), .A(n16466), .ZN(
        n16467) );
  OAI21_X1 U18662 ( .B1(n19656), .B2(n16474), .A(n16467), .ZN(P2_U2867) );
  INV_X1 U18663 ( .A(n16460), .ZN(n16468) );
  OAI21_X1 U18664 ( .B1(n15449), .B2(n16469), .A(n16468), .ZN(n16553) );
  OAI21_X1 U18665 ( .B1(n16471), .B2(n16470), .A(n16463), .ZN(n16891) );
  NOR2_X1 U18666 ( .A1(n16891), .A2(n16433), .ZN(n16472) );
  AOI21_X1 U18667 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n16433), .A(n16472), .ZN(
        n16473) );
  OAI21_X1 U18668 ( .B1(n16553), .B2(n16474), .A(n16473), .ZN(P2_U2868) );
  OR2_X1 U18669 ( .A1(n16490), .A2(n16475), .ZN(n16476) );
  NAND2_X1 U18670 ( .A1(n16477), .A2(n16476), .ZN(n18781) );
  OAI22_X1 U18671 ( .A1(n16564), .A2(n19374), .B1(n19556), .B2(n16478), .ZN(
        n16479) );
  AOI21_X1 U18672 ( .B1(n19764), .B2(BUF2_REG_29__SCAN_IN), .A(n16479), .ZN(
        n16481) );
  NAND2_X1 U18673 ( .A1(n19765), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16480) );
  OAI211_X1 U18674 ( .C1(n18781), .C2(n19549), .A(n16481), .B(n16480), .ZN(
        n16482) );
  INV_X1 U18675 ( .A(n16482), .ZN(n16483) );
  OAI21_X1 U18676 ( .B1(n16484), .B2(n19812), .A(n16483), .ZN(P2_U2890) );
  OAI22_X1 U18677 ( .A1(n16564), .A2(n19377), .B1(n19556), .B2(n16485), .ZN(
        n16489) );
  INV_X1 U18678 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n16486) );
  NOR2_X1 U18679 ( .A1(n16487), .A2(n16486), .ZN(n16488) );
  AOI211_X1 U18680 ( .C1(BUF1_REG_28__SCAN_IN), .C2(n19765), .A(n16489), .B(
        n16488), .ZN(n16493) );
  AOI21_X1 U18681 ( .B1(n16491), .B2(n16498), .A(n16490), .ZN(n18759) );
  NAND2_X1 U18682 ( .A1(n18759), .A2(n19860), .ZN(n16492) );
  OAI211_X1 U18683 ( .C1(n16494), .C2(n19812), .A(n16493), .B(n16492), .ZN(
        P2_U2891) );
  OAI22_X1 U18684 ( .A1(n16564), .A2(n19380), .B1(n19556), .B2(n16495), .ZN(
        n16496) );
  AOI21_X1 U18685 ( .B1(n19764), .B2(BUF2_REG_27__SCAN_IN), .A(n16496), .ZN(
        n16502) );
  INV_X1 U18686 ( .A(n16498), .ZN(n16499) );
  AOI21_X1 U18687 ( .B1(n16500), .B2(n16497), .A(n16499), .ZN(n18747) );
  AOI22_X1 U18688 ( .A1(n18747), .A2(n19860), .B1(n19765), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16501) );
  OAI211_X1 U18689 ( .C1(n16503), .C2(n19812), .A(n16502), .B(n16501), .ZN(
        P2_U2892) );
  NAND2_X1 U18690 ( .A1(n16504), .A2(n19862), .ZN(n16510) );
  AOI22_X1 U18691 ( .A1(n19763), .A2(n19384), .B1(n19859), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16509) );
  AOI22_X1 U18692 ( .A1(n19765), .A2(BUF1_REG_26__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n16508) );
  OR2_X1 U18693 ( .A1(n16514), .A2(n16505), .ZN(n16506) );
  AND2_X1 U18694 ( .A1(n16506), .A2(n16497), .ZN(n18733) );
  NAND2_X1 U18695 ( .A1(n18733), .A2(n19860), .ZN(n16507) );
  NAND4_X1 U18696 ( .A1(n16510), .A2(n16509), .A3(n16508), .A4(n16507), .ZN(
        P2_U2893) );
  NOR2_X1 U18697 ( .A1(n16512), .A2(n16511), .ZN(n16513) );
  OR2_X1 U18698 ( .A1(n16514), .A2(n16513), .ZN(n18724) );
  OAI22_X1 U18699 ( .A1(n18724), .A2(n19549), .B1(n19556), .B2(n16515), .ZN(
        n16516) );
  AOI21_X1 U18700 ( .B1(n19763), .B2(n16517), .A(n16516), .ZN(n16519) );
  AOI22_X1 U18701 ( .A1(n19765), .A2(BUF1_REG_25__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n16518) );
  OAI211_X1 U18702 ( .C1(n16520), .C2(n19812), .A(n16519), .B(n16518), .ZN(
        P2_U2894) );
  XNOR2_X1 U18703 ( .A(n16529), .B(n16521), .ZN(n18711) );
  INV_X1 U18704 ( .A(n18711), .ZN(n16822) );
  OAI22_X1 U18705 ( .A1(n16564), .A2(n19391), .B1(n16522), .B2(n19556), .ZN(
        n16523) );
  AOI21_X1 U18706 ( .B1(n16822), .B2(n19860), .A(n16523), .ZN(n16525) );
  AOI22_X1 U18707 ( .A1(n19765), .A2(BUF1_REG_24__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n16524) );
  OAI211_X1 U18708 ( .C1(n16526), .C2(n19812), .A(n16525), .B(n16524), .ZN(
        P2_U2895) );
  AND2_X1 U18709 ( .A1(n16844), .A2(n16527), .ZN(n16528) );
  NOR2_X1 U18710 ( .A1(n16529), .A2(n16528), .ZN(n18695) );
  INV_X1 U18711 ( .A(n18695), .ZN(n16531) );
  OAI22_X1 U18712 ( .A1(n16531), .A2(n19549), .B1(n16530), .B2(n19556), .ZN(
        n16532) );
  AOI21_X1 U18713 ( .B1(n19763), .B2(n16533), .A(n16532), .ZN(n16535) );
  AOI22_X1 U18714 ( .A1(n19765), .A2(BUF1_REG_23__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n16534) );
  OAI211_X1 U18715 ( .C1(n16536), .C2(n19812), .A(n16535), .B(n16534), .ZN(
        P2_U2896) );
  INV_X1 U18716 ( .A(n16537), .ZN(n16545) );
  INV_X1 U18717 ( .A(n16842), .ZN(n16539) );
  AOI21_X1 U18718 ( .B1(n16540), .B2(n16538), .A(n16539), .ZN(n18666) );
  INV_X1 U18719 ( .A(n18666), .ZN(n16857) );
  OAI22_X1 U18720 ( .A1(n16857), .A2(n19549), .B1(n16541), .B2(n19556), .ZN(
        n16542) );
  AOI21_X1 U18721 ( .B1(n19763), .B2(n19607), .A(n16542), .ZN(n16544) );
  AOI22_X1 U18722 ( .A1(n19765), .A2(BUF1_REG_21__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n16543) );
  OAI211_X1 U18723 ( .C1(n16545), .C2(n19812), .A(n16544), .B(n16543), .ZN(
        P2_U2898) );
  AND2_X1 U18724 ( .A1(n16901), .A2(n16546), .ZN(n16547) );
  NOR2_X1 U18725 ( .A1(n16877), .A2(n16547), .ZN(n18649) );
  NOR2_X1 U18726 ( .A1(n19556), .A2(n16548), .ZN(n16550) );
  NOR2_X1 U18727 ( .A1(n16564), .A2(n19719), .ZN(n16549) );
  AOI211_X1 U18728 ( .C1(n18649), .C2(n19860), .A(n16550), .B(n16549), .ZN(
        n16552) );
  AOI22_X1 U18729 ( .A1(n19765), .A2(BUF1_REG_19__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n16551) );
  OAI211_X1 U18730 ( .C1(n16553), .C2(n19812), .A(n16552), .B(n16551), .ZN(
        P2_U2900) );
  AOI22_X1 U18731 ( .A1(n19765), .A2(BUF1_REG_17__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n16557) );
  INV_X1 U18732 ( .A(n16554), .ZN(n16555) );
  XNOR2_X1 U18733 ( .A(n16347), .B(n16555), .ZN(n18627) );
  AOI22_X1 U18734 ( .A1(n19860), .A2(n18627), .B1(n19859), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16556) );
  OAI211_X1 U18735 ( .C1(n19816), .C2(n16564), .A(n16557), .B(n16556), .ZN(
        n16558) );
  AOI21_X1 U18736 ( .B1(n16559), .B2(n19862), .A(n16558), .ZN(n16560) );
  INV_X1 U18737 ( .A(n16560), .ZN(P2_U2902) );
  AOI22_X1 U18738 ( .A1(n19765), .A2(BUF1_REG_16__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n16563) );
  INV_X1 U18739 ( .A(n16934), .ZN(n16561) );
  AOI22_X1 U18740 ( .A1(n19860), .A2(n16561), .B1(n19859), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n16562) );
  OAI211_X1 U18741 ( .C1(n19870), .C2(n16564), .A(n16563), .B(n16562), .ZN(
        n16565) );
  INV_X1 U18742 ( .A(n16565), .ZN(n16566) );
  OAI21_X1 U18743 ( .B1(n16567), .B2(n19812), .A(n16566), .ZN(P2_U2903) );
  NAND2_X1 U18744 ( .A1(n17470), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16568) );
  OAI211_X1 U18745 ( .C1(n17479), .C2(n16570), .A(n16569), .B(n16568), .ZN(
        n16572) );
  OAI21_X1 U18746 ( .B1(n16574), .B2(n17461), .A(n16573), .ZN(P2_U2983) );
  NOR2_X1 U18747 ( .A1(n16576), .A2(n16575), .ZN(n16581) );
  INV_X1 U18748 ( .A(n16577), .ZN(n16579) );
  NAND2_X1 U18749 ( .A1(n16579), .A2(n16578), .ZN(n16580) );
  XNOR2_X1 U18750 ( .A(n16581), .B(n16580), .ZN(n16760) );
  NOR2_X1 U18751 ( .A1(n18848), .A2(n18790), .ZN(n16750) );
  AOI21_X1 U18752 ( .B1(n17470), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16750), .ZN(n16582) );
  OAI21_X1 U18753 ( .B1(n17479), .B2(n18787), .A(n16582), .ZN(n16585) );
  INV_X1 U18754 ( .A(n16620), .ZN(n16609) );
  NAND3_X1 U18755 ( .A1(n16586), .A2(n16587), .A3(n16609), .ZN(n16588) );
  NAND2_X1 U18756 ( .A1(n16588), .A2(n16589), .ZN(n16600) );
  NAND2_X1 U18757 ( .A1(n16600), .A2(n16764), .ZN(n16599) );
  INV_X1 U18758 ( .A(n16589), .ZN(n16590) );
  NAND2_X1 U18759 ( .A1(n16586), .A2(n16590), .ZN(n16601) );
  NAND2_X1 U18760 ( .A1(n16599), .A2(n16601), .ZN(n16593) );
  XNOR2_X1 U18761 ( .A(n16591), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16592) );
  XNOR2_X1 U18762 ( .A(n16593), .B(n16592), .ZN(n16781) );
  INV_X1 U18763 ( .A(n16775), .ZN(n18760) );
  AND2_X1 U18764 ( .A1(n16675), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n16772) );
  AOI21_X1 U18765 ( .B1(n17470), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16772), .ZN(n16594) );
  OAI21_X1 U18766 ( .B1(n17479), .B2(n18754), .A(n16594), .ZN(n16597) );
  NOR2_X1 U18767 ( .A1(n16776), .A2(n17463), .ZN(n16596) );
  AOI211_X1 U18768 ( .C1(n18760), .C2(n17474), .A(n16597), .B(n16596), .ZN(
        n16598) );
  OAI21_X1 U18769 ( .B1(n17461), .B2(n16781), .A(n16598), .ZN(P2_U2986) );
  INV_X1 U18770 ( .A(n16599), .ZN(n16603) );
  AOI21_X1 U18771 ( .B1(n16600), .B2(n16601), .A(n16764), .ZN(n16602) );
  OAI22_X1 U18772 ( .A1(n16603), .A2(n16602), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16601), .ZN(n16793) );
  NAND2_X1 U18773 ( .A1(n17453), .A2(n18743), .ZN(n16604) );
  NAND2_X1 U18774 ( .A1(n16675), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n16783) );
  OAI211_X1 U18775 ( .C1(n17459), .C2(n18740), .A(n16604), .B(n16783), .ZN(
        n16607) );
  OAI21_X1 U18776 ( .B1(n16613), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16605), .ZN(n16788) );
  NOR2_X1 U18777 ( .A1(n16788), .A2(n17463), .ZN(n16606) );
  AOI211_X1 U18778 ( .C1(n18748), .C2(n17474), .A(n16607), .B(n16606), .ZN(
        n16608) );
  OAI21_X1 U18779 ( .B1(n16793), .B2(n17461), .A(n16608), .ZN(P2_U2987) );
  AOI21_X1 U18780 ( .B1(n16621), .B2(n16609), .A(n16619), .ZN(n16610) );
  XOR2_X1 U18781 ( .A(n16611), .B(n16610), .Z(n16805) );
  NAND2_X1 U18782 ( .A1(n16627), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16810) );
  AOI21_X1 U18783 ( .B1(n16799), .B2(n16810), .A(n16613), .ZN(n16802) );
  NAND2_X1 U18784 ( .A1(n16675), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16794) );
  OAI21_X1 U18785 ( .B1(n17459), .B2(n16614), .A(n16794), .ZN(n16615) );
  AOI21_X1 U18786 ( .B1(n17453), .B2(n18727), .A(n16615), .ZN(n16616) );
  OAI21_X1 U18787 ( .B1(n18738), .B2(n17449), .A(n16616), .ZN(n16617) );
  AOI21_X1 U18788 ( .B1(n16802), .B2(n17473), .A(n16617), .ZN(n16618) );
  OAI21_X1 U18789 ( .B1(n16805), .B2(n17461), .A(n16618), .ZN(P2_U2988) );
  NOR2_X1 U18790 ( .A1(n16620), .A2(n16619), .ZN(n16622) );
  XOR2_X1 U18791 ( .A(n16622), .B(n16621), .Z(n16816) );
  NAND2_X1 U18792 ( .A1(n17453), .A2(n18715), .ZN(n16624) );
  NAND2_X1 U18793 ( .A1(n16675), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16806) );
  OAI211_X1 U18794 ( .C1(n17459), .C2(n16625), .A(n16624), .B(n16806), .ZN(
        n16626) );
  AOI21_X1 U18795 ( .B1(n18720), .B2(n17474), .A(n16626), .ZN(n16629) );
  INV_X1 U18796 ( .A(n16627), .ZN(n16636) );
  NAND2_X1 U18797 ( .A1(n16636), .A2(n16798), .ZN(n16811) );
  NAND3_X1 U18798 ( .A1(n16811), .A2(n17473), .A3(n16810), .ZN(n16628) );
  OAI211_X1 U18799 ( .C1(n16816), .C2(n17461), .A(n16629), .B(n16628), .ZN(
        P2_U2989) );
  NAND2_X1 U18800 ( .A1(n16632), .A2(n16631), .ZN(n16633) );
  XNOR2_X1 U18801 ( .A(n16630), .B(n16633), .ZN(n16829) );
  NOR2_X1 U18802 ( .A1(n18848), .A2(n17565), .ZN(n16821) );
  AOI21_X1 U18803 ( .B1(n17470), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16821), .ZN(n16634) );
  OAI21_X1 U18804 ( .B1(n17479), .B2(n16635), .A(n16634), .ZN(n16638) );
  OAI21_X1 U18805 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16640), .A(
        n16636), .ZN(n16817) );
  NOR2_X1 U18806 ( .A1(n16817), .A2(n17463), .ZN(n16637) );
  AOI211_X1 U18807 ( .C1(n17474), .C2(n18707), .A(n16638), .B(n16637), .ZN(
        n16639) );
  OAI21_X1 U18808 ( .B1(n17461), .B2(n16829), .A(n16639), .ZN(P2_U2990) );
  INV_X1 U18809 ( .A(n11063), .ZN(n16656) );
  NOR2_X1 U18810 ( .A1(n16656), .A2(n16847), .ZN(n16655) );
  OAI21_X1 U18811 ( .B1(n16655), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11276), .ZN(n16840) );
  NAND2_X1 U18812 ( .A1(n17453), .A2(n18691), .ZN(n16641) );
  NAND2_X1 U18813 ( .A1(n16675), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16831) );
  OAI211_X1 U18814 ( .C1(n17459), .C2(n18688), .A(n16641), .B(n16831), .ZN(
        n16642) );
  AOI21_X1 U18815 ( .B1(n18696), .B2(n17474), .A(n16642), .ZN(n16647) );
  OAI21_X1 U18816 ( .B1(n16645), .B2(n16644), .A(n16643), .ZN(n16838) );
  NAND2_X1 U18817 ( .A1(n16838), .A2(n17475), .ZN(n16646) );
  OAI211_X1 U18818 ( .C1(n16840), .C2(n17463), .A(n16647), .B(n16646), .ZN(
        P2_U2991) );
  INV_X1 U18819 ( .A(n16648), .ZN(n16649) );
  AOI21_X1 U18820 ( .B1(n16651), .B2(n16650), .A(n16649), .ZN(n16855) );
  NOR2_X1 U18821 ( .A1(n18848), .A2(n16652), .ZN(n16845) );
  AOI21_X1 U18822 ( .B1(n17470), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16845), .ZN(n16653) );
  OAI21_X1 U18823 ( .B1(n17479), .B2(n18677), .A(n16653), .ZN(n16654) );
  AOI21_X1 U18824 ( .B1(n18683), .B2(n17474), .A(n16654), .ZN(n16658) );
  INV_X1 U18825 ( .A(n16655), .ZN(n16852) );
  NAND2_X1 U18826 ( .A1(n16656), .A2(n16847), .ZN(n16851) );
  NAND3_X1 U18827 ( .A1(n16852), .A2(n17473), .A3(n16851), .ZN(n16657) );
  OAI211_X1 U18828 ( .C1(n16855), .C2(n17461), .A(n16658), .B(n16657), .ZN(
        P2_U2992) );
  NAND3_X1 U18829 ( .A1(n16729), .A2(n16728), .A3(n16740), .ZN(n16661) );
  NAND2_X1 U18830 ( .A1(n16716), .A2(n16715), .ZN(n16939) );
  INV_X1 U18831 ( .A(n16707), .ZN(n16663) );
  INV_X1 U18832 ( .A(n16664), .ZN(n16665) );
  XNOR2_X1 U18833 ( .A(n16668), .B(n16667), .ZN(n16681) );
  AOI22_X1 U18834 ( .A1(n16681), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16669), .B2(n16668), .ZN(n16673) );
  NAND2_X1 U18835 ( .A1(n16671), .A2(n16670), .ZN(n16672) );
  XNOR2_X1 U18836 ( .A(n16673), .B(n16672), .ZN(n16866) );
  INV_X1 U18837 ( .A(n16674), .ZN(n18667) );
  INV_X1 U18838 ( .A(n18671), .ZN(n16677) );
  NAND2_X1 U18839 ( .A1(n16675), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16856) );
  NAND2_X1 U18840 ( .A1(n17470), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16676) );
  OAI211_X1 U18841 ( .C1(n17479), .C2(n16677), .A(n16856), .B(n16676), .ZN(
        n16678) );
  AOI21_X1 U18842 ( .B1(n18667), .B2(n17474), .A(n16678), .ZN(n16680) );
  NAND2_X1 U18843 ( .A1(n11052), .A2(n16873), .ZN(n16683) );
  AOI21_X1 U18844 ( .B1(n16861), .B2(n16683), .A(n11063), .ZN(n16864) );
  NAND2_X1 U18845 ( .A1(n16864), .A2(n17473), .ZN(n16679) );
  OAI211_X1 U18846 ( .C1(n16866), .C2(n17461), .A(n16680), .B(n16679), .ZN(
        P2_U2993) );
  XNOR2_X1 U18847 ( .A(n16681), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16887) );
  INV_X1 U18848 ( .A(n18661), .ZN(n16880) );
  NAND2_X1 U18849 ( .A1(n16675), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n16878) );
  NAND2_X1 U18850 ( .A1(n17470), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16682) );
  OAI211_X1 U18851 ( .C1(n17479), .C2(n18656), .A(n16878), .B(n16682), .ZN(
        n16685) );
  NAND2_X1 U18852 ( .A1(n11052), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16699) );
  NOR2_X1 U18853 ( .A1(n16699), .A2(n16888), .ZN(n16696) );
  OAI21_X1 U18854 ( .B1(n16696), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16683), .ZN(n16867) );
  NOR2_X1 U18855 ( .A1(n16867), .A2(n17463), .ZN(n16684) );
  AOI211_X1 U18856 ( .C1(n17474), .C2(n16880), .A(n16685), .B(n16684), .ZN(
        n16686) );
  OAI21_X1 U18857 ( .B1(n16887), .B2(n17461), .A(n16686), .ZN(P2_U2994) );
  NAND2_X1 U18858 ( .A1(n16688), .A2(n16687), .ZN(n16692) );
  XNOR2_X1 U18859 ( .A(n16689), .B(n16907), .ZN(n16701) );
  OAI22_X1 U18860 ( .A1(n16701), .A2(n16690), .B1(n16907), .B2(n16689), .ZN(
        n16691) );
  XOR2_X1 U18861 ( .A(n16692), .B(n16691), .Z(n16898) );
  INV_X1 U18862 ( .A(n16891), .ZN(n18650) );
  NAND2_X1 U18863 ( .A1(n17453), .A2(n18644), .ZN(n16693) );
  NAND2_X1 U18864 ( .A1(n16675), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16890) );
  OAI211_X1 U18865 ( .C1(n17459), .C2(n16694), .A(n16693), .B(n16890), .ZN(
        n16695) );
  AOI21_X1 U18866 ( .B1(n18650), .B2(n17474), .A(n16695), .ZN(n16698) );
  AOI21_X1 U18867 ( .B1(n16888), .B2(n16699), .A(n16696), .ZN(n16895) );
  NAND2_X1 U18868 ( .A1(n16895), .A2(n17473), .ZN(n16697) );
  OAI211_X1 U18869 ( .C1(n16898), .C2(n17461), .A(n16698), .B(n16697), .ZN(
        P2_U2995) );
  OAI21_X1 U18870 ( .B1(n11052), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16699), .ZN(n16911) );
  XNOR2_X1 U18871 ( .A(n16701), .B(n16700), .ZN(n16899) );
  NAND2_X1 U18872 ( .A1(n16899), .A2(n17475), .ZN(n16706) );
  NAND2_X1 U18873 ( .A1(n16328), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16904) );
  NAND2_X1 U18874 ( .A1(n17470), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16702) );
  OAI211_X1 U18875 ( .C1(n17479), .C2(n18636), .A(n16904), .B(n16702), .ZN(
        n16703) );
  AOI21_X1 U18876 ( .B1(n16704), .B2(n17474), .A(n16703), .ZN(n16705) );
  OAI211_X1 U18877 ( .C1(n17463), .C2(n16911), .A(n16706), .B(n16705), .ZN(
        P2_U2996) );
  NAND2_X1 U18878 ( .A1(n16708), .A2(n16707), .ZN(n16710) );
  XOR2_X1 U18879 ( .A(n16710), .B(n16709), .Z(n16931) );
  NAND2_X1 U18880 ( .A1(n17453), .A2(n18621), .ZN(n16711) );
  NAND2_X1 U18881 ( .A1(n16675), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16925) );
  AOI211_X1 U18882 ( .C1(n16922), .C2(n16920), .A(n17463), .B(n11052), .ZN(
        n16712) );
  AOI211_X1 U18883 ( .C1(n17474), .C2(n18628), .A(n16713), .B(n16712), .ZN(
        n16714) );
  OAI21_X1 U18884 ( .B1(n16931), .B2(n17461), .A(n16714), .ZN(P2_U2997) );
  XNOR2_X1 U18885 ( .A(n16734), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16723) );
  OR2_X1 U18886 ( .A1(n16716), .A2(n16715), .ZN(n16940) );
  NAND3_X1 U18887 ( .A1(n16940), .A2(n16939), .A3(n17475), .ZN(n16722) );
  INV_X1 U18888 ( .A(n16717), .ZN(n16938) );
  NOR2_X1 U18889 ( .A1(n18848), .A2(n17557), .ZN(n16932) );
  AOI21_X1 U18890 ( .B1(n17470), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16932), .ZN(n16718) );
  OAI21_X1 U18891 ( .B1(n17479), .B2(n16719), .A(n16718), .ZN(n16720) );
  AOI21_X1 U18892 ( .B1(n16938), .B2(n17474), .A(n16720), .ZN(n16721) );
  OAI211_X1 U18893 ( .C1(n16723), .C2(n17463), .A(n16722), .B(n16721), .ZN(
        P2_U2998) );
  INV_X1 U18894 ( .A(n16744), .ZN(n16725) );
  NOR2_X1 U18895 ( .A1(n16724), .A2(n16730), .ZN(n16742) );
  OAI21_X1 U18896 ( .B1(n16725), .B2(n16742), .A(n16740), .ZN(n16963) );
  OAI21_X1 U18897 ( .B1(n16726), .B2(n16730), .A(n16728), .ZN(n16727) );
  INV_X1 U18898 ( .A(n16727), .ZN(n16962) );
  NAND2_X1 U18899 ( .A1(n16963), .A2(n16962), .ZN(n16961) );
  NAND2_X1 U18900 ( .A1(n16961), .A2(n16728), .ZN(n16733) );
  OAI21_X1 U18901 ( .B1(n16731), .B2(n16730), .A(n16729), .ZN(n16732) );
  XNOR2_X1 U18902 ( .A(n16733), .B(n16732), .ZN(n16956) );
  AOI21_X1 U18903 ( .B1(n16913), .B2(n16959), .A(n16734), .ZN(n16954) );
  NAND2_X1 U18904 ( .A1(n16675), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16947) );
  AOI21_X1 U18905 ( .B1(n17453), .B2(n18615), .A(n16735), .ZN(n16736) );
  OAI21_X1 U18906 ( .B1(n16946), .B2(n17449), .A(n16736), .ZN(n16737) );
  AOI21_X1 U18907 ( .B1(n16954), .B2(n17473), .A(n16737), .ZN(n16738) );
  OAI21_X1 U18908 ( .B1(n16956), .B2(n17461), .A(n16738), .ZN(P2_U2999) );
  NAND2_X1 U18909 ( .A1(n17034), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17443) );
  NOR2_X2 U18910 ( .A1(n17443), .A2(n18814), .ZN(n17442) );
  NAND2_X1 U18911 ( .A1(n17442), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17014) );
  NOR2_X1 U18912 ( .A1(n17014), .A2(n17002), .ZN(n17464) );
  NAND2_X1 U18913 ( .A1(n17034), .A2(n16968), .ZN(n16958) );
  OAI21_X1 U18914 ( .B1(n17464), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16958), .ZN(n16994) );
  INV_X1 U18915 ( .A(n16740), .ZN(n16741) );
  NOR2_X1 U18916 ( .A1(n16742), .A2(n16741), .ZN(n16743) );
  XNOR2_X1 U18917 ( .A(n16744), .B(n16743), .ZN(n16992) );
  NAND2_X1 U18918 ( .A1(n16675), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16985) );
  OAI21_X1 U18919 ( .B1(n17459), .B2(n16745), .A(n16985), .ZN(n16746) );
  AOI21_X1 U18920 ( .B1(n17453), .B2(n18591), .A(n16746), .ZN(n16747) );
  OAI21_X1 U18921 ( .B1(n16980), .B2(n17449), .A(n16747), .ZN(n16748) );
  AOI21_X1 U18922 ( .B1(n16992), .B2(n17475), .A(n16748), .ZN(n16749) );
  OAI21_X1 U18923 ( .B1(n16994), .B2(n17463), .A(n16749), .ZN(P2_U3001) );
  INV_X1 U18924 ( .A(n18797), .ZN(n16758) );
  AOI21_X1 U18925 ( .B1(n16751), .B2(n18852), .A(n16750), .ZN(n16755) );
  INV_X1 U18926 ( .A(n16766), .ZN(n16787) );
  NAND3_X1 U18927 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16752) );
  AOI21_X1 U18928 ( .B1(n16753), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11466), .ZN(n16754) );
  OAI21_X1 U18929 ( .B1(n16760), .B2(n18869), .A(n16759), .ZN(P2_U3016) );
  NOR3_X1 U18930 ( .A1(n16787), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16762), .ZN(n16763) );
  OAI21_X1 U18931 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17047), .A(
        n16782), .ZN(n16779) );
  NOR2_X1 U18932 ( .A1(n16764), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16765) );
  NAND2_X1 U18933 ( .A1(n16766), .A2(n16765), .ZN(n16774) );
  INV_X1 U18934 ( .A(n16774), .ZN(n16767) );
  OAI21_X1 U18935 ( .B1(n16779), .B2(n16767), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16768) );
  OAI21_X1 U18936 ( .B1(n16771), .B2(n18869), .A(n16770), .ZN(P2_U3017) );
  AOI21_X1 U18937 ( .B1(n18759), .B2(n18852), .A(n16772), .ZN(n16773) );
  OAI211_X1 U18938 ( .C1(n16775), .C2(n18849), .A(n16774), .B(n16773), .ZN(
        n16778) );
  NOR2_X1 U18939 ( .A1(n16776), .A2(n18881), .ZN(n16777) );
  AOI211_X1 U18940 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16779), .A(
        n16778), .B(n16777), .ZN(n16780) );
  OAI21_X1 U18941 ( .B1(n18869), .B2(n16781), .A(n16780), .ZN(P2_U3018) );
  INV_X1 U18942 ( .A(n16782), .ZN(n16791) );
  INV_X1 U18943 ( .A(n18747), .ZN(n16784) );
  OAI21_X1 U18944 ( .B1(n16784), .B2(n18870), .A(n16783), .ZN(n16785) );
  AOI21_X1 U18945 ( .B1(n18748), .B2(n14189), .A(n16785), .ZN(n16786) );
  OAI21_X1 U18946 ( .B1(n16787), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16786), .ZN(n16790) );
  NOR2_X1 U18947 ( .A1(n16788), .A2(n18881), .ZN(n16789) );
  AOI211_X1 U18948 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16791), .A(
        n16790), .B(n16789), .ZN(n16792) );
  OAI21_X1 U18949 ( .B1(n16793), .B2(n18869), .A(n16792), .ZN(P2_U3019) );
  INV_X1 U18950 ( .A(n16794), .ZN(n16795) );
  AOI21_X1 U18951 ( .B1(n18733), .B2(n18852), .A(n16795), .ZN(n16796) );
  OAI21_X1 U18952 ( .B1(n18738), .B2(n18849), .A(n16796), .ZN(n16801) );
  AOI211_X1 U18953 ( .C1(n16799), .C2(n16798), .A(n16797), .B(n16809), .ZN(
        n16800) );
  AOI211_X1 U18954 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n16814), .A(
        n16801), .B(n16800), .ZN(n16804) );
  NAND2_X1 U18955 ( .A1(n16802), .A2(n18825), .ZN(n16803) );
  OAI211_X1 U18956 ( .C1(n16805), .C2(n18869), .A(n16804), .B(n16803), .ZN(
        P2_U3020) );
  OAI21_X1 U18957 ( .B1(n18724), .B2(n18870), .A(n16806), .ZN(n16807) );
  AOI21_X1 U18958 ( .B1(n18720), .B2(n14189), .A(n16807), .ZN(n16808) );
  OAI21_X1 U18959 ( .B1(n16809), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16808), .ZN(n16813) );
  AND3_X1 U18960 ( .A1(n16811), .A2(n18825), .A3(n16810), .ZN(n16812) );
  AOI211_X1 U18961 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n16814), .A(
        n16813), .B(n16812), .ZN(n16815) );
  OAI21_X1 U18962 ( .B1(n18869), .B2(n16816), .A(n16815), .ZN(P2_U3021) );
  INV_X1 U18963 ( .A(n16817), .ZN(n16827) );
  NOR2_X1 U18964 ( .A1(n16819), .A2(n16818), .ZN(n16820) );
  AOI211_X1 U18965 ( .C1(n18852), .C2(n16822), .A(n16821), .B(n16820), .ZN(
        n16823) );
  OAI211_X1 U18966 ( .C1(n18849), .C2(n16825), .A(n16824), .B(n16823), .ZN(
        n16826) );
  AOI21_X1 U18967 ( .B1(n16827), .B2(n18825), .A(n16826), .ZN(n16828) );
  OAI21_X1 U18968 ( .B1(n18869), .B2(n16829), .A(n16828), .ZN(P2_U3022) );
  OAI21_X1 U18969 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16830), .ZN(n16836) );
  NAND2_X1 U18970 ( .A1(n18695), .A2(n18852), .ZN(n16832) );
  OAI211_X1 U18971 ( .C1(n16862), .C2(n16833), .A(n16832), .B(n16831), .ZN(
        n16834) );
  AOI21_X1 U18972 ( .B1(n18696), .B2(n14189), .A(n16834), .ZN(n16835) );
  OAI21_X1 U18973 ( .B1(n16848), .B2(n16836), .A(n16835), .ZN(n16837) );
  AOI21_X1 U18974 ( .B1(n16838), .B2(n18856), .A(n16837), .ZN(n16839) );
  OAI21_X1 U18975 ( .B1(n16840), .B2(n18881), .A(n16839), .ZN(P2_U3023) );
  NAND2_X1 U18976 ( .A1(n16842), .A2(n16841), .ZN(n16843) );
  AND2_X1 U18977 ( .A1(n16844), .A2(n16843), .ZN(n19547) );
  AOI21_X1 U18978 ( .B1(n19547), .B2(n18852), .A(n16845), .ZN(n16846) );
  OAI21_X1 U18979 ( .B1(n16862), .B2(n16847), .A(n16846), .ZN(n16850) );
  NOR2_X1 U18980 ( .A1(n16848), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16849) );
  AOI211_X1 U18981 ( .C1(n18683), .C2(n14189), .A(n16850), .B(n16849), .ZN(
        n16854) );
  NAND3_X1 U18982 ( .A1(n16852), .A2(n18825), .A3(n16851), .ZN(n16853) );
  OAI211_X1 U18983 ( .C1(n16855), .C2(n18869), .A(n16854), .B(n16853), .ZN(
        P2_U3024) );
  NAND3_X1 U18984 ( .A1(n16908), .A2(n16873), .A3(n16861), .ZN(n16860) );
  OAI21_X1 U18985 ( .B1(n16857), .B2(n18870), .A(n16856), .ZN(n16858) );
  AOI21_X1 U18986 ( .B1(n18667), .B2(n14189), .A(n16858), .ZN(n16859) );
  OAI211_X1 U18987 ( .C1(n16862), .C2(n16861), .A(n16860), .B(n16859), .ZN(
        n16863) );
  AOI21_X1 U18988 ( .B1(n16864), .B2(n18825), .A(n16863), .ZN(n16865) );
  OAI21_X1 U18989 ( .B1(n16866), .B2(n18869), .A(n16865), .ZN(P2_U3025) );
  INV_X1 U18990 ( .A(n16867), .ZN(n16885) );
  NAND2_X1 U18991 ( .A1(n16921), .A2(n16868), .ZN(n16914) );
  NOR2_X1 U18992 ( .A1(n16912), .A2(n16921), .ZN(n16869) );
  OR2_X1 U18993 ( .A1(n16870), .A2(n16869), .ZN(n16915) );
  NOR2_X1 U18994 ( .A1(n17047), .A2(n11476), .ZN(n16871) );
  AOI211_X1 U18995 ( .C1(n16872), .C2(n16914), .A(n16915), .B(n16871), .ZN(
        n16900) );
  INV_X1 U18996 ( .A(n16873), .ZN(n16874) );
  OAI211_X1 U18997 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n16875), .A(
        n16908), .B(n16874), .ZN(n16882) );
  OAI21_X1 U18998 ( .B1(n16877), .B2(n16876), .A(n16538), .ZN(n18657) );
  OAI21_X1 U18999 ( .B1(n18657), .B2(n18870), .A(n16878), .ZN(n16879) );
  AOI21_X1 U19000 ( .B1(n16880), .B2(n14189), .A(n16879), .ZN(n16881) );
  OAI211_X1 U19001 ( .C1(n16900), .C2(n16883), .A(n16882), .B(n16881), .ZN(
        n16884) );
  AOI21_X1 U19002 ( .B1(n16885), .B2(n18825), .A(n16884), .ZN(n16886) );
  OAI21_X1 U19003 ( .B1(n16887), .B2(n18869), .A(n16886), .ZN(P2_U3026) );
  XNOR2_X1 U19004 ( .A(n16888), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16894) );
  NOR2_X1 U19005 ( .A1(n16900), .A2(n16888), .ZN(n16893) );
  NAND2_X1 U19006 ( .A1(n18852), .A2(n18649), .ZN(n16889) );
  OAI211_X1 U19007 ( .C1(n16891), .C2(n18849), .A(n16890), .B(n16889), .ZN(
        n16892) );
  AOI211_X1 U19008 ( .C1(n16908), .C2(n16894), .A(n16893), .B(n16892), .ZN(
        n16897) );
  NAND2_X1 U19009 ( .A1(n16895), .A2(n18825), .ZN(n16896) );
  OAI211_X1 U19010 ( .C1(n16898), .C2(n18869), .A(n16897), .B(n16896), .ZN(
        P2_U3027) );
  NAND2_X1 U19011 ( .A1(n16899), .A2(n18856), .ZN(n16910) );
  NOR2_X1 U19012 ( .A1(n16900), .A2(n16907), .ZN(n16906) );
  AOI21_X1 U19013 ( .B1(n16902), .B2(n11091), .A(n11374), .ZN(n19766) );
  NAND2_X1 U19014 ( .A1(n18852), .A2(n19766), .ZN(n16903) );
  OAI211_X1 U19015 ( .C1(n18641), .C2(n18849), .A(n16904), .B(n16903), .ZN(
        n16905) );
  AOI211_X1 U19016 ( .C1(n16908), .C2(n16907), .A(n16906), .B(n16905), .ZN(
        n16909) );
  OAI211_X1 U19017 ( .C1(n16911), .C2(n18881), .A(n16910), .B(n16909), .ZN(
        P2_U3028) );
  NAND2_X1 U19018 ( .A1(n18881), .A2(n16912), .ZN(n16919) );
  NOR2_X1 U19019 ( .A1(n16914), .A2(n16913), .ZN(n16918) );
  INV_X1 U19020 ( .A(n16915), .ZN(n16916) );
  OAI21_X1 U19021 ( .B1(n16918), .B2(n16917), .A(n16916), .ZN(n16950) );
  AOI21_X1 U19022 ( .B1(n16920), .B2(n16919), .A(n16950), .ZN(n16944) );
  OAI21_X1 U19023 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17047), .A(
        n16944), .ZN(n16929) );
  INV_X1 U19024 ( .A(n17037), .ZN(n16965) );
  NAND2_X1 U19025 ( .A1(n16965), .A2(n16921), .ZN(n16952) );
  OAI21_X1 U19026 ( .B1(n16959), .B2(n18881), .A(n16952), .ZN(n16935) );
  AND3_X1 U19027 ( .A1(n16935), .A2(n16923), .A3(n16922), .ZN(n16928) );
  NAND2_X1 U19028 ( .A1(n18852), .A2(n18627), .ZN(n16924) );
  OAI211_X1 U19029 ( .C1(n16926), .C2(n18849), .A(n16925), .B(n16924), .ZN(
        n16927) );
  AOI211_X1 U19030 ( .C1(n16929), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16928), .B(n16927), .ZN(n16930) );
  OAI21_X1 U19031 ( .B1(n16931), .B2(n18869), .A(n16930), .ZN(P2_U3029) );
  INV_X1 U19032 ( .A(n16932), .ZN(n16933) );
  OAI21_X1 U19033 ( .B1(n18870), .B2(n16934), .A(n16933), .ZN(n16937) );
  AND3_X1 U19034 ( .A1(n16935), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16943), .ZN(n16936) );
  AOI211_X1 U19035 ( .C1(n16938), .C2(n14189), .A(n16937), .B(n16936), .ZN(
        n16942) );
  NAND3_X1 U19036 ( .A1(n16940), .A2(n16939), .A3(n18856), .ZN(n16941) );
  OAI211_X1 U19037 ( .C1(n16944), .C2(n16943), .A(n16942), .B(n16941), .ZN(
        P2_U3030) );
  XNOR2_X1 U19038 ( .A(n11039), .B(n16945), .ZN(n19369) );
  INV_X1 U19039 ( .A(n16946), .ZN(n18616) );
  NAND2_X1 U19040 ( .A1(n18616), .A2(n14189), .ZN(n16948) );
  OAI211_X1 U19041 ( .C1(n19369), .C2(n18870), .A(n16948), .B(n16947), .ZN(
        n16949) );
  AOI21_X1 U19042 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16950), .A(
        n16949), .ZN(n16951) );
  OAI21_X1 U19043 ( .B1(n16952), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16951), .ZN(n16953) );
  AOI21_X1 U19044 ( .B1(n16954), .B2(n18825), .A(n16953), .ZN(n16955) );
  OAI21_X1 U19045 ( .B1(n16956), .B2(n18869), .A(n16955), .ZN(P2_U3031) );
  NAND2_X1 U19046 ( .A1(n16958), .A2(n16957), .ZN(n16960) );
  AND2_X1 U19047 ( .A1(n16960), .A2(n16959), .ZN(n17472) );
  INV_X1 U19048 ( .A(n17472), .ZN(n16979) );
  OAI21_X1 U19049 ( .B1(n16963), .B2(n16962), .A(n16961), .ZN(n17476) );
  NAND2_X1 U19050 ( .A1(n17476), .A2(n18856), .ZN(n16978) );
  INV_X1 U19051 ( .A(n16967), .ZN(n16964) );
  NAND2_X1 U19052 ( .A1(n16965), .A2(n16964), .ZN(n17001) );
  NOR2_X1 U19053 ( .A1(n17001), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16966) );
  AOI211_X1 U19054 ( .C1(n16967), .C2(n18808), .A(n17043), .B(n16966), .ZN(
        n17000) );
  OAI21_X1 U19055 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17001), .A(
        n17000), .ZN(n16976) );
  INV_X1 U19056 ( .A(n16968), .ZN(n16969) );
  NOR3_X1 U19057 ( .A1(n17037), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16969), .ZN(n16975) );
  NAND2_X1 U19058 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n16328), .ZN(n16973) );
  NAND2_X1 U19059 ( .A1(n16984), .A2(n16970), .ZN(n16971) );
  AND2_X1 U19060 ( .A1(n11039), .A2(n16971), .ZN(n19370) );
  NAND2_X1 U19061 ( .A1(n18852), .A2(n19370), .ZN(n16972) );
  OAI211_X1 U19062 ( .C1(n17471), .C2(n18849), .A(n16973), .B(n16972), .ZN(
        n16974) );
  AOI211_X1 U19063 ( .C1(n16976), .C2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16975), .B(n16974), .ZN(n16977) );
  OAI211_X1 U19064 ( .C1(n16979), .C2(n18881), .A(n16978), .B(n16977), .ZN(
        P2_U3032) );
  INV_X1 U19065 ( .A(n16980), .ZN(n18592) );
  OR2_X1 U19066 ( .A1(n16982), .A2(n16981), .ZN(n16983) );
  NAND2_X1 U19067 ( .A1(n16984), .A2(n16983), .ZN(n19376) );
  OAI21_X1 U19068 ( .B1(n18870), .B2(n19376), .A(n16985), .ZN(n16986) );
  AOI21_X1 U19069 ( .B1(n18592), .B2(n14189), .A(n16986), .ZN(n16989) );
  INV_X1 U19070 ( .A(n17001), .ZN(n16987) );
  NAND3_X1 U19071 ( .A1(n16987), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n16990), .ZN(n16988) );
  OAI211_X1 U19072 ( .C1(n17000), .C2(n16990), .A(n16989), .B(n16988), .ZN(
        n16991) );
  AOI21_X1 U19073 ( .B1(n16992), .B2(n18856), .A(n16991), .ZN(n16993) );
  OAI21_X1 U19074 ( .B1(n16994), .B2(n18881), .A(n16993), .ZN(P2_U3033) );
  XNOR2_X1 U19075 ( .A(n16995), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16996) );
  XNOR2_X1 U19076 ( .A(n16659), .B(n16996), .ZN(n17462) );
  INV_X1 U19077 ( .A(n17014), .ZN(n16997) );
  NOR2_X1 U19078 ( .A1(n16997), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17465) );
  OR3_X1 U19079 ( .A1(n17465), .A2(n17464), .A3(n18881), .ZN(n17006) );
  AOI21_X1 U19080 ( .B1(n16999), .B2(n16998), .A(n16981), .ZN(n18579) );
  INV_X1 U19081 ( .A(n18579), .ZN(n19379) );
  OAI22_X1 U19082 ( .A1(n18870), .A2(n19379), .B1(n13071), .B2(n18848), .ZN(
        n17004) );
  AOI21_X1 U19083 ( .B1(n17002), .B2(n17001), .A(n17000), .ZN(n17003) );
  AOI211_X1 U19084 ( .C1(n18580), .C2(n14189), .A(n17004), .B(n17003), .ZN(
        n17005) );
  OAI211_X1 U19085 ( .C1(n17462), .C2(n18869), .A(n17006), .B(n17005), .ZN(
        P2_U3034) );
  NAND2_X1 U19086 ( .A1(n17008), .A2(n17007), .ZN(n17013) );
  INV_X1 U19087 ( .A(n17009), .ZN(n17011) );
  AND2_X1 U19088 ( .A1(n17011), .A2(n17010), .ZN(n17012) );
  XNOR2_X1 U19089 ( .A(n17013), .B(n17012), .ZN(n17454) );
  OAI21_X1 U19090 ( .B1(n17442), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17014), .ZN(n17455) );
  OR2_X1 U19091 ( .A1(n17455), .A2(n18881), .ZN(n17027) );
  AOI21_X1 U19092 ( .B1(n17020), .B2(n18808), .A(n17043), .ZN(n18815) );
  NOR2_X1 U19093 ( .A1(n17020), .A2(n17037), .ZN(n17015) );
  NAND2_X1 U19094 ( .A1(n17015), .A2(n18814), .ZN(n18813) );
  INV_X1 U19095 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17016) );
  AOI21_X1 U19096 ( .B1(n18815), .B2(n18813), .A(n17016), .ZN(n17025) );
  OR2_X1 U19097 ( .A1(n17018), .A2(n17017), .ZN(n17019) );
  NAND2_X1 U19098 ( .A1(n17019), .A2(n16998), .ZN(n19382) );
  NAND2_X1 U19099 ( .A1(n14189), .A2(n18570), .ZN(n17023) );
  NOR4_X1 U19100 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18814), .A3(
        n17020), .A4(n17037), .ZN(n17021) );
  AOI21_X1 U19101 ( .B1(n16328), .B2(P2_REIP_REG_11__SCAN_IN), .A(n17021), 
        .ZN(n17022) );
  OAI211_X1 U19102 ( .C1(n19382), .C2(n18870), .A(n17023), .B(n17022), .ZN(
        n17024) );
  NOR2_X1 U19103 ( .A1(n17025), .A2(n17024), .ZN(n17026) );
  OAI211_X1 U19104 ( .C1(n17454), .C2(n18869), .A(n17027), .B(n17026), .ZN(
        P2_U3035) );
  NAND2_X1 U19105 ( .A1(n17028), .A2(n17029), .ZN(n17033) );
  INV_X1 U19106 ( .A(n17029), .ZN(n17444) );
  OAI21_X1 U19107 ( .B1(n17031), .B2(n17444), .A(n17030), .ZN(n17032) );
  NAND2_X1 U19108 ( .A1(n17033), .A2(n17032), .ZN(n17436) );
  OAI21_X1 U19109 ( .B1(n17034), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17443), .ZN(n17437) );
  OR2_X1 U19110 ( .A1(n17437), .A2(n18881), .ZN(n17045) );
  OR2_X1 U19111 ( .A1(n17035), .A2(n18530), .ZN(n17036) );
  NAND2_X1 U19112 ( .A1(n17036), .A2(n18555), .ZN(n19389) );
  NAND2_X1 U19113 ( .A1(n14189), .A2(n18544), .ZN(n17041) );
  NOR2_X1 U19114 ( .A1(n13061), .A2(n18848), .ZN(n17039) );
  NOR2_X1 U19115 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17037), .ZN(
        n17038) );
  NOR2_X1 U19116 ( .A1(n17039), .A2(n17038), .ZN(n17040) );
  OAI211_X1 U19117 ( .C1(n19389), .C2(n18870), .A(n17041), .B(n17040), .ZN(
        n17042) );
  AOI21_X1 U19118 ( .B1(n17043), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17042), .ZN(n17044) );
  OAI211_X1 U19119 ( .C1(n17436), .C2(n18869), .A(n17045), .B(n17044), .ZN(
        P2_U3037) );
  NOR2_X1 U19120 ( .A1(n17046), .A2(n18869), .ZN(n17050) );
  AOI211_X1 U19121 ( .C1(n17065), .C2(n17048), .A(n18864), .B(n17047), .ZN(
        n17049) );
  AOI211_X1 U19122 ( .C1(n18825), .C2(n17051), .A(n17050), .B(n17049), .ZN(
        n17056) );
  AOI22_X1 U19123 ( .A1(n18470), .A2(n14189), .B1(n18852), .B2(n19809), .ZN(
        n17055) );
  NAND2_X1 U19124 ( .A1(n17052), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17053) );
  NAND4_X1 U19125 ( .A1(n17056), .A2(n17055), .A3(n17054), .A4(n17053), .ZN(
        P2_U3045) );
  INV_X1 U19126 ( .A(n17071), .ZN(n17060) );
  OAI21_X1 U19127 ( .B1(n17057), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n18890), 
        .ZN(n17059) );
  AOI22_X1 U19128 ( .A1(n17060), .A2(n17059), .B1(n17058), .B2(n18897), .ZN(
        n17062) );
  NAND2_X1 U19129 ( .A1(n17073), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17061) );
  OAI21_X1 U19130 ( .B1(n17062), .B2(n17073), .A(n17061), .ZN(P2_U3601) );
  OAI21_X1 U19131 ( .B1(n18462), .B2(n17064), .A(n17063), .ZN(n18476) );
  OAI21_X1 U19132 ( .B1(n11029), .B2(n17065), .A(n18476), .ZN(n17070) );
  INV_X1 U19133 ( .A(n17070), .ZN(n17066) );
  AOI222_X1 U19134 ( .A1(n17067), .A2(n17387), .B1(n17066), .B2(n17071), .C1(
        n18471), .C2(n18897), .ZN(n17069) );
  NAND2_X1 U19135 ( .A1(n17073), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17068) );
  OAI21_X1 U19136 ( .B1(n17069), .B2(n17073), .A(n17068), .ZN(P2_U3600) );
  AOI222_X1 U19137 ( .A1(n17072), .A2(n17387), .B1(n17071), .B2(n17070), .C1(
        n18897), .C2(n17488), .ZN(n17074) );
  MUX2_X1 U19138 ( .A(n17074), .B(n11409), .S(n17073), .Z(n17075) );
  INV_X1 U19139 ( .A(n17075), .ZN(P2_U3599) );
  NOR2_X1 U19140 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17076), .ZN(
        n18955) );
  INV_X1 U19141 ( .A(n18356), .ZN(n17089) );
  OAI211_X1 U19142 ( .C1(n17076), .C2(n18353), .A(n21398), .B(n17089), .ZN(
        n17078) );
  NAND2_X1 U19143 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18939) );
  INV_X1 U19144 ( .A(n18306), .ZN(n18254) );
  OAI21_X1 U19145 ( .B1(n17972), .B2(n18254), .A(n21426), .ZN(n17077) );
  AOI211_X1 U19146 ( .C1(n18939), .C2(n17077), .A(n18356), .B(n18942), .ZN(
        n18354) );
  OAI22_X1 U19147 ( .A1(n18955), .A2(n17078), .B1(n18354), .B2(n21398), .ZN(
        P3_U2865) );
  INV_X1 U19148 ( .A(n21670), .ZN(n17082) );
  INV_X1 U19149 ( .A(n12287), .ZN(n17080) );
  NAND4_X1 U19150 ( .A1(n17082), .A2(n17081), .A3(n17080), .A4(n17079), .ZN(
        n17083) );
  OAI21_X1 U19151 ( .B1(n21829), .B2(n17084), .A(n17083), .ZN(P1_U3468) );
  INV_X1 U19152 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17085) );
  OAI21_X1 U19153 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n21862), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18418) );
  NAND2_X1 U19154 ( .A1(n11798), .A2(n18418), .ZN(n17087) );
  INV_X1 U19155 ( .A(n17087), .ZN(n21858) );
  INV_X1 U19156 ( .A(BS16), .ZN(n17228) );
  INV_X1 U19157 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21909) );
  NAND2_X1 U19158 ( .A1(n21909), .A2(n21862), .ZN(n21860) );
  AOI21_X1 U19159 ( .B1(n17228), .B2(n21860), .A(n17086), .ZN(n21854) );
  AOI21_X1 U19160 ( .B1(n17085), .B2(n17086), .A(n21854), .ZN(P3_U3280) );
  AND2_X1 U19161 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17086), .ZN(P3_U3028) );
  AND2_X1 U19162 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17086), .ZN(P3_U3027) );
  AND2_X1 U19163 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17086), .ZN(P3_U3026) );
  AND2_X1 U19164 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17086), .ZN(P3_U3025) );
  AND2_X1 U19165 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17086), .ZN(P3_U3024) );
  AND2_X1 U19166 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17086), .ZN(P3_U3023) );
  AND2_X1 U19167 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17086), .ZN(P3_U3022) );
  AND2_X1 U19168 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17086), .ZN(P3_U3021) );
  AND2_X1 U19169 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17086), .ZN(
        P3_U3020) );
  AND2_X1 U19170 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17086), .ZN(
        P3_U3019) );
  AND2_X1 U19171 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17086), .ZN(
        P3_U3018) );
  AND2_X1 U19172 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17086), .ZN(
        P3_U3017) );
  AND2_X1 U19173 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17086), .ZN(
        P3_U3016) );
  AND2_X1 U19174 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17087), .ZN(
        P3_U3015) );
  AND2_X1 U19175 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17087), .ZN(
        P3_U3014) );
  AND2_X1 U19176 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17087), .ZN(
        P3_U3013) );
  AND2_X1 U19177 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17087), .ZN(
        P3_U3012) );
  AND2_X1 U19178 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17087), .ZN(
        P3_U3011) );
  AND2_X1 U19179 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17087), .ZN(
        P3_U3010) );
  AND2_X1 U19180 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17087), .ZN(
        P3_U3009) );
  AND2_X1 U19181 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17087), .ZN(
        P3_U3008) );
  AND2_X1 U19182 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17087), .ZN(
        P3_U3007) );
  AND2_X1 U19183 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17087), .ZN(
        P3_U3006) );
  AND2_X1 U19184 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17087), .ZN(
        P3_U3005) );
  AND2_X1 U19185 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17087), .ZN(
        P3_U3004) );
  AND2_X1 U19186 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17087), .ZN(
        P3_U3003) );
  AND2_X1 U19187 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17087), .ZN(
        P3_U3002) );
  AND2_X1 U19188 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17086), .ZN(
        P3_U3001) );
  AND2_X1 U19189 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17086), .ZN(
        P3_U3000) );
  AND2_X1 U19190 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17087), .ZN(
        P3_U2999) );
  AOI21_X1 U19191 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17088)
         );
  NOR4_X1 U19192 ( .A1(n18347), .A2(n21438), .A3(n21907), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21378) );
  AOI211_X1 U19193 ( .C1(n18306), .C2(n17088), .A(n21424), .B(n21378), .ZN(
        P3_U2998) );
  NOR2_X1 U19194 ( .A1(n17090), .A2(n17089), .ZN(P3_U2867) );
  NAND2_X1 U19195 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18086), .ZN(n20317) );
  INV_X2 U19196 ( .A(n20317), .ZN(n18415) );
  NOR2_X4 U19197 ( .A1(n18415), .A2(n18399), .ZN(n18410) );
  AND2_X1 U19198 ( .A1(n18410), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U19199 ( .A(n20369), .ZN(n20316) );
  OAI21_X1 U19200 ( .B1(n17969), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n20316), 
        .ZN(n17093) );
  OAI21_X1 U19201 ( .B1(n20314), .B2(n20316), .A(n17093), .ZN(P3_U3298) );
  NOR2_X1 U19202 ( .A1(n17969), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n17095)
         );
  OAI21_X1 U19203 ( .B1(n20369), .B2(n17095), .A(n17094), .ZN(P3_U3299) );
  INV_X1 U19204 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n17096) );
  NOR2_X1 U19205 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17096), .ZN(n21889) );
  AOI21_X1 U19206 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21889), .A(n17541), 
        .ZN(n17097) );
  INV_X1 U19207 ( .A(n17097), .ZN(n21853) );
  INV_X1 U19208 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17113) );
  INV_X1 U19209 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21890) );
  NAND2_X1 U19210 ( .A1(n21890), .A2(n17096), .ZN(n21885) );
  AOI21_X1 U19211 ( .B1(n17228), .B2(n21885), .A(n17098), .ZN(n21850) );
  AOI21_X1 U19212 ( .B1(n17098), .B2(n17113), .A(n21850), .ZN(P2_U3591) );
  AND2_X1 U19213 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17098), .ZN(P2_U3208) );
  AND2_X1 U19214 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17098), .ZN(P2_U3207) );
  AND2_X1 U19215 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17098), .ZN(P2_U3206) );
  AND2_X1 U19216 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17098), .ZN(P2_U3205) );
  AND2_X1 U19217 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17098), .ZN(P2_U3204) );
  AND2_X1 U19218 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17098), .ZN(P2_U3203) );
  AND2_X1 U19219 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17098), .ZN(P2_U3202) );
  AND2_X1 U19220 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17098), .ZN(P2_U3201) );
  AND2_X1 U19221 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17098), .ZN(
        P2_U3200) );
  AND2_X1 U19222 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17098), .ZN(
        P2_U3199) );
  AND2_X1 U19223 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17098), .ZN(
        P2_U3198) );
  AND2_X1 U19224 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17098), .ZN(
        P2_U3197) );
  AND2_X1 U19225 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17098), .ZN(
        P2_U3196) );
  AND2_X1 U19226 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17098), .ZN(
        P2_U3195) );
  AND2_X1 U19227 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17098), .ZN(
        P2_U3194) );
  AND2_X1 U19228 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17097), .ZN(
        P2_U3193) );
  AND2_X1 U19229 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17097), .ZN(
        P2_U3192) );
  AND2_X1 U19230 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17097), .ZN(
        P2_U3191) );
  AND2_X1 U19231 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17097), .ZN(
        P2_U3190) );
  AND2_X1 U19232 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17097), .ZN(
        P2_U3189) );
  AND2_X1 U19233 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17097), .ZN(
        P2_U3188) );
  AND2_X1 U19234 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17097), .ZN(
        P2_U3187) );
  AND2_X1 U19235 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17097), .ZN(
        P2_U3186) );
  AND2_X1 U19236 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17097), .ZN(
        P2_U3185) );
  AND2_X1 U19237 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17097), .ZN(
        P2_U3184) );
  AND2_X1 U19238 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17097), .ZN(
        P2_U3183) );
  AND2_X1 U19239 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17097), .ZN(
        P2_U3182) );
  AND2_X1 U19240 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17098), .ZN(
        P2_U3181) );
  AND2_X1 U19241 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17098), .ZN(
        P2_U3180) );
  AND2_X1 U19242 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17098), .ZN(
        P2_U3179) );
  OAI221_X1 U19243 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(
        P2_STATEBS16_REG_SCAN_IN), .C1(n14841), .C2(n18899), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n17100) );
  AOI21_X1 U19244 ( .B1(n17100), .B2(n19473), .A(n17099), .ZN(P2_U3178) );
  OAI221_X1 U19245 ( .B1(n18912), .B2(n18893), .C1(n17101), .C2(n18893), .A(
        n19869), .ZN(n17497) );
  NOR2_X1 U19246 ( .A1(n17102), .A2(n17497), .ZN(P2_U3047) );
  AND2_X1 U19247 ( .A1(n17529), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19248 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17106) );
  NOR4_X1 U19249 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17105) );
  NOR4_X1 U19250 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17104) );
  NOR4_X1 U19251 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17103) );
  NAND4_X1 U19252 ( .A1(n17106), .A2(n17105), .A3(n17104), .A4(n17103), .ZN(
        n17112) );
  NOR4_X1 U19253 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17110) );
  AOI211_X1 U19254 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17109) );
  NOR4_X1 U19255 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17108) );
  NOR4_X1 U19256 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17107) );
  NAND4_X1 U19257 ( .A1(n17110), .A2(n17109), .A3(n17108), .A4(n17107), .ZN(
        n17111) );
  NOR2_X1 U19258 ( .A1(n17112), .A2(n17111), .ZN(n17508) );
  INV_X1 U19259 ( .A(n17508), .ZN(n17506) );
  NOR2_X1 U19260 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17506), .ZN(n17500) );
  INV_X1 U19261 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21852) );
  NAND3_X1 U19262 ( .A1(n17501), .A2(n21852), .A3(n17113), .ZN(n17505) );
  INV_X1 U19263 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U19264 ( .A1(n17500), .A2(n17505), .B1(n17506), .B2(n17114), .ZN(
        P2_U2821) );
  INV_X1 U19265 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U19266 ( .A1(n17500), .A2(n17501), .B1(n17506), .B2(n17115), .ZN(
        P2_U2820) );
  INV_X1 U19267 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17116) );
  INV_X1 U19268 ( .A(n21865), .ZN(n17157) );
  INV_X1 U19269 ( .A(n22398), .ZN(n20100) );
  CLKBUF_X1 U19270 ( .A(n20100), .Z(n22395) );
  OAI21_X1 U19271 ( .B1(n17157), .B2(n12216), .A(n22395), .ZN(n17117) );
  NAND2_X1 U19272 ( .A1(n21873), .A2(n12216), .ZN(n20242) );
  AOI21_X1 U19273 ( .B1(n17228), .B2(n20242), .A(n21848), .ZN(n21847) );
  AOI21_X1 U19274 ( .B1(n17116), .B2(n21848), .A(n21847), .ZN(P1_U3464) );
  AND2_X1 U19275 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21848), .ZN(P1_U3193) );
  AND2_X1 U19276 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21848), .ZN(P1_U3192) );
  AND2_X1 U19277 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21848), .ZN(P1_U3191) );
  AND2_X1 U19278 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n17117), .ZN(P1_U3190) );
  AND2_X1 U19279 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n17117), .ZN(P1_U3189) );
  AND2_X1 U19280 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n17117), .ZN(P1_U3188) );
  AND2_X1 U19281 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n17117), .ZN(P1_U3187) );
  AND2_X1 U19282 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n17117), .ZN(P1_U3186) );
  AND2_X1 U19283 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n17117), .ZN(
        P1_U3185) );
  AND2_X1 U19284 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n17117), .ZN(
        P1_U3184) );
  AND2_X1 U19285 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n17117), .ZN(
        P1_U3183) );
  AND2_X1 U19286 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n17117), .ZN(
        P1_U3182) );
  AND2_X1 U19287 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n17117), .ZN(
        P1_U3181) );
  AND2_X1 U19288 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n17117), .ZN(
        P1_U3180) );
  AND2_X1 U19289 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n17117), .ZN(
        P1_U3179) );
  AND2_X1 U19290 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n17117), .ZN(
        P1_U3178) );
  AND2_X1 U19291 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21848), .ZN(
        P1_U3177) );
  AND2_X1 U19292 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21848), .ZN(
        P1_U3176) );
  AND2_X1 U19293 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21848), .ZN(
        P1_U3175) );
  AND2_X1 U19294 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21848), .ZN(
        P1_U3174) );
  AND2_X1 U19295 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21848), .ZN(
        P1_U3173) );
  AND2_X1 U19296 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21848), .ZN(
        P1_U3172) );
  AND2_X1 U19297 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21848), .ZN(
        P1_U3171) );
  AND2_X1 U19298 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n17117), .ZN(
        P1_U3170) );
  AND2_X1 U19299 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21848), .ZN(
        P1_U3169) );
  AND2_X1 U19300 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21848), .ZN(
        P1_U3168) );
  AND2_X1 U19301 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21848), .ZN(
        P1_U3167) );
  AND2_X1 U19302 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21848), .ZN(
        P1_U3166) );
  AND2_X1 U19303 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21848), .ZN(
        P1_U3165) );
  AND2_X1 U19304 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21848), .ZN(
        P1_U3164) );
  INV_X1 U19305 ( .A(n17128), .ZN(n17126) );
  AOI21_X1 U19306 ( .B1(n17118), .B2(n11008), .A(n22029), .ZN(n17119) );
  AND2_X1 U19307 ( .A1(n17120), .A2(n17119), .ZN(n17123) );
  OAI22_X1 U19308 ( .A1(n17122), .A2(n17121), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17123), .ZN(n17125) );
  NAND2_X1 U19309 ( .A1(n17123), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n17124) );
  OAI211_X1 U19310 ( .C1(n17126), .C2(n22018), .A(n17125), .B(n17124), .ZN(
        n17127) );
  OAI21_X1 U19311 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17128), .A(
        n17127), .ZN(n17132) );
  NAND2_X1 U19312 ( .A1(n17129), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17131) );
  INV_X1 U19313 ( .A(n17129), .ZN(n17130) );
  AOI22_X1 U19314 ( .A1(n17132), .A2(n17131), .B1(n17130), .B2(n12225), .ZN(
        n17141) );
  INV_X1 U19315 ( .A(n17133), .ZN(n17138) );
  AOI21_X1 U19316 ( .B1(n21823), .B2(n17135), .A(n17134), .ZN(n17137) );
  NOR4_X1 U19317 ( .A1(n17139), .A2(n17138), .A3(n17137), .A4(n17136), .ZN(
        n17140) );
  OAI21_X1 U19318 ( .B1(n17141), .B2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n17140), .ZN(n17142) );
  INV_X1 U19319 ( .A(n17142), .ZN(n21845) );
  NOR2_X1 U19320 ( .A1(n21875), .A2(n17143), .ZN(n17145) );
  AND3_X1 U19321 ( .A1(n17146), .A2(n17145), .A3(n17144), .ZN(n17147) );
  AOI221_X1 U19322 ( .B1(n17149), .B2(n17148), .C1(n21455), .C2(n17148), .A(
        n17147), .ZN(n17151) );
  OAI221_X1 U19323 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n21845), 
        .A(n17151), .ZN(n21831) );
  OAI211_X1 U19324 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21455), .A(n17150), 
        .B(n21831), .ZN(n21841) );
  OAI221_X1 U19325 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n21832), .C2(n21455), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21833) );
  AOI21_X1 U19326 ( .B1(n21833), .B2(n17152), .A(n17151), .ZN(n17153) );
  AOI21_X1 U19327 ( .B1(n17154), .B2(n21841), .A(n17153), .ZN(P1_U3162) );
  NOR2_X1 U19328 ( .A1(n17156), .A2(n17155), .ZN(P1_U3032) );
  AND2_X1 U19329 ( .A1(n20060), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19330 ( .A1(n17157), .A2(n12216), .ZN(n17159) );
  INV_X1 U19331 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17158) );
  AOI21_X1 U19332 ( .B1(n17159), .B2(n17158), .A(n22398), .ZN(P1_U2802) );
  OAI22_X1 U19333 ( .A1(n17161), .A2(keyinput_59), .B1(n17260), .B2(
        keyinput_60), .ZN(n17160) );
  AOI221_X1 U19334 ( .B1(n17161), .B2(keyinput_59), .C1(keyinput_60), .C2(
        n17260), .A(n17160), .ZN(n17255) );
  OAI22_X1 U19335 ( .A1(n16065), .A2(keyinput_57), .B1(n16058), .B2(
        keyinput_56), .ZN(n17162) );
  AOI221_X1 U19336 ( .B1(n16065), .B2(keyinput_57), .C1(keyinput_56), .C2(
        n16058), .A(n17162), .ZN(n17252) );
  INV_X1 U19337 ( .A(keyinput_55), .ZN(n17250) );
  INV_X1 U19338 ( .A(keyinput_54), .ZN(n17248) );
  INV_X1 U19339 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U19340 ( .A1(n17263), .A2(keyinput_51), .B1(n17264), .B2(
        keyinput_52), .ZN(n17163) );
  OAI221_X1 U19341 ( .B1(n17263), .B2(keyinput_51), .C1(n17264), .C2(
        keyinput_52), .A(n17163), .ZN(n17246) );
  INV_X1 U19342 ( .A(keyinput_50), .ZN(n17243) );
  INV_X1 U19343 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20121) );
  INV_X1 U19344 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20125) );
  OAI22_X1 U19345 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_46), .B1(
        P1_W_R_N_REG_SCAN_IN), .B2(keyinput_47), .ZN(n17164) );
  AOI221_X1 U19346 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_46), .C1(
        keyinput_47), .C2(P1_W_R_N_REG_SCAN_IN), .A(n17164), .ZN(n17170) );
  OAI22_X1 U19347 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_42), .B1(
        P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_43), .ZN(n17165) );
  AOI221_X1 U19348 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_42), .C1(
        keyinput_43), .C2(P1_REQUESTPENDING_REG_SCAN_IN), .A(n17165), .ZN(
        n17169) );
  OAI22_X1 U19349 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(keyinput_44), .B1(
        P1_MORE_REG_SCAN_IN), .B2(keyinput_45), .ZN(n17166) );
  AOI221_X1 U19350 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_44), .C1(
        keyinput_45), .C2(P1_MORE_REG_SCAN_IN), .A(n17166), .ZN(n17168) );
  INV_X1 U19351 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20128) );
  XOR2_X1 U19352 ( .A(n20128), .B(keyinput_48), .Z(n17167) );
  NAND4_X1 U19353 ( .A1(n17170), .A2(n17169), .A3(n17168), .A4(n17167), .ZN(
        n17240) );
  OAI22_X1 U19354 ( .A1(n17172), .A2(keyinput_40), .B1(P1_ADS_N_REG_SCAN_IN), 
        .B2(keyinput_39), .ZN(n17171) );
  AOI221_X1 U19355 ( .B1(n17172), .B2(keyinput_40), .C1(keyinput_39), .C2(
        P1_ADS_N_REG_SCAN_IN), .A(n17171), .ZN(n17237) );
  INV_X1 U19356 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n17344) );
  INV_X1 U19357 ( .A(keyinput_38), .ZN(n17235) );
  INV_X1 U19358 ( .A(READY2), .ZN(n17342) );
  INV_X1 U19359 ( .A(keyinput_37), .ZN(n17233) );
  INV_X1 U19360 ( .A(HOLD), .ZN(n21908) );
  INV_X1 U19361 ( .A(keyinput_33), .ZN(n17226) );
  AOI22_X1 U19362 ( .A1(DATAI_1_), .A2(keyinput_31), .B1(DATAI_2_), .B2(
        keyinput_30), .ZN(n17173) );
  OAI221_X1 U19363 ( .B1(DATAI_1_), .B2(keyinput_31), .C1(DATAI_2_), .C2(
        keyinput_30), .A(n17173), .ZN(n17223) );
  INV_X1 U19364 ( .A(DATAI_3_), .ZN(n17328) );
  INV_X1 U19365 ( .A(keyinput_29), .ZN(n17221) );
  INV_X1 U19366 ( .A(DATAI_6_), .ZN(n17276) );
  OAI22_X1 U19367 ( .A1(n17276), .A2(keyinput_26), .B1(keyinput_28), .B2(
        DATAI_4_), .ZN(n17174) );
  AOI221_X1 U19368 ( .B1(n17276), .B2(keyinput_26), .C1(DATAI_4_), .C2(
        keyinput_28), .A(n17174), .ZN(n17218) );
  INV_X1 U19369 ( .A(DATAI_7_), .ZN(n17322) );
  INV_X1 U19370 ( .A(keyinput_25), .ZN(n17216) );
  INV_X1 U19371 ( .A(DATAI_14_), .ZN(n17278) );
  INV_X1 U19372 ( .A(DATAI_13_), .ZN(n17176) );
  OAI22_X1 U19373 ( .A1(n17278), .A2(keyinput_18), .B1(n17176), .B2(
        keyinput_19), .ZN(n17175) );
  AOI221_X1 U19374 ( .B1(n17278), .B2(keyinput_18), .C1(keyinput_19), .C2(
        n17176), .A(n17175), .ZN(n17214) );
  OAI22_X1 U19375 ( .A1(DATAI_12_), .A2(keyinput_20), .B1(DATAI_15_), .B2(
        keyinput_17), .ZN(n17177) );
  AOI221_X1 U19376 ( .B1(DATAI_12_), .B2(keyinput_20), .C1(keyinput_17), .C2(
        DATAI_15_), .A(n17177), .ZN(n17213) );
  INV_X1 U19377 ( .A(DATAI_8_), .ZN(n17179) );
  OAI22_X1 U19378 ( .A1(n17179), .A2(keyinput_24), .B1(keyinput_22), .B2(
        DATAI_10_), .ZN(n17178) );
  AOI221_X1 U19379 ( .B1(n17179), .B2(keyinput_24), .C1(DATAI_10_), .C2(
        keyinput_22), .A(n17178), .ZN(n17183) );
  INV_X1 U19380 ( .A(DATAI_9_), .ZN(n17287) );
  OAI22_X1 U19381 ( .A1(n17287), .A2(keyinput_23), .B1(n17181), .B2(
        keyinput_16), .ZN(n17180) );
  AOI221_X1 U19382 ( .B1(n17287), .B2(keyinput_23), .C1(keyinput_16), .C2(
        n17181), .A(n17180), .ZN(n17182) );
  OAI211_X1 U19383 ( .C1(DATAI_11_), .C2(keyinput_21), .A(n17183), .B(n17182), 
        .ZN(n17184) );
  AOI21_X1 U19384 ( .B1(DATAI_11_), .B2(keyinput_21), .A(n17184), .ZN(n17212)
         );
  INV_X1 U19385 ( .A(keyinput_15), .ZN(n17210) );
  OAI22_X1 U19386 ( .A1(n17289), .A2(keyinput_12), .B1(n17186), .B2(
        keyinput_13), .ZN(n17185) );
  AOI221_X1 U19387 ( .B1(n17289), .B2(keyinput_12), .C1(keyinput_13), .C2(
        n17186), .A(n17185), .ZN(n17206) );
  INV_X1 U19388 ( .A(keyinput_11), .ZN(n17204) );
  INV_X1 U19389 ( .A(keyinput_10), .ZN(n17202) );
  OAI22_X1 U19390 ( .A1(DATAI_31_), .A2(keyinput_1), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_0), .ZN(n17187) );
  AOI221_X1 U19391 ( .B1(DATAI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P1_MEMORYFETCH_REG_SCAN_IN), .A(n17187), .ZN(n17190) );
  XNOR2_X1 U19392 ( .A(n17188), .B(keyinput_2), .ZN(n17189) );
  AOI22_X1 U19393 ( .A1(n17190), .A2(n17189), .B1(keyinput_4), .B2(n17192), 
        .ZN(n17191) );
  OAI21_X1 U19394 ( .B1(keyinput_4), .B2(n17192), .A(n17191), .ZN(n17200) );
  AOI22_X1 U19395 ( .A1(DATAI_27_), .A2(keyinput_5), .B1(n17194), .B2(
        keyinput_3), .ZN(n17193) );
  OAI221_X1 U19396 ( .B1(DATAI_27_), .B2(keyinput_5), .C1(n17194), .C2(
        keyinput_3), .A(n17193), .ZN(n17199) );
  OAI22_X1 U19397 ( .A1(n17299), .A2(keyinput_9), .B1(keyinput_8), .B2(
        DATAI_24_), .ZN(n17195) );
  AOI221_X1 U19398 ( .B1(n17299), .B2(keyinput_9), .C1(DATAI_24_), .C2(
        keyinput_8), .A(n17195), .ZN(n17198) );
  OAI22_X1 U19399 ( .A1(DATAI_26_), .A2(keyinput_6), .B1(keyinput_7), .B2(
        DATAI_25_), .ZN(n17196) );
  AOI221_X1 U19400 ( .B1(DATAI_26_), .B2(keyinput_6), .C1(DATAI_25_), .C2(
        keyinput_7), .A(n17196), .ZN(n17197) );
  OAI211_X1 U19401 ( .C1(n17200), .C2(n17199), .A(n17198), .B(n17197), .ZN(
        n17201) );
  OAI221_X1 U19402 ( .B1(DATAI_22_), .B2(n17202), .C1(n17307), .C2(keyinput_10), .A(n17201), .ZN(n17203) );
  OAI221_X1 U19403 ( .B1(DATAI_21_), .B2(keyinput_11), .C1(n17309), .C2(n17204), .A(n17203), .ZN(n17205) );
  AOI22_X1 U19404 ( .A1(keyinput_14), .A2(n17208), .B1(n17206), .B2(n17205), 
        .ZN(n17207) );
  OAI21_X1 U19405 ( .B1(n17208), .B2(keyinput_14), .A(n17207), .ZN(n17209) );
  OAI221_X1 U19406 ( .B1(DATAI_17_), .B2(keyinput_15), .C1(n17315), .C2(n17210), .A(n17209), .ZN(n17211) );
  NAND4_X1 U19407 ( .A1(n17214), .A2(n17213), .A3(n17212), .A4(n17211), .ZN(
        n17215) );
  OAI221_X1 U19408 ( .B1(DATAI_7_), .B2(keyinput_25), .C1(n17322), .C2(n17216), 
        .A(n17215), .ZN(n17217) );
  OAI211_X1 U19409 ( .C1(DATAI_5_), .C2(keyinput_27), .A(n17218), .B(n17217), 
        .ZN(n17219) );
  AOI21_X1 U19410 ( .B1(DATAI_5_), .B2(keyinput_27), .A(n17219), .ZN(n17220)
         );
  AOI221_X1 U19411 ( .B1(DATAI_3_), .B2(keyinput_29), .C1(n17328), .C2(n17221), 
        .A(n17220), .ZN(n17222) );
  OAI22_X1 U19412 ( .A1(n17223), .A2(n17222), .B1(keyinput_32), .B2(DATAI_0_), 
        .ZN(n17224) );
  AOI21_X1 U19413 ( .B1(keyinput_32), .B2(DATAI_0_), .A(n17224), .ZN(n17225)
         );
  AOI221_X1 U19414 ( .B1(HOLD), .B2(keyinput_33), .C1(n21908), .C2(n17226), 
        .A(n17225), .ZN(n17230) );
  AOI22_X1 U19415 ( .A1(NA), .A2(keyinput_34), .B1(n17228), .B2(keyinput_35), 
        .ZN(n17227) );
  OAI221_X1 U19416 ( .B1(NA), .B2(keyinput_34), .C1(n17228), .C2(keyinput_35), 
        .A(n17227), .ZN(n17229) );
  AOI211_X1 U19417 ( .C1(READY1), .C2(keyinput_36), .A(n17230), .B(n17229), 
        .ZN(n17231) );
  OAI21_X1 U19418 ( .B1(READY1), .B2(keyinput_36), .A(n17231), .ZN(n17232) );
  OAI221_X1 U19419 ( .B1(READY2), .B2(keyinput_37), .C1(n17342), .C2(n17233), 
        .A(n17232), .ZN(n17234) );
  OAI221_X1 U19420 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_38), .C1(
        n17344), .C2(n17235), .A(n17234), .ZN(n17236) );
  OAI211_X1 U19421 ( .C1(n22396), .C2(keyinput_41), .A(n17237), .B(n17236), 
        .ZN(n17238) );
  AOI21_X1 U19422 ( .B1(n22396), .B2(keyinput_41), .A(n17238), .ZN(n17239) );
  OAI22_X1 U19423 ( .A1(keyinput_49), .A2(n20125), .B1(n17240), .B2(n17239), 
        .ZN(n17241) );
  AOI21_X1 U19424 ( .B1(keyinput_49), .B2(n20125), .A(n17241), .ZN(n17242) );
  AOI221_X1 U19425 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n17243), .C1(
        n20121), .C2(keyinput_50), .A(n17242), .ZN(n17245) );
  NAND2_X1 U19426 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_53), .ZN(n17244) );
  OAI221_X1 U19427 ( .B1(n17246), .B2(n17245), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(keyinput_53), .A(n17244), .ZN(n17247) );
  OAI221_X1 U19428 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_54), .C1(
        n17359), .C2(n17248), .A(n17247), .ZN(n17249) );
  OAI221_X1 U19429 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_55), .C1(
        n17362), .C2(n17250), .A(n17249), .ZN(n17251) );
  AOI22_X1 U19430 ( .A1(keyinput_58), .A2(n17367), .B1(n17252), .B2(n17251), 
        .ZN(n17253) );
  OAI21_X1 U19431 ( .B1(n17367), .B2(keyinput_58), .A(n17253), .ZN(n17254) );
  AOI22_X1 U19432 ( .A1(n17255), .A2(n17254), .B1(keyinput_61), .B2(n21803), 
        .ZN(n17256) );
  OAI21_X1 U19433 ( .B1(keyinput_61), .B2(n21803), .A(n17256), .ZN(n17374) );
  AOI22_X1 U19434 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_62), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_63), .ZN(n17257) );
  OAI221_X1 U19435 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_62), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_63), .A(n17257), .ZN(n17373) );
  OAI22_X1 U19436 ( .A1(n21807), .A2(keyinput_126), .B1(n21803), .B2(
        keyinput_125), .ZN(n17258) );
  AOI221_X1 U19437 ( .B1(n21807), .B2(keyinput_126), .C1(keyinput_125), .C2(
        n21803), .A(n17258), .ZN(n17372) );
  AOI22_X1 U19438 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_123), .B1(
        n17260), .B2(keyinput_124), .ZN(n17259) );
  OAI221_X1 U19439 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_123), .C1(
        n17260), .C2(keyinput_124), .A(n17259), .ZN(n17369) );
  AOI22_X1 U19440 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(keyinput_120), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(keyinput_121), .ZN(n17261) );
  OAI221_X1 U19441 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput_120), .C1(
        P1_REIP_REG_26__SCAN_IN), .C2(keyinput_121), .A(n17261), .ZN(n17365)
         );
  INV_X1 U19442 ( .A(keyinput_119), .ZN(n17363) );
  INV_X1 U19443 ( .A(keyinput_118), .ZN(n17360) );
  AOI22_X1 U19444 ( .A1(n17264), .A2(keyinput_116), .B1(keyinput_115), .B2(
        n17263), .ZN(n17262) );
  OAI221_X1 U19445 ( .B1(n17264), .B2(keyinput_116), .C1(n17263), .C2(
        keyinput_115), .A(n17262), .ZN(n17355) );
  INV_X1 U19446 ( .A(keyinput_114), .ZN(n17353) );
  OAI22_X1 U19447 ( .A1(n22050), .A2(keyinput_108), .B1(n21823), .B2(
        keyinput_110), .ZN(n17265) );
  AOI221_X1 U19448 ( .B1(n22050), .B2(keyinput_108), .C1(keyinput_110), .C2(
        n21823), .A(n17265), .ZN(n17271) );
  OAI22_X1 U19449 ( .A1(n20128), .A2(keyinput_112), .B1(keyinput_109), .B2(
        P1_MORE_REG_SCAN_IN), .ZN(n17266) );
  AOI221_X1 U19450 ( .B1(n20128), .B2(keyinput_112), .C1(P1_MORE_REG_SCAN_IN), 
        .C2(keyinput_109), .A(n17266), .ZN(n17270) );
  INV_X1 U19451 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20241) );
  OAI22_X1 U19452 ( .A1(n20241), .A2(keyinput_106), .B1(keyinput_107), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n17267) );
  AOI221_X1 U19453 ( .B1(n20241), .B2(keyinput_106), .C1(
        P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_107), .A(n17267), .ZN(
        n17269) );
  XNOR2_X1 U19454 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_111), .ZN(n17268) );
  NAND4_X1 U19455 ( .A1(n17271), .A2(n17270), .A3(n17269), .A4(n17268), .ZN(
        n17350) );
  OAI22_X1 U19456 ( .A1(n22396), .A2(keyinput_105), .B1(keyinput_104), .B2(
        P1_CODEFETCH_REG_SCAN_IN), .ZN(n17272) );
  AOI221_X1 U19457 ( .B1(n22396), .B2(keyinput_105), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_104), .A(n17272), .ZN(n17347)
         );
  INV_X1 U19458 ( .A(keyinput_102), .ZN(n17345) );
  INV_X1 U19459 ( .A(keyinput_101), .ZN(n17341) );
  INV_X1 U19460 ( .A(keyinput_97), .ZN(n17334) );
  INV_X1 U19461 ( .A(DATAI_1_), .ZN(n17274) );
  AOI22_X1 U19462 ( .A1(DATAI_2_), .A2(keyinput_94), .B1(n17274), .B2(
        keyinput_95), .ZN(n17273) );
  OAI221_X1 U19463 ( .B1(DATAI_2_), .B2(keyinput_94), .C1(n17274), .C2(
        keyinput_95), .A(n17273), .ZN(n17331) );
  INV_X1 U19464 ( .A(keyinput_93), .ZN(n17329) );
  OAI22_X1 U19465 ( .A1(n17276), .A2(keyinput_90), .B1(DATAI_5_), .B2(
        keyinput_91), .ZN(n17275) );
  AOI221_X1 U19466 ( .B1(n17276), .B2(keyinput_90), .C1(keyinput_91), .C2(
        DATAI_5_), .A(n17275), .ZN(n17325) );
  INV_X1 U19467 ( .A(keyinput_89), .ZN(n17323) );
  OAI22_X1 U19468 ( .A1(n17278), .A2(keyinput_82), .B1(keyinput_84), .B2(
        DATAI_12_), .ZN(n17277) );
  AOI221_X1 U19469 ( .B1(n17278), .B2(keyinput_82), .C1(DATAI_12_), .C2(
        keyinput_84), .A(n17277), .ZN(n17320) );
  OAI22_X1 U19470 ( .A1(DATAI_13_), .A2(keyinput_83), .B1(DATAI_15_), .B2(
        keyinput_81), .ZN(n17279) );
  AOI221_X1 U19471 ( .B1(DATAI_13_), .B2(keyinput_83), .C1(keyinput_81), .C2(
        DATAI_15_), .A(n17279), .ZN(n17319) );
  INV_X1 U19472 ( .A(DATAI_10_), .ZN(n17282) );
  INV_X1 U19473 ( .A(DATAI_11_), .ZN(n17281) );
  AOI22_X1 U19474 ( .A1(n17282), .A2(keyinput_86), .B1(n17281), .B2(
        keyinput_85), .ZN(n17280) );
  OAI221_X1 U19475 ( .B1(n17282), .B2(keyinput_86), .C1(n17281), .C2(
        keyinput_85), .A(n17280), .ZN(n17286) );
  OAI22_X1 U19476 ( .A1(DATAI_8_), .A2(keyinput_88), .B1(keyinput_80), .B2(
        DATAI_16_), .ZN(n17283) );
  AOI221_X1 U19477 ( .B1(DATAI_8_), .B2(keyinput_88), .C1(DATAI_16_), .C2(
        keyinput_80), .A(n17283), .ZN(n17284) );
  OAI21_X1 U19478 ( .B1(keyinput_87), .B2(n17287), .A(n17284), .ZN(n17285) );
  AOI211_X1 U19479 ( .C1(keyinput_87), .C2(n17287), .A(n17286), .B(n17285), 
        .ZN(n17318) );
  INV_X1 U19480 ( .A(keyinput_79), .ZN(n17316) );
  AOI22_X1 U19481 ( .A1(DATAI_19_), .A2(keyinput_77), .B1(n17289), .B2(
        keyinput_76), .ZN(n17288) );
  OAI221_X1 U19482 ( .B1(DATAI_19_), .B2(keyinput_77), .C1(n17289), .C2(
        keyinput_76), .A(n17288), .ZN(n17313) );
  INV_X1 U19483 ( .A(keyinput_75), .ZN(n17310) );
  INV_X1 U19484 ( .A(keyinput_74), .ZN(n17306) );
  XOR2_X1 U19485 ( .A(n17290), .B(keyinput_65), .Z(n17293) );
  AOI22_X1 U19486 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_64), .B1(
        DATAI_30_), .B2(keyinput_66), .ZN(n17291) );
  OAI221_X1 U19487 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_64), .C1(
        DATAI_30_), .C2(keyinput_66), .A(n17291), .ZN(n17292) );
  OAI22_X1 U19488 ( .A1(n17293), .A2(n17292), .B1(n17295), .B2(keyinput_69), 
        .ZN(n17294) );
  AOI21_X1 U19489 ( .B1(n17295), .B2(keyinput_69), .A(n17294), .ZN(n17304) );
  OAI22_X1 U19490 ( .A1(DATAI_29_), .A2(keyinput_67), .B1(keyinput_68), .B2(
        DATAI_28_), .ZN(n17296) );
  AOI221_X1 U19491 ( .B1(DATAI_29_), .B2(keyinput_67), .C1(DATAI_28_), .C2(
        keyinput_68), .A(n17296), .ZN(n17303) );
  AOI22_X1 U19492 ( .A1(n17299), .A2(keyinput_73), .B1(n17298), .B2(
        keyinput_71), .ZN(n17297) );
  OAI221_X1 U19493 ( .B1(n17299), .B2(keyinput_73), .C1(n17298), .C2(
        keyinput_71), .A(n17297), .ZN(n17302) );
  AOI22_X1 U19494 ( .A1(DATAI_24_), .A2(keyinput_72), .B1(DATAI_26_), .B2(
        keyinput_70), .ZN(n17300) );
  OAI221_X1 U19495 ( .B1(DATAI_24_), .B2(keyinput_72), .C1(DATAI_26_), .C2(
        keyinput_70), .A(n17300), .ZN(n17301) );
  AOI211_X1 U19496 ( .C1(n17304), .C2(n17303), .A(n17302), .B(n17301), .ZN(
        n17305) );
  AOI221_X1 U19497 ( .B1(DATAI_22_), .B2(keyinput_74), .C1(n17307), .C2(n17306), .A(n17305), .ZN(n17308) );
  AOI221_X1 U19498 ( .B1(DATAI_21_), .B2(n17310), .C1(n17309), .C2(keyinput_75), .A(n17308), .ZN(n17312) );
  NAND2_X1 U19499 ( .A1(DATAI_18_), .A2(keyinput_78), .ZN(n17311) );
  OAI221_X1 U19500 ( .B1(n17313), .B2(n17312), .C1(DATAI_18_), .C2(keyinput_78), .A(n17311), .ZN(n17314) );
  OAI221_X1 U19501 ( .B1(DATAI_17_), .B2(n17316), .C1(n17315), .C2(keyinput_79), .A(n17314), .ZN(n17317) );
  NAND4_X1 U19502 ( .A1(n17320), .A2(n17319), .A3(n17318), .A4(n17317), .ZN(
        n17321) );
  OAI221_X1 U19503 ( .B1(DATAI_7_), .B2(n17323), .C1(n17322), .C2(keyinput_89), 
        .A(n17321), .ZN(n17324) );
  OAI211_X1 U19504 ( .C1(DATAI_4_), .C2(keyinput_92), .A(n17325), .B(n17324), 
        .ZN(n17326) );
  AOI21_X1 U19505 ( .B1(DATAI_4_), .B2(keyinput_92), .A(n17326), .ZN(n17327)
         );
  AOI221_X1 U19506 ( .B1(DATAI_3_), .B2(n17329), .C1(n17328), .C2(keyinput_93), 
        .A(n17327), .ZN(n17330) );
  OAI22_X1 U19507 ( .A1(n17331), .A2(n17330), .B1(keyinput_96), .B2(DATAI_0_), 
        .ZN(n17332) );
  AOI21_X1 U19508 ( .B1(keyinput_96), .B2(DATAI_0_), .A(n17332), .ZN(n17333)
         );
  AOI221_X1 U19509 ( .B1(HOLD), .B2(keyinput_97), .C1(n21908), .C2(n17334), 
        .A(n17333), .ZN(n17338) );
  INV_X1 U19510 ( .A(READY1), .ZN(n17336) );
  INV_X1 U19511 ( .A(NA), .ZN(n21911) );
  AOI22_X1 U19512 ( .A1(n17336), .A2(keyinput_100), .B1(keyinput_98), .B2(
        n21911), .ZN(n17335) );
  OAI221_X1 U19513 ( .B1(n17336), .B2(keyinput_100), .C1(n21911), .C2(
        keyinput_98), .A(n17335), .ZN(n17337) );
  AOI211_X1 U19514 ( .C1(BS16), .C2(keyinput_99), .A(n17338), .B(n17337), .ZN(
        n17339) );
  OAI21_X1 U19515 ( .B1(BS16), .B2(keyinput_99), .A(n17339), .ZN(n17340) );
  OAI221_X1 U19516 ( .B1(READY2), .B2(keyinput_101), .C1(n17342), .C2(n17341), 
        .A(n17340), .ZN(n17343) );
  OAI221_X1 U19517 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(n17345), .C1(n17344), 
        .C2(keyinput_102), .A(n17343), .ZN(n17346) );
  OAI211_X1 U19518 ( .C1(P1_ADS_N_REG_SCAN_IN), .C2(keyinput_103), .A(n17347), 
        .B(n17346), .ZN(n17348) );
  AOI21_X1 U19519 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_103), .A(n17348), 
        .ZN(n17349) );
  OAI22_X1 U19520 ( .A1(keyinput_113), .A2(n20125), .B1(n17350), .B2(n17349), 
        .ZN(n17351) );
  AOI21_X1 U19521 ( .B1(keyinput_113), .B2(n20125), .A(n17351), .ZN(n17352) );
  AOI221_X1 U19522 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_114), 
        .C1(n20121), .C2(n17353), .A(n17352), .ZN(n17354) );
  OAI22_X1 U19523 ( .A1(keyinput_117), .A2(n17357), .B1(n17355), .B2(n17354), 
        .ZN(n17356) );
  AOI21_X1 U19524 ( .B1(keyinput_117), .B2(n17357), .A(n17356), .ZN(n17358) );
  AOI221_X1 U19525 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n17360), .C1(n17359), 
        .C2(keyinput_118), .A(n17358), .ZN(n17361) );
  AOI221_X1 U19526 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n17363), .C1(n17362), 
        .C2(keyinput_119), .A(n17361), .ZN(n17364) );
  OAI22_X1 U19527 ( .A1(keyinput_122), .A2(n17367), .B1(n17365), .B2(n17364), 
        .ZN(n17366) );
  AOI21_X1 U19528 ( .B1(keyinput_122), .B2(n17367), .A(n17366), .ZN(n17368) );
  OAI22_X1 U19529 ( .A1(n17369), .A2(n17368), .B1(P1_REIP_REG_20__SCAN_IN), 
        .B2(keyinput_127), .ZN(n17370) );
  AOI21_X1 U19530 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_127), .A(n17370), .ZN(n17371) );
  OAI211_X1 U19531 ( .C1(n17374), .C2(n17373), .A(n17372), .B(n17371), .ZN(
        n17386) );
  AOI22_X1 U19532 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19875), .ZN(n19852) );
  NOR2_X1 U19533 ( .A1(n19495), .A2(n19528), .ZN(n19959) );
  OAI21_X1 U19534 ( .B1(n17377), .B2(n19959), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17375) );
  OR2_X1 U19535 ( .A1(n19497), .A2(n19528), .ZN(n17379) );
  NAND2_X1 U19536 ( .A1(n17375), .A2(n17379), .ZN(n19960) );
  NOR2_X2 U19537 ( .A1(n15667), .A2(n19871), .ZN(n19853) );
  AOI22_X1 U19538 ( .A1(n19960), .A2(n17376), .B1(n19853), .B2(n19959), .ZN(
        n17384) );
  INV_X1 U19539 ( .A(n17377), .ZN(n17378) );
  AOI21_X1 U19540 ( .B1(n17378), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n17382) );
  OAI21_X1 U19541 ( .B1(n19846), .B2(n19961), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n17380) );
  NAND3_X1 U19542 ( .A1(n17380), .A2(n19508), .A3(n17379), .ZN(n17381) );
  OAI211_X1 U19543 ( .C1(n19959), .C2(n17382), .A(n17381), .B(n19475), .ZN(
        n19962) );
  AOI22_X1 U19544 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19875), .ZN(n19842) );
  AOI22_X1 U19545 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n19854), .ZN(n17383) );
  OAI211_X1 U19546 ( .C1(n19852), .C2(n19965), .A(n17384), .B(n17383), .ZN(
        n17385) );
  XNOR2_X1 U19547 ( .A(n17386), .B(n17385), .ZN(P2_U3065) );
  INV_X1 U19548 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17542) );
  INV_X1 U19549 ( .A(n17387), .ZN(n18883) );
  OAI22_X1 U19550 ( .A1(n17388), .A2(n17542), .B1(n18883), .B2(n18891), .ZN(
        P2_U2816) );
  AOI22_X1 U19551 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n16328), .B1(n17453), 
        .B2(n17389), .ZN(n17399) );
  XNOR2_X1 U19552 ( .A(n17390), .B(n18860), .ZN(n17402) );
  XNOR2_X1 U19553 ( .A(n17402), .B(n17391), .ZN(n18857) );
  CLKBUF_X1 U19554 ( .A(n17392), .Z(n17395) );
  XNOR2_X1 U19555 ( .A(n17393), .B(n18860), .ZN(n17394) );
  XNOR2_X1 U19556 ( .A(n17395), .B(n17394), .ZN(n18854) );
  INV_X1 U19557 ( .A(n18854), .ZN(n17396) );
  AOI222_X1 U19558 ( .A1(n18857), .A2(n17475), .B1(n17397), .B2(n17474), .C1(
        n17473), .C2(n17396), .ZN(n17398) );
  OAI211_X1 U19559 ( .C1(n17400), .C2(n17459), .A(n17399), .B(n17398), .ZN(
        P2_U3011) );
  AOI22_X1 U19560 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17470), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n16328), .ZN(n17408) );
  AOI22_X1 U19561 ( .A1(n17402), .A2(n17401), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17390), .ZN(n17404) );
  XNOR2_X1 U19562 ( .A(n18482), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17403) );
  XNOR2_X1 U19563 ( .A(n17404), .B(n17403), .ZN(n18841) );
  INV_X1 U19564 ( .A(n18484), .ZN(n18837) );
  XNOR2_X1 U19565 ( .A(n17405), .B(n18844), .ZN(n18839) );
  INV_X1 U19566 ( .A(n18839), .ZN(n17406) );
  AOI222_X1 U19567 ( .A1(n18841), .A2(n17475), .B1(n17474), .B2(n18837), .C1(
        n17473), .C2(n17406), .ZN(n17407) );
  OAI211_X1 U19568 ( .C1(n17479), .C2(n18487), .A(n17408), .B(n17407), .ZN(
        P2_U3010) );
  AOI22_X1 U19569 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n16675), .B1(n17453), 
        .B2(n18501), .ZN(n17413) );
  OAI22_X1 U19570 ( .A1(n17463), .A2(n17410), .B1(n17409), .B2(n17461), .ZN(
        n17411) );
  AOI21_X1 U19571 ( .B1(n17474), .B2(n18503), .A(n17411), .ZN(n17412) );
  OAI211_X1 U19572 ( .C1(n17414), .C2(n17459), .A(n17413), .B(n17412), .ZN(
        P2_U3009) );
  AOI22_X1 U19573 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17470), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n16675), .ZN(n17422) );
  NAND3_X1 U19574 ( .A1(n17416), .A2(n17473), .A3(n17415), .ZN(n17418) );
  NAND2_X1 U19575 ( .A1(n18514), .A2(n17474), .ZN(n17417) );
  OAI211_X1 U19576 ( .C1(n17461), .C2(n17419), .A(n17418), .B(n17417), .ZN(
        n17420) );
  INV_X1 U19577 ( .A(n17420), .ZN(n17421) );
  OAI211_X1 U19578 ( .C1(n17479), .C2(n18511), .A(n17422), .B(n17421), .ZN(
        P2_U3008) );
  AOI22_X1 U19579 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17470), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n16328), .ZN(n17435) );
  NOR2_X1 U19580 ( .A1(n17424), .A2(n17423), .ZN(n17429) );
  INV_X1 U19581 ( .A(n17425), .ZN(n17427) );
  NOR2_X1 U19582 ( .A1(n17427), .A2(n17426), .ZN(n17428) );
  XNOR2_X1 U19583 ( .A(n17429), .B(n17428), .ZN(n18827) );
  INV_X1 U19584 ( .A(n18538), .ZN(n18826) );
  OAI21_X1 U19585 ( .B1(n17432), .B2(n17431), .A(n17430), .ZN(n17433) );
  INV_X1 U19586 ( .A(n17433), .ZN(n18824) );
  AOI222_X1 U19587 ( .A1(n18827), .A2(n17475), .B1(n17474), .B2(n18826), .C1(
        n17473), .C2(n18824), .ZN(n17434) );
  OAI211_X1 U19588 ( .C1(n17479), .C2(n18533), .A(n17435), .B(n17434), .ZN(
        P2_U3006) );
  AOI22_X1 U19589 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n16328), .B1(n17453), 
        .B2(n18540), .ZN(n17440) );
  OAI22_X1 U19590 ( .A1(n17437), .A2(n17463), .B1(n17461), .B2(n17436), .ZN(
        n17438) );
  AOI21_X1 U19591 ( .B1(n17474), .B2(n18544), .A(n17438), .ZN(n17439) );
  OAI211_X1 U19592 ( .C1(n17441), .C2(n17459), .A(n17440), .B(n17439), .ZN(
        P2_U3005) );
  AOI22_X1 U19593 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17470), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n16675), .ZN(n17452) );
  AOI21_X1 U19594 ( .B1(n18814), .B2(n17443), .A(n17442), .ZN(n18819) );
  NOR2_X1 U19595 ( .A1(n17028), .A2(n17444), .ZN(n17448) );
  NAND2_X1 U19596 ( .A1(n17446), .A2(n17445), .ZN(n17447) );
  XNOR2_X1 U19597 ( .A(n17448), .B(n17447), .ZN(n18822) );
  OAI22_X1 U19598 ( .A1(n18822), .A2(n17461), .B1(n17449), .B2(n18817), .ZN(
        n17450) );
  AOI21_X1 U19599 ( .B1(n18819), .B2(n17473), .A(n17450), .ZN(n17451) );
  OAI211_X1 U19600 ( .C1(n17479), .C2(n18558), .A(n17452), .B(n17451), .ZN(
        P2_U3004) );
  AOI22_X1 U19601 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n16675), .B1(n17453), 
        .B2(n18568), .ZN(n17458) );
  OAI22_X1 U19602 ( .A1(n17455), .A2(n17463), .B1(n17454), .B2(n17461), .ZN(
        n17456) );
  AOI21_X1 U19603 ( .B1(n17474), .B2(n18570), .A(n17456), .ZN(n17457) );
  OAI211_X1 U19604 ( .C1(n17460), .C2(n17459), .A(n17458), .B(n17457), .ZN(
        P2_U3003) );
  AOI22_X1 U19605 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17470), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n16328), .ZN(n17469) );
  NOR2_X1 U19606 ( .A1(n17462), .A2(n17461), .ZN(n17467) );
  NOR3_X1 U19607 ( .A1(n17465), .A2(n17464), .A3(n17463), .ZN(n17466) );
  AOI211_X1 U19608 ( .C1(n17474), .C2(n18580), .A(n17467), .B(n17466), .ZN(
        n17468) );
  OAI211_X1 U19609 ( .C1(n17479), .C2(n18574), .A(n17469), .B(n17468), .ZN(
        P2_U3002) );
  AOI22_X1 U19610 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17470), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n16675), .ZN(n17478) );
  INV_X1 U19611 ( .A(n17471), .ZN(n18600) );
  AOI222_X1 U19612 ( .A1(n17476), .A2(n17475), .B1(n17474), .B2(n18600), .C1(
        n17473), .C2(n17472), .ZN(n17477) );
  OAI211_X1 U19613 ( .C1(n17479), .C2(n18595), .A(n17478), .B(n17477), .ZN(
        P2_U3000) );
  INV_X1 U19614 ( .A(n17497), .ZN(n17499) );
  OAI22_X1 U19615 ( .A1(n17481), .A2(n17480), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19472), .ZN(n17482) );
  AOI21_X1 U19616 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n17483), .A(n17482), 
        .ZN(n17484) );
  AOI22_X1 U19617 ( .A1(n17499), .A2(n17485), .B1(n17484), .B2(n17497), .ZN(
        P2_U3605) );
  NAND2_X1 U19618 ( .A1(n19489), .A2(n19508), .ZN(n17486) );
  NAND2_X1 U19619 ( .A1(n17486), .A2(n18883), .ZN(n17496) );
  AOI222_X1 U19620 ( .A1(n17496), .A2(n17488), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19608), .C1(n19508), .C2(n17487), .ZN(n17489) );
  AOI22_X1 U19621 ( .A1(n17499), .A2(n17490), .B1(n17489), .B2(n17497), .ZN(
        P2_U3603) );
  AND2_X1 U19622 ( .A1(n19508), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17494) );
  INV_X1 U19623 ( .A(n17494), .ZN(n17491) );
  NAND2_X1 U19624 ( .A1(n19420), .A2(n17491), .ZN(n17492) );
  AOI22_X1 U19625 ( .A1(n17496), .A2(n17492), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19809), .ZN(n17493) );
  AOI22_X1 U19626 ( .A1(n17499), .A2(n19488), .B1(n17493), .B2(n17497), .ZN(
        P2_U3604) );
  INV_X1 U19627 ( .A(n19499), .ZN(n19509) );
  OAI21_X1 U19628 ( .B1(n19509), .B2(n19420), .A(n19455), .ZN(n17495) );
  AOI222_X1 U19629 ( .A1(n17496), .A2(n19614), .B1(n17495), .B2(n17494), .C1(
        n19712), .C2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U19630 ( .A1(n17499), .A2(n19432), .B1(n17498), .B2(n17497), .ZN(
        P2_U3602) );
  NAND2_X1 U19631 ( .A1(n17500), .A2(n21852), .ZN(n17504) );
  OAI21_X1 U19632 ( .B1(n17501), .B2(n18464), .A(n17508), .ZN(n17502) );
  OAI21_X1 U19633 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17508), .A(n17502), 
        .ZN(n17503) );
  OAI221_X1 U19634 ( .B1(n17504), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17504), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17503), .ZN(P2_U2822) );
  INV_X1 U19635 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17507) );
  OAI221_X1 U19636 ( .B1(n17508), .B2(n17507), .C1(n17506), .C2(n17505), .A(
        n17504), .ZN(P2_U2823) );
  OAI22_X1 U19637 ( .A1(n17572), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n21882), .ZN(n17509) );
  INV_X1 U19638 ( .A(n17509), .ZN(P2_U3611) );
  INV_X1 U19639 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17510) );
  AOI22_X1 U19640 ( .A1(n21882), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17510), 
        .B2(n17572), .ZN(P2_U3608) );
  AOI21_X1 U19641 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n21853), .ZN(n17511) );
  INV_X1 U19642 ( .A(n17511), .ZN(P2_U2815) );
  AOI22_X1 U19643 ( .A1(n17538), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17513) );
  OAI21_X1 U19644 ( .B1(n17514), .B2(n17540), .A(n17513), .ZN(P2_U2951) );
  INV_X1 U19645 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17516) );
  AOI22_X1 U19646 ( .A1(n17538), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17515) );
  OAI21_X1 U19647 ( .B1(n17516), .B2(n17540), .A(n17515), .ZN(P2_U2950) );
  INV_X1 U19648 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17518) );
  AOI22_X1 U19649 ( .A1(n17538), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17517) );
  OAI21_X1 U19650 ( .B1(n17518), .B2(n17540), .A(n17517), .ZN(P2_U2949) );
  INV_X1 U19651 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17520) );
  AOI22_X1 U19652 ( .A1(n17530), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17519) );
  OAI21_X1 U19653 ( .B1(n17520), .B2(n17540), .A(n17519), .ZN(P2_U2948) );
  INV_X1 U19654 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17522) );
  AOI22_X1 U19655 ( .A1(n17538), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U19656 ( .B1(n17522), .B2(n17540), .A(n17521), .ZN(P2_U2947) );
  INV_X1 U19657 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U19658 ( .A1(n17530), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17523) );
  OAI21_X1 U19659 ( .B1(n17524), .B2(n17540), .A(n17523), .ZN(P2_U2946) );
  INV_X1 U19660 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19557) );
  AOI22_X1 U19661 ( .A1(n17530), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17525) );
  OAI21_X1 U19662 ( .B1(n19557), .B2(n17540), .A(n17525), .ZN(P2_U2945) );
  INV_X1 U19663 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19395) );
  AOI22_X1 U19664 ( .A1(n17530), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17526) );
  OAI21_X1 U19665 ( .B1(n19395), .B2(n17540), .A(n17526), .ZN(P2_U2944) );
  INV_X1 U19666 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19392) );
  AOI22_X1 U19667 ( .A1(n17530), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17527) );
  OAI21_X1 U19668 ( .B1(n19392), .B2(n17540), .A(n17527), .ZN(P2_U2943) );
  INV_X1 U19669 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19388) );
  AOI22_X1 U19670 ( .A1(n17538), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17528) );
  OAI21_X1 U19671 ( .B1(n19388), .B2(n17540), .A(n17528), .ZN(P2_U2942) );
  AOI22_X1 U19672 ( .A1(n17530), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17531) );
  OAI21_X1 U19673 ( .B1(n17532), .B2(n17540), .A(n17531), .ZN(P2_U2941) );
  INV_X1 U19674 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19381) );
  AOI22_X1 U19675 ( .A1(n17538), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U19676 ( .B1(n19381), .B2(n17540), .A(n17533), .ZN(P2_U2940) );
  INV_X1 U19677 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19378) );
  AOI22_X1 U19678 ( .A1(n17538), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17534) );
  OAI21_X1 U19679 ( .B1(n19378), .B2(n17540), .A(n17534), .ZN(P2_U2939) );
  INV_X1 U19680 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19375) );
  AOI22_X1 U19681 ( .A1(n17538), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U19682 ( .B1(n19375), .B2(n17540), .A(n17535), .ZN(P2_U2938) );
  INV_X1 U19683 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19372) );
  AOI22_X1 U19684 ( .A1(n17538), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17536) );
  OAI21_X1 U19685 ( .B1(n19372), .B2(n17540), .A(n17536), .ZN(P2_U2937) );
  AOI22_X1 U19686 ( .A1(n17538), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17537), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17539) );
  OAI21_X1 U19687 ( .B1(n14281), .B2(n17540), .A(n17539), .ZN(P2_U2936) );
  INV_X1 U19688 ( .A(n17541), .ZN(n21884) );
  AOI22_X1 U19689 ( .A1(n21882), .A2(n17542), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n17572), .ZN(n17543) );
  OAI21_X1 U19690 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n21884), .A(n17543), 
        .ZN(P2_U2817) );
  NOR2_X2 U19691 ( .A1(n21890), .A2(n17572), .ZN(n21888) );
  INV_X1 U19692 ( .A(n17563), .ZN(n17569) );
  OAI222_X1 U19693 ( .A1(n17567), .A2(n18464), .B1(n17544), .B2(n21882), .C1(
        n14336), .C2(n17569), .ZN(P2_U3212) );
  AOI222_X1 U19694 ( .A1(n21888), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_3__SCAN_IN), 
        .C2(n17563), .ZN(n17545) );
  INV_X1 U19695 ( .A(n17545), .ZN(P2_U3213) );
  AOI222_X1 U19696 ( .A1(n21888), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_4__SCAN_IN), 
        .C2(n17563), .ZN(n17546) );
  INV_X1 U19697 ( .A(n17546), .ZN(P2_U3214) );
  AOI222_X1 U19698 ( .A1(n17563), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_4__SCAN_IN), 
        .C2(n21888), .ZN(n17547) );
  INV_X1 U19699 ( .A(n17547), .ZN(P2_U3215) );
  AOI222_X1 U19700 ( .A1(n17563), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_5__SCAN_IN), 
        .C2(n21888), .ZN(n17548) );
  INV_X1 U19701 ( .A(n17548), .ZN(P2_U3216) );
  AOI222_X1 U19702 ( .A1(n17563), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_6__SCAN_IN), 
        .C2(n21888), .ZN(n17549) );
  INV_X1 U19703 ( .A(n17549), .ZN(P2_U3217) );
  AOI222_X1 U19704 ( .A1(n17563), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_7__SCAN_IN), 
        .C2(n21888), .ZN(n17550) );
  INV_X1 U19705 ( .A(n17550), .ZN(P2_U3218) );
  INV_X1 U19706 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19994) );
  INV_X1 U19707 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n17551) );
  OAI222_X1 U19708 ( .A1(n17569), .A2(n13061), .B1(n19994), .B2(n21882), .C1(
        n17551), .C2(n17567), .ZN(P2_U3219) );
  INV_X1 U19709 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19996) );
  INV_X1 U19710 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n17552) );
  OAI222_X1 U19711 ( .A1(n17567), .A2(n13061), .B1(n19996), .B2(n21882), .C1(
        n17552), .C2(n17569), .ZN(P2_U3220) );
  INV_X1 U19712 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19998) );
  OAI222_X1 U19713 ( .A1(n17567), .A2(n17552), .B1(n19998), .B2(n21882), .C1(
        n13069), .C2(n17569), .ZN(P2_U3221) );
  INV_X1 U19714 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20000) );
  OAI222_X1 U19715 ( .A1(n17567), .A2(n13069), .B1(n20000), .B2(n21882), .C1(
        n13071), .C2(n17569), .ZN(P2_U3222) );
  AOI222_X1 U19716 ( .A1(n21888), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_ADDRESS_REG_11__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_13__SCAN_IN), 
        .C2(n17563), .ZN(n17553) );
  INV_X1 U19717 ( .A(n17553), .ZN(P2_U3223) );
  AOI222_X1 U19718 ( .A1(n21888), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_ADDRESS_REG_12__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_14__SCAN_IN), 
        .C2(n17563), .ZN(n17554) );
  INV_X1 U19719 ( .A(n17554), .ZN(P2_U3224) );
  AOI222_X1 U19720 ( .A1(n21888), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_ADDRESS_REG_13__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_15__SCAN_IN), 
        .C2(n17563), .ZN(n17555) );
  INV_X1 U19721 ( .A(n17555), .ZN(P2_U3225) );
  INV_X1 U19722 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20005) );
  OAI222_X1 U19723 ( .A1(n17567), .A2(n17556), .B1(n20005), .B2(n21882), .C1(
        n17557), .C2(n17569), .ZN(P2_U3226) );
  INV_X1 U19724 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20007) );
  OAI222_X1 U19725 ( .A1(n17567), .A2(n17557), .B1(n20007), .B2(n21882), .C1(
        n13091), .C2(n17569), .ZN(P2_U3227) );
  INV_X1 U19726 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20009) );
  OAI222_X1 U19727 ( .A1(n17567), .A2(n13091), .B1(n20009), .B2(n21882), .C1(
        n17558), .C2(n17569), .ZN(P2_U3228) );
  INV_X1 U19728 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20011) );
  OAI222_X1 U19729 ( .A1(n17569), .A2(n18647), .B1(n20011), .B2(n21882), .C1(
        n17558), .C2(n17567), .ZN(P2_U3229) );
  AOI222_X1 U19730 ( .A1(n21888), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_ADDRESS_REG_18__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_20__SCAN_IN), 
        .C2(n17563), .ZN(n17559) );
  INV_X1 U19731 ( .A(n17559), .ZN(P2_U3230) );
  AOI222_X1 U19732 ( .A1(n17563), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_ADDRESS_REG_19__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_20__SCAN_IN), 
        .C2(n21888), .ZN(n17560) );
  INV_X1 U19733 ( .A(n17560), .ZN(P2_U3231) );
  AOI222_X1 U19734 ( .A1(n17563), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_ADDRESS_REG_20__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_21__SCAN_IN), 
        .C2(n21888), .ZN(n17561) );
  INV_X1 U19735 ( .A(n17561), .ZN(P2_U3232) );
  AOI222_X1 U19736 ( .A1(n17563), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_ADDRESS_REG_21__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_22__SCAN_IN), 
        .C2(n21888), .ZN(n17562) );
  INV_X1 U19737 ( .A(n17562), .ZN(P2_U3233) );
  AOI222_X1 U19738 ( .A1(n17563), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_ADDRESS_REG_22__SCAN_IN), .B2(n17572), .C1(P2_REIP_REG_23__SCAN_IN), 
        .C2(n21888), .ZN(n17564) );
  INV_X1 U19739 ( .A(n17564), .ZN(P2_U3234) );
  INV_X1 U19740 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20019) );
  OAI222_X1 U19741 ( .A1(n17569), .A2(n18717), .B1(n20019), .B2(n21882), .C1(
        n17565), .C2(n17567), .ZN(P2_U3235) );
  INV_X1 U19742 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20021) );
  OAI222_X1 U19743 ( .A1(n17567), .A2(n18717), .B1(n20021), .B2(n21882), .C1(
        n17566), .C2(n17569), .ZN(P2_U3236) );
  INV_X1 U19744 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20023) );
  OAI222_X1 U19745 ( .A1(n17569), .A2(n18739), .B1(n20023), .B2(n21882), .C1(
        n17566), .C2(n17567), .ZN(P2_U3237) );
  INV_X1 U19746 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20025) );
  OAI222_X1 U19747 ( .A1(n17567), .A2(n18739), .B1(n20025), .B2(n21882), .C1(
        n13130), .C2(n17569), .ZN(P2_U3238) );
  INV_X1 U19748 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20027) );
  OAI222_X1 U19749 ( .A1(n17567), .A2(n13130), .B1(n20027), .B2(n21882), .C1(
        n18764), .C2(n17569), .ZN(P2_U3239) );
  INV_X1 U19750 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20030) );
  OAI222_X1 U19751 ( .A1(n17567), .A2(n18764), .B1(n20030), .B2(n21882), .C1(
        n18790), .C2(n17569), .ZN(P2_U3240) );
  INV_X1 U19752 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20032) );
  OAI222_X1 U19753 ( .A1(n17569), .A2(n17568), .B1(n20032), .B2(n21882), .C1(
        n18790), .C2(n17567), .ZN(P2_U3241) );
  OAI22_X1 U19754 ( .A1(n17572), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n21882), .ZN(n17570) );
  INV_X1 U19755 ( .A(n17570), .ZN(P2_U3588) );
  OAI22_X1 U19756 ( .A1(n17572), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n21882), .ZN(n17571) );
  INV_X1 U19757 ( .A(n17571), .ZN(P2_U3587) );
  MUX2_X1 U19758 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n17572), .Z(P2_U3586) );
  OAI22_X1 U19759 ( .A1(n17572), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n21882), .ZN(n17573) );
  INV_X1 U19760 ( .A(n17573), .ZN(P2_U3585) );
  INV_X1 U19761 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17967) );
  INV_X1 U19762 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20372) );
  NOR3_X1 U19763 ( .A1(n20388), .A2(n17967), .A3(n20372), .ZN(n17579) );
  NAND3_X1 U19764 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17579), .ZN(n17608) );
  INV_X1 U19765 ( .A(n17608), .ZN(n17600) );
  NOR2_X1 U19766 ( .A1(n21385), .A2(n17574), .ZN(n17578) );
  NOR3_X1 U19767 ( .A1(n20809), .A2(n17576), .A3(n17575), .ZN(n17577) );
  NOR3_X1 U19768 ( .A1(n19220), .A2(n20370), .A3(n20777), .ZN(n17968) );
  NOR2_X1 U19769 ( .A1(n20809), .A2(n17962), .ZN(n17964) );
  AND2_X1 U19770 ( .A1(n17600), .A2(n17964), .ZN(n17605) );
  NAND2_X1 U19771 ( .A1(n17579), .A2(n17964), .ZN(n17583) );
  INV_X1 U19772 ( .A(n17583), .ZN(n17585) );
  AOI22_X1 U19773 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17935), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(n17585), .ZN(n17580) );
  OAI22_X1 U19774 ( .A1(n17605), .A2(n17580), .B1(n17891), .B2(n17935), .ZN(
        P3_U2699) );
  NAND3_X1 U19775 ( .A1(n17583), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17935), .ZN(
        n17581) );
  OAI221_X1 U19776 ( .B1(n17583), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17935), 
        .C2(n17582), .A(n17581), .ZN(P3_U2700) );
  NOR2_X1 U19777 ( .A1(n17967), .A2(n20372), .ZN(n17584) );
  AOI21_X1 U19778 ( .B1(n17968), .B2(n17584), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17586) );
  AOI221_X1 U19779 ( .B1(n17586), .B2(n17935), .C1(n17905), .C2(n17965), .A(
        n17585), .ZN(P3_U2701) );
  NAND4_X1 U19780 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n17600), .ZN(n17720) );
  NOR3_X1 U19781 ( .A1(n20470), .A2(n17962), .A3(n17720), .ZN(n17715) );
  NOR2_X1 U19782 ( .A1(n17962), .A2(n17720), .ZN(n17601) );
  OAI21_X1 U19783 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17601), .A(n17935), .ZN(
        n17599) );
  AOI22_X1 U19784 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17597) );
  AOI22_X1 U19785 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17596) );
  AOI22_X1 U19786 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17587) );
  OAI21_X1 U19787 ( .B1(n17690), .B2(n17770), .A(n17587), .ZN(n17594) );
  AOI22_X1 U19788 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17592) );
  AOI22_X1 U19789 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17591) );
  AOI22_X1 U19790 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17590) );
  AOI22_X1 U19791 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17589) );
  NAND4_X1 U19792 ( .A1(n17592), .A2(n17591), .A3(n17590), .A4(n17589), .ZN(
        n17593) );
  AOI211_X1 U19793 ( .C1(n17803), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17594), .B(n17593), .ZN(n17595) );
  NAND3_X1 U19794 ( .A1(n17597), .A2(n17596), .A3(n17595), .ZN(n20960) );
  INV_X1 U19795 ( .A(n20960), .ZN(n17598) );
  OAI22_X1 U19796 ( .A1(n17715), .A2(n17599), .B1(n17598), .B2(n17935), .ZN(
        P3_U2695) );
  NAND3_X1 U19797 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17968), .A3(n17600), .ZN(
        n17609) );
  NOR2_X1 U19798 ( .A1(n20446), .A2(n17609), .ZN(n17603) );
  INV_X1 U19799 ( .A(n17601), .ZN(n17602) );
  OAI221_X1 U19800 ( .B1(n17603), .B2(P3_EBX_REG_7__SCAN_IN), .C1(n20959), 
        .C2(n17962), .A(n17602), .ZN(n17604) );
  OAI21_X1 U19801 ( .B1(n17782), .B2(n17935), .A(n17604), .ZN(P3_U2696) );
  NAND3_X1 U19802 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17935), .A3(n17609), .ZN(
        n17607) );
  NAND3_X1 U19803 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17605), .A3(n20446), .ZN(
        n17606) );
  OAI211_X1 U19804 ( .C1(n17935), .C2(n17815), .A(n17607), .B(n17606), .ZN(
        P3_U2697) );
  INV_X1 U19805 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17830) );
  NOR2_X1 U19806 ( .A1(n17962), .A2(n17608), .ZN(n17610) );
  OAI211_X1 U19807 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17610), .A(n17609), .B(
        n17935), .ZN(n17611) );
  OAI21_X1 U19808 ( .B1(n17935), .B2(n17830), .A(n17611), .ZN(P3_U2698) );
  NAND3_X1 U19809 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .ZN(n17719) );
  NAND2_X1 U19810 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17715), .ZN(n17714) );
  NAND2_X1 U19811 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17702), .ZN(n17687) );
  NAND2_X1 U19812 ( .A1(n20959), .A2(n17637), .ZN(n17661) );
  OR2_X1 U19813 ( .A1(n17719), .A2(n17661), .ZN(n17623) );
  AOI22_X1 U19814 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17615) );
  AOI22_X1 U19815 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U19816 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17613) );
  AOI22_X1 U19817 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17612) );
  NAND4_X1 U19818 ( .A1(n17615), .A2(n17614), .A3(n17613), .A4(n17612), .ZN(
        n17621) );
  AOI22_X1 U19819 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17619) );
  AOI22_X1 U19820 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17618) );
  AOI22_X1 U19821 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17617) );
  AOI22_X1 U19822 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17616) );
  NAND4_X1 U19823 ( .A1(n17619), .A2(n17618), .A3(n17617), .A4(n17616), .ZN(
        n17620) );
  NOR2_X1 U19824 ( .A1(n17621), .A2(n17620), .ZN(n20945) );
  NAND3_X1 U19825 ( .A1(n17623), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17935), 
        .ZN(n17622) );
  OAI221_X1 U19826 ( .B1(n17623), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17935), 
        .C2(n20945), .A(n17622), .ZN(P3_U2687) );
  INV_X1 U19827 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17662) );
  NOR2_X1 U19828 ( .A1(n20562), .A2(n17662), .ZN(n17624) );
  AOI21_X1 U19829 ( .B1(n17624), .B2(n17637), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n17636) );
  OAI21_X1 U19830 ( .B1(n17719), .B2(n17661), .A(n17935), .ZN(n17635) );
  AOI22_X1 U19831 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17628) );
  AOI22_X1 U19832 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17627) );
  AOI22_X1 U19833 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17626) );
  AOI22_X1 U19834 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17625) );
  NAND4_X1 U19835 ( .A1(n17628), .A2(n17627), .A3(n17626), .A4(n17625), .ZN(
        n17634) );
  AOI22_X1 U19836 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11537), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17632) );
  AOI22_X1 U19837 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17631) );
  AOI22_X1 U19838 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17630) );
  AOI22_X1 U19839 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17629) );
  NAND4_X1 U19840 ( .A1(n17632), .A2(n17631), .A3(n17630), .A4(n17629), .ZN(
        n17633) );
  NOR2_X1 U19841 ( .A1(n17634), .A2(n17633), .ZN(n20957) );
  OAI22_X1 U19842 ( .A1(n17636), .A2(n17635), .B1(n20957), .B2(n17935), .ZN(
        P3_U2688) );
  INV_X1 U19843 ( .A(n17637), .ZN(n17660) );
  NAND2_X1 U19844 ( .A1(n17935), .A2(n17660), .ZN(n17676) );
  AOI22_X1 U19845 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17647) );
  AOI22_X1 U19846 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17646) );
  AOI22_X1 U19847 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17638) );
  OAI21_X1 U19848 ( .B1(n17690), .B2(n17830), .A(n17638), .ZN(n17644) );
  AOI22_X1 U19849 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17642) );
  AOI22_X1 U19850 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17641) );
  AOI22_X1 U19851 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17640) );
  AOI22_X1 U19852 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17639) );
  NAND4_X1 U19853 ( .A1(n17642), .A2(n17641), .A3(n17640), .A4(n17639), .ZN(
        n17643) );
  AOI211_X1 U19854 ( .C1(n10992), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n17644), .B(n17643), .ZN(n17645) );
  NAND3_X1 U19855 ( .A1(n17647), .A2(n17646), .A3(n17645), .ZN(n20788) );
  NAND2_X1 U19856 ( .A1(n17965), .A2(n20788), .ZN(n17648) );
  OAI221_X1 U19857 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17661), .C1(n17662), 
        .C2(n17676), .A(n17648), .ZN(P3_U2690) );
  AOI22_X1 U19858 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17653) );
  AOI22_X1 U19859 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11621), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17652) );
  AOI22_X1 U19860 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17651) );
  AOI22_X1 U19861 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17650) );
  NAND4_X1 U19862 ( .A1(n17653), .A2(n17652), .A3(n17651), .A4(n17650), .ZN(
        n17659) );
  AOI22_X1 U19863 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17881), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17657) );
  AOI22_X1 U19864 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17656) );
  AOI22_X1 U19865 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17655) );
  AOI22_X1 U19866 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17771), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17654) );
  NAND4_X1 U19867 ( .A1(n17657), .A2(n17656), .A3(n17655), .A4(n17654), .ZN(
        n17658) );
  NOR2_X1 U19868 ( .A1(n17659), .A2(n17658), .ZN(n20951) );
  OAI211_X1 U19869 ( .C1(n17662), .C2(n17660), .A(P3_EBX_REG_14__SCAN_IN), .B(
        n17935), .ZN(n17664) );
  OR3_X1 U19870 ( .A1(n17662), .A2(n17661), .A3(P3_EBX_REG_14__SCAN_IN), .ZN(
        n17663) );
  OAI211_X1 U19871 ( .C1(n20951), .C2(n17935), .A(n17664), .B(n17663), .ZN(
        P3_U2689) );
  AOI22_X1 U19872 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17674) );
  AOI22_X1 U19873 ( .A1(n17771), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17673) );
  AOI22_X1 U19874 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17665) );
  OAI21_X1 U19875 ( .B1(n17690), .B2(n17891), .A(n17665), .ZN(n17671) );
  AOI22_X1 U19876 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10992), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17669) );
  AOI22_X1 U19877 ( .A1(n17951), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11621), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17668) );
  AOI22_X1 U19878 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17667) );
  AOI22_X1 U19879 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17666) );
  NAND4_X1 U19880 ( .A1(n17669), .A2(n17668), .A3(n17667), .A4(n17666), .ZN(
        n17670) );
  AOI211_X1 U19881 ( .C1(n10996), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n17671), .B(n17670), .ZN(n17672) );
  NAND3_X1 U19882 ( .A1(n17674), .A2(n17673), .A3(n17672), .ZN(n20792) );
  NAND2_X1 U19883 ( .A1(n17965), .A2(n20792), .ZN(n17675) );
  OAI221_X1 U19884 ( .B1(n17676), .B2(n20530), .C1(n17676), .C2(n17687), .A(
        n17675), .ZN(P3_U2691) );
  AOI22_X1 U19885 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11621), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17680) );
  AOI22_X1 U19886 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17679) );
  AOI22_X1 U19887 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17678) );
  AOI22_X1 U19888 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17677) );
  NAND4_X1 U19889 ( .A1(n17680), .A2(n17679), .A3(n17678), .A4(n17677), .ZN(
        n17686) );
  AOI22_X1 U19890 ( .A1(n17951), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17684) );
  AOI22_X1 U19891 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17683) );
  AOI22_X1 U19892 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17771), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17682) );
  AOI22_X1 U19893 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17681) );
  NAND4_X1 U19894 ( .A1(n17684), .A2(n17683), .A3(n17682), .A4(n17681), .ZN(
        n17685) );
  NOR2_X1 U19895 ( .A1(n17686), .A2(n17685), .ZN(n20796) );
  OAI21_X1 U19896 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17702), .A(n17687), .ZN(
        n17688) );
  AOI22_X1 U19897 ( .A1(n17965), .A2(n20796), .B1(n17688), .B2(n17935), .ZN(
        P3_U2692) );
  AOI22_X1 U19898 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17699) );
  AOI22_X1 U19899 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17698) );
  AOI22_X1 U19900 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17689) );
  OAI21_X1 U19901 ( .B1(n17690), .B2(n17905), .A(n17689), .ZN(n17696) );
  AOI22_X1 U19902 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17771), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17694) );
  AOI22_X1 U19903 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11621), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17693) );
  AOI22_X1 U19904 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17692) );
  AOI22_X1 U19905 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17691) );
  NAND4_X1 U19906 ( .A1(n17694), .A2(n17693), .A3(n17692), .A4(n17691), .ZN(
        n17695) );
  AOI211_X1 U19907 ( .C1(n17951), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n17696), .B(n17695), .ZN(n17697) );
  NAND3_X1 U19908 ( .A1(n17699), .A2(n17698), .A3(n17697), .ZN(n20800) );
  INV_X1 U19909 ( .A(n20800), .ZN(n17703) );
  INV_X1 U19910 ( .A(n17714), .ZN(n17700) );
  OAI21_X1 U19911 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17700), .A(n17935), .ZN(
        n17701) );
  OAI22_X1 U19912 ( .A1(n17703), .A2(n17935), .B1(n17702), .B2(n17701), .ZN(
        P3_U2693) );
  AOI22_X1 U19913 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17927), .B1(
        n17771), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17707) );
  AOI22_X1 U19914 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17881), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U19915 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17942), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17943), .ZN(n17705) );
  AOI22_X1 U19916 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11632), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17941), .ZN(n17704) );
  NAND4_X1 U19917 ( .A1(n17707), .A2(n17706), .A3(n17705), .A4(n17704), .ZN(
        n17713) );
  AOI22_X1 U19918 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17950), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17711) );
  AOI22_X1 U19919 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17803), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17710) );
  AOI22_X1 U19920 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17949), .ZN(n17709) );
  AOI22_X1 U19921 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17708) );
  NAND4_X1 U19922 ( .A1(n17711), .A2(n17710), .A3(n17709), .A4(n17708), .ZN(
        n17712) );
  NOR2_X1 U19923 ( .A1(n17713), .A2(n17712), .ZN(n20805) );
  OAI21_X1 U19924 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17715), .A(n17714), .ZN(
        n17716) );
  AOI22_X1 U19925 ( .A1(n17965), .A2(n20805), .B1(n17716), .B2(n17935), .ZN(
        P3_U2694) );
  INV_X1 U19926 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20737) );
  INV_X1 U19927 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20685) );
  NOR4_X1 U19928 ( .A1(n20737), .A2(n20701), .A3(n20685), .A4(n20677), .ZN(
        n17722) );
  INV_X1 U19929 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n20708) );
  INV_X1 U19930 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20635) );
  INV_X1 U19931 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20608) );
  NOR3_X1 U19932 ( .A1(n20592), .A2(n20530), .A3(n20493), .ZN(n17717) );
  NAND4_X1 U19933 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(n17717), .ZN(n17718) );
  NOR3_X1 U19934 ( .A1(n17720), .A2(n17719), .A3(n17718), .ZN(n17959) );
  NAND2_X1 U19935 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17959), .ZN(n17958) );
  NAND2_X1 U19936 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17918), .ZN(n17921) );
  NAND2_X1 U19937 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17937), .ZN(n17840) );
  NOR4_X1 U19938 ( .A1(n20728), .A2(n20708), .A3(n20635), .A4(n17840), .ZN(
        n17721) );
  NAND4_X1 U19939 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17722), .A4(n17721), .ZN(n17725) );
  NOR2_X1 U19940 ( .A1(n20747), .A2(n17725), .ZN(n17828) );
  NAND2_X1 U19941 ( .A1(n17935), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17724) );
  NAND2_X1 U19942 ( .A1(n17828), .A2(n20959), .ZN(n17723) );
  OAI22_X1 U19943 ( .A1(n17828), .A2(n17724), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17723), .ZN(P3_U2672) );
  NAND2_X1 U19944 ( .A1(n20747), .A2(n17725), .ZN(n17726) );
  NAND2_X1 U19945 ( .A1(n17726), .A2(n17935), .ZN(n17827) );
  AOI22_X1 U19946 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17731) );
  AOI22_X1 U19947 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17771), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17730) );
  AOI22_X1 U19948 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17729) );
  AOI22_X1 U19949 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17728) );
  NAND4_X1 U19950 ( .A1(n17731), .A2(n17730), .A3(n17729), .A4(n17728), .ZN(
        n17738) );
  AOI22_X1 U19951 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17736) );
  AOI22_X1 U19952 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17881), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17735) );
  AOI22_X1 U19953 ( .A1(n17949), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17734) );
  AOI22_X1 U19954 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17733) );
  NAND4_X1 U19955 ( .A1(n17736), .A2(n17735), .A3(n17734), .A4(n17733), .ZN(
        n17737) );
  NOR2_X1 U19956 ( .A1(n17738), .A2(n17737), .ZN(n17826) );
  AOI22_X1 U19957 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17742) );
  AOI22_X1 U19958 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17741) );
  AOI22_X1 U19959 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17740) );
  AOI22_X1 U19960 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17739) );
  NAND4_X1 U19961 ( .A1(n17742), .A2(n17741), .A3(n17740), .A4(n17739), .ZN(
        n17748) );
  AOI22_X1 U19962 ( .A1(n11547), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U19963 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17771), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17745) );
  AOI22_X1 U19964 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17744) );
  AOI22_X1 U19965 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17743) );
  NAND4_X1 U19966 ( .A1(n17746), .A2(n17745), .A3(n17744), .A4(n17743), .ZN(
        n17747) );
  NOR2_X1 U19967 ( .A1(n17748), .A2(n17747), .ZN(n17851) );
  AOI22_X1 U19968 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17752) );
  AOI22_X1 U19969 ( .A1(n17951), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17771), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U19970 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17750) );
  AOI22_X1 U19971 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17749) );
  NAND4_X1 U19972 ( .A1(n17752), .A2(n17751), .A3(n17750), .A4(n17749), .ZN(
        n17758) );
  AOI22_X1 U19973 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17756) );
  AOI22_X1 U19974 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17755) );
  AOI22_X1 U19975 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17754) );
  AOI22_X1 U19976 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17753) );
  NAND4_X1 U19977 ( .A1(n17756), .A2(n17755), .A3(n17754), .A4(n17753), .ZN(
        n17757) );
  NOR2_X1 U19978 ( .A1(n17758), .A2(n17757), .ZN(n17857) );
  AOI22_X1 U19979 ( .A1(n17771), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n11547), .ZN(n17762) );
  AOI22_X1 U19980 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17927), .ZN(n17761) );
  AOI22_X1 U19981 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17942), .ZN(n17760) );
  AOI22_X1 U19982 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17943), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17759) );
  NAND4_X1 U19983 ( .A1(n17762), .A2(n17761), .A3(n17760), .A4(n17759), .ZN(
        n17768) );
  AOI22_X1 U19984 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17928), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17766) );
  AOI22_X1 U19985 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17949), .B1(
        n17783), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17765) );
  AOI22_X1 U19986 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17938), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17764) );
  AOI22_X1 U19987 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17763) );
  NAND4_X1 U19988 ( .A1(n17766), .A2(n17765), .A3(n17764), .A4(n17763), .ZN(
        n17767) );
  NOR2_X1 U19989 ( .A1(n17768), .A2(n17767), .ZN(n17867) );
  AOI22_X1 U19990 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17780) );
  AOI22_X1 U19991 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17779) );
  AOI22_X1 U19992 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17769) );
  OAI21_X1 U19993 ( .B1(n17816), .B2(n17770), .A(n17769), .ZN(n17777) );
  AOI22_X1 U19994 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17775) );
  AOI22_X1 U19995 ( .A1(n17771), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17774) );
  AOI22_X1 U19996 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17773) );
  AOI22_X1 U19997 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17772) );
  NAND4_X1 U19998 ( .A1(n17775), .A2(n17774), .A3(n17773), .A4(n17772), .ZN(
        n17776) );
  AOI211_X1 U19999 ( .C1(n17914), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17777), .B(n17776), .ZN(n17778) );
  NAND3_X1 U20000 ( .A1(n17780), .A2(n17779), .A3(n17778), .ZN(n17873) );
  AOI22_X1 U20001 ( .A1(n11547), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17792) );
  AOI22_X1 U20002 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17791) );
  AOI22_X1 U20003 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17781) );
  OAI21_X1 U20004 ( .B1(n17906), .B2(n17782), .A(n17781), .ZN(n17789) );
  AOI22_X1 U20005 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17783), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U20006 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17786) );
  AOI22_X1 U20007 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17785) );
  AOI22_X1 U20008 ( .A1(n17943), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17784) );
  NAND4_X1 U20009 ( .A1(n17787), .A2(n17786), .A3(n17785), .A4(n17784), .ZN(
        n17788) );
  AOI211_X1 U20010 ( .C1(n10996), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n17789), .B(n17788), .ZN(n17790) );
  NAND3_X1 U20011 ( .A1(n17792), .A2(n17791), .A3(n17790), .ZN(n17874) );
  NAND2_X1 U20012 ( .A1(n17873), .A2(n17874), .ZN(n17872) );
  NOR2_X1 U20013 ( .A1(n17867), .A2(n17872), .ZN(n17866) );
  AOI22_X1 U20014 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17802) );
  AOI22_X1 U20015 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17801) );
  AOI22_X1 U20016 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17793) );
  OAI21_X1 U20017 ( .B1(n17816), .B2(n17905), .A(n17793), .ZN(n17799) );
  AOI22_X1 U20018 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17797) );
  AOI22_X1 U20019 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17796) );
  AOI22_X1 U20020 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17795) );
  AOI22_X1 U20021 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17794) );
  NAND4_X1 U20022 ( .A1(n17797), .A2(n17796), .A3(n17795), .A4(n17794), .ZN(
        n17798) );
  AOI211_X1 U20023 ( .C1(n17914), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17799), .B(n17798), .ZN(n17800) );
  NAND3_X1 U20024 ( .A1(n17802), .A2(n17801), .A3(n17800), .ZN(n17862) );
  NAND2_X1 U20025 ( .A1(n17866), .A2(n17862), .ZN(n17861) );
  NOR2_X1 U20026 ( .A1(n17857), .A2(n17861), .ZN(n17856) );
  AOI22_X1 U20027 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10992), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17813) );
  AOI22_X1 U20028 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17812) );
  AOI22_X1 U20029 ( .A1(n17949), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17804) );
  OAI21_X1 U20030 ( .B1(n17816), .B2(n17891), .A(n17804), .ZN(n17810) );
  AOI22_X1 U20031 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17808) );
  AOI22_X1 U20032 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17807) );
  AOI22_X1 U20033 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17943), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17806) );
  AOI22_X1 U20034 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17805) );
  NAND4_X1 U20035 ( .A1(n17808), .A2(n17807), .A3(n17806), .A4(n17805), .ZN(
        n17809) );
  AOI211_X1 U20036 ( .C1(n17783), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17810), .B(n17809), .ZN(n17811) );
  NAND3_X1 U20037 ( .A1(n17813), .A2(n17812), .A3(n17811), .ZN(n17842) );
  NAND2_X1 U20038 ( .A1(n17856), .A2(n17842), .ZN(n17850) );
  NOR2_X1 U20039 ( .A1(n17851), .A2(n17850), .ZN(n17849) );
  AOI22_X1 U20040 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U20041 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17824) );
  AOI22_X1 U20042 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17928), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17814) );
  OAI21_X1 U20043 ( .B1(n17816), .B2(n17815), .A(n17814), .ZN(n17822) );
  AOI22_X1 U20044 ( .A1(n17949), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17820) );
  AOI22_X1 U20045 ( .A1(n17939), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17819) );
  AOI22_X1 U20046 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17818) );
  AOI22_X1 U20047 ( .A1(n17943), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17817) );
  NAND4_X1 U20048 ( .A1(n17820), .A2(n17819), .A3(n17818), .A4(n17817), .ZN(
        n17821) );
  AOI211_X1 U20049 ( .C1(n17783), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17822), .B(n17821), .ZN(n17823) );
  NAND3_X1 U20050 ( .A1(n17825), .A2(n17824), .A3(n17823), .ZN(n17846) );
  NAND2_X1 U20051 ( .A1(n17849), .A2(n17846), .ZN(n17845) );
  XNOR2_X1 U20052 ( .A(n17826), .B(n17845), .ZN(n20899) );
  OAI22_X1 U20053 ( .A1(n17828), .A2(n17827), .B1(n20899), .B2(n17935), .ZN(
        P3_U2673) );
  NAND2_X1 U20054 ( .A1(n17935), .A2(n17840), .ZN(n17901) );
  AOI22_X1 U20055 ( .A1(n11537), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11621), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17839) );
  AOI22_X1 U20056 ( .A1(n17914), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17838) );
  AOI22_X1 U20057 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17829) );
  OAI21_X1 U20058 ( .B1(n17906), .B2(n17830), .A(n17829), .ZN(n17836) );
  AOI22_X1 U20059 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17834) );
  AOI22_X1 U20060 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U20061 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17943), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17832) );
  AOI22_X1 U20062 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17831) );
  NAND4_X1 U20063 ( .A1(n17834), .A2(n17833), .A3(n17832), .A4(n17831), .ZN(
        n17835) );
  AOI211_X1 U20064 ( .C1(n17783), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n17836), .B(n17835), .ZN(n17837) );
  NAND3_X1 U20065 ( .A1(n17839), .A2(n17838), .A3(n17837), .ZN(n20842) );
  NOR2_X1 U20066 ( .A1(n20809), .A2(n17840), .ZN(n17843) );
  AOI22_X1 U20067 ( .A1(n17965), .A2(n20842), .B1(n17843), .B2(n20635), .ZN(
        n17841) );
  OAI21_X1 U20068 ( .B1(n20635), .B2(n17901), .A(n17841), .ZN(P3_U2682) );
  OAI21_X1 U20069 ( .B1(n17856), .B2(n17842), .A(n17850), .ZN(n20919) );
  NAND2_X1 U20070 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17843), .ZN(n17889) );
  NAND2_X1 U20071 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17871), .ZN(n17865) );
  NAND2_X1 U20072 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17870), .ZN(n17855) );
  NAND2_X1 U20073 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17860), .ZN(n17854) );
  OAI211_X1 U20074 ( .C1(n17860), .C2(P3_EBX_REG_27__SCAN_IN), .A(n17935), .B(
        n17854), .ZN(n17844) );
  OAI21_X1 U20075 ( .B1(n17935), .B2(n20919), .A(n17844), .ZN(P3_U2676) );
  NAND3_X1 U20076 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17860), .ZN(n17848) );
  OAI21_X1 U20077 ( .B1(n17849), .B2(n17846), .A(n17845), .ZN(n20908) );
  NAND3_X1 U20078 ( .A1(n17848), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17935), 
        .ZN(n17847) );
  OAI221_X1 U20079 ( .B1(n17848), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17935), 
        .C2(n20908), .A(n17847), .ZN(P3_U2674) );
  AND2_X1 U20080 ( .A1(n17935), .A2(n17848), .ZN(n17852) );
  AOI21_X1 U20081 ( .B1(n17851), .B2(n17850), .A(n17849), .ZN(n20909) );
  AOI22_X1 U20082 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17852), .B1(n20909), 
        .B2(n17965), .ZN(n17853) );
  OAI21_X1 U20083 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17854), .A(n17853), .ZN(
        P3_U2675) );
  INV_X1 U20084 ( .A(n17855), .ZN(n17864) );
  AOI21_X1 U20085 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17935), .A(n17864), .ZN(
        n17859) );
  AOI21_X1 U20086 ( .B1(n17857), .B2(n17861), .A(n17856), .ZN(n20890) );
  INV_X1 U20087 ( .A(n20890), .ZN(n17858) );
  OAI22_X1 U20088 ( .A1(n17860), .A2(n17859), .B1(n17858), .B2(n17935), .ZN(
        P3_U2677) );
  AOI21_X1 U20089 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17935), .A(n17870), .ZN(
        n17863) );
  OAI21_X1 U20090 ( .B1(n17866), .B2(n17862), .A(n17861), .ZN(n20889) );
  OAI22_X1 U20091 ( .A1(n17864), .A2(n17863), .B1(n20889), .B2(n17935), .ZN(
        P3_U2678) );
  INV_X1 U20092 ( .A(n17865), .ZN(n17876) );
  AOI21_X1 U20093 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17935), .A(n17876), .ZN(
        n17869) );
  AOI21_X1 U20094 ( .B1(n17867), .B2(n17872), .A(n17866), .ZN(n20920) );
  INV_X1 U20095 ( .A(n20920), .ZN(n17868) );
  OAI22_X1 U20096 ( .A1(n17870), .A2(n17869), .B1(n17935), .B2(n17868), .ZN(
        P3_U2679) );
  AOI21_X1 U20097 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17935), .A(n17871), .ZN(
        n17875) );
  OAI21_X1 U20098 ( .B1(n17874), .B2(n17873), .A(n17872), .ZN(n20932) );
  OAI22_X1 U20099 ( .A1(n17876), .A2(n17875), .B1(n17935), .B2(n20932), .ZN(
        P3_U2680) );
  AOI22_X1 U20100 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17880) );
  AOI22_X1 U20101 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17879) );
  AOI22_X1 U20102 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17878) );
  AOI22_X1 U20103 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17943), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17877) );
  NAND4_X1 U20104 ( .A1(n17880), .A2(n17879), .A3(n17878), .A4(n17877), .ZN(
        n17887) );
  AOI22_X1 U20105 ( .A1(n17881), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17885) );
  AOI22_X1 U20106 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17884) );
  AOI22_X1 U20107 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17883) );
  AOI22_X1 U20108 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17882) );
  NAND4_X1 U20109 ( .A1(n17885), .A2(n17884), .A3(n17883), .A4(n17882), .ZN(
        n17886) );
  NOR2_X1 U20110 ( .A1(n17887), .A2(n17886), .ZN(n20854) );
  NAND3_X1 U20111 ( .A1(n17889), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17935), 
        .ZN(n17888) );
  OAI221_X1 U20112 ( .B1(n17889), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17935), 
        .C2(n20854), .A(n17888), .ZN(P3_U2681) );
  AOI22_X1 U20113 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11654), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17900) );
  AOI22_X1 U20114 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17899) );
  AOI22_X1 U20115 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17890) );
  OAI21_X1 U20116 ( .B1(n17906), .B2(n17891), .A(n17890), .ZN(n17897) );
  AOI22_X1 U20117 ( .A1(n17951), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17895) );
  AOI22_X1 U20118 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17894) );
  AOI22_X1 U20119 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17727), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17893) );
  AOI22_X1 U20120 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17892) );
  NAND4_X1 U20121 ( .A1(n17895), .A2(n17894), .A3(n17893), .A4(n17892), .ZN(
        n17896) );
  AOI211_X1 U20122 ( .C1(n10992), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n17897), .B(n17896), .ZN(n17898) );
  NAND3_X1 U20123 ( .A1(n17900), .A2(n17899), .A3(n17898), .ZN(n20849) );
  INV_X1 U20124 ( .A(n20849), .ZN(n17903) );
  NOR2_X1 U20125 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17937), .ZN(n17902) );
  OAI22_X1 U20126 ( .A1(n17903), .A2(n17935), .B1(n17902), .B2(n17901), .ZN(
        P3_U2683) );
  AOI22_X1 U20127 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17917) );
  AOI22_X1 U20128 ( .A1(n17951), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17927), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17916) );
  AOI22_X1 U20129 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17904) );
  OAI21_X1 U20130 ( .B1(n17906), .B2(n17905), .A(n17904), .ZN(n17913) );
  AOI22_X1 U20131 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17907), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17911) );
  AOI22_X1 U20132 ( .A1(n17803), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17910) );
  AOI22_X1 U20133 ( .A1(n21008), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17942), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17909) );
  AOI22_X1 U20134 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17941), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17908) );
  NAND4_X1 U20135 ( .A1(n17911), .A2(n17910), .A3(n17909), .A4(n17908), .ZN(
        n17912) );
  AOI211_X1 U20136 ( .C1(n17914), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17913), .B(n17912), .ZN(n17915) );
  NAND3_X1 U20137 ( .A1(n17917), .A2(n17916), .A3(n17915), .ZN(n20871) );
  INV_X1 U20138 ( .A(n20871), .ZN(n17920) );
  OAI21_X1 U20139 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17918), .A(n17921), .ZN(
        n17919) );
  AOI22_X1 U20140 ( .A1(n17965), .A2(n17920), .B1(n17919), .B2(n17935), .ZN(
        P3_U2685) );
  AOI21_X1 U20141 ( .B1(n20608), .B2(n17921), .A(n17965), .ZN(n17922) );
  INV_X1 U20142 ( .A(n17922), .ZN(n17936) );
  AOI22_X1 U20143 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17926) );
  AOI22_X1 U20144 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17925) );
  AOI22_X1 U20145 ( .A1(n11632), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17942), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17924) );
  AOI22_X1 U20146 ( .A1(n17941), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n21008), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17923) );
  NAND4_X1 U20147 ( .A1(n17926), .A2(n17925), .A3(n17924), .A4(n17923), .ZN(
        n17934) );
  AOI22_X1 U20148 ( .A1(n17938), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17927), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17932) );
  AOI22_X1 U20149 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11537), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17931) );
  AOI22_X1 U20150 ( .A1(n17950), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11547), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17930) );
  AOI22_X1 U20151 ( .A1(n17928), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17949), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17929) );
  NAND4_X1 U20152 ( .A1(n17932), .A2(n17931), .A3(n17930), .A4(n17929), .ZN(
        n17933) );
  NOR2_X1 U20153 ( .A1(n17934), .A2(n17933), .ZN(n20870) );
  OAI22_X1 U20154 ( .A1(n17937), .A2(n17936), .B1(n20870), .B2(n17935), .ZN(
        P3_U2684) );
  AOI22_X1 U20155 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17907), .B1(
        n17938), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17947) );
  AOI22_X1 U20156 ( .A1(n17940), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17939), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17946) );
  AOI22_X1 U20157 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11632), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17941), .ZN(n17945) );
  AOI22_X1 U20158 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17943), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17942), .ZN(n17944) );
  NAND4_X1 U20159 ( .A1(n17947), .A2(n17946), .A3(n17945), .A4(n17944), .ZN(
        n17957) );
  AOI22_X1 U20160 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17928), .ZN(n17955) );
  AOI22_X1 U20161 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17949), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17954) );
  AOI22_X1 U20162 ( .A1(n10992), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17950), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17953) );
  AOI22_X1 U20163 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11537), .B1(
        n17951), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17952) );
  NAND4_X1 U20164 ( .A1(n17955), .A2(n17954), .A3(n17953), .A4(n17952), .ZN(
        n17956) );
  NOR2_X1 U20165 ( .A1(n17957), .A2(n17956), .ZN(n20883) );
  OAI211_X1 U20166 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n17959), .A(n17964), .B(
        n17958), .ZN(n17961) );
  NAND2_X1 U20167 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17962), .ZN(n17960) );
  OAI211_X1 U20168 ( .C1(n20883), .C2(n17935), .A(n17961), .B(n17960), .ZN(
        P3_U2686) );
  AOI21_X1 U20169 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n20389), .ZN(n20371) );
  AOI222_X1 U20170 ( .A1(n17964), .A2(n20371), .B1(P3_EBX_REG_1__SCAN_IN), 
        .B2(n17962), .C1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .C2(n17965), .ZN(
        n17963) );
  INV_X1 U20171 ( .A(n17963), .ZN(P3_U2702) );
  AOI22_X1 U20172 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17965), .B1(
        n17964), .B2(n17967), .ZN(n17966) );
  OAI21_X1 U20173 ( .B1(n17968), .B2(n17967), .A(n17966), .ZN(P3_U2703) );
  INV_X1 U20174 ( .A(n17969), .ZN(n17971) );
  OAI21_X1 U20175 ( .B1(n21403), .B2(n20322), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17970) );
  OAI21_X1 U20176 ( .B1(n17971), .B2(n21438), .A(n17970), .ZN(P3_U2634) );
  OAI21_X1 U20177 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n17973), .A(n17972), .ZN(
        n21436) );
  OAI21_X1 U20178 ( .B1(n20319), .B2(n18356), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17974) );
  OAI221_X1 U20179 ( .B1(n18356), .B2(n21436), .C1(n18356), .C2(n17975), .A(
        n17974), .ZN(P3_U2863) );
  INV_X1 U20180 ( .A(n21314), .ZN(n21310) );
  OAI22_X1 U20181 ( .A1(n21192), .A2(n18351), .B1(n21177), .B2(n11041), .ZN(
        n18022) );
  AOI21_X1 U20182 ( .B1(n18184), .B2(n21310), .A(n18022), .ZN(n18189) );
  INV_X1 U20183 ( .A(n18132), .ZN(n18129) );
  AND3_X1 U20184 ( .A1(n11268), .A2(n18129), .A3(n17976), .ZN(n17979) );
  OAI21_X1 U20185 ( .B1(n17976), .B2(n18306), .A(n18345), .ZN(n18192) );
  AOI211_X1 U20186 ( .C1(n18086), .C2(n17977), .A(n17979), .B(n18192), .ZN(
        n17978) );
  INV_X1 U20187 ( .A(n17978), .ZN(n17992) );
  INV_X1 U20188 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21326) );
  OAI22_X1 U20189 ( .A1(n21329), .A2(n21326), .B1(n20603), .B2(n18180), .ZN(
        n17980) );
  AOI211_X1 U20190 ( .C1(n17992), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17980), .B(n17979), .ZN(n17984) );
  OAI21_X1 U20191 ( .B1(n18258), .B2(n17985), .A(n17981), .ZN(n17982) );
  XNOR2_X1 U20192 ( .A(n17982), .B(n17988), .ZN(n21324) );
  NOR2_X1 U20193 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21310), .ZN(
        n21323) );
  AOI22_X1 U20194 ( .A1(n18261), .A2(n21324), .B1(n18184), .B2(n21323), .ZN(
        n17983) );
  OAI211_X1 U20195 ( .C1(n18189), .C2(n17985), .A(n17984), .B(n17983), .ZN(
        P3_U2812) );
  NAND2_X1 U20196 ( .A1(n17986), .A2(n18184), .ZN(n18123) );
  NOR2_X1 U20197 ( .A1(n17987), .A2(n21300), .ZN(n21034) );
  NAND2_X1 U20198 ( .A1(n21177), .A2(n21034), .ZN(n21292) );
  NAND2_X1 U20199 ( .A1(n21192), .A2(n21034), .ZN(n21291) );
  AOI22_X1 U20200 ( .A1(n18262), .A2(n21292), .B1(n18275), .B2(n21291), .ZN(
        n18083) );
  AND2_X1 U20201 ( .A1(n18072), .A2(n17988), .ZN(n18063) );
  NOR2_X1 U20202 ( .A1(n18063), .A2(n18071), .ZN(n17990) );
  XOR2_X1 U20203 ( .A(n17990), .B(n21300), .Z(n21298) );
  NOR2_X1 U20204 ( .A1(n18132), .A2(n17991), .ZN(n17993) );
  MUX2_X1 U20205 ( .A(n17993), .B(n17992), .S(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .Z(n17995) );
  INV_X1 U20206 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20622) );
  OAI22_X1 U20207 ( .A1(n21329), .A2(n20622), .B1(n20617), .B2(n18180), .ZN(
        n17994) );
  AOI211_X1 U20208 ( .C1(n18261), .C2(n21298), .A(n17995), .B(n17994), .ZN(
        n17996) );
  OAI221_X1 U20209 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18123), 
        .C1(n21300), .C2(n18083), .A(n17996), .ZN(P3_U2811) );
  NAND2_X1 U20210 ( .A1(n18196), .A2(n18004), .ZN(n21186) );
  NOR2_X1 U20211 ( .A1(n18132), .A2(n17997), .ZN(n18016) );
  INV_X1 U20212 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17999) );
  NOR2_X1 U20213 ( .A1(n17997), .A2(n20374), .ZN(n18198) );
  AOI21_X1 U20214 ( .B1(n18254), .B2(n17997), .A(n18318), .ZN(n18200) );
  OAI21_X1 U20215 ( .B1(n18198), .B2(n18346), .A(n18200), .ZN(n18014) );
  INV_X1 U20216 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20579) );
  NAND2_X1 U20217 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18198), .ZN(
        n20581) );
  OAI21_X1 U20218 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18198), .A(
        n20581), .ZN(n20570) );
  OAI22_X1 U20219 ( .A1(n21329), .A2(n20579), .B1(n18180), .B2(n20570), .ZN(
        n17998) );
  AOI221_X1 U20220 ( .B1(n18016), .B2(n17999), .C1(n18014), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17998), .ZN(n18009) );
  NAND2_X1 U20221 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18000) );
  NOR3_X1 U20222 ( .A1(n11717), .A2(n18258), .A3(n18000), .ZN(n18235) );
  NAND2_X1 U20223 ( .A1(n21163), .A2(n18235), .ZN(n18206) );
  NAND2_X1 U20224 ( .A1(n18002), .A2(n18001), .ZN(n18207) );
  AOI22_X1 U20225 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18206), .B1(
        n18207), .B2(n18205), .ZN(n18003) );
  XOR2_X1 U20226 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18003), .Z(
        n21189) );
  INV_X1 U20227 ( .A(n21135), .ZN(n18005) );
  OAI21_X1 U20228 ( .B1(n18006), .B2(n18005), .A(n18004), .ZN(n18007) );
  AOI22_X1 U20229 ( .A1(n18261), .A2(n21189), .B1(n18022), .B2(n18007), .ZN(
        n18008) );
  OAI211_X1 U20230 ( .C1(n18351), .C2(n21186), .A(n18009), .B(n18008), .ZN(
        P3_U2815) );
  AOI22_X1 U20231 ( .A1(n13191), .A2(n21338), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18258), .ZN(n18010) );
  XOR2_X1 U20232 ( .A(n18011), .B(n18010), .Z(n21340) );
  INV_X1 U20233 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18013) );
  AOI21_X1 U20234 ( .B1(n18013), .B2(n20581), .A(n18012), .ZN(n20583) );
  AOI22_X1 U20235 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18014), .B1(
        n18171), .B2(n20583), .ZN(n18018) );
  OAI211_X1 U20236 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18016), .B(n18015), .ZN(n18017) );
  OAI211_X1 U20237 ( .C1(n21342), .C2(n21329), .A(n18018), .B(n18017), .ZN(
        n18019) );
  AOI21_X1 U20238 ( .B1(n18261), .B2(n21340), .A(n18019), .ZN(n18020) );
  INV_X1 U20239 ( .A(n18020), .ZN(n18021) );
  AOI221_X1 U20240 ( .B1(n21338), .B2(n18184), .C1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18022), .A(n18021), .ZN(
        n18023) );
  INV_X1 U20241 ( .A(n18023), .ZN(P3_U2814) );
  NOR2_X1 U20242 ( .A1(n18029), .A2(n20374), .ZN(n18025) );
  AOI21_X1 U20243 ( .B1(n18254), .B2(n18029), .A(n18318), .ZN(n18024) );
  OAI21_X1 U20244 ( .B1(n18025), .B2(n18346), .A(n18024), .ZN(n18040) );
  INV_X1 U20245 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18030) );
  INV_X1 U20246 ( .A(n18025), .ZN(n18214) );
  NOR2_X1 U20247 ( .A1(n18030), .A2(n18214), .ZN(n20541) );
  AOI21_X1 U20248 ( .B1(n18030), .B2(n18214), .A(n20541), .ZN(n20527) );
  AOI22_X1 U20249 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18040), .B1(
        n18171), .B2(n20527), .ZN(n18034) );
  INV_X1 U20250 ( .A(n21130), .ZN(n21142) );
  NOR2_X1 U20251 ( .A1(n21142), .A2(n18220), .ZN(n21154) );
  NAND2_X1 U20252 ( .A1(n18258), .A2(n18026), .ZN(n18043) );
  OAI221_X1 U20253 ( .B1(n18258), .B2(n18027), .C1(n18258), .C2(n21154), .A(
        n18043), .ZN(n18028) );
  XOR2_X1 U20254 ( .A(n11751), .B(n18028), .Z(n21155) );
  NOR2_X1 U20255 ( .A1(n18132), .A2(n18029), .ZN(n18036) );
  AOI22_X1 U20256 ( .A1(n21155), .A2(n18261), .B1(n18036), .B2(n18030), .ZN(
        n18033) );
  NAND2_X1 U20257 ( .A1(n10995), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21156) );
  INV_X1 U20258 ( .A(n18247), .ZN(n18217) );
  OAI22_X1 U20259 ( .A1(n18351), .A2(n21132), .B1(n11041), .B2(n21135), .ZN(
        n18031) );
  INV_X1 U20260 ( .A(n18031), .ZN(n18246) );
  OAI21_X1 U20261 ( .B1(n21152), .B2(n18247), .A(n18246), .ZN(n18045) );
  OAI221_X1 U20262 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21154), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18217), .A(n18045), .ZN(
        n18032) );
  NAND4_X1 U20263 ( .A1(n18034), .A2(n18033), .A3(n21156), .A4(n18032), .ZN(
        P3_U2818) );
  OR2_X1 U20264 ( .A1(n18041), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n21350) );
  NAND2_X1 U20265 ( .A1(n18199), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20556) );
  OAI21_X1 U20266 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n20541), .A(
        n20556), .ZN(n20542) );
  OAI211_X1 U20267 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18036), .B(n18035), .ZN(n18038) );
  NAND2_X1 U20268 ( .A1(n10995), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18037) );
  OAI211_X1 U20269 ( .C1(n18180), .C2(n20542), .A(n18038), .B(n18037), .ZN(
        n18039) );
  AOI21_X1 U20270 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18040), .A(
        n18039), .ZN(n18047) );
  OAI22_X1 U20271 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n13191), .B1(
        n18221), .B2(n18041), .ZN(n18042) );
  NAND2_X1 U20272 ( .A1(n18043), .A2(n18042), .ZN(n18044) );
  XNOR2_X1 U20273 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18044), .ZN(
        n21344) );
  AOI22_X1 U20274 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18045), .B1(
        n18261), .B2(n21344), .ZN(n18046) );
  OAI211_X1 U20275 ( .C1(n18247), .C2(n21350), .A(n18047), .B(n18046), .ZN(
        P3_U2817) );
  AOI22_X1 U20276 ( .A1(n18275), .A2(n21038), .B1(n18262), .B2(n21039), .ZN(
        n18070) );
  OAI21_X1 U20277 ( .B1(n18051), .B2(n18050), .A(n11764), .ZN(n18094) );
  XOR2_X1 U20278 ( .A(n18095), .B(n18094), .Z(n21201) );
  INV_X1 U20279 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18052) );
  NAND2_X1 U20280 ( .A1(n11100), .A2(n18129), .ZN(n18059) );
  AOI221_X1 U20281 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n18052), .C2(n20636), .A(
        n18059), .ZN(n18057) );
  OAI21_X1 U20282 ( .B1(n11100), .B2(n18306), .A(n18345), .ZN(n18053) );
  AOI21_X1 U20283 ( .B1(n18086), .B2(n18054), .A(n18053), .ZN(n18074) );
  OAI21_X1 U20284 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18181), .A(
        n18074), .ZN(n18062) );
  AOI22_X1 U20285 ( .A1(n10995), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18062), .ZN(n18055) );
  OAI21_X1 U20286 ( .B1(n20651), .B2(n18180), .A(n18055), .ZN(n18056) );
  AOI211_X1 U20287 ( .C1(n21201), .C2(n18261), .A(n18057), .B(n18056), .ZN(
        n18058) );
  OAI221_X1 U20288 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18157), 
        .C1(n18095), .C2(n18070), .A(n18058), .ZN(P3_U2808) );
  INV_X1 U20289 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18069) );
  NAND2_X1 U20290 ( .A1(n10995), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n21045) );
  INV_X1 U20291 ( .A(n21045), .ZN(n18061) );
  OAI22_X1 U20292 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18059), .B1(
        n18180), .B2(n20641), .ZN(n18060) );
  AOI211_X1 U20293 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n18062), .A(
        n18061), .B(n18060), .ZN(n18068) );
  NOR2_X1 U20294 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18064) );
  AOI22_X1 U20295 ( .A1(n21042), .A2(n18071), .B1(n18064), .B2(n18063), .ZN(
        n18065) );
  XOR2_X1 U20296 ( .A(n18069), .B(n18065), .Z(n21033) );
  AND2_X1 U20297 ( .A1(n18069), .A2(n21042), .ZN(n21032) );
  INV_X1 U20298 ( .A(n18123), .ZN(n18066) );
  AOI22_X1 U20299 ( .A1(n18261), .A2(n21033), .B1(n21032), .B2(n18066), .ZN(
        n18067) );
  OAI211_X1 U20300 ( .C1(n18070), .C2(n18069), .A(n18068), .B(n18067), .ZN(
        P3_U2809) );
  OAI221_X1 U20301 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18072), 
        .C1(n21300), .C2(n18071), .A(n11764), .ZN(n18073) );
  XOR2_X1 U20302 ( .A(n18082), .B(n18073), .Z(n21304) );
  NAND2_X1 U20303 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18082), .ZN(
        n21309) );
  INV_X1 U20304 ( .A(n20627), .ZN(n18078) );
  AOI221_X1 U20305 ( .B1(n18076), .B2(n18075), .C1(n18333), .C2(n18075), .A(
        n18074), .ZN(n18077) );
  AOI221_X1 U20306 ( .B1(n18171), .B2(n18078), .C1(n18152), .C2(n18078), .A(
        n18077), .ZN(n18079) );
  NAND2_X1 U20307 ( .A1(n10995), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21306) );
  OAI211_X1 U20308 ( .C1(n21309), .C2(n18123), .A(n18079), .B(n21306), .ZN(
        n18080) );
  AOI21_X1 U20309 ( .B1(n18261), .B2(n21304), .A(n18080), .ZN(n18081) );
  OAI21_X1 U20310 ( .B1(n18083), .B2(n18082), .A(n18081), .ZN(P3_U2810) );
  AOI22_X1 U20311 ( .A1(n18275), .A2(n18091), .B1(n18262), .B2(n21272), .ZN(
        n18117) );
  OAI21_X1 U20312 ( .B1(n18103), .B2(n18333), .A(n18345), .ZN(n18084) );
  AOI21_X1 U20313 ( .B1(n18086), .B2(n18085), .A(n18084), .ZN(n18102) );
  AOI221_X1 U20314 ( .B1(n18088), .B2(n18087), .C1(n18333), .C2(n18087), .A(
        n18102), .ZN(n18090) );
  AOI21_X1 U20315 ( .B1(n18180), .B2(n18181), .A(n20666), .ZN(n18089) );
  AOI211_X1 U20316 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n10995), .A(n18090), 
        .B(n18089), .ZN(n18100) );
  NAND2_X1 U20317 ( .A1(n18262), .A2(n21272), .ZN(n18093) );
  NAND2_X1 U20318 ( .A1(n18275), .A2(n18091), .ZN(n18092) );
  OAI22_X1 U20319 ( .A1(n21039), .A2(n18093), .B1(n21038), .B2(n18092), .ZN(
        n18098) );
  AOI221_X1 U20320 ( .B1(n18258), .B2(n18096), .C1(n18095), .C2(n18096), .A(
        n18094), .ZN(n18097) );
  XOR2_X1 U20321 ( .A(n18097), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n21277) );
  AOI22_X1 U20322 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18098), .B1(
        n18261), .B2(n21277), .ZN(n18099) );
  OAI211_X1 U20323 ( .C1(n18117), .C2(n21280), .A(n18100), .B(n18099), .ZN(
        P3_U2807) );
  XOR2_X1 U20324 ( .A(n21205), .B(n18101), .Z(n21210) );
  OAI21_X1 U20325 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18181), .A(
        n18102), .ZN(n18116) );
  INV_X1 U20326 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n20686) );
  NAND2_X1 U20327 ( .A1(n18103), .A2(n18129), .ZN(n18114) );
  AOI221_X1 U20328 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n20686), .C2(n18104), .A(
        n18114), .ZN(n18106) );
  INV_X1 U20329 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20689) );
  OAI22_X1 U20330 ( .A1(n21329), .A2(n20689), .B1(n20692), .B2(n18180), .ZN(
        n18105) );
  AOI211_X1 U20331 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18116), .A(
        n18106), .B(n18105), .ZN(n18111) );
  XOR2_X1 U20332 ( .A(n18107), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n21211) );
  INV_X1 U20333 ( .A(n18108), .ZN(n18159) );
  OAI21_X1 U20334 ( .B1(n18258), .B2(n18159), .A(n18158), .ZN(n18109) );
  XOR2_X1 U20335 ( .A(n18109), .B(n21205), .Z(n21214) );
  AOI22_X1 U20336 ( .A1(n18262), .A2(n21211), .B1(n18261), .B2(n21214), .ZN(
        n18110) );
  OAI211_X1 U20337 ( .C1(n18351), .C2(n21210), .A(n18111), .B(n18110), .ZN(
        P3_U2805) );
  NAND3_X1 U20338 ( .A1(n18113), .A2(n18112), .A3(n21283), .ZN(n21290) );
  NOR2_X1 U20339 ( .A1(n21329), .A2(n20671), .ZN(n21287) );
  OAI22_X1 U20340 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18114), .B1(
        n18180), .B2(n20676), .ZN(n18115) );
  AOI211_X1 U20341 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n18116), .A(
        n21287), .B(n18115), .ZN(n18122) );
  INV_X1 U20342 ( .A(n18117), .ZN(n18120) );
  OAI21_X1 U20343 ( .B1(n18119), .B2(n21283), .A(n18118), .ZN(n21288) );
  AOI22_X1 U20344 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18120), .B1(
        n18261), .B2(n21288), .ZN(n18121) );
  OAI211_X1 U20345 ( .C1(n18123), .C2(n21290), .A(n18122), .B(n18121), .ZN(
        P3_U2806) );
  AOI211_X1 U20346 ( .C1(n18126), .C2(n18125), .A(n18124), .B(n18187), .ZN(
        n18136) );
  OAI22_X1 U20347 ( .A1(n18346), .A2(n18127), .B1(n18306), .B2(n11101), .ZN(
        n18128) );
  OR2_X1 U20348 ( .A1(n18128), .A2(n18318), .ZN(n18156) );
  AOI21_X1 U20349 ( .B1(n18152), .B2(n18150), .A(n18156), .ZN(n18149) );
  NAND3_X1 U20350 ( .A1(n11101), .A2(n11261), .A3(n18129), .ZN(n18144) );
  AOI21_X1 U20351 ( .B1(n18149), .B2(n18144), .A(n18130), .ZN(n18135) );
  NOR3_X1 U20352 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18132), .A3(
        n18131), .ZN(n18134) );
  OAI22_X1 U20353 ( .A1(n21329), .A2(n20720), .B1(n20726), .B2(n18180), .ZN(
        n18133) );
  NOR4_X1 U20354 ( .A1(n18136), .A2(n18135), .A3(n18134), .A4(n18133), .ZN(
        n18142) );
  AOI22_X1 U20355 ( .A1(n18275), .A2(n18137), .B1(n18262), .B2(n21234), .ZN(
        n18165) );
  NAND2_X1 U20356 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18165), .ZN(
        n18146) );
  OAI211_X1 U20357 ( .C1(n18262), .C2(n18275), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18146), .ZN(n18141) );
  NAND3_X1 U20358 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18166), .A3(
        n18139), .ZN(n18140) );
  NAND3_X1 U20359 ( .A1(n18142), .A2(n18141), .A3(n18140), .ZN(P3_U2802) );
  XOR2_X1 U20360 ( .A(n13191), .B(n18143), .Z(n21230) );
  NAND2_X1 U20361 ( .A1(n10995), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21240) );
  OAI211_X1 U20362 ( .C1(n18180), .C2(n20714), .A(n18144), .B(n21240), .ZN(
        n18145) );
  AOI21_X1 U20363 ( .B1(n18261), .B2(n21230), .A(n18145), .ZN(n18148) );
  OAI21_X1 U20364 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18166), .A(
        n18146), .ZN(n18147) );
  OAI211_X1 U20365 ( .C1(n18149), .C2(n11261), .A(n18148), .B(n18147), .ZN(
        P3_U2803) );
  OAI21_X1 U20366 ( .B1(n18151), .B2(n18333), .A(n18150), .ZN(n18155) );
  AOI21_X1 U20367 ( .B1(n18180), .B2(n18181), .A(n20699), .ZN(n18154) );
  NAND2_X1 U20368 ( .A1(n10995), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n21227) );
  INV_X1 U20369 ( .A(n21227), .ZN(n18153) );
  AOI211_X1 U20370 ( .C1(n18156), .C2(n18155), .A(n18154), .B(n18153), .ZN(
        n18164) );
  NOR2_X1 U20371 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18157), .ZN(
        n18161) );
  OAI221_X1 U20372 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18258), 
        .C1(n21205), .C2(n18159), .A(n18158), .ZN(n18160) );
  XOR2_X1 U20373 ( .A(n21229), .B(n18160), .Z(n21226) );
  AOI22_X1 U20374 ( .A1(n18162), .A2(n18161), .B1(n18261), .B2(n21226), .ZN(
        n18163) );
  OAI211_X1 U20375 ( .C1(n18165), .C2(n21229), .A(n18164), .B(n18163), .ZN(
        P3_U2804) );
  NAND2_X1 U20376 ( .A1(n18169), .A2(n18168), .ZN(n18170) );
  XOR2_X1 U20377 ( .A(n18170), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n21258) );
  AOI22_X1 U20378 ( .A1(n10995), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n20757), 
        .B2(n18171), .ZN(n18172) );
  OAI221_X1 U20379 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18174), .C1(
        n11259), .C2(n18173), .A(n18172), .ZN(n18175) );
  AOI21_X1 U20380 ( .B1(n18261), .B2(n21258), .A(n18175), .ZN(n18176) );
  OAI221_X1 U20381 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18179), 
        .C1(n18178), .C2(n18177), .A(n18176), .ZN(P3_U2800) );
  OAI21_X1 U20382 ( .B1(n18183), .B2(n18333), .A(n18182), .ZN(n18191) );
  AOI21_X1 U20383 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18184), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18188) );
  AOI21_X1 U20384 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18186), .A(
        n18185), .ZN(n21334) );
  OAI22_X1 U20385 ( .A1(n18189), .A2(n18188), .B1(n21334), .B2(n18187), .ZN(
        n18190) );
  AOI21_X1 U20386 ( .B1(n18192), .B2(n18191), .A(n18190), .ZN(n18194) );
  NAND2_X1 U20387 ( .A1(n10995), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18193) );
  OAI211_X1 U20388 ( .C1(n18342), .C2(n18195), .A(n18194), .B(n18193), .ZN(
        P3_U2813) );
  AOI21_X1 U20389 ( .B1(n18205), .B2(n18197), .A(n18196), .ZN(n21171) );
  NOR2_X1 U20390 ( .A1(n21329), .A2(n18431), .ZN(n18203) );
  INV_X1 U20391 ( .A(n20556), .ZN(n20537) );
  INV_X1 U20392 ( .A(n18198), .ZN(n20567) );
  OAI21_X1 U20393 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n20537), .A(
        n20567), .ZN(n20558) );
  AOI21_X1 U20394 ( .B1(n18199), .B2(n19264), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18201) );
  OAI22_X1 U20395 ( .A1(n18342), .A2(n20558), .B1(n18201), .B2(n18200), .ZN(
        n18202) );
  AOI211_X1 U20396 ( .C1(n21171), .C2(n18275), .A(n18203), .B(n18202), .ZN(
        n18210) );
  AOI21_X1 U20397 ( .B1(n18205), .B2(n18204), .A(n21188), .ZN(n21170) );
  NAND2_X1 U20398 ( .A1(n18207), .A2(n18206), .ZN(n18208) );
  XOR2_X1 U20399 ( .A(n18208), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n21173) );
  AOI22_X1 U20400 ( .A1(n18262), .A2(n21170), .B1(n18261), .B2(n21173), .ZN(
        n18209) );
  NAND2_X1 U20401 ( .A1(n18210), .A2(n18209), .ZN(P3_U2816) );
  NOR2_X1 U20402 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18211), .ZN(
        n18236) );
  AOI22_X1 U20403 ( .A1(n21130), .A2(n18235), .B1(n18226), .B2(n18236), .ZN(
        n18212) );
  XOR2_X1 U20404 ( .A(n18220), .B(n18212), .Z(n21144) );
  NOR2_X1 U20405 ( .A1(n18318), .A2(n18254), .ZN(n18341) );
  INV_X1 U20406 ( .A(n18341), .ZN(n18238) );
  NAND2_X1 U20407 ( .A1(n18213), .A2(n19264), .ZN(n18228) );
  NAND2_X1 U20408 ( .A1(n18238), .A2(n18228), .ZN(n18231) );
  AOI22_X1 U20409 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18231), .B1(
        n18228), .B2(n11265), .ZN(n18216) );
  INV_X1 U20410 ( .A(n18213), .ZN(n20522) );
  NOR2_X1 U20411 ( .A1(n20522), .A2(n20374), .ZN(n18227) );
  OAI21_X1 U20412 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18227), .A(
        n18214), .ZN(n20511) );
  OAI22_X1 U20413 ( .A1(n18342), .A2(n20511), .B1(n21329), .B2(n21146), .ZN(
        n18215) );
  AOI211_X1 U20414 ( .C1(n18261), .C2(n21144), .A(n18216), .B(n18215), .ZN(
        n18219) );
  INV_X1 U20415 ( .A(n21154), .ZN(n21134) );
  OAI211_X1 U20416 ( .C1(n21130), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n21134), .B(n18217), .ZN(n18218) );
  OAI211_X1 U20417 ( .C1(n18246), .C2(n18220), .A(n18219), .B(n18218), .ZN(
        P3_U2819) );
  INV_X1 U20418 ( .A(n18221), .ZN(n18223) );
  AOI21_X1 U20419 ( .B1(n18258), .B2(n21376), .A(n18235), .ZN(n18222) );
  AOI21_X1 U20420 ( .B1(n21376), .B2(n18223), .A(n18222), .ZN(n18225) );
  AOI221_X1 U20421 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18235), .C1(
        n21376), .C2(n18236), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18224) );
  AOI21_X1 U20422 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18225), .A(
        n18224), .ZN(n21352) );
  NOR3_X1 U20423 ( .A1(n21130), .A2(n18226), .A3(n18247), .ZN(n18233) );
  NAND3_X1 U20424 ( .A1(n18285), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n19264), .ZN(n18267) );
  NOR2_X1 U20425 ( .A1(n20481), .A2(n18267), .ZN(n18242) );
  INV_X1 U20426 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18255) );
  INV_X1 U20427 ( .A(n20482), .ZN(n18251) );
  NAND3_X1 U20428 ( .A1(n18251), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18266) );
  NOR2_X1 U20429 ( .A1(n18255), .A2(n18266), .ZN(n18250) );
  NAND2_X1 U20430 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18250), .ZN(
        n18240) );
  AOI21_X1 U20431 ( .B1(n20496), .B2(n18240), .A(n18227), .ZN(n20505) );
  AOI22_X1 U20432 ( .A1(n18242), .A2(n18228), .B1(n20505), .B2(n18321), .ZN(
        n18230) );
  NAND2_X1 U20433 ( .A1(n10995), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18229) );
  OAI211_X1 U20434 ( .C1(n20496), .C2(n18231), .A(n18230), .B(n18229), .ZN(
        n18232) );
  AOI211_X1 U20435 ( .C1(n21352), .C2(n18261), .A(n18233), .B(n18232), .ZN(
        n18234) );
  OAI21_X1 U20436 ( .B1(n18246), .B2(n21351), .A(n18234), .ZN(P3_U2820) );
  NOR2_X1 U20437 ( .A1(n18236), .A2(n18235), .ZN(n18237) );
  XOR2_X1 U20438 ( .A(n18237), .B(n21376), .Z(n21372) );
  INV_X1 U20439 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18427) );
  NOR2_X1 U20440 ( .A1(n21329), .A2(n18427), .ZN(n18244) );
  INV_X1 U20441 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20457) );
  NOR2_X1 U20442 ( .A1(n18255), .A2(n20457), .ZN(n18252) );
  INV_X1 U20443 ( .A(n18267), .ZN(n18239) );
  AOI22_X1 U20444 ( .A1(n18252), .A2(n18239), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18238), .ZN(n18241) );
  OAI21_X1 U20445 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18250), .A(
        n18240), .ZN(n20486) );
  OAI22_X1 U20446 ( .A1(n18242), .A2(n18241), .B1(n18342), .B2(n20486), .ZN(
        n18243) );
  AOI211_X1 U20447 ( .C1(n18261), .C2(n21372), .A(n18244), .B(n18243), .ZN(
        n18245) );
  OAI221_X1 U20448 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18247), .C1(
        n21376), .C2(n18246), .A(n18245), .ZN(P3_U2821) );
  OAI21_X1 U20449 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18249), .A(
        n18248), .ZN(n21129) );
  AOI21_X1 U20450 ( .B1(n18255), .B2(n18266), .A(n18250), .ZN(n20467) );
  NAND2_X1 U20451 ( .A1(n18251), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18253) );
  AOI211_X1 U20452 ( .C1(n18255), .C2(n18253), .A(n18252), .B(n18333), .ZN(
        n18257) );
  AOI21_X1 U20453 ( .B1(n18254), .B2(n20482), .A(n18318), .ZN(n18278) );
  OAI22_X1 U20454 ( .A1(n21329), .A2(n20484), .B1(n18255), .B2(n18278), .ZN(
        n18256) );
  AOI211_X1 U20455 ( .C1(n20467), .C2(n18321), .A(n18257), .B(n18256), .ZN(
        n18265) );
  AOI22_X1 U20456 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18258), .B1(
        n13191), .B2(n21122), .ZN(n18259) );
  XOR2_X1 U20457 ( .A(n18260), .B(n18259), .Z(n18263) );
  INV_X1 U20458 ( .A(n18263), .ZN(n21125) );
  AOI22_X1 U20459 ( .A1(n18263), .A2(n18262), .B1(n18261), .B2(n21125), .ZN(
        n18264) );
  OAI211_X1 U20460 ( .C1(n18351), .C2(n21129), .A(n18265), .B(n18264), .ZN(
        P3_U2822) );
  NOR2_X1 U20461 ( .A1(n20482), .A2(n20374), .ZN(n18286) );
  OAI21_X1 U20462 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18286), .A(
        n18266), .ZN(n20452) );
  OAI22_X1 U20463 ( .A1(n18342), .A2(n20452), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18267), .ZN(n18268) );
  AOI21_X1 U20464 ( .B1(n10995), .B2(P3_REIP_REG_7__SCAN_IN), .A(n18268), .ZN(
        n18277) );
  AOI21_X1 U20465 ( .B1(n21116), .B2(n18270), .A(n18269), .ZN(n21109) );
  AOI21_X1 U20466 ( .B1(n18273), .B2(n18272), .A(n18271), .ZN(n18274) );
  XOR2_X1 U20467 ( .A(n18274), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n21108) );
  AOI22_X1 U20468 ( .A1(n18339), .A2(n21109), .B1(n18275), .B2(n21108), .ZN(
        n18276) );
  OAI211_X1 U20469 ( .C1(n20457), .C2(n18278), .A(n18277), .B(n18276), .ZN(
        P3_U2823) );
  OAI21_X1 U20470 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18280), .A(
        n18279), .ZN(n21107) );
  AOI21_X1 U20471 ( .B1(n11111), .B2(n18282), .A(n18281), .ZN(n21105) );
  NAND2_X1 U20472 ( .A1(n18285), .A2(n19264), .ZN(n18283) );
  OAI22_X1 U20473 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18283), .B1(
        n21329), .B2(n21102), .ZN(n18284) );
  AOI21_X1 U20474 ( .B1(n18339), .B2(n21105), .A(n18284), .ZN(n18288) );
  AOI21_X1 U20475 ( .B1(n19264), .B2(n18285), .A(n18341), .ZN(n18299) );
  INV_X1 U20476 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20440) );
  NAND2_X1 U20477 ( .A1(n18285), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18289) );
  AOI21_X1 U20478 ( .B1(n20440), .B2(n18289), .A(n18286), .ZN(n20439) );
  AOI22_X1 U20479 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18299), .B1(
        n20439), .B2(n18321), .ZN(n18287) );
  OAI211_X1 U20480 ( .C1(n18351), .C2(n21107), .A(n18288), .B(n18287), .ZN(
        P3_U2824) );
  NOR2_X1 U20481 ( .A1(n20406), .A2(n20374), .ZN(n18308) );
  OAI21_X1 U20482 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18308), .A(
        n18289), .ZN(n20426) );
  OAI21_X1 U20483 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18290), .A(
        n21084), .ZN(n18295) );
  OAI211_X1 U20484 ( .C1(n18293), .C2(n18292), .A(n21384), .B(n18291), .ZN(
        n18294) );
  OAI21_X1 U20485 ( .B1(n18296), .B2(n18295), .A(n18294), .ZN(n21097) );
  OAI21_X1 U20486 ( .B1(n18318), .B2(n20406), .A(n18297), .ZN(n18298) );
  AOI22_X1 U20487 ( .A1(n21443), .A2(n21097), .B1(n18299), .B2(n18298), .ZN(
        n18300) );
  NAND2_X1 U20488 ( .A1(n10995), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21098) );
  OAI211_X1 U20489 ( .C1(n18342), .C2(n20426), .A(n18300), .B(n21098), .ZN(
        P3_U2825) );
  OAI21_X1 U20490 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18302), .A(
        n18301), .ZN(n21086) );
  AOI21_X1 U20491 ( .B1(n11119), .B2(n18304), .A(n18303), .ZN(n21085) );
  NOR2_X1 U20492 ( .A1(n21329), .A2(n20408), .ZN(n21087) );
  INV_X1 U20493 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20424) );
  AND3_X1 U20494 ( .A1(n20424), .A2(n18307), .A3(n19264), .ZN(n18305) );
  AOI211_X1 U20495 ( .C1(n18339), .C2(n21085), .A(n21087), .B(n18305), .ZN(
        n18310) );
  OAI21_X1 U20496 ( .B1(n18307), .B2(n18306), .A(n18345), .ZN(n18320) );
  NAND2_X1 U20497 ( .A1(n18307), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18317) );
  AOI21_X1 U20498 ( .B1(n20424), .B2(n18317), .A(n18308), .ZN(n20412) );
  AOI22_X1 U20499 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18320), .B1(
        n20412), .B2(n18321), .ZN(n18309) );
  OAI211_X1 U20500 ( .C1(n18351), .C2(n21086), .A(n18310), .B(n18309), .ZN(
        P3_U2826) );
  OAI21_X1 U20501 ( .B1(n18313), .B2(n18312), .A(n18311), .ZN(n21080) );
  AOI21_X1 U20502 ( .B1(n18316), .B2(n18315), .A(n18314), .ZN(n21077) );
  AOI22_X1 U20503 ( .A1(n10995), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18339), 
        .B2(n21077), .ZN(n18323) );
  NAND2_X1 U20504 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18327) );
  INV_X1 U20505 ( .A(n18317), .ZN(n20411) );
  AOI21_X1 U20506 ( .B1(n20401), .B2(n18327), .A(n20411), .ZN(n20394) );
  OAI21_X1 U20507 ( .B1(n18318), .B2(n20378), .A(n20401), .ZN(n18319) );
  AOI22_X1 U20508 ( .A1(n20394), .A2(n18321), .B1(n18320), .B2(n18319), .ZN(
        n18322) );
  OAI211_X1 U20509 ( .C1(n18351), .C2(n21080), .A(n18323), .B(n18322), .ZN(
        P3_U2827) );
  AOI21_X1 U20510 ( .B1(n18326), .B2(n18325), .A(n18324), .ZN(n21063) );
  INV_X1 U20511 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20386) );
  NOR2_X1 U20512 ( .A1(n21329), .A2(n20386), .ZN(n21067) );
  OAI21_X1 U20513 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n18327), .ZN(n20383) );
  OAI21_X1 U20514 ( .B1(n18330), .B2(n18329), .A(n18328), .ZN(n21066) );
  OAI22_X1 U20515 ( .A1(n18342), .A2(n20383), .B1(n18351), .B2(n21066), .ZN(
        n18331) );
  AOI211_X1 U20516 ( .C1(n18339), .C2(n21063), .A(n21067), .B(n18331), .ZN(
        n18332) );
  OAI221_X1 U20517 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18333), .C1(
        n20378), .C2(n18345), .A(n18332), .ZN(P3_U2828) );
  AOI21_X1 U20518 ( .B1(n18335), .B2(n18344), .A(n18334), .ZN(n21055) );
  AOI21_X1 U20519 ( .B1(n18337), .B2(n18343), .A(n18336), .ZN(n21059) );
  INV_X1 U20520 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20385) );
  OAI22_X1 U20521 ( .A1(n21059), .A2(n18351), .B1(n21329), .B2(n20385), .ZN(
        n18338) );
  AOI21_X1 U20522 ( .B1(n18339), .B2(n21055), .A(n18338), .ZN(n18340) );
  OAI221_X1 U20523 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18342), .C1(
        n20374), .C2(n18341), .A(n18340), .ZN(P3_U2829) );
  NAND2_X1 U20524 ( .A1(n18344), .A2(n18343), .ZN(n21049) );
  INV_X1 U20525 ( .A(n21049), .ZN(n21048) );
  NAND3_X1 U20526 ( .A1(n18347), .A2(n18346), .A3(n18345), .ZN(n18348) );
  AOI22_X1 U20527 ( .A1(n10995), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18348), .ZN(n18349) );
  OAI221_X1 U20528 ( .B1(n21048), .B2(n18351), .C1(n21049), .C2(n18350), .A(
        n18349), .ZN(P3_U2830) );
  NOR2_X1 U20529 ( .A1(n18939), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18970) );
  NAND2_X1 U20530 ( .A1(n21398), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18961) );
  NOR2_X1 U20531 ( .A1(n21398), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18982) );
  INV_X1 U20532 ( .A(n18982), .ZN(n18981) );
  AOI21_X1 U20533 ( .B1(n18961), .B2(n18981), .A(n18976), .ZN(n18352) );
  AOI21_X1 U20534 ( .B1(n18970), .B2(n18353), .A(n18352), .ZN(n18355) );
  OAI22_X1 U20535 ( .A1(n18356), .A2(n18355), .B1(n18354), .B2(n18975), .ZN(
        P3_U2866) );
  NOR4_X1 U20536 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18360) );
  NOR4_X1 U20537 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18359) );
  NOR4_X1 U20538 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18358) );
  NOR4_X1 U20539 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18357) );
  NAND4_X1 U20540 ( .A1(n18360), .A2(n18359), .A3(n18358), .A4(n18357), .ZN(
        n18366) );
  NOR4_X1 U20541 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18364) );
  AOI211_X1 U20542 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18363) );
  NOR4_X1 U20543 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18362) );
  NOR4_X1 U20544 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18361) );
  NAND4_X1 U20545 ( .A1(n18364), .A2(n18363), .A3(n18362), .A4(n18361), .ZN(
        n18365) );
  NOR2_X1 U20546 ( .A1(n18366), .A2(n18365), .ZN(n18378) );
  INV_X1 U20547 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18368) );
  OAI21_X1 U20548 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18378), .ZN(n18367) );
  OAI21_X1 U20549 ( .B1(n18378), .B2(n18368), .A(n18367), .ZN(P3_U3293) );
  INV_X1 U20550 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18371) );
  AOI21_X1 U20551 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18369) );
  OAI221_X1 U20552 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18369), .C1(n20385), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18378), .ZN(n18370) );
  OAI21_X1 U20553 ( .B1(n18378), .B2(n18371), .A(n18370), .ZN(P3_U3292) );
  INV_X1 U20554 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18373) );
  NOR3_X1 U20555 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18374) );
  OAI21_X1 U20556 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18374), .A(n18378), .ZN(
        n18372) );
  OAI21_X1 U20557 ( .B1(n18378), .B2(n18373), .A(n18372), .ZN(P3_U2638) );
  INV_X1 U20558 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21857) );
  AOI21_X1 U20559 ( .B1(n20385), .B2(n21857), .A(n18374), .ZN(n18377) );
  INV_X1 U20560 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18376) );
  INV_X1 U20561 ( .A(n18378), .ZN(n18375) );
  AOI22_X1 U20562 ( .A1(n18378), .A2(n18377), .B1(n18376), .B2(n18375), .ZN(
        P3_U2639) );
  OAI22_X1 U20563 ( .A1(n11798), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n21864), .ZN(n18379) );
  INV_X1 U20564 ( .A(n18379), .ZN(P3_U3297) );
  INV_X1 U20565 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18380) );
  AOI22_X1 U20566 ( .A1(n21864), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18380), 
        .B2(n11798), .ZN(P3_U3294) );
  AOI21_X1 U20567 ( .B1(n21909), .B2(n21861), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18381) );
  AOI22_X1 U20568 ( .A1(n21864), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18381), 
        .B2(n11798), .ZN(P3_U2635) );
  INV_X1 U20569 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20976) );
  AOI22_X1 U20570 ( .A1(n18415), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18382) );
  OAI21_X1 U20571 ( .B1(n20976), .B2(n18398), .A(n18382), .ZN(P3_U2767) );
  INV_X1 U20572 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20345) );
  AOI22_X1 U20573 ( .A1(n18415), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18383) );
  OAI21_X1 U20574 ( .B1(n20345), .B2(n18398), .A(n18383), .ZN(P3_U2766) );
  INV_X1 U20575 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20774) );
  AOI22_X1 U20576 ( .A1(n18415), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18384) );
  OAI21_X1 U20577 ( .B1(n20774), .B2(n18398), .A(n18384), .ZN(P3_U2765) );
  INV_X1 U20578 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20775) );
  AOI22_X1 U20579 ( .A1(n18415), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18385) );
  OAI21_X1 U20580 ( .B1(n20775), .B2(n18398), .A(n18385), .ZN(P3_U2764) );
  INV_X1 U20581 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20824) );
  AOI22_X1 U20582 ( .A1(n18415), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18386) );
  OAI21_X1 U20583 ( .B1(n20824), .B2(n18398), .A(n18386), .ZN(P3_U2763) );
  INV_X1 U20584 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20772) );
  AOI22_X1 U20585 ( .A1(n18415), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18387) );
  OAI21_X1 U20586 ( .B1(n20772), .B2(n18398), .A(n18387), .ZN(P3_U2762) );
  INV_X1 U20587 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20811) );
  AOI22_X1 U20588 ( .A1(n18415), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18388) );
  OAI21_X1 U20589 ( .B1(n20811), .B2(n18398), .A(n18388), .ZN(P3_U2761) );
  INV_X1 U20590 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20773) );
  AOI22_X1 U20591 ( .A1(n18415), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18389) );
  OAI21_X1 U20592 ( .B1(n20773), .B2(n18398), .A(n18389), .ZN(P3_U2760) );
  INV_X1 U20593 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20963) );
  AOI22_X1 U20594 ( .A1(n18415), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18390) );
  OAI21_X1 U20595 ( .B1(n20963), .B2(n18398), .A(n18390), .ZN(P3_U2759) );
  INV_X1 U20596 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20783) );
  AOI22_X1 U20597 ( .A1(n18415), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18391) );
  OAI21_X1 U20598 ( .B1(n20783), .B2(n18398), .A(n18391), .ZN(P3_U2758) );
  INV_X1 U20599 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20802) );
  AOI22_X1 U20600 ( .A1(n18415), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18392) );
  OAI21_X1 U20601 ( .B1(n20802), .B2(n18398), .A(n18392), .ZN(P3_U2757) );
  INV_X1 U20602 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20356) );
  AOI22_X1 U20603 ( .A1(n18415), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18393) );
  OAI21_X1 U20604 ( .B1(n20356), .B2(n18398), .A(n18393), .ZN(P3_U2756) );
  INV_X1 U20605 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20359) );
  AOI22_X1 U20606 ( .A1(n18415), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18394) );
  OAI21_X1 U20607 ( .B1(n20359), .B2(n18398), .A(n18394), .ZN(P3_U2755) );
  INV_X1 U20608 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20361) );
  AOI22_X1 U20609 ( .A1(n18415), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18395) );
  OAI21_X1 U20610 ( .B1(n20361), .B2(n18398), .A(n18395), .ZN(P3_U2754) );
  INV_X1 U20611 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20947) );
  AOI22_X1 U20612 ( .A1(n18415), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18396) );
  OAI21_X1 U20613 ( .B1(n20947), .B2(n18398), .A(n18396), .ZN(P3_U2753) );
  INV_X1 U20614 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20367) );
  AOI22_X1 U20615 ( .A1(n18415), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18397) );
  OAI21_X1 U20616 ( .B1(n20367), .B2(n18398), .A(n18397), .ZN(P3_U2752) );
  INV_X1 U20617 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20941) );
  AOI22_X1 U20618 ( .A1(n18415), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18400) );
  OAI21_X1 U20619 ( .B1(n20941), .B2(n18417), .A(n18400), .ZN(P3_U2751) );
  INV_X1 U20620 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20878) );
  AOI22_X1 U20621 ( .A1(n18415), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18401) );
  OAI21_X1 U20622 ( .B1(n20878), .B2(n18417), .A(n18401), .ZN(P3_U2750) );
  INV_X1 U20623 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20859) );
  AOI22_X1 U20624 ( .A1(n18415), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18402) );
  OAI21_X1 U20625 ( .B1(n20859), .B2(n18417), .A(n18402), .ZN(P3_U2749) );
  INV_X1 U20626 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20861) );
  AOI22_X1 U20627 ( .A1(n18415), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18403) );
  OAI21_X1 U20628 ( .B1(n20861), .B2(n18417), .A(n18403), .ZN(P3_U2748) );
  INV_X1 U20629 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20860) );
  AOI22_X1 U20630 ( .A1(n18415), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18404) );
  OAI21_X1 U20631 ( .B1(n20860), .B2(n18417), .A(n18404), .ZN(P3_U2747) );
  INV_X1 U20632 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20858) );
  AOI22_X1 U20633 ( .A1(n18415), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18405) );
  OAI21_X1 U20634 ( .B1(n20858), .B2(n18417), .A(n18405), .ZN(P3_U2746) );
  INV_X1 U20635 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20862) );
  AOI22_X1 U20636 ( .A1(n18415), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18406) );
  OAI21_X1 U20637 ( .B1(n20862), .B2(n18417), .A(n18406), .ZN(P3_U2745) );
  INV_X1 U20638 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20930) );
  AOI22_X1 U20639 ( .A1(n18415), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18407) );
  OAI21_X1 U20640 ( .B1(n20930), .B2(n18417), .A(n18407), .ZN(P3_U2744) );
  INV_X1 U20641 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20922) );
  AOI22_X1 U20642 ( .A1(n18415), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18408) );
  OAI21_X1 U20643 ( .B1(n20922), .B2(n18417), .A(n18408), .ZN(P3_U2743) );
  INV_X1 U20644 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20885) );
  AOI22_X1 U20645 ( .A1(n18415), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18409) );
  OAI21_X1 U20646 ( .B1(n20885), .B2(n18417), .A(n18409), .ZN(P3_U2742) );
  INV_X1 U20647 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20336) );
  AOI22_X1 U20648 ( .A1(n18415), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18411) );
  OAI21_X1 U20649 ( .B1(n20336), .B2(n18417), .A(n18411), .ZN(P3_U2741) );
  INV_X1 U20650 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20915) );
  AOI22_X1 U20651 ( .A1(n18415), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18412) );
  OAI21_X1 U20652 ( .B1(n20915), .B2(n18417), .A(n18412), .ZN(P3_U2740) );
  INV_X1 U20653 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20339) );
  AOI22_X1 U20654 ( .A1(n18415), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18413) );
  OAI21_X1 U20655 ( .B1(n20339), .B2(n18417), .A(n18413), .ZN(P3_U2739) );
  INV_X1 U20656 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20341) );
  AOI22_X1 U20657 ( .A1(n18415), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18414) );
  OAI21_X1 U20658 ( .B1(n20341), .B2(n18417), .A(n18414), .ZN(P3_U2738) );
  INV_X1 U20659 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20903) );
  AOI22_X1 U20660 ( .A1(n18415), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18410), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18416) );
  OAI21_X1 U20661 ( .B1(n20903), .B2(n18417), .A(n18416), .ZN(P3_U2737) );
  NOR2_X1 U20662 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18418), .ZN(n18419) );
  NOR2_X1 U20663 ( .A1(n21864), .A2(n18419), .ZN(P3_U2633) );
  NOR2_X1 U20664 ( .A1(n11798), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18436) );
  AOI22_X1 U20665 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18438), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n11798), .ZN(n18420) );
  OAI21_X1 U20666 ( .B1(n20386), .B2(n18443), .A(n18420), .ZN(P3_U3032) );
  AOI22_X1 U20667 ( .A1(n18436), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n11798), .ZN(n18421) );
  OAI21_X1 U20668 ( .B1(n18444), .B2(n20386), .A(n18421), .ZN(P3_U3033) );
  AOI22_X1 U20669 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n18438), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n11798), .ZN(n18422) );
  OAI21_X1 U20670 ( .B1(n20408), .B2(n18443), .A(n18422), .ZN(P3_U3034) );
  AOI22_X1 U20671 ( .A1(n18436), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n11798), .ZN(n18423) );
  OAI21_X1 U20672 ( .B1(n18444), .B2(n20408), .A(n18423), .ZN(P3_U3035) );
  AOI22_X1 U20673 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18438), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n11798), .ZN(n18424) );
  OAI21_X1 U20674 ( .B1(n21102), .B2(n18443), .A(n18424), .ZN(P3_U3036) );
  AOI22_X1 U20675 ( .A1(n18436), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n11798), .ZN(n18425) );
  OAI21_X1 U20676 ( .B1(n18444), .B2(n21102), .A(n18425), .ZN(P3_U3037) );
  AOI22_X1 U20677 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n18438), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n11798), .ZN(n18426) );
  OAI21_X1 U20678 ( .B1(n20484), .B2(n18443), .A(n18426), .ZN(P3_U3038) );
  INV_X1 U20679 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19995) );
  OAI222_X1 U20680 ( .A1(n18443), .A2(n18427), .B1(n19995), .B2(n21864), .C1(
        n20484), .C2(n18444), .ZN(P3_U3039) );
  INV_X1 U20681 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19997) );
  OAI222_X1 U20682 ( .A1(n18443), .A2(n18428), .B1(n19997), .B2(n21864), .C1(
        n18427), .C2(n18444), .ZN(P3_U3040) );
  INV_X1 U20683 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19999) );
  OAI222_X1 U20684 ( .A1(n18443), .A2(n21146), .B1(n19999), .B2(n21864), .C1(
        n18428), .C2(n18444), .ZN(P3_U3041) );
  INV_X1 U20685 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20529) );
  INV_X1 U20686 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20001) );
  OAI222_X1 U20687 ( .A1(n18443), .A2(n20529), .B1(n20001), .B2(n21864), .C1(
        n21146), .C2(n18444), .ZN(P3_U3042) );
  AOI22_X1 U20688 ( .A1(n18436), .A2(P3_REIP_REG_13__SCAN_IN), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n11798), .ZN(n18429) );
  OAI21_X1 U20689 ( .B1(n18444), .B2(n20529), .A(n18429), .ZN(P3_U3043) );
  AOI22_X1 U20690 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n18438), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n11798), .ZN(n18430) );
  OAI21_X1 U20691 ( .B1(n18431), .B2(n18443), .A(n18430), .ZN(P3_U3044) );
  AOI222_X1 U20692 ( .A1(n18436), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n11798), .C1(P3_REIP_REG_14__SCAN_IN), 
        .C2(n18438), .ZN(n18432) );
  INV_X1 U20693 ( .A(n18432), .ZN(P3_U3045) );
  INV_X1 U20694 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20006) );
  OAI222_X1 U20695 ( .A1(n18443), .A2(n21342), .B1(n20006), .B2(n21864), .C1(
        n20579), .C2(n18444), .ZN(P3_U3046) );
  INV_X1 U20696 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20008) );
  OAI222_X1 U20697 ( .A1(n18443), .A2(n18433), .B1(n20008), .B2(n21864), .C1(
        n21342), .C2(n18444), .ZN(P3_U3047) );
  INV_X1 U20698 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20010) );
  OAI222_X1 U20699 ( .A1(n18433), .A2(n18444), .B1(n20010), .B2(n21864), .C1(
        n21326), .C2(n18443), .ZN(P3_U3048) );
  INV_X1 U20700 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20012) );
  OAI222_X1 U20701 ( .A1(n21326), .A2(n18444), .B1(n20012), .B2(n21864), .C1(
        n20622), .C2(n18443), .ZN(P3_U3049) );
  AOI22_X1 U20702 ( .A1(n18436), .A2(P3_REIP_REG_20__SCAN_IN), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n11798), .ZN(n18434) );
  OAI21_X1 U20703 ( .B1(n18444), .B2(n20622), .A(n18434), .ZN(P3_U3050) );
  INV_X1 U20704 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20646) );
  AOI22_X1 U20705 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18438), .B1(
        P3_ADDRESS_REG_19__SCAN_IN), .B2(n11798), .ZN(n18435) );
  OAI21_X1 U20706 ( .B1(n20646), .B2(n18443), .A(n18435), .ZN(P3_U3051) );
  INV_X1 U20707 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20645) );
  INV_X1 U20708 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20016) );
  OAI222_X1 U20709 ( .A1(n18443), .A2(n20645), .B1(n20016), .B2(n21864), .C1(
        n20646), .C2(n18444), .ZN(P3_U3052) );
  AOI22_X1 U20710 ( .A1(n18436), .A2(P3_REIP_REG_23__SCAN_IN), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n11798), .ZN(n18437) );
  OAI21_X1 U20711 ( .B1(n18444), .B2(n20645), .A(n18437), .ZN(P3_U3053) );
  AOI22_X1 U20712 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n18438), .B1(
        P3_ADDRESS_REG_22__SCAN_IN), .B2(n11798), .ZN(n18439) );
  OAI21_X1 U20713 ( .B1(n20671), .B2(n18443), .A(n18439), .ZN(P3_U3054) );
  INV_X1 U20714 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20020) );
  OAI222_X1 U20715 ( .A1(n20671), .A2(n18444), .B1(n20020), .B2(n21864), .C1(
        n20689), .C2(n18443), .ZN(P3_U3055) );
  INV_X1 U20716 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18440) );
  INV_X1 U20717 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20022) );
  OAI222_X1 U20718 ( .A1(n18443), .A2(n18440), .B1(n20022), .B2(n21864), .C1(
        n20689), .C2(n18444), .ZN(P3_U3056) );
  INV_X1 U20719 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20024) );
  OAI222_X1 U20720 ( .A1(n18443), .A2(n18441), .B1(n20024), .B2(n21864), .C1(
        n18440), .C2(n18444), .ZN(P3_U3057) );
  INV_X1 U20721 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20026) );
  OAI222_X1 U20722 ( .A1(n18443), .A2(n20720), .B1(n20026), .B2(n21864), .C1(
        n18441), .C2(n18444), .ZN(P3_U3058) );
  INV_X1 U20723 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20028) );
  OAI222_X1 U20724 ( .A1(n20720), .A2(n18444), .B1(n20028), .B2(n21864), .C1(
        n18442), .C2(n18443), .ZN(P3_U3059) );
  INV_X1 U20725 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20031) );
  OAI222_X1 U20726 ( .A1(n18443), .A2(n20750), .B1(n20031), .B2(n21864), .C1(
        n18442), .C2(n18444), .ZN(P3_U3060) );
  INV_X1 U20727 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20033) );
  INV_X1 U20728 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20752) );
  OAI222_X1 U20729 ( .A1(n20750), .A2(n18444), .B1(n20033), .B2(n21864), .C1(
        n20752), .C2(n18443), .ZN(P3_U3061) );
  OAI22_X1 U20730 ( .A1(n11798), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n21864), .ZN(n18445) );
  INV_X1 U20731 ( .A(n18445), .ZN(P3_U3277) );
  OAI22_X1 U20732 ( .A1(n11798), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n21864), .ZN(n18446) );
  INV_X1 U20733 ( .A(n18446), .ZN(P3_U3276) );
  OAI22_X1 U20734 ( .A1(n11798), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n21864), .ZN(n18447) );
  INV_X1 U20735 ( .A(n18447), .ZN(P3_U3275) );
  OAI22_X1 U20736 ( .A1(n11798), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n21864), .ZN(n18448) );
  INV_X1 U20737 ( .A(n18448), .ZN(P3_U3274) );
  NOR4_X1 U20738 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18451)
         );
  INV_X1 U20739 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18449) );
  NOR4_X1 U20740 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18449), .ZN(n18450) );
  INV_X2 U20741 ( .A(n19261), .ZN(U215) );
  NAND3_X1 U20742 ( .A1(n18451), .A2(n18450), .A3(U215), .ZN(U213) );
  NAND2_X1 U20743 ( .A1(n18452), .A2(n18796), .ZN(n18458) );
  INV_X1 U20744 ( .A(n18802), .ZN(n19864) );
  AOI22_X1 U20745 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(n18774), .B1(n18795), .B2(
        n19864), .ZN(n18457) );
  INV_X1 U20746 ( .A(n18453), .ZN(n18454) );
  NAND2_X1 U20747 ( .A1(n18776), .A2(n18454), .ZN(n18456) );
  NAND2_X1 U20748 ( .A1(n18755), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18455) );
  NAND4_X1 U20749 ( .A1(n18458), .A2(n18457), .A3(n18456), .A4(n18455), .ZN(
        n18459) );
  AOI21_X1 U20750 ( .B1(n19865), .B2(n18472), .A(n18459), .ZN(n18461) );
  NAND2_X1 U20751 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18794), .ZN(
        n18460) );
  OAI211_X1 U20752 ( .C1(n18462), .C2(n18888), .A(n18461), .B(n18460), .ZN(
        P2_U2855) );
  AOI22_X1 U20753 ( .A1(n18774), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18794), .ZN(n18463) );
  OAI21_X1 U20754 ( .B1(n18791), .B2(n18464), .A(n18463), .ZN(n18465) );
  AOI21_X1 U20755 ( .B1(n18776), .B2(n18466), .A(n18465), .ZN(n18467) );
  OAI21_X1 U20756 ( .B1(n18780), .B2(n18468), .A(n18467), .ZN(n18469) );
  AOI21_X1 U20757 ( .B1(n18470), .B2(n18796), .A(n18469), .ZN(n18475) );
  NOR2_X1 U20758 ( .A1(n18888), .A2(n11029), .ZN(n18614) );
  AOI22_X1 U20759 ( .A1(n18614), .A2(n18473), .B1(n18472), .B2(n18471), .ZN(
        n18474) );
  OAI211_X1 U20760 ( .C1(n18888), .C2(n18476), .A(n18475), .B(n18474), .ZN(
        P2_U2854) );
  AOI22_X1 U20761 ( .A1(n18774), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18794), .ZN(n18495) );
  NAND2_X1 U20762 ( .A1(n18478), .A2(n18477), .ZN(n18481) );
  INV_X1 U20763 ( .A(n18479), .ZN(n18480) );
  NAND2_X1 U20764 ( .A1(n18481), .A2(n18480), .ZN(n19663) );
  OAI22_X1 U20765 ( .A1(n18482), .A2(n18800), .B1(n18780), .B2(n19663), .ZN(
        n18483) );
  AOI211_X1 U20766 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n18755), .A(n16328), .B(
        n18483), .ZN(n18494) );
  OAI22_X1 U20767 ( .A1(n19665), .A2(n18485), .B1(n18484), .B2(n18737), .ZN(
        n18486) );
  INV_X1 U20768 ( .A(n18486), .ZN(n18493) );
  INV_X1 U20769 ( .A(n18487), .ZN(n18491) );
  NOR2_X1 U20770 ( .A1(n18783), .A2(n18488), .ZN(n18490) );
  AOI21_X1 U20771 ( .B1(n18491), .B2(n18490), .A(n18888), .ZN(n18489) );
  OAI21_X1 U20772 ( .B1(n18491), .B2(n18490), .A(n18489), .ZN(n18492) );
  NAND4_X1 U20773 ( .A1(n18495), .A2(n18494), .A3(n18493), .A4(n18492), .ZN(
        P2_U2851) );
  AOI22_X1 U20774 ( .A1(n18774), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18794), .ZN(n18496) );
  OAI21_X1 U20775 ( .B1(n18497), .B2(n18800), .A(n18496), .ZN(n18498) );
  AOI211_X1 U20776 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18755), .A(n16328), .B(
        n18498), .ZN(n18505) );
  NAND2_X1 U20777 ( .A1(n11029), .A2(n18499), .ZN(n18500) );
  XNOR2_X1 U20778 ( .A(n18501), .B(n18500), .ZN(n18502) );
  AOI22_X1 U20779 ( .A1(n18796), .A2(n18503), .B1(n18784), .B2(n18502), .ZN(
        n18504) );
  OAI211_X1 U20780 ( .C1(n18780), .C2(n19619), .A(n18505), .B(n18504), .ZN(
        P2_U2850) );
  OAI21_X1 U20781 ( .B1(n13049), .B2(n18791), .A(n18848), .ZN(n18509) );
  OAI22_X1 U20782 ( .A1(n18800), .A2(n18507), .B1(n18506), .B2(n18788), .ZN(
        n18508) );
  AOI211_X1 U20783 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18794), .A(
        n18509), .B(n18508), .ZN(n18516) );
  NOR2_X1 U20784 ( .A1(n18783), .A2(n18510), .ZN(n18512) );
  XNOR2_X1 U20785 ( .A(n18512), .B(n18511), .ZN(n18513) );
  AOI22_X1 U20786 ( .A1(n18796), .A2(n18514), .B1(n18784), .B2(n18513), .ZN(
        n18515) );
  OAI211_X1 U20787 ( .C1(n18780), .C2(n19558), .A(n18516), .B(n18515), .ZN(
        P2_U2849) );
  NAND2_X1 U20788 ( .A1(n11029), .A2(n18517), .ZN(n18519) );
  XOR2_X1 U20789 ( .A(n18519), .B(n18518), .Z(n18526) );
  AOI22_X1 U20790 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18794), .B1(
        n18520), .B2(n18776), .ZN(n18521) );
  OAI211_X1 U20791 ( .C1(n18788), .C2(n14508), .A(n18521), .B(n18848), .ZN(
        n18523) );
  OAI22_X1 U20792 ( .A1(n18791), .A2(n13056), .B1(n18780), .B2(n19396), .ZN(
        n18522) );
  AOI211_X1 U20793 ( .C1(n18524), .C2(n18796), .A(n18523), .B(n18522), .ZN(
        n18525) );
  OAI21_X1 U20794 ( .B1(n18526), .B2(n18888), .A(n18525), .ZN(P2_U2848) );
  AOI22_X1 U20795 ( .A1(n18774), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18794), .ZN(n18527) );
  OAI21_X1 U20796 ( .B1(n18528), .B2(n18800), .A(n18527), .ZN(n18529) );
  AOI211_X1 U20797 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n18755), .A(n16328), .B(
        n18529), .ZN(n18537) );
  AOI21_X1 U20798 ( .B1(n18531), .B2(n15306), .A(n18530), .ZN(n19390) );
  NOR2_X1 U20799 ( .A1(n18783), .A2(n18532), .ZN(n18534) );
  XNOR2_X1 U20800 ( .A(n18534), .B(n18533), .ZN(n18535) );
  AOI22_X1 U20801 ( .A1(n18795), .A2(n19390), .B1(n18784), .B2(n18535), .ZN(
        n18536) );
  OAI211_X1 U20802 ( .C1(n18737), .C2(n18538), .A(n18537), .B(n18536), .ZN(
        P2_U2847) );
  NAND2_X1 U20803 ( .A1(n11029), .A2(n18539), .ZN(n18541) );
  XOR2_X1 U20804 ( .A(n18541), .B(n18540), .Z(n18549) );
  AOI22_X1 U20805 ( .A1(n18542), .A2(n18776), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n18774), .ZN(n18543) );
  OAI211_X1 U20806 ( .C1(n13061), .C2(n18791), .A(n18543), .B(n18848), .ZN(
        n18547) );
  INV_X1 U20807 ( .A(n18544), .ZN(n18545) );
  OAI22_X1 U20808 ( .A1(n18545), .A2(n18737), .B1(n19389), .B2(n18780), .ZN(
        n18546) );
  AOI211_X1 U20809 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18794), .A(
        n18547), .B(n18546), .ZN(n18548) );
  OAI21_X1 U20810 ( .B1(n18549), .B2(n18888), .A(n18548), .ZN(P2_U2846) );
  NAND2_X1 U20811 ( .A1(n18550), .A2(n18776), .ZN(n18552) );
  NAND2_X1 U20812 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18794), .ZN(
        n18551) );
  OAI211_X1 U20813 ( .C1(n18553), .C2(n18788), .A(n18552), .B(n18551), .ZN(
        n18554) );
  AOI211_X1 U20814 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n18755), .A(n16675), 
        .B(n18554), .ZN(n18562) );
  AOI21_X1 U20815 ( .B1(n18556), .B2(n18555), .A(n17017), .ZN(n19383) );
  NOR2_X1 U20816 ( .A1(n18783), .A2(n18557), .ZN(n18559) );
  XNOR2_X1 U20817 ( .A(n18559), .B(n18558), .ZN(n18560) );
  AOI22_X1 U20818 ( .A1(n19383), .A2(n18795), .B1(n18784), .B2(n18560), .ZN(
        n18561) );
  OAI211_X1 U20819 ( .C1(n18817), .C2(n18737), .A(n18562), .B(n18561), .ZN(
        P2_U2845) );
  AOI22_X1 U20820 ( .A1(n18774), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18794), .ZN(n18563) );
  OAI21_X1 U20821 ( .B1(n18564), .B2(n18800), .A(n18563), .ZN(n18565) );
  AOI211_X1 U20822 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n18755), .A(n16328), 
        .B(n18565), .ZN(n18572) );
  NAND2_X1 U20823 ( .A1(n11029), .A2(n18566), .ZN(n18567) );
  XNOR2_X1 U20824 ( .A(n18568), .B(n18567), .ZN(n18569) );
  AOI22_X1 U20825 ( .A1(n18570), .A2(n18796), .B1(n18784), .B2(n18569), .ZN(
        n18571) );
  OAI211_X1 U20826 ( .C1(n19382), .C2(n18780), .A(n18572), .B(n18571), .ZN(
        P2_U2844) );
  NOR2_X1 U20827 ( .A1(n18783), .A2(n18573), .ZN(n18575) );
  XOR2_X1 U20828 ( .A(n18575), .B(n18574), .Z(n18583) );
  AOI22_X1 U20829 ( .A1(n18576), .A2(n18776), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n18774), .ZN(n18577) );
  OAI211_X1 U20830 ( .C1(n13071), .C2(n18791), .A(n18577), .B(n18848), .ZN(
        n18578) );
  AOI21_X1 U20831 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18794), .A(
        n18578), .ZN(n18582) );
  AOI22_X1 U20832 ( .A1(n18580), .A2(n18796), .B1(n18579), .B2(n18795), .ZN(
        n18581) );
  OAI211_X1 U20833 ( .C1(n18888), .C2(n18583), .A(n18582), .B(n18581), .ZN(
        P2_U2843) );
  AOI22_X1 U20834 ( .A1(n18774), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18794), .ZN(n18588) );
  OR2_X1 U20835 ( .A1(n18783), .A2(n18584), .ZN(n18596) );
  AOI211_X1 U20836 ( .C1(n18585), .C2(n18591), .A(n18888), .B(n18596), .ZN(
        n18586) );
  INV_X1 U20837 ( .A(n18586), .ZN(n18587) );
  OAI211_X1 U20838 ( .C1(n18800), .C2(n18589), .A(n18588), .B(n18587), .ZN(
        n18590) );
  AOI211_X1 U20839 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18755), .A(n16328), 
        .B(n18590), .ZN(n18594) );
  AOI22_X1 U20840 ( .A1(n18592), .A2(n18796), .B1(n18591), .B2(n18614), .ZN(
        n18593) );
  OAI211_X1 U20841 ( .C1(n19376), .C2(n18780), .A(n18594), .B(n18593), .ZN(
        P2_U2842) );
  XNOR2_X1 U20842 ( .A(n18596), .B(n18595), .ZN(n18603) );
  AOI22_X1 U20843 ( .A1(n18774), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18794), .ZN(n18597) );
  OAI21_X1 U20844 ( .B1(n18598), .B2(n18800), .A(n18597), .ZN(n18599) );
  AOI211_X1 U20845 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18755), .A(n16328), 
        .B(n18599), .ZN(n18602) );
  AOI22_X1 U20846 ( .A1(n18600), .A2(n18796), .B1(n19370), .B2(n18795), .ZN(
        n18601) );
  OAI211_X1 U20847 ( .C1(n18888), .C2(n18603), .A(n18602), .B(n18601), .ZN(
        P2_U2841) );
  OAI22_X1 U20848 ( .A1(n18788), .A2(n18605), .B1(n18765), .B2(n18604), .ZN(
        n18606) );
  INV_X1 U20849 ( .A(n18606), .ZN(n18611) );
  AOI211_X1 U20850 ( .C1(n18608), .C2(n18615), .A(n18888), .B(n18607), .ZN(
        n18609) );
  INV_X1 U20851 ( .A(n18609), .ZN(n18610) );
  OAI211_X1 U20852 ( .C1(n18800), .C2(n18612), .A(n18611), .B(n18610), .ZN(
        n18613) );
  AOI211_X1 U20853 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18755), .A(n16675), 
        .B(n18613), .ZN(n18618) );
  AOI22_X1 U20854 ( .A1(n18616), .A2(n18796), .B1(n18615), .B2(n18614), .ZN(
        n18617) );
  OAI211_X1 U20855 ( .C1(n19369), .C2(n18780), .A(n18618), .B(n18617), .ZN(
        P2_U2840) );
  NAND2_X1 U20856 ( .A1(n11029), .A2(n18619), .ZN(n18620) );
  XOR2_X1 U20857 ( .A(n18621), .B(n18620), .Z(n18631) );
  OAI21_X1 U20858 ( .B1(n18765), .B2(n18622), .A(n18848), .ZN(n18623) );
  AOI21_X1 U20859 ( .B1(n18774), .B2(P2_EBX_REG_17__SCAN_IN), .A(n18623), .ZN(
        n18624) );
  OAI21_X1 U20860 ( .B1(n18791), .B2(n13091), .A(n18624), .ZN(n18625) );
  AOI21_X1 U20861 ( .B1(n18626), .B2(n18776), .A(n18625), .ZN(n18630) );
  AOI22_X1 U20862 ( .A1(n18628), .A2(n18796), .B1(n18627), .B2(n18795), .ZN(
        n18629) );
  OAI211_X1 U20863 ( .C1(n18888), .C2(n18631), .A(n18630), .B(n18629), .ZN(
        P2_U2838) );
  AOI22_X1 U20864 ( .A1(n18774), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18794), .ZN(n18632) );
  OAI21_X1 U20865 ( .B1(n18633), .B2(n18800), .A(n18632), .ZN(n18634) );
  AOI211_X1 U20866 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18755), .A(n16675), 
        .B(n18634), .ZN(n18640) );
  NOR2_X1 U20867 ( .A1(n18783), .A2(n18635), .ZN(n18637) );
  XNOR2_X1 U20868 ( .A(n18637), .B(n18636), .ZN(n18638) );
  AOI22_X1 U20869 ( .A1(n19766), .A2(n18795), .B1(n18784), .B2(n18638), .ZN(
        n18639) );
  OAI211_X1 U20870 ( .C1(n18641), .C2(n18737), .A(n18640), .B(n18639), .ZN(
        P2_U2837) );
  NAND2_X1 U20871 ( .A1(n11029), .A2(n18642), .ZN(n18643) );
  XOR2_X1 U20872 ( .A(n18644), .B(n18643), .Z(n18653) );
  AOI22_X1 U20873 ( .A1(n18645), .A2(n18776), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n18774), .ZN(n18646) );
  OAI211_X1 U20874 ( .C1(n18647), .C2(n18791), .A(n18646), .B(n18848), .ZN(
        n18648) );
  AOI21_X1 U20875 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18794), .A(
        n18648), .ZN(n18652) );
  AOI22_X1 U20876 ( .A1(n18650), .A2(n18796), .B1(n18649), .B2(n18795), .ZN(
        n18651) );
  OAI211_X1 U20877 ( .C1(n18888), .C2(n18653), .A(n18652), .B(n18651), .ZN(
        P2_U2836) );
  NOR2_X1 U20878 ( .A1(n18783), .A2(n18654), .ZN(n18655) );
  XOR2_X1 U20879 ( .A(n18656), .B(n18655), .Z(n18664) );
  INV_X1 U20880 ( .A(n18657), .ZN(n19657) );
  AOI22_X1 U20881 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18794), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18755), .ZN(n18660) );
  AOI22_X1 U20882 ( .A1(n18658), .A2(n18776), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n18774), .ZN(n18659) );
  OAI211_X1 U20883 ( .C1(n18661), .C2(n18737), .A(n18660), .B(n18659), .ZN(
        n18662) );
  AOI21_X1 U20884 ( .B1(n19657), .B2(n18795), .A(n18662), .ZN(n18663) );
  OAI21_X1 U20885 ( .B1(n18888), .B2(n18664), .A(n18663), .ZN(P2_U2835) );
  AOI22_X1 U20886 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18794), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18755), .ZN(n18675) );
  AOI22_X1 U20887 ( .A1(n18665), .A2(n18776), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n18774), .ZN(n18674) );
  AOI22_X1 U20888 ( .A1(n18667), .A2(n18796), .B1(n18666), .B2(n18795), .ZN(
        n18673) );
  AND2_X1 U20889 ( .A1(n11029), .A2(n18668), .ZN(n18670) );
  AOI21_X1 U20890 ( .B1(n18671), .B2(n18670), .A(n18888), .ZN(n18669) );
  OAI21_X1 U20891 ( .B1(n18671), .B2(n18670), .A(n18669), .ZN(n18672) );
  NAND4_X1 U20892 ( .A1(n18675), .A2(n18674), .A3(n18673), .A4(n18672), .ZN(
        P2_U2834) );
  NOR2_X1 U20893 ( .A1(n18783), .A2(n18676), .ZN(n18678) );
  XOR2_X1 U20894 ( .A(n18678), .B(n18677), .Z(n18686) );
  AOI22_X1 U20895 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18794), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18755), .ZN(n18679) );
  OAI21_X1 U20896 ( .B1(n18788), .B2(n18680), .A(n18679), .ZN(n18681) );
  AOI21_X1 U20897 ( .B1(n18682), .B2(n18776), .A(n18681), .ZN(n18685) );
  AOI22_X1 U20898 ( .A1(n18683), .A2(n18796), .B1(n19547), .B2(n18795), .ZN(
        n18684) );
  OAI211_X1 U20899 ( .C1(n18888), .C2(n18686), .A(n18685), .B(n18684), .ZN(
        P2_U2833) );
  OAI22_X1 U20900 ( .A1(n18688), .A2(n18765), .B1(n18687), .B2(n18791), .ZN(
        n18694) );
  AND2_X1 U20901 ( .A1(n11029), .A2(n18689), .ZN(n18692) );
  OAI21_X1 U20902 ( .B1(n18691), .B2(n18692), .A(n18784), .ZN(n18690) );
  AOI21_X1 U20903 ( .B1(n18692), .B2(n18691), .A(n18690), .ZN(n18693) );
  AOI211_X1 U20904 ( .C1(n18774), .C2(P2_EBX_REG_23__SCAN_IN), .A(n18694), .B(
        n18693), .ZN(n18698) );
  AOI22_X1 U20905 ( .A1(n18696), .A2(n18796), .B1(n18695), .B2(n18795), .ZN(
        n18697) );
  OAI211_X1 U20906 ( .C1(n18699), .C2(n18800), .A(n18698), .B(n18697), .ZN(
        P2_U2832) );
  AOI22_X1 U20907 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18794), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18755), .ZN(n18700) );
  INV_X1 U20908 ( .A(n18700), .ZN(n18706) );
  NOR2_X1 U20909 ( .A1(n18783), .A2(n18701), .ZN(n18704) );
  OAI21_X1 U20910 ( .B1(n18703), .B2(n18704), .A(n18784), .ZN(n18702) );
  AOI21_X1 U20911 ( .B1(n18704), .B2(n18703), .A(n18702), .ZN(n18705) );
  AOI211_X1 U20912 ( .C1(n18774), .C2(P2_EBX_REG_24__SCAN_IN), .A(n18706), .B(
        n18705), .ZN(n18710) );
  AOI22_X1 U20913 ( .A1(n18708), .A2(n18776), .B1(n18707), .B2(n18796), .ZN(
        n18709) );
  OAI211_X1 U20914 ( .C1(n18711), .C2(n18780), .A(n18710), .B(n18709), .ZN(
        P2_U2831) );
  AND2_X1 U20915 ( .A1(n11029), .A2(n18712), .ZN(n18714) );
  OAI21_X1 U20916 ( .B1(n18715), .B2(n18714), .A(n18784), .ZN(n18713) );
  AOI21_X1 U20917 ( .B1(n18715), .B2(n18714), .A(n18713), .ZN(n18719) );
  INV_X1 U20918 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n18716) );
  OAI22_X1 U20919 ( .A1(n18791), .A2(n18717), .B1(n18716), .B2(n18788), .ZN(
        n18718) );
  AOI211_X1 U20920 ( .C1(n18794), .C2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n18719), .B(n18718), .ZN(n18723) );
  AOI22_X1 U20921 ( .A1(n18721), .A2(n18776), .B1(n18720), .B2(n18796), .ZN(
        n18722) );
  OAI211_X1 U20922 ( .C1(n18724), .C2(n18780), .A(n18723), .B(n18722), .ZN(
        P2_U2830) );
  NOR2_X1 U20923 ( .A1(n18783), .A2(n18725), .ZN(n18728) );
  OAI21_X1 U20924 ( .B1(n18727), .B2(n18728), .A(n18784), .ZN(n18726) );
  AOI21_X1 U20925 ( .B1(n18728), .B2(n18727), .A(n18726), .ZN(n18732) );
  AOI22_X1 U20926 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18794), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18755), .ZN(n18729) );
  OAI21_X1 U20927 ( .B1(n18788), .B2(n18730), .A(n18729), .ZN(n18731) );
  NOR2_X1 U20928 ( .A1(n18732), .A2(n18731), .ZN(n18736) );
  AOI22_X1 U20929 ( .A1(n18734), .A2(n18776), .B1(n18733), .B2(n18795), .ZN(
        n18735) );
  OAI211_X1 U20930 ( .C1(n18738), .C2(n18737), .A(n18736), .B(n18735), .ZN(
        P2_U2829) );
  OAI22_X1 U20931 ( .A1(n18740), .A2(n18765), .B1(n18739), .B2(n18791), .ZN(
        n18746) );
  AND2_X1 U20932 ( .A1(n11029), .A2(n18741), .ZN(n18744) );
  OAI21_X1 U20933 ( .B1(n18743), .B2(n18744), .A(n18784), .ZN(n18742) );
  AOI21_X1 U20934 ( .B1(n18744), .B2(n18743), .A(n18742), .ZN(n18745) );
  AOI211_X1 U20935 ( .C1(n18774), .C2(P2_EBX_REG_27__SCAN_IN), .A(n18746), .B(
        n18745), .ZN(n18750) );
  AOI22_X1 U20936 ( .A1(n18748), .A2(n18796), .B1(n18747), .B2(n18795), .ZN(
        n18749) );
  OAI211_X1 U20937 ( .C1(n18751), .C2(n18800), .A(n18750), .B(n18749), .ZN(
        P2_U2828) );
  NOR2_X1 U20938 ( .A1(n18783), .A2(n18752), .ZN(n18753) );
  XOR2_X1 U20939 ( .A(n18754), .B(n18753), .Z(n18757) );
  AOI22_X1 U20940 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18794), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18755), .ZN(n18756) );
  OAI21_X1 U20941 ( .B1(n18888), .B2(n18757), .A(n18756), .ZN(n18758) );
  AOI21_X1 U20942 ( .B1(n18774), .B2(P2_EBX_REG_28__SCAN_IN), .A(n18758), .ZN(
        n18762) );
  AOI22_X1 U20943 ( .A1(n18760), .A2(n18796), .B1(n18759), .B2(n18795), .ZN(
        n18761) );
  OAI211_X1 U20944 ( .C1(n18763), .C2(n18800), .A(n18762), .B(n18761), .ZN(
        P2_U2827) );
  OAI22_X1 U20945 ( .A1(n18766), .A2(n18765), .B1(n18764), .B2(n18791), .ZN(
        n18773) );
  AND2_X1 U20946 ( .A1(n11029), .A2(n18767), .ZN(n18771) );
  OAI21_X1 U20947 ( .B1(n18770), .B2(n18771), .A(n18784), .ZN(n18769) );
  AOI21_X1 U20948 ( .B1(n18771), .B2(n18770), .A(n18769), .ZN(n18772) );
  AOI211_X1 U20949 ( .C1(n18774), .C2(P2_EBX_REG_29__SCAN_IN), .A(n18773), .B(
        n18772), .ZN(n18779) );
  AOI22_X1 U20950 ( .A1(n18777), .A2(n18776), .B1(n18775), .B2(n18796), .ZN(
        n18778) );
  OAI211_X1 U20951 ( .C1(n18781), .C2(n18780), .A(n18779), .B(n18778), .ZN(
        P2_U2826) );
  OR2_X1 U20952 ( .A1(n18783), .A2(n18782), .ZN(n18786) );
  OAI21_X1 U20953 ( .B1(n18787), .B2(n18786), .A(n18784), .ZN(n18785) );
  AOI21_X1 U20954 ( .B1(n18787), .B2(n18786), .A(n18785), .ZN(n18793) );
  OAI22_X1 U20955 ( .A1(n18791), .A2(n18790), .B1(n18789), .B2(n18788), .ZN(
        n18792) );
  AOI211_X1 U20956 ( .C1(n18794), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n18793), .B(n18792), .ZN(n18799) );
  AOI22_X1 U20957 ( .A1(n18797), .A2(n18796), .B1(n16751), .B2(n18795), .ZN(
        n18798) );
  OAI211_X1 U20958 ( .C1(n18801), .C2(n18800), .A(n18799), .B(n18798), .ZN(
        P2_U2825) );
  OAI22_X1 U20959 ( .A1(n18869), .A2(n18803), .B1(n18870), .B2(n18802), .ZN(
        n18807) );
  OAI22_X1 U20960 ( .A1(n18805), .A2(n18849), .B1(n17048), .B2(n18804), .ZN(
        n18806) );
  AOI211_X1 U20961 ( .C1(n17048), .C2(n18808), .A(n18807), .B(n18806), .ZN(
        n18810) );
  OAI211_X1 U20962 ( .C1(n18811), .C2(n18881), .A(n18810), .B(n18809), .ZN(
        P2_U3046) );
  NAND2_X1 U20963 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n16675), .ZN(n18812) );
  OAI211_X1 U20964 ( .C1(n18815), .C2(n18814), .A(n18813), .B(n18812), .ZN(
        n18816) );
  AOI21_X1 U20965 ( .B1(n18852), .B2(n19383), .A(n18816), .ZN(n18821) );
  INV_X1 U20966 ( .A(n18817), .ZN(n18818) );
  AOI22_X1 U20967 ( .A1(n18819), .A2(n18825), .B1(n14189), .B2(n18818), .ZN(
        n18820) );
  OAI211_X1 U20968 ( .C1(n18822), .C2(n18869), .A(n18821), .B(n18820), .ZN(
        P2_U3036) );
  AOI22_X1 U20969 ( .A1(n18823), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n18852), .B2(n19390), .ZN(n18833) );
  AOI222_X1 U20970 ( .A1(n18827), .A2(n18856), .B1(n14189), .B2(n18826), .C1(
        n18825), .C2(n18824), .ZN(n18832) );
  NAND2_X1 U20971 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16328), .ZN(n18831) );
  OAI211_X1 U20972 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18829), .B(n18828), .ZN(n18830) );
  NAND4_X1 U20973 ( .A1(n18833), .A2(n18832), .A3(n18831), .A4(n18830), .ZN(
        P2_U3038) );
  INV_X1 U20974 ( .A(n18834), .ZN(n18843) );
  OAI22_X1 U20975 ( .A1(n18870), .A2(n19663), .B1(n18848), .B2(n18835), .ZN(
        n18836) );
  AOI21_X1 U20976 ( .B1(n18837), .B2(n14189), .A(n18836), .ZN(n18838) );
  OAI21_X1 U20977 ( .B1(n18839), .B2(n18881), .A(n18838), .ZN(n18840) );
  AOI21_X1 U20978 ( .B1(n18856), .B2(n18841), .A(n18840), .ZN(n18842) );
  OAI221_X1 U20979 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18845), .C1(
        n18844), .C2(n18843), .A(n18842), .ZN(P2_U3042) );
  NAND2_X1 U20980 ( .A1(n18847), .A2(n18846), .ZN(n18861) );
  OAI22_X1 U20981 ( .A1(n18850), .A2(n18849), .B1(n16366), .B2(n18848), .ZN(
        n18851) );
  AOI21_X1 U20982 ( .B1(n19712), .B2(n18852), .A(n18851), .ZN(n18853) );
  OAI21_X1 U20983 ( .B1(n18854), .B2(n18881), .A(n18853), .ZN(n18855) );
  AOI21_X1 U20984 ( .B1(n18857), .B2(n18856), .A(n18855), .ZN(n18858) );
  OAI221_X1 U20985 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18861), .C1(
        n18860), .C2(n18859), .A(n18858), .ZN(P2_U3043) );
  AOI21_X1 U20986 ( .B1(n18863), .B2(n14189), .A(n18862), .ZN(n18867) );
  NAND2_X1 U20987 ( .A1(n18865), .A2(n18864), .ZN(n18866) );
  OAI211_X1 U20988 ( .C1(n18869), .C2(n18868), .A(n18867), .B(n18866), .ZN(
        n18873) );
  INV_X1 U20989 ( .A(n19608), .ZN(n18871) );
  NOR2_X1 U20990 ( .A1(n18871), .A2(n18870), .ZN(n18872) );
  AOI211_X1 U20991 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n18874), .A(
        n18873), .B(n18872), .ZN(n18879) );
  OAI21_X1 U20992 ( .B1(n18877), .B2(n18876), .A(n18875), .ZN(n18878) );
  OAI211_X1 U20993 ( .C1(n18881), .C2(n18880), .A(n18879), .B(n18878), .ZN(
        P2_U3044) );
  NAND2_X1 U20994 ( .A1(n18896), .A2(n18882), .ZN(n18898) );
  NAND2_X1 U20995 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18899), .ZN(n18884) );
  OAI21_X1 U20996 ( .B1(n18884), .B2(n18883), .A(n18904), .ZN(n18887) );
  NAND2_X1 U20997 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21883), .ZN(n18885) );
  AOI21_X1 U20998 ( .B1(n18891), .B2(n18898), .A(n18885), .ZN(n18886) );
  AOI21_X1 U20999 ( .B1(n18898), .B2(n18887), .A(n18886), .ZN(n18889) );
  NAND2_X1 U21000 ( .A1(n18889), .A2(n18888), .ZN(P2_U3177) );
  AOI21_X1 U21001 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n18890), .A(n21883), 
        .ZN(n18892) );
  OAI22_X1 U21002 ( .A1(n18894), .A2(n18893), .B1(n18892), .B2(n18891), .ZN(
        n18895) );
  AOI21_X1 U21003 ( .B1(n18896), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n18895), 
        .ZN(n18903) );
  NOR2_X1 U21004 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18897), .ZN(n18901) );
  OAI22_X1 U21005 ( .A1(n18901), .A2(n18900), .B1(n18899), .B2(n18898), .ZN(
        n18902) );
  OAI211_X1 U21006 ( .C1(n18905), .C2(n18904), .A(n18903), .B(n18902), .ZN(
        P2_U3176) );
  NAND2_X1 U21007 ( .A1(n18907), .A2(n18906), .ZN(n18910) );
  NAND2_X1 U21008 ( .A1(n18910), .A2(P2_MORE_REG_SCAN_IN), .ZN(n18908) );
  OAI21_X1 U21009 ( .B1(n18910), .B2(n18909), .A(n18908), .ZN(P2_U3609) );
  INV_X1 U21010 ( .A(n18910), .ZN(n18913) );
  OAI21_X1 U21011 ( .B1(n18913), .B2(n18912), .A(n18911), .ZN(P2_U2819) );
  INV_X1 U21012 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20310) );
  INV_X1 U21013 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n20898) );
  AOI22_X1 U21014 ( .A1(n19261), .A2(n20310), .B1(n20898), .B2(U215), .ZN(U282) );
  OAI22_X1 U21015 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19261), .ZN(n18914) );
  INV_X1 U21016 ( .A(n18914), .ZN(U281) );
  OAI22_X1 U21017 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19261), .ZN(n18915) );
  INV_X1 U21018 ( .A(n18915), .ZN(U280) );
  OAI22_X1 U21019 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19261), .ZN(n18916) );
  INV_X1 U21020 ( .A(n18916), .ZN(U279) );
  OAI22_X1 U21021 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19261), .ZN(n18917) );
  INV_X1 U21022 ( .A(n18917), .ZN(U278) );
  OAI22_X1 U21023 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19261), .ZN(n18918) );
  INV_X1 U21024 ( .A(n18918), .ZN(U277) );
  OAI22_X1 U21025 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19261), .ZN(n18919) );
  INV_X1 U21026 ( .A(n18919), .ZN(U276) );
  OAI22_X1 U21027 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19261), .ZN(n18920) );
  INV_X1 U21028 ( .A(n18920), .ZN(U275) );
  OAI22_X1 U21029 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19261), .ZN(n18921) );
  INV_X1 U21030 ( .A(n18921), .ZN(U274) );
  OAI22_X1 U21031 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19261), .ZN(n18922) );
  INV_X1 U21032 ( .A(n18922), .ZN(U273) );
  OAI22_X1 U21033 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19261), .ZN(n18923) );
  INV_X1 U21034 ( .A(n18923), .ZN(U272) );
  OAI22_X1 U21035 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19261), .ZN(n18924) );
  INV_X1 U21036 ( .A(n18924), .ZN(U271) );
  OAI22_X1 U21037 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18937), .ZN(n18925) );
  INV_X1 U21038 ( .A(n18925), .ZN(U270) );
  OAI22_X1 U21039 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19261), .ZN(n18926) );
  INV_X1 U21040 ( .A(n18926), .ZN(U269) );
  OAI22_X1 U21041 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18937), .ZN(n18927) );
  INV_X1 U21042 ( .A(n18927), .ZN(U268) );
  OAI22_X1 U21043 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19261), .ZN(n18928) );
  INV_X1 U21044 ( .A(n18928), .ZN(U267) );
  OAI22_X1 U21045 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18937), .ZN(n18929) );
  INV_X1 U21046 ( .A(n18929), .ZN(U266) );
  OAI22_X1 U21047 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19261), .ZN(n18930) );
  INV_X1 U21048 ( .A(n18930), .ZN(U265) );
  OAI22_X1 U21049 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n18937), .ZN(n18931) );
  INV_X1 U21050 ( .A(n18931), .ZN(U264) );
  OAI22_X1 U21051 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n18937), .ZN(n18932) );
  INV_X1 U21052 ( .A(n18932), .ZN(U263) );
  OAI22_X1 U21053 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n18937), .ZN(n18933) );
  INV_X1 U21054 ( .A(n18933), .ZN(U262) );
  OAI22_X1 U21055 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n18937), .ZN(n18934) );
  INV_X1 U21056 ( .A(n18934), .ZN(U261) );
  OAI22_X1 U21057 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n18937), .ZN(n18935) );
  INV_X1 U21058 ( .A(n18935), .ZN(U260) );
  OAI22_X1 U21059 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18937), .ZN(n18936) );
  INV_X1 U21060 ( .A(n18936), .ZN(U259) );
  OAI22_X1 U21061 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n18937), .ZN(n18938) );
  INV_X1 U21062 ( .A(n18938), .ZN(U258) );
  NOR2_X1 U21063 ( .A1(n18975), .A2(n18939), .ZN(n19004) );
  NAND2_X1 U21064 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19004), .ZN(
        n19345) );
  NOR2_X1 U21065 ( .A1(n18941), .A2(n18940), .ZN(n19055) );
  NAND2_X1 U21066 ( .A1(n19055), .A2(n20809), .ZN(n19015) );
  NOR3_X1 U21067 ( .A1(n21398), .A2(n18975), .A3(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18947) );
  NAND2_X1 U21068 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18947), .ZN(
        n19271) );
  INV_X1 U21069 ( .A(n19271), .ZN(n19357) );
  AND2_X1 U21070 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19264), .ZN(n19008) );
  INV_X1 U21071 ( .A(n18992), .ZN(n21418) );
  AND2_X1 U21072 ( .A1(n21418), .A2(n19004), .ZN(n19266) );
  INV_X1 U21073 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20934) );
  NOR2_X2 U21074 ( .A1(n20934), .A2(n19176), .ZN(n19007) );
  AOI22_X1 U21075 ( .A1(n19357), .A2(n19008), .B1(n19266), .B2(n19007), .ZN(
        n18944) );
  NOR2_X1 U21076 ( .A1(n18942), .A2(n19176), .ZN(n18962) );
  AOI22_X1 U21077 ( .A1(n19264), .A2(n18947), .B1(n19004), .B2(n18962), .ZN(
        n19268) );
  NAND2_X1 U21078 ( .A1(n18980), .A2(n18947), .ZN(n19182) );
  INV_X1 U21079 ( .A(n19182), .ZN(n19283) );
  NOR2_X2 U21080 ( .A1(n20898), .A2(n18333), .ZN(n19012) );
  AOI22_X1 U21081 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19268), .B1(
        n19283), .B2(n19012), .ZN(n18943) );
  OAI211_X1 U21082 ( .C1(n19345), .C2(n19015), .A(n18944), .B(n18943), .ZN(
        P3_U2995) );
  NAND2_X1 U21083 ( .A1(n19004), .A2(n18980), .ZN(n19364) );
  NOR2_X1 U21084 ( .A1(n21388), .A2(n18961), .ZN(n18953) );
  NAND2_X1 U21085 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18953), .ZN(
        n19281) );
  INV_X1 U21086 ( .A(n19281), .ZN(n19290) );
  NAND2_X1 U21087 ( .A1(n19271), .A2(n19364), .ZN(n19011) );
  AND2_X1 U21088 ( .A1(n21418), .A2(n19011), .ZN(n19272) );
  AOI22_X1 U21089 ( .A1(n19012), .A2(n19290), .B1(n19007), .B2(n19272), .ZN(
        n18946) );
  NAND2_X1 U21090 ( .A1(n19182), .A2(n19281), .ZN(n18950) );
  AOI21_X1 U21091 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19176), .ZN(n19010) );
  AOI22_X1 U21092 ( .A1(n19264), .A2(n18950), .B1(n19010), .B2(n19011), .ZN(
        n19274) );
  AOI22_X1 U21093 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19274), .B1(
        n19283), .B2(n19008), .ZN(n18945) );
  OAI211_X1 U21094 ( .C1(n19015), .C2(n19364), .A(n18946), .B(n18945), .ZN(
        P3_U2987) );
  AND2_X1 U21095 ( .A1(n21418), .A2(n18947), .ZN(n19277) );
  AOI22_X1 U21096 ( .A1(n19008), .A2(n19290), .B1(n19007), .B2(n19277), .ZN(
        n18949) );
  AOI22_X1 U21097 ( .A1(n19264), .A2(n18953), .B1(n18962), .B2(n18947), .ZN(
        n19278) );
  NAND2_X1 U21098 ( .A1(n18980), .A2(n18953), .ZN(n19229) );
  INV_X1 U21099 ( .A(n19229), .ZN(n19294) );
  AOI22_X1 U21100 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19278), .B1(
        n19012), .B2(n19294), .ZN(n18948) );
  OAI211_X1 U21101 ( .C1(n19015), .C2(n19271), .A(n18949), .B(n18948), .ZN(
        P3_U2979) );
  AND2_X1 U21102 ( .A1(n21418), .A2(n18950), .ZN(n19282) );
  AOI22_X1 U21103 ( .A1(n19008), .A2(n19294), .B1(n19007), .B2(n19282), .ZN(
        n18952) );
  NAND2_X1 U21104 ( .A1(n21388), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18986) );
  NOR2_X2 U21105 ( .A1(n18961), .A2(n18986), .ZN(n19300) );
  INV_X1 U21106 ( .A(n19300), .ZN(n19287) );
  NAND2_X1 U21107 ( .A1(n19229), .A2(n19287), .ZN(n18958) );
  AOI22_X1 U21108 ( .A1(n19264), .A2(n18958), .B1(n19010), .B2(n18950), .ZN(
        n19284) );
  AOI22_X1 U21109 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19284), .B1(
        n19012), .B2(n19300), .ZN(n18951) );
  OAI211_X1 U21110 ( .C1(n19182), .C2(n19015), .A(n18952), .B(n18951), .ZN(
        P3_U2971) );
  INV_X1 U21111 ( .A(n18953), .ZN(n18954) );
  NOR2_X1 U21112 ( .A1(n18992), .A2(n18954), .ZN(n19288) );
  AOI22_X1 U21113 ( .A1(n19008), .A2(n19300), .B1(n19007), .B2(n19288), .ZN(
        n18957) );
  INV_X1 U21114 ( .A(n18961), .ZN(n18963) );
  NAND2_X1 U21115 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21387) );
  AOI211_X1 U21116 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(n21387), .A(n18955), 
        .B(n19176), .ZN(n18993) );
  NAND2_X1 U21117 ( .A1(n18963), .A2(n18993), .ZN(n19289) );
  NAND2_X1 U21118 ( .A1(n21388), .A2(n18980), .ZN(n21391) );
  NOR2_X2 U21119 ( .A1(n21391), .A2(n18961), .ZN(n19306) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19289), .B1(
        n19012), .B2(n19306), .ZN(n18956) );
  OAI211_X1 U21121 ( .C1(n19015), .C2(n19281), .A(n18957), .B(n18956), .ZN(
        P3_U2963) );
  NAND2_X1 U21122 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18970), .ZN(
        n19191) );
  INV_X1 U21123 ( .A(n19191), .ZN(n19311) );
  AND2_X1 U21124 ( .A1(n21418), .A2(n18958), .ZN(n19293) );
  AOI22_X1 U21125 ( .A1(n19012), .A2(n19311), .B1(n19007), .B2(n19293), .ZN(
        n18960) );
  NAND2_X1 U21126 ( .A1(n19298), .A2(n19191), .ZN(n18967) );
  AOI22_X1 U21127 ( .A1(n19264), .A2(n18967), .B1(n19010), .B2(n18958), .ZN(
        n19295) );
  AOI22_X1 U21128 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19295), .B1(
        n19008), .B2(n19306), .ZN(n18959) );
  OAI211_X1 U21129 ( .C1(n19015), .C2(n19229), .A(n18960), .B(n18959), .ZN(
        P3_U2955) );
  NAND2_X1 U21130 ( .A1(n18980), .A2(n18970), .ZN(n19304) );
  INV_X1 U21131 ( .A(n19304), .ZN(n19317) );
  NAND2_X1 U21132 ( .A1(n21388), .A2(n21418), .ZN(n19001) );
  NOR2_X1 U21133 ( .A1(n18961), .A2(n19001), .ZN(n19299) );
  AOI22_X1 U21134 ( .A1(n19012), .A2(n19317), .B1(n19007), .B2(n19299), .ZN(
        n18965) );
  AND2_X1 U21135 ( .A1(n21388), .A2(n18962), .ZN(n19003) );
  AOI22_X1 U21136 ( .A1(n19264), .A2(n18970), .B1(n18963), .B2(n19003), .ZN(
        n19301) );
  AOI22_X1 U21137 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19301), .B1(
        n19008), .B2(n19311), .ZN(n18964) );
  OAI211_X1 U21138 ( .C1(n19015), .C2(n19287), .A(n18965), .B(n18964), .ZN(
        P3_U2947) );
  INV_X1 U21139 ( .A(n18986), .ZN(n18966) );
  NAND2_X1 U21140 ( .A1(n18966), .A2(n18982), .ZN(n19315) );
  INV_X1 U21141 ( .A(n19315), .ZN(n19323) );
  AND2_X1 U21142 ( .A1(n21418), .A2(n18967), .ZN(n19305) );
  AOI22_X1 U21143 ( .A1(n19012), .A2(n19323), .B1(n19007), .B2(n19305), .ZN(
        n18969) );
  NAND2_X1 U21144 ( .A1(n19304), .A2(n19315), .ZN(n18974) );
  AOI22_X1 U21145 ( .A1(n19264), .A2(n18974), .B1(n19010), .B2(n18967), .ZN(
        n19307) );
  AOI22_X1 U21146 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19307), .B1(
        n19008), .B2(n19317), .ZN(n18968) );
  OAI211_X1 U21147 ( .C1(n19015), .C2(n19298), .A(n18969), .B(n18968), .ZN(
        P3_U2939) );
  NAND2_X1 U21148 ( .A1(n18993), .A2(n18982), .ZN(n19312) );
  INV_X1 U21149 ( .A(n18970), .ZN(n18971) );
  NOR2_X1 U21150 ( .A1(n18992), .A2(n18971), .ZN(n19310) );
  AOI22_X1 U21151 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19312), .B1(
        n19007), .B2(n19310), .ZN(n18973) );
  NOR2_X2 U21152 ( .A1(n21391), .A2(n18981), .ZN(n19329) );
  AOI22_X1 U21153 ( .A1(n19012), .A2(n19329), .B1(n19008), .B2(n19323), .ZN(
        n18972) );
  OAI211_X1 U21154 ( .C1(n19015), .C2(n19191), .A(n18973), .B(n18972), .ZN(
        P3_U2931) );
  AND2_X1 U21155 ( .A1(n21418), .A2(n18974), .ZN(n19316) );
  AOI22_X1 U21156 ( .A1(n19008), .A2(n19329), .B1(n19007), .B2(n19316), .ZN(
        n18979) );
  NAND2_X1 U21157 ( .A1(n21398), .A2(n18975), .ZN(n19000) );
  NOR2_X1 U21158 ( .A1(n21388), .A2(n19000), .ZN(n18990) );
  NAND2_X1 U21159 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18990), .ZN(
        n19327) );
  NAND2_X1 U21160 ( .A1(n19321), .A2(n19327), .ZN(n18987) );
  INV_X1 U21161 ( .A(n18987), .ZN(n18985) );
  OAI22_X1 U21162 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19315), .B1(n18985), 
        .B2(n18976), .ZN(n18977) );
  OAI21_X1 U21163 ( .B1(n19317), .B2(n18977), .A(n19265), .ZN(n19318) );
  INV_X1 U21164 ( .A(n19327), .ZN(n19335) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19318), .B1(
        n19012), .B2(n19335), .ZN(n18978) );
  OAI211_X1 U21166 ( .C1(n19015), .C2(n19304), .A(n18979), .B(n18978), .ZN(
        P3_U2923) );
  NAND2_X1 U21167 ( .A1(n18980), .A2(n18990), .ZN(n19244) );
  NOR2_X1 U21168 ( .A1(n19001), .A2(n18981), .ZN(n19322) );
  AOI22_X1 U21169 ( .A1(n19012), .A2(n19341), .B1(n19007), .B2(n19322), .ZN(
        n18984) );
  AOI22_X1 U21170 ( .A1(n19264), .A2(n18990), .B1(n19003), .B2(n18982), .ZN(
        n19324) );
  AOI22_X1 U21171 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19324), .B1(
        n19008), .B2(n19335), .ZN(n18983) );
  OAI211_X1 U21172 ( .C1(n19015), .C2(n19315), .A(n18984), .B(n18983), .ZN(
        P3_U2915) );
  NOR2_X1 U21173 ( .A1(n18992), .A2(n18985), .ZN(n19328) );
  AOI22_X1 U21174 ( .A1(n19008), .A2(n19341), .B1(n19007), .B2(n19328), .ZN(
        n18989) );
  NOR2_X2 U21175 ( .A1(n18986), .A2(n19000), .ZN(n19349) );
  INV_X1 U21176 ( .A(n19349), .ZN(n19333) );
  NAND2_X1 U21177 ( .A1(n19244), .A2(n19333), .ZN(n18996) );
  AOI22_X1 U21178 ( .A1(n19264), .A2(n18996), .B1(n19010), .B2(n18987), .ZN(
        n19330) );
  AOI22_X1 U21179 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19330), .B1(
        n19012), .B2(n19349), .ZN(n18988) );
  OAI211_X1 U21180 ( .C1(n19015), .C2(n19321), .A(n18989), .B(n18988), .ZN(
        P3_U2907) );
  INV_X1 U21181 ( .A(n18990), .ZN(n18991) );
  NOR2_X1 U21182 ( .A1(n18992), .A2(n18991), .ZN(n19334) );
  AOI22_X1 U21183 ( .A1(n19008), .A2(n19349), .B1(n19007), .B2(n19334), .ZN(
        n18995) );
  INV_X1 U21184 ( .A(n19000), .ZN(n19002) );
  NAND2_X1 U21185 ( .A1(n18993), .A2(n19002), .ZN(n19336) );
  NOR2_X2 U21186 ( .A1(n21391), .A2(n19000), .ZN(n19359) );
  AOI22_X1 U21187 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19336), .B1(
        n19012), .B2(n19359), .ZN(n18994) );
  OAI211_X1 U21188 ( .C1(n19015), .C2(n19327), .A(n18995), .B(n18994), .ZN(
        P3_U2899) );
  AND2_X1 U21189 ( .A1(n21418), .A2(n18996), .ZN(n19340) );
  AOI22_X1 U21190 ( .A1(n19008), .A2(n19359), .B1(n19007), .B2(n19340), .ZN(
        n18999) );
  OAI21_X1 U21191 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19333), .A(n19244), 
        .ZN(n18997) );
  NAND2_X1 U21192 ( .A1(n19345), .A2(n19339), .ZN(n19009) );
  AOI22_X1 U21193 ( .A1(n19265), .A2(n18997), .B1(n19264), .B2(n19009), .ZN(
        n19342) );
  INV_X1 U21194 ( .A(n19345), .ZN(n19348) );
  AOI22_X1 U21195 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19342), .B1(
        n19012), .B2(n19348), .ZN(n18998) );
  OAI211_X1 U21196 ( .C1(n19015), .C2(n19244), .A(n18999), .B(n18998), .ZN(
        P3_U2891) );
  INV_X1 U21197 ( .A(n19364), .ZN(n19273) );
  NOR2_X1 U21198 ( .A1(n19001), .A2(n19000), .ZN(n19346) );
  AOI22_X1 U21199 ( .A1(n19012), .A2(n19273), .B1(n19007), .B2(n19346), .ZN(
        n19006) );
  AOI22_X1 U21200 ( .A1(n19264), .A2(n19004), .B1(n19003), .B2(n19002), .ZN(
        n19350) );
  AOI22_X1 U21201 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19350), .B1(
        n19348), .B2(n19008), .ZN(n19005) );
  OAI211_X1 U21202 ( .C1(n19015), .C2(n19333), .A(n19006), .B(n19005), .ZN(
        P3_U2883) );
  AND2_X1 U21203 ( .A1(n21418), .A2(n19009), .ZN(n19355) );
  AOI22_X1 U21204 ( .A1(n19008), .A2(n19273), .B1(n19007), .B2(n19355), .ZN(
        n19014) );
  AOI22_X1 U21205 ( .A1(n19264), .A2(n19011), .B1(n19010), .B2(n19009), .ZN(
        n19360) );
  AOI22_X1 U21206 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19360), .B1(
        n19012), .B2(n19357), .ZN(n19013) );
  OAI211_X1 U21207 ( .C1(n19015), .C2(n19339), .A(n19014), .B(n19013), .ZN(
        P3_U2875) );
  OAI22_X1 U21208 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19261), .ZN(n19016) );
  INV_X1 U21209 ( .A(n19016), .ZN(U257) );
  NAND2_X1 U21210 ( .A1(n19055), .A2(n19017), .ZN(n19053) );
  NOR2_X2 U21211 ( .A1(n15699), .A2(n18333), .ZN(n19049) );
  NOR2_X2 U21212 ( .A1(n20865), .A2(n19176), .ZN(n19048) );
  AOI22_X1 U21213 ( .A1(n19283), .A2(n19049), .B1(n19266), .B2(n19048), .ZN(
        n19019) );
  INV_X1 U21214 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n20853) );
  NOR2_X2 U21215 ( .A1(n20853), .A2(n18333), .ZN(n19050) );
  AOI22_X1 U21216 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19268), .B1(
        n19357), .B2(n19050), .ZN(n19018) );
  OAI211_X1 U21217 ( .C1(n19345), .C2(n19053), .A(n19019), .B(n19018), .ZN(
        P3_U2994) );
  AOI22_X1 U21218 ( .A1(n19283), .A2(n19050), .B1(n19272), .B2(n19048), .ZN(
        n19021) );
  AOI22_X1 U21219 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19274), .B1(
        n19290), .B2(n19049), .ZN(n19020) );
  OAI211_X1 U21220 ( .C1(n19364), .C2(n19053), .A(n19021), .B(n19020), .ZN(
        P3_U2986) );
  AOI22_X1 U21221 ( .A1(n19290), .A2(n19050), .B1(n19277), .B2(n19048), .ZN(
        n19023) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19278), .B1(
        n19294), .B2(n19049), .ZN(n19022) );
  OAI211_X1 U21223 ( .C1(n19271), .C2(n19053), .A(n19023), .B(n19022), .ZN(
        P3_U2978) );
  AOI22_X1 U21224 ( .A1(n19300), .A2(n19049), .B1(n19282), .B2(n19048), .ZN(
        n19025) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19284), .B1(
        n19294), .B2(n19050), .ZN(n19024) );
  OAI211_X1 U21226 ( .C1(n19182), .C2(n19053), .A(n19025), .B(n19024), .ZN(
        P3_U2970) );
  AOI22_X1 U21227 ( .A1(n19306), .A2(n19049), .B1(n19288), .B2(n19048), .ZN(
        n19027) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19289), .B1(
        n19300), .B2(n19050), .ZN(n19026) );
  OAI211_X1 U21229 ( .C1(n19281), .C2(n19053), .A(n19027), .B(n19026), .ZN(
        P3_U2962) );
  AOI22_X1 U21230 ( .A1(n19306), .A2(n19050), .B1(n19293), .B2(n19048), .ZN(
        n19029) );
  AOI22_X1 U21231 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19295), .B1(
        n19311), .B2(n19049), .ZN(n19028) );
  OAI211_X1 U21232 ( .C1(n19229), .C2(n19053), .A(n19029), .B(n19028), .ZN(
        P3_U2954) );
  AOI22_X1 U21233 ( .A1(n19299), .A2(n19048), .B1(n19317), .B2(n19049), .ZN(
        n19031) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19301), .B1(
        n19311), .B2(n19050), .ZN(n19030) );
  OAI211_X1 U21235 ( .C1(n19287), .C2(n19053), .A(n19031), .B(n19030), .ZN(
        P3_U2946) );
  AOI22_X1 U21236 ( .A1(n19323), .A2(n19049), .B1(n19305), .B2(n19048), .ZN(
        n19033) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19307), .B1(
        n19317), .B2(n19050), .ZN(n19032) );
  OAI211_X1 U21238 ( .C1(n19298), .C2(n19053), .A(n19033), .B(n19032), .ZN(
        P3_U2938) );
  AOI22_X1 U21239 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19312), .B1(
        n19310), .B2(n19048), .ZN(n19035) );
  AOI22_X1 U21240 ( .A1(n19323), .A2(n19050), .B1(n19329), .B2(n19049), .ZN(
        n19034) );
  OAI211_X1 U21241 ( .C1(n19191), .C2(n19053), .A(n19035), .B(n19034), .ZN(
        P3_U2930) );
  AOI22_X1 U21242 ( .A1(n19329), .A2(n19050), .B1(n19316), .B2(n19048), .ZN(
        n19037) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19318), .B1(
        n19335), .B2(n19049), .ZN(n19036) );
  OAI211_X1 U21244 ( .C1(n19304), .C2(n19053), .A(n19037), .B(n19036), .ZN(
        P3_U2922) );
  AOI22_X1 U21245 ( .A1(n19335), .A2(n19050), .B1(n19322), .B2(n19048), .ZN(
        n19039) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19324), .B1(
        n19341), .B2(n19049), .ZN(n19038) );
  OAI211_X1 U21247 ( .C1(n19315), .C2(n19053), .A(n19039), .B(n19038), .ZN(
        P3_U2914) );
  AOI22_X1 U21248 ( .A1(n19341), .A2(n19050), .B1(n19328), .B2(n19048), .ZN(
        n19041) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19330), .B1(
        n19349), .B2(n19049), .ZN(n19040) );
  OAI211_X1 U21250 ( .C1(n19321), .C2(n19053), .A(n19041), .B(n19040), .ZN(
        P3_U2906) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19336), .B1(
        n19334), .B2(n19048), .ZN(n19043) );
  AOI22_X1 U21252 ( .A1(n19349), .A2(n19050), .B1(n19359), .B2(n19049), .ZN(
        n19042) );
  OAI211_X1 U21253 ( .C1(n19327), .C2(n19053), .A(n19043), .B(n19042), .ZN(
        P3_U2898) );
  AOI22_X1 U21254 ( .A1(n19348), .A2(n19049), .B1(n19340), .B2(n19048), .ZN(
        n19045) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19342), .B1(
        n19359), .B2(n19050), .ZN(n19044) );
  OAI211_X1 U21256 ( .C1(n19244), .C2(n19053), .A(n19045), .B(n19044), .ZN(
        P3_U2890) );
  AOI22_X1 U21257 ( .A1(n19273), .A2(n19049), .B1(n19346), .B2(n19048), .ZN(
        n19047) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19350), .B1(
        n19348), .B2(n19050), .ZN(n19046) );
  OAI211_X1 U21259 ( .C1(n19333), .C2(n19053), .A(n19047), .B(n19046), .ZN(
        P3_U2882) );
  AOI22_X1 U21260 ( .A1(n19357), .A2(n19049), .B1(n19355), .B2(n19048), .ZN(
        n19052) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19360), .B1(
        n19273), .B2(n19050), .ZN(n19051) );
  OAI211_X1 U21262 ( .C1(n19339), .C2(n19053), .A(n19052), .B(n19051), .ZN(
        P3_U2874) );
  OAI22_X1 U21263 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19261), .ZN(n19054) );
  INV_X1 U21264 ( .A(n19054), .ZN(U256) );
  NAND2_X1 U21265 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n19264), .ZN(n19085) );
  NAND2_X1 U21266 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19264), .ZN(n19093) );
  INV_X1 U21267 ( .A(n19093), .ZN(n19082) );
  INV_X1 U21268 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20848) );
  NOR2_X2 U21269 ( .A1(n20848), .A2(n19176), .ZN(n19088) );
  AOI22_X1 U21270 ( .A1(n19283), .A2(n19082), .B1(n19266), .B2(n19088), .ZN(
        n19057) );
  INV_X1 U21271 ( .A(n19055), .ZN(n19267) );
  NOR2_X2 U21272 ( .A1(n20840), .A2(n19267), .ZN(n19090) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19268), .B1(
        n19348), .B2(n19090), .ZN(n19056) );
  OAI211_X1 U21274 ( .C1(n19271), .C2(n19085), .A(n19057), .B(n19056), .ZN(
        P3_U2993) );
  INV_X1 U21275 ( .A(n19085), .ZN(n19089) );
  AOI22_X1 U21276 ( .A1(n19283), .A2(n19089), .B1(n19272), .B2(n19088), .ZN(
        n19059) );
  AOI22_X1 U21277 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19090), .ZN(n19058) );
  OAI211_X1 U21278 ( .C1(n19281), .C2(n19093), .A(n19059), .B(n19058), .ZN(
        P3_U2985) );
  AOI22_X1 U21279 ( .A1(n19290), .A2(n19089), .B1(n19277), .B2(n19088), .ZN(
        n19061) );
  AOI22_X1 U21280 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19278), .B1(
        n19357), .B2(n19090), .ZN(n19060) );
  OAI211_X1 U21281 ( .C1(n19229), .C2(n19093), .A(n19061), .B(n19060), .ZN(
        P3_U2977) );
  AOI22_X1 U21282 ( .A1(n19300), .A2(n19082), .B1(n19282), .B2(n19088), .ZN(
        n19063) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19090), .ZN(n19062) );
  OAI211_X1 U21284 ( .C1(n19229), .C2(n19085), .A(n19063), .B(n19062), .ZN(
        P3_U2969) );
  AOI22_X1 U21285 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19289), .B1(
        n19288), .B2(n19088), .ZN(n19065) );
  AOI22_X1 U21286 ( .A1(n19290), .A2(n19090), .B1(n19300), .B2(n19089), .ZN(
        n19064) );
  OAI211_X1 U21287 ( .C1(n19298), .C2(n19093), .A(n19065), .B(n19064), .ZN(
        P3_U2961) );
  AOI22_X1 U21288 ( .A1(n19311), .A2(n19082), .B1(n19293), .B2(n19088), .ZN(
        n19067) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19295), .B1(
        n19294), .B2(n19090), .ZN(n19066) );
  OAI211_X1 U21290 ( .C1(n19298), .C2(n19085), .A(n19067), .B(n19066), .ZN(
        P3_U2953) );
  AOI22_X1 U21291 ( .A1(n19299), .A2(n19088), .B1(n19317), .B2(n19082), .ZN(
        n19069) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19301), .B1(
        n19300), .B2(n19090), .ZN(n19068) );
  OAI211_X1 U21293 ( .C1(n19191), .C2(n19085), .A(n19069), .B(n19068), .ZN(
        P3_U2945) );
  AOI22_X1 U21294 ( .A1(n19323), .A2(n19082), .B1(n19305), .B2(n19088), .ZN(
        n19071) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19307), .B1(
        n19306), .B2(n19090), .ZN(n19070) );
  OAI211_X1 U21296 ( .C1(n19304), .C2(n19085), .A(n19071), .B(n19070), .ZN(
        P3_U2937) );
  AOI22_X1 U21297 ( .A1(n19323), .A2(n19089), .B1(n19310), .B2(n19088), .ZN(
        n19073) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19090), .ZN(n19072) );
  OAI211_X1 U21299 ( .C1(n19321), .C2(n19093), .A(n19073), .B(n19072), .ZN(
        P3_U2929) );
  AOI22_X1 U21300 ( .A1(n19335), .A2(n19082), .B1(n19316), .B2(n19088), .ZN(
        n19075) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19318), .B1(
        n19317), .B2(n19090), .ZN(n19074) );
  OAI211_X1 U21302 ( .C1(n19321), .C2(n19085), .A(n19075), .B(n19074), .ZN(
        P3_U2921) );
  AOI22_X1 U21303 ( .A1(n19341), .A2(n19082), .B1(n19322), .B2(n19088), .ZN(
        n19077) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19090), .ZN(n19076) );
  OAI211_X1 U21305 ( .C1(n19327), .C2(n19085), .A(n19077), .B(n19076), .ZN(
        P3_U2913) );
  AOI22_X1 U21306 ( .A1(n19341), .A2(n19089), .B1(n19328), .B2(n19088), .ZN(
        n19079) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19090), .ZN(n19078) );
  OAI211_X1 U21308 ( .C1(n19333), .C2(n19093), .A(n19079), .B(n19078), .ZN(
        P3_U2905) );
  AOI22_X1 U21309 ( .A1(n19349), .A2(n19089), .B1(n19334), .B2(n19088), .ZN(
        n19081) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19336), .B1(
        n19335), .B2(n19090), .ZN(n19080) );
  OAI211_X1 U21311 ( .C1(n19339), .C2(n19093), .A(n19081), .B(n19080), .ZN(
        P3_U2897) );
  AOI22_X1 U21312 ( .A1(n19348), .A2(n19082), .B1(n19340), .B2(n19088), .ZN(
        n19084) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19090), .ZN(n19083) );
  OAI211_X1 U21314 ( .C1(n19339), .C2(n19085), .A(n19084), .B(n19083), .ZN(
        P3_U2889) );
  AOI22_X1 U21315 ( .A1(n19348), .A2(n19089), .B1(n19346), .B2(n19088), .ZN(
        n19087) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19090), .ZN(n19086) );
  OAI211_X1 U21317 ( .C1(n19364), .C2(n19093), .A(n19087), .B(n19086), .ZN(
        P3_U2881) );
  AOI22_X1 U21318 ( .A1(n19273), .A2(n19089), .B1(n19355), .B2(n19088), .ZN(
        n19092) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19090), .ZN(n19091) );
  OAI211_X1 U21320 ( .C1(n19271), .C2(n19093), .A(n19092), .B(n19091), .ZN(
        P3_U2873) );
  OAI22_X1 U21321 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19261), .ZN(n19094) );
  INV_X1 U21322 ( .A(n19094), .ZN(U255) );
  NOR2_X1 U21323 ( .A1(n16486), .A2(n18333), .ZN(n19122) );
  NAND2_X1 U21324 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n19264), .ZN(n19125) );
  INV_X1 U21325 ( .A(n19125), .ZN(n19129) );
  NOR2_X2 U21326 ( .A1(n20829), .A2(n19176), .ZN(n19128) );
  AOI22_X1 U21327 ( .A1(n19357), .A2(n19129), .B1(n19266), .B2(n19128), .ZN(
        n19097) );
  NOR2_X2 U21328 ( .A1(n19095), .A2(n19267), .ZN(n19130) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19268), .B1(
        n19348), .B2(n19130), .ZN(n19096) );
  OAI211_X1 U21330 ( .C1(n19182), .C2(n19133), .A(n19097), .B(n19096), .ZN(
        P3_U2992) );
  AOI22_X1 U21331 ( .A1(n19290), .A2(n19122), .B1(n19272), .B2(n19128), .ZN(
        n19099) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19130), .ZN(n19098) );
  OAI211_X1 U21333 ( .C1(n19182), .C2(n19125), .A(n19099), .B(n19098), .ZN(
        P3_U2984) );
  AOI22_X1 U21334 ( .A1(n19294), .A2(n19122), .B1(n19277), .B2(n19128), .ZN(
        n19101) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19278), .B1(
        n19357), .B2(n19130), .ZN(n19100) );
  OAI211_X1 U21336 ( .C1(n19281), .C2(n19125), .A(n19101), .B(n19100), .ZN(
        P3_U2976) );
  AOI22_X1 U21337 ( .A1(n19294), .A2(n19129), .B1(n19282), .B2(n19128), .ZN(
        n19103) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19130), .ZN(n19102) );
  OAI211_X1 U21339 ( .C1(n19287), .C2(n19133), .A(n19103), .B(n19102), .ZN(
        P3_U2968) );
  AOI22_X1 U21340 ( .A1(n19300), .A2(n19129), .B1(n19288), .B2(n19128), .ZN(
        n19105) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19289), .B1(
        n19290), .B2(n19130), .ZN(n19104) );
  OAI211_X1 U21342 ( .C1(n19298), .C2(n19133), .A(n19105), .B(n19104), .ZN(
        P3_U2960) );
  AOI22_X1 U21343 ( .A1(n19306), .A2(n19129), .B1(n19293), .B2(n19128), .ZN(
        n19107) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19295), .B1(
        n19294), .B2(n19130), .ZN(n19106) );
  OAI211_X1 U21345 ( .C1(n19191), .C2(n19133), .A(n19107), .B(n19106), .ZN(
        P3_U2952) );
  AOI22_X1 U21346 ( .A1(n19311), .A2(n19129), .B1(n19299), .B2(n19128), .ZN(
        n19109) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19301), .B1(
        n19300), .B2(n19130), .ZN(n19108) );
  OAI211_X1 U21348 ( .C1(n19304), .C2(n19133), .A(n19109), .B(n19108), .ZN(
        P3_U2944) );
  AOI22_X1 U21349 ( .A1(n19317), .A2(n19129), .B1(n19305), .B2(n19128), .ZN(
        n19111) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19307), .B1(
        n19306), .B2(n19130), .ZN(n19110) );
  OAI211_X1 U21351 ( .C1(n19315), .C2(n19133), .A(n19111), .B(n19110), .ZN(
        P3_U2936) );
  AOI22_X1 U21352 ( .A1(n19329), .A2(n19122), .B1(n19310), .B2(n19128), .ZN(
        n19113) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19130), .ZN(n19112) );
  OAI211_X1 U21354 ( .C1(n19315), .C2(n19125), .A(n19113), .B(n19112), .ZN(
        P3_U2928) );
  AOI22_X1 U21355 ( .A1(n19329), .A2(n19129), .B1(n19316), .B2(n19128), .ZN(
        n19115) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19318), .B1(
        n19317), .B2(n19130), .ZN(n19114) );
  OAI211_X1 U21357 ( .C1(n19327), .C2(n19133), .A(n19115), .B(n19114), .ZN(
        P3_U2920) );
  AOI22_X1 U21358 ( .A1(n19335), .A2(n19129), .B1(n19322), .B2(n19128), .ZN(
        n19117) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19130), .ZN(n19116) );
  OAI211_X1 U21360 ( .C1(n19244), .C2(n19133), .A(n19117), .B(n19116), .ZN(
        P3_U2912) );
  AOI22_X1 U21361 ( .A1(n19341), .A2(n19129), .B1(n19328), .B2(n19128), .ZN(
        n19119) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19130), .ZN(n19118) );
  OAI211_X1 U21363 ( .C1(n19333), .C2(n19133), .A(n19119), .B(n19118), .ZN(
        P3_U2904) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19336), .B1(
        n19334), .B2(n19128), .ZN(n19121) );
  AOI22_X1 U21365 ( .A1(n19335), .A2(n19130), .B1(n19359), .B2(n19122), .ZN(
        n19120) );
  OAI211_X1 U21366 ( .C1(n19333), .C2(n19125), .A(n19121), .B(n19120), .ZN(
        P3_U2896) );
  AOI22_X1 U21367 ( .A1(n19348), .A2(n19122), .B1(n19340), .B2(n19128), .ZN(
        n19124) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19130), .ZN(n19123) );
  OAI211_X1 U21369 ( .C1(n19339), .C2(n19125), .A(n19124), .B(n19123), .ZN(
        P3_U2888) );
  AOI22_X1 U21370 ( .A1(n19348), .A2(n19129), .B1(n19346), .B2(n19128), .ZN(
        n19127) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19130), .ZN(n19126) );
  OAI211_X1 U21372 ( .C1(n19364), .C2(n19133), .A(n19127), .B(n19126), .ZN(
        P3_U2880) );
  AOI22_X1 U21373 ( .A1(n19273), .A2(n19129), .B1(n19355), .B2(n19128), .ZN(
        n19132) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19130), .ZN(n19131) );
  OAI211_X1 U21375 ( .C1(n19271), .C2(n19133), .A(n19132), .B(n19131), .ZN(
        P3_U2872) );
  OAI22_X1 U21376 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19261), .ZN(n19134) );
  INV_X1 U21377 ( .A(n19134), .ZN(U254) );
  NAND2_X1 U21378 ( .A1(n19264), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19167) );
  NAND2_X1 U21379 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19264), .ZN(n19173) );
  INV_X1 U21380 ( .A(n19173), .ZN(n19164) );
  INV_X1 U21381 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n20833) );
  NOR2_X2 U21382 ( .A1(n19176), .A2(n20833), .ZN(n19168) );
  AOI22_X1 U21383 ( .A1(n19283), .A2(n19164), .B1(n19266), .B2(n19168), .ZN(
        n19137) );
  NOR2_X2 U21384 ( .A1(n19135), .A2(n19267), .ZN(n19170) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19268), .B1(
        n19348), .B2(n19170), .ZN(n19136) );
  OAI211_X1 U21386 ( .C1(n19271), .C2(n19167), .A(n19137), .B(n19136), .ZN(
        P3_U2991) );
  AOI22_X1 U21387 ( .A1(n19290), .A2(n19164), .B1(n19272), .B2(n19168), .ZN(
        n19139) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19170), .ZN(n19138) );
  OAI211_X1 U21389 ( .C1(n19182), .C2(n19167), .A(n19139), .B(n19138), .ZN(
        P3_U2983) );
  INV_X1 U21390 ( .A(n19167), .ZN(n19169) );
  AOI22_X1 U21391 ( .A1(n19290), .A2(n19169), .B1(n19277), .B2(n19168), .ZN(
        n19141) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19278), .B1(
        n19357), .B2(n19170), .ZN(n19140) );
  OAI211_X1 U21393 ( .C1(n19229), .C2(n19173), .A(n19141), .B(n19140), .ZN(
        P3_U2975) );
  AOI22_X1 U21394 ( .A1(n19300), .A2(n19164), .B1(n19282), .B2(n19168), .ZN(
        n19143) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19170), .ZN(n19142) );
  OAI211_X1 U21396 ( .C1(n19229), .C2(n19167), .A(n19143), .B(n19142), .ZN(
        P3_U2967) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19289), .B1(
        n19288), .B2(n19168), .ZN(n19145) );
  AOI22_X1 U21398 ( .A1(n19290), .A2(n19170), .B1(n19300), .B2(n19169), .ZN(
        n19144) );
  OAI211_X1 U21399 ( .C1(n19298), .C2(n19173), .A(n19145), .B(n19144), .ZN(
        P3_U2959) );
  AOI22_X1 U21400 ( .A1(n19311), .A2(n19164), .B1(n19293), .B2(n19168), .ZN(
        n19147) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19295), .B1(
        n19294), .B2(n19170), .ZN(n19146) );
  OAI211_X1 U21402 ( .C1(n19298), .C2(n19167), .A(n19147), .B(n19146), .ZN(
        P3_U2951) );
  AOI22_X1 U21403 ( .A1(n19299), .A2(n19168), .B1(n19317), .B2(n19164), .ZN(
        n19149) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19301), .B1(
        n19300), .B2(n19170), .ZN(n19148) );
  OAI211_X1 U21405 ( .C1(n19191), .C2(n19167), .A(n19149), .B(n19148), .ZN(
        P3_U2943) );
  AOI22_X1 U21406 ( .A1(n19323), .A2(n19164), .B1(n19305), .B2(n19168), .ZN(
        n19151) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19307), .B1(
        n19306), .B2(n19170), .ZN(n19150) );
  OAI211_X1 U21408 ( .C1(n19304), .C2(n19167), .A(n19151), .B(n19150), .ZN(
        P3_U2935) );
  AOI22_X1 U21409 ( .A1(n19323), .A2(n19169), .B1(n19310), .B2(n19168), .ZN(
        n19153) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19170), .ZN(n19152) );
  OAI211_X1 U21411 ( .C1(n19321), .C2(n19173), .A(n19153), .B(n19152), .ZN(
        P3_U2927) );
  AOI22_X1 U21412 ( .A1(n19329), .A2(n19169), .B1(n19316), .B2(n19168), .ZN(
        n19155) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19318), .B1(
        n19317), .B2(n19170), .ZN(n19154) );
  OAI211_X1 U21414 ( .C1(n19327), .C2(n19173), .A(n19155), .B(n19154), .ZN(
        P3_U2919) );
  AOI22_X1 U21415 ( .A1(n19335), .A2(n19169), .B1(n19322), .B2(n19168), .ZN(
        n19157) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19170), .ZN(n19156) );
  OAI211_X1 U21417 ( .C1(n19244), .C2(n19173), .A(n19157), .B(n19156), .ZN(
        P3_U2911) );
  AOI22_X1 U21418 ( .A1(n19341), .A2(n19169), .B1(n19328), .B2(n19168), .ZN(
        n19159) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19170), .ZN(n19158) );
  OAI211_X1 U21420 ( .C1(n19333), .C2(n19173), .A(n19159), .B(n19158), .ZN(
        P3_U2903) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19336), .B1(
        n19334), .B2(n19168), .ZN(n19161) );
  AOI22_X1 U21422 ( .A1(n19335), .A2(n19170), .B1(n19349), .B2(n19169), .ZN(
        n19160) );
  OAI211_X1 U21423 ( .C1(n19339), .C2(n19173), .A(n19161), .B(n19160), .ZN(
        P3_U2895) );
  AOI22_X1 U21424 ( .A1(n19359), .A2(n19169), .B1(n19340), .B2(n19168), .ZN(
        n19163) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19170), .ZN(n19162) );
  OAI211_X1 U21426 ( .C1(n19345), .C2(n19173), .A(n19163), .B(n19162), .ZN(
        P3_U2887) );
  AOI22_X1 U21427 ( .A1(n19273), .A2(n19164), .B1(n19346), .B2(n19168), .ZN(
        n19166) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19170), .ZN(n19165) );
  OAI211_X1 U21429 ( .C1(n19345), .C2(n19167), .A(n19166), .B(n19165), .ZN(
        P3_U2879) );
  AOI22_X1 U21430 ( .A1(n19273), .A2(n19169), .B1(n19355), .B2(n19168), .ZN(
        n19172) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19170), .ZN(n19171) );
  OAI211_X1 U21432 ( .C1(n19271), .C2(n19173), .A(n19172), .B(n19171), .ZN(
        P3_U2871) );
  OAI22_X1 U21433 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19261), .ZN(n19174) );
  INV_X1 U21434 ( .A(n19174), .ZN(U253) );
  INV_X1 U21435 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19175) );
  NOR2_X1 U21436 ( .A1(n18333), .A2(n19175), .ZN(n19204) );
  INV_X1 U21437 ( .A(n19204), .ZN(n19217) );
  NAND2_X1 U21438 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19264), .ZN(n19207) );
  INV_X1 U21439 ( .A(n19207), .ZN(n19213) );
  INV_X1 U21440 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n20876) );
  NOR2_X2 U21441 ( .A1(n19176), .A2(n20876), .ZN(n19212) );
  AOI22_X1 U21442 ( .A1(n19283), .A2(n19213), .B1(n19266), .B2(n19212), .ZN(
        n19179) );
  NOR2_X2 U21443 ( .A1(n19177), .A2(n19267), .ZN(n19214) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19268), .B1(
        n19348), .B2(n19214), .ZN(n19178) );
  OAI211_X1 U21445 ( .C1(n19271), .C2(n19217), .A(n19179), .B(n19178), .ZN(
        P3_U2990) );
  AOI22_X1 U21446 ( .A1(n19290), .A2(n19213), .B1(n19272), .B2(n19212), .ZN(
        n19181) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19214), .ZN(n19180) );
  OAI211_X1 U21448 ( .C1(n19182), .C2(n19217), .A(n19181), .B(n19180), .ZN(
        P3_U2982) );
  AOI22_X1 U21449 ( .A1(n19294), .A2(n19213), .B1(n19277), .B2(n19212), .ZN(
        n19184) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19278), .B1(
        n19357), .B2(n19214), .ZN(n19183) );
  OAI211_X1 U21451 ( .C1(n19281), .C2(n19217), .A(n19184), .B(n19183), .ZN(
        P3_U2974) );
  AOI22_X1 U21452 ( .A1(n19300), .A2(n19213), .B1(n19282), .B2(n19212), .ZN(
        n19186) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19214), .ZN(n19185) );
  OAI211_X1 U21454 ( .C1(n19229), .C2(n19217), .A(n19186), .B(n19185), .ZN(
        P3_U2966) );
  AOI22_X1 U21455 ( .A1(n19300), .A2(n19204), .B1(n19288), .B2(n19212), .ZN(
        n19188) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19289), .B1(
        n19290), .B2(n19214), .ZN(n19187) );
  OAI211_X1 U21457 ( .C1(n19298), .C2(n19207), .A(n19188), .B(n19187), .ZN(
        P3_U2958) );
  AOI22_X1 U21458 ( .A1(n19306), .A2(n19204), .B1(n19293), .B2(n19212), .ZN(
        n19190) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19295), .B1(
        n19294), .B2(n19214), .ZN(n19189) );
  OAI211_X1 U21460 ( .C1(n19191), .C2(n19207), .A(n19190), .B(n19189), .ZN(
        P3_U2950) );
  AOI22_X1 U21461 ( .A1(n19311), .A2(n19204), .B1(n19299), .B2(n19212), .ZN(
        n19193) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19301), .B1(
        n19300), .B2(n19214), .ZN(n19192) );
  OAI211_X1 U21463 ( .C1(n19304), .C2(n19207), .A(n19193), .B(n19192), .ZN(
        P3_U2942) );
  AOI22_X1 U21464 ( .A1(n19323), .A2(n19213), .B1(n19305), .B2(n19212), .ZN(
        n19195) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19307), .B1(
        n19306), .B2(n19214), .ZN(n19194) );
  OAI211_X1 U21466 ( .C1(n19304), .C2(n19217), .A(n19195), .B(n19194), .ZN(
        P3_U2934) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19312), .B1(
        n19310), .B2(n19212), .ZN(n19197) );
  AOI22_X1 U21468 ( .A1(n19311), .A2(n19214), .B1(n19323), .B2(n19204), .ZN(
        n19196) );
  OAI211_X1 U21469 ( .C1(n19321), .C2(n19207), .A(n19197), .B(n19196), .ZN(
        P3_U2926) );
  AOI22_X1 U21470 ( .A1(n19329), .A2(n19204), .B1(n19316), .B2(n19212), .ZN(
        n19199) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19318), .B1(
        n19317), .B2(n19214), .ZN(n19198) );
  OAI211_X1 U21472 ( .C1(n19327), .C2(n19207), .A(n19199), .B(n19198), .ZN(
        P3_U2918) );
  AOI22_X1 U21473 ( .A1(n19335), .A2(n19204), .B1(n19322), .B2(n19212), .ZN(
        n19201) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19214), .ZN(n19200) );
  OAI211_X1 U21475 ( .C1(n19244), .C2(n19207), .A(n19201), .B(n19200), .ZN(
        P3_U2910) );
  AOI22_X1 U21476 ( .A1(n19349), .A2(n19213), .B1(n19328), .B2(n19212), .ZN(
        n19203) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19214), .ZN(n19202) );
  OAI211_X1 U21478 ( .C1(n19244), .C2(n19217), .A(n19203), .B(n19202), .ZN(
        P3_U2902) );
  AOI22_X1 U21479 ( .A1(n19349), .A2(n19204), .B1(n19334), .B2(n19212), .ZN(
        n19206) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19336), .B1(
        n19335), .B2(n19214), .ZN(n19205) );
  OAI211_X1 U21481 ( .C1(n19339), .C2(n19207), .A(n19206), .B(n19205), .ZN(
        P3_U2894) );
  AOI22_X1 U21482 ( .A1(n19348), .A2(n19213), .B1(n19340), .B2(n19212), .ZN(
        n19209) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19214), .ZN(n19208) );
  OAI211_X1 U21484 ( .C1(n19339), .C2(n19217), .A(n19209), .B(n19208), .ZN(
        P3_U2886) );
  AOI22_X1 U21485 ( .A1(n19273), .A2(n19213), .B1(n19346), .B2(n19212), .ZN(
        n19211) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19214), .ZN(n19210) );
  OAI211_X1 U21487 ( .C1(n19345), .C2(n19217), .A(n19211), .B(n19210), .ZN(
        P3_U2878) );
  AOI22_X1 U21488 ( .A1(n19357), .A2(n19213), .B1(n19355), .B2(n19212), .ZN(
        n19216) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19214), .ZN(n19215) );
  OAI211_X1 U21490 ( .C1(n19364), .C2(n19217), .A(n19216), .B(n19215), .ZN(
        P3_U2870) );
  OAI22_X1 U21491 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19261), .ZN(n19218) );
  INV_X1 U21492 ( .A(n19218), .ZN(U252) );
  INV_X1 U21493 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19219) );
  NOR2_X1 U21494 ( .A1(n18333), .A2(n19219), .ZN(n19256) );
  INV_X1 U21495 ( .A(n19256), .ZN(n19254) );
  NAND2_X1 U21496 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19264), .ZN(n19260) );
  INV_X1 U21497 ( .A(n19260), .ZN(n19251) );
  AND2_X1 U21498 ( .A1(n19265), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19255) );
  AOI22_X1 U21499 ( .A1(n19283), .A2(n19251), .B1(n19266), .B2(n19255), .ZN(
        n19222) );
  NOR2_X2 U21500 ( .A1(n19220), .A2(n19267), .ZN(n19257) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19268), .B1(
        n19348), .B2(n19257), .ZN(n19221) );
  OAI211_X1 U21502 ( .C1(n19271), .C2(n19254), .A(n19222), .B(n19221), .ZN(
        P3_U2989) );
  AOI22_X1 U21503 ( .A1(n19283), .A2(n19256), .B1(n19272), .B2(n19255), .ZN(
        n19224) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19257), .ZN(n19223) );
  OAI211_X1 U21505 ( .C1(n19281), .C2(n19260), .A(n19224), .B(n19223), .ZN(
        P3_U2981) );
  AOI22_X1 U21506 ( .A1(n19294), .A2(n19251), .B1(n19277), .B2(n19255), .ZN(
        n19226) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19278), .B1(
        n19357), .B2(n19257), .ZN(n19225) );
  OAI211_X1 U21508 ( .C1(n19281), .C2(n19254), .A(n19226), .B(n19225), .ZN(
        P3_U2973) );
  AOI22_X1 U21509 ( .A1(n19300), .A2(n19251), .B1(n19282), .B2(n19255), .ZN(
        n19228) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19257), .ZN(n19227) );
  OAI211_X1 U21511 ( .C1(n19229), .C2(n19254), .A(n19228), .B(n19227), .ZN(
        P3_U2965) );
  AOI22_X1 U21512 ( .A1(n19306), .A2(n19251), .B1(n19288), .B2(n19255), .ZN(
        n19231) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19289), .B1(
        n19290), .B2(n19257), .ZN(n19230) );
  OAI211_X1 U21514 ( .C1(n19287), .C2(n19254), .A(n19231), .B(n19230), .ZN(
        P3_U2957) );
  AOI22_X1 U21515 ( .A1(n19311), .A2(n19251), .B1(n19293), .B2(n19255), .ZN(
        n19233) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19295), .B1(
        n19294), .B2(n19257), .ZN(n19232) );
  OAI211_X1 U21517 ( .C1(n19298), .C2(n19254), .A(n19233), .B(n19232), .ZN(
        P3_U2949) );
  AOI22_X1 U21518 ( .A1(n19311), .A2(n19256), .B1(n19299), .B2(n19255), .ZN(
        n19235) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19301), .B1(
        n19300), .B2(n19257), .ZN(n19234) );
  OAI211_X1 U21520 ( .C1(n19304), .C2(n19260), .A(n19235), .B(n19234), .ZN(
        P3_U2941) );
  AOI22_X1 U21521 ( .A1(n19323), .A2(n19251), .B1(n19305), .B2(n19255), .ZN(
        n19237) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19307), .B1(
        n19306), .B2(n19257), .ZN(n19236) );
  OAI211_X1 U21523 ( .C1(n19304), .C2(n19254), .A(n19237), .B(n19236), .ZN(
        P3_U2933) );
  AOI22_X1 U21524 ( .A1(n19323), .A2(n19256), .B1(n19310), .B2(n19255), .ZN(
        n19239) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19257), .ZN(n19238) );
  OAI211_X1 U21526 ( .C1(n19321), .C2(n19260), .A(n19239), .B(n19238), .ZN(
        P3_U2925) );
  AOI22_X1 U21527 ( .A1(n19329), .A2(n19256), .B1(n19316), .B2(n19255), .ZN(
        n19241) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19318), .B1(
        n19317), .B2(n19257), .ZN(n19240) );
  OAI211_X1 U21529 ( .C1(n19327), .C2(n19260), .A(n19241), .B(n19240), .ZN(
        P3_U2917) );
  AOI22_X1 U21530 ( .A1(n19335), .A2(n19256), .B1(n19322), .B2(n19255), .ZN(
        n19243) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19257), .ZN(n19242) );
  OAI211_X1 U21532 ( .C1(n19244), .C2(n19260), .A(n19243), .B(n19242), .ZN(
        P3_U2909) );
  AOI22_X1 U21533 ( .A1(n19341), .A2(n19256), .B1(n19328), .B2(n19255), .ZN(
        n19246) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19257), .ZN(n19245) );
  OAI211_X1 U21535 ( .C1(n19333), .C2(n19260), .A(n19246), .B(n19245), .ZN(
        P3_U2901) );
  AOI22_X1 U21536 ( .A1(n19349), .A2(n19256), .B1(n19334), .B2(n19255), .ZN(
        n19248) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19336), .B1(
        n19335), .B2(n19257), .ZN(n19247) );
  OAI211_X1 U21538 ( .C1(n19339), .C2(n19260), .A(n19248), .B(n19247), .ZN(
        P3_U2893) );
  AOI22_X1 U21539 ( .A1(n19348), .A2(n19251), .B1(n19340), .B2(n19255), .ZN(
        n19250) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19257), .ZN(n19249) );
  OAI211_X1 U21541 ( .C1(n19339), .C2(n19254), .A(n19250), .B(n19249), .ZN(
        P3_U2885) );
  AOI22_X1 U21542 ( .A1(n19273), .A2(n19251), .B1(n19346), .B2(n19255), .ZN(
        n19253) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19257), .ZN(n19252) );
  OAI211_X1 U21544 ( .C1(n19345), .C2(n19254), .A(n19253), .B(n19252), .ZN(
        P3_U2877) );
  AOI22_X1 U21545 ( .A1(n19273), .A2(n19256), .B1(n19355), .B2(n19255), .ZN(
        n19259) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19257), .ZN(n19258) );
  OAI211_X1 U21547 ( .C1(n19271), .C2(n19260), .A(n19259), .B(n19258), .ZN(
        P3_U2869) );
  OAI22_X1 U21548 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19261), .ZN(n19263) );
  INV_X1 U21549 ( .A(n19263), .ZN(U251) );
  NAND2_X1 U21550 ( .A1(n19264), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19363) );
  NAND2_X1 U21551 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19264), .ZN(n19353) );
  INV_X1 U21552 ( .A(n19353), .ZN(n19356) );
  AND2_X1 U21553 ( .A1(n19265), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19354) );
  AOI22_X1 U21554 ( .A1(n19283), .A2(n19356), .B1(n19266), .B2(n19354), .ZN(
        n19270) );
  NOR2_X2 U21555 ( .A1(n20370), .A2(n19267), .ZN(n19358) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19268), .B1(
        n19348), .B2(n19358), .ZN(n19269) );
  OAI211_X1 U21557 ( .C1(n19271), .C2(n19363), .A(n19270), .B(n19269), .ZN(
        P3_U2988) );
  INV_X1 U21558 ( .A(n19363), .ZN(n19347) );
  AOI22_X1 U21559 ( .A1(n19283), .A2(n19347), .B1(n19272), .B2(n19354), .ZN(
        n19276) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19358), .ZN(n19275) );
  OAI211_X1 U21561 ( .C1(n19281), .C2(n19353), .A(n19276), .B(n19275), .ZN(
        P3_U2980) );
  AOI22_X1 U21562 ( .A1(n19294), .A2(n19356), .B1(n19277), .B2(n19354), .ZN(
        n19280) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19278), .B1(
        n19357), .B2(n19358), .ZN(n19279) );
  OAI211_X1 U21564 ( .C1(n19281), .C2(n19363), .A(n19280), .B(n19279), .ZN(
        P3_U2972) );
  AOI22_X1 U21565 ( .A1(n19294), .A2(n19347), .B1(n19282), .B2(n19354), .ZN(
        n19286) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19284), .B1(
        n19283), .B2(n19358), .ZN(n19285) );
  OAI211_X1 U21567 ( .C1(n19287), .C2(n19353), .A(n19286), .B(n19285), .ZN(
        P3_U2964) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19289), .B1(
        n19288), .B2(n19354), .ZN(n19292) );
  AOI22_X1 U21569 ( .A1(n19290), .A2(n19358), .B1(n19300), .B2(n19347), .ZN(
        n19291) );
  OAI211_X1 U21570 ( .C1(n19298), .C2(n19353), .A(n19292), .B(n19291), .ZN(
        P3_U2956) );
  AOI22_X1 U21571 ( .A1(n19311), .A2(n19356), .B1(n19293), .B2(n19354), .ZN(
        n19297) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19295), .B1(
        n19294), .B2(n19358), .ZN(n19296) );
  OAI211_X1 U21573 ( .C1(n19298), .C2(n19363), .A(n19297), .B(n19296), .ZN(
        P3_U2948) );
  AOI22_X1 U21574 ( .A1(n19311), .A2(n19347), .B1(n19299), .B2(n19354), .ZN(
        n19303) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19301), .B1(
        n19300), .B2(n19358), .ZN(n19302) );
  OAI211_X1 U21576 ( .C1(n19304), .C2(n19353), .A(n19303), .B(n19302), .ZN(
        P3_U2940) );
  AOI22_X1 U21577 ( .A1(n19317), .A2(n19347), .B1(n19305), .B2(n19354), .ZN(
        n19309) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19307), .B1(
        n19306), .B2(n19358), .ZN(n19308) );
  OAI211_X1 U21579 ( .C1(n19315), .C2(n19353), .A(n19309), .B(n19308), .ZN(
        P3_U2932) );
  AOI22_X1 U21580 ( .A1(n19329), .A2(n19356), .B1(n19310), .B2(n19354), .ZN(
        n19314) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19312), .B1(
        n19311), .B2(n19358), .ZN(n19313) );
  OAI211_X1 U21582 ( .C1(n19315), .C2(n19363), .A(n19314), .B(n19313), .ZN(
        P3_U2924) );
  AOI22_X1 U21583 ( .A1(n19335), .A2(n19356), .B1(n19316), .B2(n19354), .ZN(
        n19320) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19318), .B1(
        n19317), .B2(n19358), .ZN(n19319) );
  OAI211_X1 U21585 ( .C1(n19321), .C2(n19363), .A(n19320), .B(n19319), .ZN(
        P3_U2916) );
  AOI22_X1 U21586 ( .A1(n19341), .A2(n19356), .B1(n19322), .B2(n19354), .ZN(
        n19326) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19358), .ZN(n19325) );
  OAI211_X1 U21588 ( .C1(n19327), .C2(n19363), .A(n19326), .B(n19325), .ZN(
        P3_U2908) );
  AOI22_X1 U21589 ( .A1(n19341), .A2(n19347), .B1(n19328), .B2(n19354), .ZN(
        n19332) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19358), .ZN(n19331) );
  OAI211_X1 U21591 ( .C1(n19333), .C2(n19353), .A(n19332), .B(n19331), .ZN(
        P3_U2900) );
  AOI22_X1 U21592 ( .A1(n19349), .A2(n19347), .B1(n19334), .B2(n19354), .ZN(
        n19338) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19336), .B1(
        n19335), .B2(n19358), .ZN(n19337) );
  OAI211_X1 U21594 ( .C1(n19339), .C2(n19353), .A(n19338), .B(n19337), .ZN(
        P3_U2892) );
  AOI22_X1 U21595 ( .A1(n19359), .A2(n19347), .B1(n19340), .B2(n19354), .ZN(
        n19344) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19342), .B1(
        n19341), .B2(n19358), .ZN(n19343) );
  OAI211_X1 U21597 ( .C1(n19345), .C2(n19353), .A(n19344), .B(n19343), .ZN(
        P3_U2884) );
  AOI22_X1 U21598 ( .A1(n19348), .A2(n19347), .B1(n19346), .B2(n19354), .ZN(
        n19352) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19358), .ZN(n19351) );
  OAI211_X1 U21600 ( .C1(n19364), .C2(n19353), .A(n19352), .B(n19351), .ZN(
        P3_U2876) );
  AOI22_X1 U21601 ( .A1(n19357), .A2(n19356), .B1(n19355), .B2(n19354), .ZN(
        n19362) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19358), .ZN(n19361) );
  OAI211_X1 U21603 ( .C1(n19364), .C2(n19363), .A(n19362), .B(n19361), .ZN(
        P3_U2868) );
  INV_X1 U21604 ( .A(n16341), .ZN(n19365) );
  AOI22_X1 U21605 ( .A1(n19365), .A2(n19860), .B1(n19764), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19367) );
  AOI22_X1 U21606 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19859), .B1(n19765), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19366) );
  NAND2_X1 U21607 ( .A1(n19367), .A2(n19366), .ZN(P2_U2888) );
  OAI222_X1 U21608 ( .A1(n19369), .A2(n19620), .B1(n14281), .B2(n19556), .C1(
        n19368), .C2(n19868), .ZN(P2_U2904) );
  INV_X1 U21609 ( .A(n19370), .ZN(n19373) );
  OAI222_X1 U21610 ( .A1(n19373), .A2(n19620), .B1(n19372), .B2(n19556), .C1(
        n19868), .C2(n19371), .ZN(P2_U2905) );
  OAI222_X1 U21611 ( .A1(n19376), .A2(n19620), .B1(n19375), .B2(n19556), .C1(
        n19868), .C2(n19374), .ZN(P2_U2906) );
  OAI222_X1 U21612 ( .A1(n19379), .A2(n19620), .B1(n19378), .B2(n19556), .C1(
        n19868), .C2(n19377), .ZN(P2_U2907) );
  OAI222_X1 U21613 ( .A1(n19382), .A2(n19620), .B1(n19381), .B2(n19556), .C1(
        n19868), .C2(n19380), .ZN(P2_U2908) );
  INV_X1 U21614 ( .A(n19383), .ZN(n19386) );
  AOI22_X1 U21615 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19859), .B1(n19384), 
        .B2(n19606), .ZN(n19385) );
  OAI21_X1 U21616 ( .B1(n19620), .B2(n19386), .A(n19385), .ZN(P2_U2909) );
  OAI222_X1 U21617 ( .A1(n19389), .A2(n19620), .B1(n19388), .B2(n19556), .C1(
        n19868), .C2(n19387), .ZN(P2_U2910) );
  INV_X1 U21618 ( .A(n19390), .ZN(n19393) );
  OAI222_X1 U21619 ( .A1(n19393), .A2(n19620), .B1(n19392), .B2(n19556), .C1(
        n19868), .C2(n19391), .ZN(P2_U2911) );
  OAI222_X1 U21620 ( .A1(n19396), .A2(n19620), .B1(n19395), .B2(n19556), .C1(
        n19868), .C2(n19394), .ZN(P2_U2912) );
  INV_X1 U21621 ( .A(n19421), .ZN(n19397) );
  NAND2_X1 U21622 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19415), .ZN(
        n19399) );
  INV_X1 U21623 ( .A(n19400), .ZN(n19873) );
  OAI21_X1 U21624 ( .B1(n12843), .B2(n19873), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19398) );
  OAI21_X1 U21625 ( .B1(n19399), .B2(n19532), .A(n19398), .ZN(n19874) );
  AOI22_X1 U21626 ( .A1(n19874), .A2(n14988), .B1(n19873), .B2(n19531), .ZN(
        n19405) );
  INV_X1 U21627 ( .A(n19511), .ZN(n19409) );
  NAND2_X1 U21628 ( .A1(n19409), .A2(n19400), .ZN(n19403) );
  OAI22_X1 U21629 ( .A1(n19421), .A2(n19489), .B1(n19408), .B2(n19488), .ZN(
        n19402) );
  AOI21_X1 U21630 ( .B1(n19535), .B2(n19400), .A(n19869), .ZN(n19401) );
  OAI211_X1 U21631 ( .C1(n12843), .C2(n19403), .A(n19402), .B(n19401), .ZN(
        n19877) );
  AOI22_X1 U21632 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19877), .B1(
        n19975), .B2(n19521), .ZN(n19404) );
  OAI211_X1 U21633 ( .C1(n19426), .C2(n19886), .A(n19405), .B(n19404), .ZN(
        P2_U3175) );
  NOR2_X1 U21634 ( .A1(n19408), .A2(n19495), .ZN(n19880) );
  OAI21_X1 U21635 ( .B1(n19406), .B2(n19880), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19407) );
  OAI21_X1 U21636 ( .B1(n19408), .B2(n19497), .A(n19407), .ZN(n19881) );
  AOI22_X1 U21637 ( .A1(n19881), .A2(n14988), .B1(n19880), .B2(n19531), .ZN(
        n19413) );
  NOR2_X1 U21638 ( .A1(n19408), .A2(n19529), .ZN(n19887) );
  INV_X1 U21639 ( .A(n19887), .ZN(n19419) );
  OAI221_X1 U21640 ( .B1(n14662), .B2(n19886), .C1(n14662), .C2(n19893), .A(
        n19419), .ZN(n19411) );
  AOI21_X1 U21641 ( .B1(n12850), .B2(n19409), .A(n19535), .ZN(n19410) );
  AOI22_X1 U21642 ( .A1(n19411), .A2(n19410), .B1(n19880), .B2(n19475), .ZN(
        n19883) );
  AOI22_X1 U21643 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19543), .ZN(n19412) );
  OAI211_X1 U21644 ( .C1(n19546), .C2(n19886), .A(n19413), .B(n19412), .ZN(
        P2_U3167) );
  NAND2_X1 U21645 ( .A1(n19415), .A2(n19488), .ZN(n19428) );
  OAI21_X1 U21646 ( .B1(n19417), .B2(n19887), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19416) );
  OAI21_X1 U21647 ( .B1(n19428), .B2(n19532), .A(n19416), .ZN(n19888) );
  AOI22_X1 U21648 ( .A1(n19888), .A2(n14988), .B1(n19531), .B2(n19887), .ZN(
        n19425) );
  NOR3_X1 U21649 ( .A1(n19417), .A2(n19887), .A3(n19511), .ZN(n19418) );
  AOI211_X1 U21650 ( .C1(n19535), .C2(n19419), .A(n19869), .B(n19418), .ZN(
        n19423) );
  NAND2_X1 U21651 ( .A1(n19420), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19538) );
  OAI21_X1 U21652 ( .B1(n19421), .B2(n19538), .A(n19428), .ZN(n19422) );
  NAND2_X1 U21653 ( .A1(n19423), .A2(n19422), .ZN(n19890) );
  AOI22_X1 U21654 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19890), .B1(
        n19882), .B2(n19521), .ZN(n19424) );
  OAI211_X1 U21655 ( .C1(n19426), .C2(n19899), .A(n19425), .B(n19424), .ZN(
        P2_U3159) );
  INV_X1 U21656 ( .A(n19427), .ZN(n19430) );
  NOR2_X1 U21657 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19428), .ZN(
        n19894) );
  OAI21_X1 U21658 ( .B1(n12841), .B2(n19894), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19429) );
  OAI21_X1 U21659 ( .B1(n19433), .B2(n19430), .A(n19429), .ZN(n19895) );
  AOI22_X1 U21660 ( .A1(n19895), .A2(n14988), .B1(n19894), .B2(n19531), .ZN(
        n19439) );
  OAI21_X1 U21661 ( .B1(n19902), .B2(n19889), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19431) );
  OAI21_X1 U21662 ( .B1(n19433), .B2(n19432), .A(n19431), .ZN(n19437) );
  INV_X1 U21663 ( .A(n19894), .ZN(n19435) );
  NOR3_X1 U21664 ( .A1(n12841), .A2(n19894), .A3(n19511), .ZN(n19434) );
  AOI211_X1 U21665 ( .C1(n19535), .C2(n19435), .A(n19869), .B(n19434), .ZN(
        n19436) );
  NAND2_X1 U21666 ( .A1(n19437), .A2(n19436), .ZN(n19896) );
  AOI22_X1 U21667 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19896), .B1(
        n19902), .B2(n19543), .ZN(n19438) );
  OAI211_X1 U21668 ( .C1(n19546), .C2(n19899), .A(n19439), .B(n19438), .ZN(
        P2_U3151) );
  NOR2_X1 U21669 ( .A1(n19495), .A2(n19454), .ZN(n19907) );
  AOI22_X1 U21670 ( .A1(n19915), .A2(n19543), .B1(n19531), .B2(n19907), .ZN(
        n19451) );
  OAI21_X1 U21671 ( .B1(n19915), .B2(n19908), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19441) );
  NAND2_X1 U21672 ( .A1(n19441), .A2(n19508), .ZN(n19449) );
  AND2_X1 U21673 ( .A1(n19442), .A2(n19456), .ZN(n19445) );
  INV_X1 U21674 ( .A(n19907), .ZN(n19573) );
  OAI211_X1 U21675 ( .C1(n19443), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19573), 
        .B(n19532), .ZN(n19444) );
  OAI211_X1 U21676 ( .C1(n19449), .C2(n19445), .A(n19475), .B(n19444), .ZN(
        n19910) );
  INV_X1 U21677 ( .A(n19445), .ZN(n19448) );
  OAI21_X1 U21678 ( .B1(n19446), .B2(n19907), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19447) );
  AOI22_X1 U21679 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19910), .B1(
        n14988), .B2(n19909), .ZN(n19450) );
  OAI211_X1 U21680 ( .C1(n19546), .C2(n19906), .A(n19451), .B(n19450), .ZN(
        P2_U3135) );
  INV_X1 U21681 ( .A(n19925), .ZN(n19831) );
  NOR2_X1 U21682 ( .A1(n19529), .A2(n19454), .ZN(n19914) );
  AOI22_X1 U21683 ( .A1(n19831), .A2(n19543), .B1(n19531), .B2(n19914), .ZN(
        n19466) );
  OAI21_X1 U21684 ( .B1(n19455), .B2(n19538), .A(n19508), .ZN(n19464) );
  NAND2_X1 U21685 ( .A1(n19456), .A2(n19488), .ZN(n19469) );
  INV_X1 U21686 ( .A(n19469), .ZN(n19461) );
  INV_X1 U21687 ( .A(n19914), .ZN(n19457) );
  AOI21_X1 U21688 ( .B1(n19457), .B2(n19532), .A(n19869), .ZN(n19460) );
  NOR2_X1 U21689 ( .A1(n19458), .A2(n19535), .ZN(n19459) );
  OAI22_X1 U21690 ( .A1(n19464), .A2(n19461), .B1(n19460), .B2(n19459), .ZN(
        n19917) );
  OAI21_X1 U21691 ( .B1(n19462), .B2(n19914), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19463) );
  OAI21_X1 U21692 ( .B1(n19464), .B2(n19469), .A(n19463), .ZN(n19916) );
  AOI22_X1 U21693 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n14988), .ZN(n19465) );
  OAI211_X1 U21694 ( .C1(n19546), .C2(n19913), .A(n19466), .B(n19465), .ZN(
        P2_U3127) );
  INV_X1 U21695 ( .A(n19467), .ZN(n19468) );
  NOR2_X1 U21696 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19469), .ZN(
        n19920) );
  AOI22_X1 U21697 ( .A1(n19928), .A2(n19543), .B1(n19531), .B2(n19920), .ZN(
        n19482) );
  NAND2_X1 U21698 ( .A1(n19925), .A2(n19837), .ZN(n19470) );
  AOI21_X1 U21699 ( .B1(n19470), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19532), 
        .ZN(n19477) );
  NAND2_X1 U21700 ( .A1(n19471), .A2(n19483), .ZN(n19487) );
  OAI21_X1 U21701 ( .B1(n19478), .B2(n19473), .A(n19472), .ZN(n19474) );
  AOI21_X1 U21702 ( .B1(n19477), .B2(n19487), .A(n19474), .ZN(n19476) );
  OAI21_X1 U21703 ( .B1(n19920), .B2(n19476), .A(n19475), .ZN(n19922) );
  INV_X1 U21704 ( .A(n19487), .ZN(n19926) );
  OAI21_X1 U21705 ( .B1(n19926), .B2(n19920), .A(n19477), .ZN(n19480) );
  OAI21_X1 U21706 ( .B1(n19478), .B2(n19920), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19479) );
  NAND2_X1 U21707 ( .A1(n19480), .A2(n19479), .ZN(n19921) );
  AOI22_X1 U21708 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n14988), .ZN(n19481) );
  OAI211_X1 U21709 ( .C1(n19546), .C2(n19925), .A(n19482), .B(n19481), .ZN(
        P2_U3119) );
  NAND2_X1 U21710 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19483), .ZN(
        n19485) );
  OAI21_X1 U21711 ( .B1(n12829), .B2(n19926), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19484) );
  OAI21_X1 U21712 ( .B1(n19485), .B2(n19532), .A(n19484), .ZN(n19927) );
  AOI22_X1 U21713 ( .A1(n19927), .A2(n14988), .B1(n19531), .B2(n19926), .ZN(
        n19494) );
  NOR3_X1 U21714 ( .A1(n12829), .A2(n19926), .A3(n19511), .ZN(n19486) );
  AOI211_X1 U21715 ( .C1(n19535), .C2(n19487), .A(n19869), .B(n19486), .ZN(
        n19491) );
  OAI22_X1 U21716 ( .A1(n19509), .A2(n19489), .B1(n19510), .B2(n19488), .ZN(
        n19490) );
  NAND2_X1 U21717 ( .A1(n19491), .A2(n19490), .ZN(n19929) );
  INV_X1 U21718 ( .A(n19937), .ZN(n19834) );
  AOI22_X1 U21719 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19929), .B1(
        n19834), .B2(n19543), .ZN(n19493) );
  OAI211_X1 U21720 ( .C1(n19546), .C2(n19837), .A(n19494), .B(n19493), .ZN(
        P2_U3111) );
  NOR2_X1 U21721 ( .A1(n19495), .A2(n19510), .ZN(n19932) );
  OAI21_X1 U21722 ( .B1(n12830), .B2(n19932), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19496) );
  OAI21_X1 U21723 ( .B1(n19510), .B2(n19497), .A(n19496), .ZN(n19933) );
  AOI22_X1 U21724 ( .A1(n19933), .A2(n14988), .B1(n19932), .B2(n19531), .ZN(
        n19507) );
  AOI21_X1 U21725 ( .B1(n19937), .B2(n19743), .A(n14662), .ZN(n19505) );
  NOR2_X1 U21726 ( .A1(n19500), .A2(n19510), .ZN(n19504) );
  INV_X1 U21727 ( .A(n19932), .ZN(n19502) );
  NOR3_X1 U21728 ( .A1(n12830), .A2(n19932), .A3(n19511), .ZN(n19501) );
  AOI211_X1 U21729 ( .C1(n19535), .C2(n19502), .A(n19869), .B(n19501), .ZN(
        n19503) );
  AOI22_X1 U21730 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19934), .B1(
        n19939), .B2(n19543), .ZN(n19506) );
  OAI211_X1 U21731 ( .C1(n19546), .C2(n19937), .A(n19507), .B(n19506), .ZN(
        P2_U3103) );
  NOR2_X1 U21732 ( .A1(n19529), .A2(n19510), .ZN(n19938) );
  AOI22_X1 U21733 ( .A1(n19946), .A2(n19543), .B1(n19531), .B2(n19938), .ZN(
        n19520) );
  OAI21_X1 U21734 ( .B1(n19509), .B2(n19538), .A(n19508), .ZN(n19518) );
  NOR2_X1 U21735 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19510), .ZN(
        n19515) );
  INV_X1 U21736 ( .A(n19938), .ZN(n19513) );
  NOR3_X1 U21737 ( .A1(n12831), .A2(n19938), .A3(n19511), .ZN(n19512) );
  AOI211_X1 U21738 ( .C1(n19535), .C2(n19513), .A(n19869), .B(n19512), .ZN(
        n19514) );
  OAI21_X1 U21739 ( .B1(n19518), .B2(n19515), .A(n19514), .ZN(n19941) );
  INV_X1 U21740 ( .A(n19515), .ZN(n19517) );
  OAI21_X1 U21741 ( .B1(n12831), .B2(n19938), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19516) );
  OAI21_X1 U21742 ( .B1(n19518), .B2(n19517), .A(n19516), .ZN(n19940) );
  AOI22_X1 U21743 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19941), .B1(
        n14988), .B2(n19940), .ZN(n19519) );
  OAI211_X1 U21744 ( .C1(n19546), .C2(n19743), .A(n19520), .B(n19519), .ZN(
        P2_U3095) );
  AOI22_X1 U21745 ( .A1(n19846), .A2(n19543), .B1(n19531), .B2(n19952), .ZN(
        n19523) );
  AOI22_X1 U21746 ( .A1(n14988), .A2(n19954), .B1(n19953), .B2(n19521), .ZN(
        n19522) );
  OAI211_X1 U21747 ( .C1(n19525), .C2(n19524), .A(n19523), .B(n19522), .ZN(
        P2_U3079) );
  AOI22_X1 U21748 ( .A1(n19960), .A2(n14988), .B1(n19531), .B2(n19959), .ZN(
        n19527) );
  AOI22_X1 U21749 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n19543), .ZN(n19526) );
  OAI211_X1 U21750 ( .C1(n19546), .C2(n19965), .A(n19527), .B(n19526), .ZN(
        P2_U3071) );
  NOR2_X1 U21751 ( .A1(n19529), .A2(n19528), .ZN(n19966) );
  OAI21_X1 U21752 ( .B1(n19534), .B2(n19966), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19530) );
  OAI21_X1 U21753 ( .B1(n19537), .B2(n19532), .A(n19530), .ZN(n19967) );
  AOI22_X1 U21754 ( .A1(n19967), .A2(n14988), .B1(n19531), .B2(n19966), .ZN(
        n19545) );
  INV_X1 U21755 ( .A(n19966), .ZN(n19533) );
  AOI21_X1 U21756 ( .B1(n19533), .B2(n19532), .A(n19869), .ZN(n19542) );
  INV_X1 U21757 ( .A(n19534), .ZN(n19536) );
  NOR2_X1 U21758 ( .A1(n19536), .A2(n19535), .ZN(n19541) );
  OAI21_X1 U21759 ( .B1(n19539), .B2(n19538), .A(n19537), .ZN(n19540) );
  OAI21_X1 U21760 ( .B1(n19542), .B2(n19541), .A(n19540), .ZN(n19968) );
  AOI22_X1 U21761 ( .A1(n19968), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n19978), .B2(n19543), .ZN(n19544) );
  OAI211_X1 U21762 ( .C1(n19546), .C2(n19971), .A(n19545), .B(n19544), .ZN(
        P2_U3063) );
  AOI22_X1 U21763 ( .A1(n19763), .A2(n19555), .B1(n19859), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n19554) );
  AOI22_X1 U21764 ( .A1(n19765), .A2(BUF1_REG_22__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n19553) );
  INV_X1 U21765 ( .A(n19547), .ZN(n19548) );
  OAI22_X1 U21766 ( .A1(n19550), .A2(n19812), .B1(n19549), .B2(n19548), .ZN(
        n19551) );
  INV_X1 U21767 ( .A(n19551), .ZN(n19552) );
  NAND3_X1 U21768 ( .A1(n19554), .A2(n19553), .A3(n19552), .ZN(P2_U2897) );
  INV_X1 U21769 ( .A(n19555), .ZN(n19561) );
  OAI222_X1 U21770 ( .A1(n19558), .A2(n19620), .B1(n19557), .B2(n19556), .C1(
        n19868), .C2(n19561), .ZN(P2_U2913) );
  OAI22_X1 U21771 ( .A1(n20306), .A2(n19560), .B1(n15699), .B2(n19559), .ZN(
        n19600) );
  NOR2_X2 U21772 ( .A1(n19561), .A2(n19869), .ZN(n19602) );
  NOR2_X2 U21773 ( .A1(n19562), .A2(n19871), .ZN(n19599) );
  AOI22_X1 U21774 ( .A1(n19874), .A2(n19602), .B1(n19873), .B2(n19599), .ZN(
        n19564) );
  AOI22_X1 U21775 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19875), .ZN(n19598) );
  INV_X1 U21776 ( .A(n19598), .ZN(n19601) );
  AOI22_X1 U21777 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19877), .B1(
        n19975), .B2(n19601), .ZN(n19563) );
  OAI211_X1 U21778 ( .C1(n19593), .C2(n19886), .A(n19564), .B(n19563), .ZN(
        P2_U3174) );
  AOI22_X1 U21779 ( .A1(n19881), .A2(n19602), .B1(n19880), .B2(n19599), .ZN(
        n19566) );
  AOI22_X1 U21780 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19600), .ZN(n19565) );
  OAI211_X1 U21781 ( .C1(n19598), .C2(n19886), .A(n19566), .B(n19565), .ZN(
        P2_U3166) );
  AOI22_X1 U21782 ( .A1(n19888), .A2(n19602), .B1(n19599), .B2(n19887), .ZN(
        n19568) );
  AOI22_X1 U21783 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19600), .ZN(n19567) );
  OAI211_X1 U21784 ( .C1(n19598), .C2(n19893), .A(n19568), .B(n19567), .ZN(
        P2_U3158) );
  AOI22_X1 U21785 ( .A1(n19895), .A2(n19602), .B1(n19894), .B2(n19599), .ZN(
        n19570) );
  AOI22_X1 U21786 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19896), .B1(
        n19902), .B2(n19600), .ZN(n19569) );
  OAI211_X1 U21787 ( .C1(n19598), .C2(n19899), .A(n19570), .B(n19569), .ZN(
        P2_U3150) );
  AOI22_X1 U21788 ( .A1(n19901), .A2(n19602), .B1(n19900), .B2(n19599), .ZN(
        n19572) );
  AOI22_X1 U21789 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19903), .B1(
        n19601), .B2(n19902), .ZN(n19571) );
  OAI211_X1 U21790 ( .C1(n19593), .C2(n19906), .A(n19572), .B(n19571), .ZN(
        P2_U3142) );
  INV_X1 U21791 ( .A(n19599), .ZN(n19574) );
  OAI22_X1 U21792 ( .A1(n19913), .A2(n19593), .B1(n19574), .B2(n19573), .ZN(
        n19575) );
  INV_X1 U21793 ( .A(n19575), .ZN(n19577) );
  AOI22_X1 U21794 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19910), .B1(
        n19602), .B2(n19909), .ZN(n19576) );
  OAI211_X1 U21795 ( .C1(n19598), .C2(n19906), .A(n19577), .B(n19576), .ZN(
        P2_U3134) );
  AOI22_X1 U21796 ( .A1(n19915), .A2(n19601), .B1(n19599), .B2(n19914), .ZN(
        n19579) );
  AOI22_X1 U21797 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19602), .ZN(n19578) );
  OAI211_X1 U21798 ( .C1(n19593), .C2(n19925), .A(n19579), .B(n19578), .ZN(
        P2_U3126) );
  AOI22_X1 U21799 ( .A1(n19831), .A2(n19601), .B1(n19599), .B2(n19920), .ZN(
        n19581) );
  AOI22_X1 U21800 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19602), .ZN(n19580) );
  OAI211_X1 U21801 ( .C1(n19593), .C2(n19837), .A(n19581), .B(n19580), .ZN(
        P2_U3118) );
  AOI22_X1 U21802 ( .A1(n19927), .A2(n19602), .B1(n19926), .B2(n19599), .ZN(
        n19583) );
  AOI22_X1 U21803 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19929), .B1(
        n19928), .B2(n19601), .ZN(n19582) );
  OAI211_X1 U21804 ( .C1(n19593), .C2(n19937), .A(n19583), .B(n19582), .ZN(
        P2_U3110) );
  AOI22_X1 U21805 ( .A1(n19933), .A2(n19602), .B1(n19932), .B2(n19599), .ZN(
        n19585) );
  AOI22_X1 U21806 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19934), .B1(
        n19939), .B2(n19600), .ZN(n19584) );
  OAI211_X1 U21807 ( .C1(n19598), .C2(n19937), .A(n19585), .B(n19584), .ZN(
        P2_U3102) );
  AOI22_X1 U21808 ( .A1(n19601), .A2(n19939), .B1(n19938), .B2(n19599), .ZN(
        n19587) );
  AOI22_X1 U21809 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19941), .B1(
        n19602), .B2(n19940), .ZN(n19586) );
  OAI211_X1 U21810 ( .C1(n19593), .C2(n19944), .A(n19587), .B(n19586), .ZN(
        P2_U3094) );
  INV_X1 U21811 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n19590) );
  AOI22_X1 U21812 ( .A1(n19601), .A2(n19946), .B1(n19945), .B2(n19599), .ZN(
        n19589) );
  AOI22_X1 U21813 ( .A1(n19602), .A2(n19947), .B1(n19953), .B2(n19600), .ZN(
        n19588) );
  OAI211_X1 U21814 ( .C1(n19951), .C2(n19590), .A(n19589), .B(n19588), .ZN(
        P2_U3086) );
  AOI22_X1 U21815 ( .A1(n19601), .A2(n19953), .B1(n19952), .B2(n19599), .ZN(
        n19592) );
  AOI22_X1 U21816 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19955), .B1(
        n19602), .B2(n19954), .ZN(n19591) );
  OAI211_X1 U21817 ( .C1(n19593), .C2(n19965), .A(n19592), .B(n19591), .ZN(
        P2_U3078) );
  AOI22_X1 U21818 ( .A1(n19960), .A2(n19602), .B1(n19599), .B2(n19959), .ZN(
        n19595) );
  AOI22_X1 U21819 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n19600), .ZN(n19594) );
  OAI211_X1 U21820 ( .C1(n19598), .C2(n19965), .A(n19595), .B(n19594), .ZN(
        P2_U3070) );
  AOI22_X1 U21821 ( .A1(n19967), .A2(n19602), .B1(n19599), .B2(n19966), .ZN(
        n19597) );
  AOI22_X1 U21822 ( .A1(n19968), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n19978), .B2(n19600), .ZN(n19596) );
  OAI211_X1 U21823 ( .C1(n19598), .C2(n19971), .A(n19597), .B(n19596), .ZN(
        P2_U3062) );
  AOI22_X1 U21824 ( .A1(n19975), .A2(n19600), .B1(n19974), .B2(n19599), .ZN(
        n19604) );
  AOI22_X1 U21825 ( .A1(n19602), .A2(n19979), .B1(n19978), .B2(n19601), .ZN(
        n19603) );
  OAI211_X1 U21826 ( .C1(n19984), .C2(n19605), .A(n19604), .B(n19603), .ZN(
        P2_U3054) );
  AOI22_X1 U21827 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19859), .B1(n19607), .B2(
        n19606), .ZN(n19618) );
  NAND2_X1 U21828 ( .A1(n19609), .A2(n19608), .ZN(n19610) );
  OAI21_X1 U21829 ( .B1(n19612), .B2(n19611), .A(n19610), .ZN(n19714) );
  XOR2_X1 U21830 ( .A(n19712), .B(n19613), .Z(n19715) );
  NOR2_X1 U21831 ( .A1(n19714), .A2(n19715), .ZN(n19713) );
  NOR2_X1 U21832 ( .A1(n19614), .A2(n19712), .ZN(n19615) );
  OAI21_X1 U21833 ( .B1(n19713), .B2(n19615), .A(n19663), .ZN(n19666) );
  INV_X1 U21834 ( .A(n19665), .ZN(n19616) );
  NAND3_X1 U21835 ( .A1(n19666), .A2(n19616), .A3(n19862), .ZN(n19617) );
  OAI211_X1 U21836 ( .C1(n19620), .C2(n19619), .A(n19618), .B(n19617), .ZN(
        P2_U2914) );
  AOI22_X1 U21837 ( .A1(n19874), .A2(n19651), .B1(n19873), .B2(n19650), .ZN(
        n19622) );
  AOI22_X1 U21838 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19877), .B1(
        n19975), .B2(n19644), .ZN(n19621) );
  OAI211_X1 U21839 ( .C1(n19635), .C2(n19886), .A(n19622), .B(n19621), .ZN(
        P2_U3173) );
  AOI22_X1 U21840 ( .A1(n19881), .A2(n19651), .B1(n19880), .B2(n19650), .ZN(
        n19624) );
  AOI22_X1 U21841 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19652), .ZN(n19623) );
  OAI211_X1 U21842 ( .C1(n19655), .C2(n19886), .A(n19624), .B(n19623), .ZN(
        P2_U3165) );
  AOI22_X1 U21843 ( .A1(n19888), .A2(n19651), .B1(n19650), .B2(n19887), .ZN(
        n19626) );
  AOI22_X1 U21844 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19652), .ZN(n19625) );
  OAI211_X1 U21845 ( .C1(n19655), .C2(n19893), .A(n19626), .B(n19625), .ZN(
        P2_U3157) );
  AOI22_X1 U21846 ( .A1(n19895), .A2(n19651), .B1(n19894), .B2(n19650), .ZN(
        n19628) );
  AOI22_X1 U21847 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19896), .B1(
        n19902), .B2(n19652), .ZN(n19627) );
  OAI211_X1 U21848 ( .C1(n19655), .C2(n19899), .A(n19628), .B(n19627), .ZN(
        P2_U3149) );
  AOI22_X1 U21849 ( .A1(n19901), .A2(n19651), .B1(n19650), .B2(n19900), .ZN(
        n19630) );
  AOI22_X1 U21850 ( .A1(n19644), .A2(n19902), .B1(n19903), .B2(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n19629) );
  OAI211_X1 U21851 ( .C1(n19635), .C2(n19906), .A(n19630), .B(n19629), .ZN(
        P2_U3141) );
  AOI22_X1 U21852 ( .A1(n19915), .A2(n19652), .B1(n19650), .B2(n19907), .ZN(
        n19632) );
  AOI22_X1 U21853 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19910), .B1(
        n19651), .B2(n19909), .ZN(n19631) );
  OAI211_X1 U21854 ( .C1(n19655), .C2(n19906), .A(n19632), .B(n19631), .ZN(
        P2_U3133) );
  AOI22_X1 U21855 ( .A1(n19915), .A2(n19644), .B1(n19650), .B2(n19914), .ZN(
        n19634) );
  AOI22_X1 U21856 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19651), .ZN(n19633) );
  OAI211_X1 U21857 ( .C1(n19635), .C2(n19925), .A(n19634), .B(n19633), .ZN(
        P2_U3125) );
  AOI22_X1 U21858 ( .A1(n19928), .A2(n19652), .B1(n19650), .B2(n19920), .ZN(
        n19637) );
  AOI22_X1 U21859 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19651), .ZN(n19636) );
  OAI211_X1 U21860 ( .C1(n19655), .C2(n19925), .A(n19637), .B(n19636), .ZN(
        P2_U3117) );
  AOI22_X1 U21861 ( .A1(n19927), .A2(n19651), .B1(n19650), .B2(n19926), .ZN(
        n19639) );
  AOI22_X1 U21862 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19929), .B1(
        n19834), .B2(n19652), .ZN(n19638) );
  OAI211_X1 U21863 ( .C1(n19655), .C2(n19837), .A(n19639), .B(n19638), .ZN(
        P2_U3109) );
  AOI22_X1 U21864 ( .A1(n19933), .A2(n19651), .B1(n19932), .B2(n19650), .ZN(
        n19641) );
  AOI22_X1 U21865 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19934), .B1(
        n19939), .B2(n19652), .ZN(n19640) );
  OAI211_X1 U21866 ( .C1(n19655), .C2(n19937), .A(n19641), .B(n19640), .ZN(
        P2_U3101) );
  AOI22_X1 U21867 ( .A1(n19946), .A2(n19652), .B1(n19650), .B2(n19938), .ZN(
        n19643) );
  AOI22_X1 U21868 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19941), .B1(
        n19651), .B2(n19940), .ZN(n19642) );
  OAI211_X1 U21869 ( .C1(n19655), .C2(n19743), .A(n19643), .B(n19642), .ZN(
        P2_U3093) );
  INV_X1 U21870 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n19647) );
  AOI22_X1 U21871 ( .A1(n19644), .A2(n19946), .B1(n19945), .B2(n19650), .ZN(
        n19646) );
  AOI22_X1 U21872 ( .A1(n19651), .A2(n19947), .B1(n19953), .B2(n19652), .ZN(
        n19645) );
  OAI211_X1 U21873 ( .C1(n19951), .C2(n19647), .A(n19646), .B(n19645), .ZN(
        P2_U3085) );
  AOI22_X1 U21874 ( .A1(n19960), .A2(n19651), .B1(n19650), .B2(n19959), .ZN(
        n19649) );
  AOI22_X1 U21875 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n19652), .ZN(n19648) );
  OAI211_X1 U21876 ( .C1(n19655), .C2(n19965), .A(n19649), .B(n19648), .ZN(
        P2_U3069) );
  AOI22_X1 U21877 ( .A1(n19967), .A2(n19651), .B1(n19650), .B2(n19966), .ZN(
        n19654) );
  AOI22_X1 U21878 ( .A1(n19968), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n19978), .B2(n19652), .ZN(n19653) );
  OAI211_X1 U21879 ( .C1(n19655), .C2(n19971), .A(n19654), .B(n19653), .ZN(
        P2_U3061) );
  AOI22_X1 U21880 ( .A1(n19763), .A2(n19662), .B1(n19859), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n19661) );
  AOI22_X1 U21881 ( .A1(n19765), .A2(BUF1_REG_20__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n19660) );
  INV_X1 U21882 ( .A(n19656), .ZN(n19658) );
  AOI22_X1 U21883 ( .A1(n19658), .A2(n19862), .B1(n19860), .B2(n19657), .ZN(
        n19659) );
  NAND3_X1 U21884 ( .A1(n19661), .A2(n19660), .A3(n19659), .ZN(P2_U2899) );
  INV_X1 U21885 ( .A(n19662), .ZN(n19670) );
  INV_X1 U21886 ( .A(n19663), .ZN(n19664) );
  AOI22_X1 U21887 ( .A1(n19860), .A2(n19664), .B1(n19859), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19669) );
  XNOR2_X1 U21888 ( .A(n19666), .B(n19665), .ZN(n19667) );
  NAND2_X1 U21889 ( .A1(n19667), .A2(n19862), .ZN(n19668) );
  OAI211_X1 U21890 ( .C1(n19670), .C2(n19868), .A(n19669), .B(n19668), .ZN(
        P2_U2915) );
  AOI22_X1 U21891 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19875), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19876), .ZN(n19699) );
  NOR2_X2 U21892 ( .A1(n19670), .A2(n19869), .ZN(n19708) );
  AOI22_X1 U21893 ( .A1(n19874), .A2(n19708), .B1(n19873), .B2(n19705), .ZN(
        n19673) );
  AOI22_X1 U21894 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19875), .ZN(n19704) );
  INV_X1 U21895 ( .A(n19704), .ZN(n19707) );
  AOI22_X1 U21896 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19877), .B1(
        n19975), .B2(n19707), .ZN(n19672) );
  OAI211_X1 U21897 ( .C1(n19699), .C2(n19886), .A(n19673), .B(n19672), .ZN(
        P2_U3172) );
  AOI22_X1 U21898 ( .A1(n19881), .A2(n19708), .B1(n19880), .B2(n19705), .ZN(
        n19675) );
  AOI22_X1 U21899 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19706), .ZN(n19674) );
  OAI211_X1 U21900 ( .C1(n19704), .C2(n19886), .A(n19675), .B(n19674), .ZN(
        P2_U3164) );
  AOI22_X1 U21901 ( .A1(n19888), .A2(n19708), .B1(n11124), .B2(n19887), .ZN(
        n19677) );
  AOI22_X1 U21902 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19890), .B1(
        n19882), .B2(n19707), .ZN(n19676) );
  OAI211_X1 U21903 ( .C1(n19699), .C2(n19899), .A(n19677), .B(n19676), .ZN(
        P2_U3156) );
  AOI22_X1 U21904 ( .A1(n19895), .A2(n19708), .B1(n19894), .B2(n19705), .ZN(
        n19679) );
  AOI22_X1 U21905 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19896), .B1(
        n19902), .B2(n19706), .ZN(n19678) );
  OAI211_X1 U21906 ( .C1(n19704), .C2(n19899), .A(n19679), .B(n19678), .ZN(
        P2_U3148) );
  AOI22_X1 U21907 ( .A1(n19901), .A2(n19708), .B1(n19900), .B2(n19705), .ZN(
        n19681) );
  AOI22_X1 U21908 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19903), .B1(
        n19707), .B2(n19902), .ZN(n19680) );
  OAI211_X1 U21909 ( .C1(n19699), .C2(n19906), .A(n19681), .B(n19680), .ZN(
        P2_U3140) );
  AOI22_X1 U21910 ( .A1(n19908), .A2(n19707), .B1(n11123), .B2(n19907), .ZN(
        n19683) );
  AOI22_X1 U21911 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19910), .B1(
        n19708), .B2(n19909), .ZN(n19682) );
  OAI211_X1 U21912 ( .C1(n19699), .C2(n19913), .A(n19683), .B(n19682), .ZN(
        P2_U3132) );
  AOI22_X1 U21913 ( .A1(n19915), .A2(n19707), .B1(n11124), .B2(n19914), .ZN(
        n19685) );
  AOI22_X1 U21914 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19708), .ZN(n19684) );
  OAI211_X1 U21915 ( .C1(n19699), .C2(n19925), .A(n19685), .B(n19684), .ZN(
        P2_U3124) );
  AOI22_X1 U21916 ( .A1(n19706), .A2(n19928), .B1(n11123), .B2(n19920), .ZN(
        n19687) );
  AOI22_X1 U21917 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19708), .ZN(n19686) );
  OAI211_X1 U21918 ( .C1(n19704), .C2(n19925), .A(n19687), .B(n19686), .ZN(
        P2_U3116) );
  AOI22_X1 U21919 ( .A1(n19927), .A2(n19708), .B1(n19926), .B2(n19705), .ZN(
        n19689) );
  AOI22_X1 U21920 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19929), .B1(
        n19834), .B2(n19706), .ZN(n19688) );
  OAI211_X1 U21921 ( .C1(n19704), .C2(n19837), .A(n19689), .B(n19688), .ZN(
        P2_U3108) );
  AOI22_X1 U21922 ( .A1(n19933), .A2(n19708), .B1(n19932), .B2(n11123), .ZN(
        n19691) );
  AOI22_X1 U21923 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19934), .B1(
        n19939), .B2(n19706), .ZN(n19690) );
  OAI211_X1 U21924 ( .C1(n19704), .C2(n19937), .A(n19691), .B(n19690), .ZN(
        P2_U3100) );
  AOI22_X1 U21925 ( .A1(n19707), .A2(n19939), .B1(n19938), .B2(n11123), .ZN(
        n19693) );
  AOI22_X1 U21926 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19941), .B1(
        n19708), .B2(n19940), .ZN(n19692) );
  OAI211_X1 U21927 ( .C1(n19699), .C2(n19944), .A(n19693), .B(n19692), .ZN(
        P2_U3092) );
  INV_X1 U21928 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n19696) );
  AOI22_X1 U21929 ( .A1(n19707), .A2(n19946), .B1(n19945), .B2(n11123), .ZN(
        n19695) );
  AOI22_X1 U21930 ( .A1(n19708), .A2(n19947), .B1(n19953), .B2(n19706), .ZN(
        n19694) );
  OAI211_X1 U21931 ( .C1(n19951), .C2(n19696), .A(n19695), .B(n19694), .ZN(
        P2_U3084) );
  AOI22_X1 U21932 ( .A1(n19707), .A2(n19953), .B1(n19952), .B2(n11124), .ZN(
        n19698) );
  AOI22_X1 U21933 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19955), .B1(
        n19708), .B2(n19954), .ZN(n19697) );
  OAI211_X1 U21934 ( .C1(n19699), .C2(n19965), .A(n19698), .B(n19697), .ZN(
        P2_U3076) );
  AOI22_X1 U21935 ( .A1(n19960), .A2(n19708), .B1(n11123), .B2(n19959), .ZN(
        n19701) );
  AOI22_X1 U21936 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n19706), .ZN(n19700) );
  OAI211_X1 U21937 ( .C1(n19704), .C2(n19965), .A(n19701), .B(n19700), .ZN(
        P2_U3068) );
  AOI22_X1 U21938 ( .A1(n19967), .A2(n19708), .B1(n11124), .B2(n19966), .ZN(
        n19703) );
  AOI22_X1 U21939 ( .A1(n19968), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n19706), .B2(n19978), .ZN(n19702) );
  OAI211_X1 U21940 ( .C1(n19704), .C2(n19971), .A(n19703), .B(n19702), .ZN(
        P2_U3060) );
  AOI22_X1 U21941 ( .A1(n19706), .A2(n19975), .B1(n19974), .B2(n11124), .ZN(
        n19710) );
  AOI22_X1 U21942 ( .A1(n19708), .A2(n19979), .B1(n19978), .B2(n19707), .ZN(
        n19709) );
  OAI211_X1 U21943 ( .C1(n19984), .C2(n19711), .A(n19710), .B(n19709), .ZN(
        P2_U3052) );
  AOI22_X1 U21944 ( .A1(n19712), .A2(n19860), .B1(n19859), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19718) );
  AOI21_X1 U21945 ( .B1(n19715), .B2(n19714), .A(n19713), .ZN(n19716) );
  OR2_X1 U21946 ( .A1(n19716), .A2(n19812), .ZN(n19717) );
  OAI211_X1 U21947 ( .C1(n19719), .C2(n19868), .A(n19718), .B(n19717), .ZN(
        P2_U2916) );
  AOI22_X1 U21948 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19875), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19876), .ZN(n19749) );
  NOR2_X2 U21949 ( .A1(n19719), .A2(n19869), .ZN(n19758) );
  NOR2_X2 U21950 ( .A1(n19720), .A2(n19871), .ZN(n19755) );
  AOI22_X1 U21951 ( .A1(n19874), .A2(n19758), .B1(n19873), .B2(n19755), .ZN(
        n19722) );
  AOI22_X2 U21952 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19875), .ZN(n19754) );
  INV_X1 U21953 ( .A(n19754), .ZN(n19757) );
  AOI22_X1 U21954 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19877), .B1(
        n19975), .B2(n19757), .ZN(n19721) );
  OAI211_X1 U21955 ( .C1(n19749), .C2(n19886), .A(n19722), .B(n19721), .ZN(
        P2_U3171) );
  AOI22_X1 U21956 ( .A1(n19881), .A2(n19758), .B1(n19880), .B2(n19755), .ZN(
        n19724) );
  AOI22_X1 U21957 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19756), .ZN(n19723) );
  OAI211_X1 U21958 ( .C1(n19754), .C2(n19886), .A(n19724), .B(n19723), .ZN(
        P2_U3163) );
  AOI22_X1 U21959 ( .A1(n19888), .A2(n19758), .B1(n19755), .B2(n19887), .ZN(
        n19726) );
  AOI22_X1 U21960 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19756), .ZN(n19725) );
  OAI211_X1 U21961 ( .C1(n19754), .C2(n19893), .A(n19726), .B(n19725), .ZN(
        P2_U3155) );
  AOI22_X1 U21962 ( .A1(n19895), .A2(n19758), .B1(n19894), .B2(n19755), .ZN(
        n19728) );
  AOI22_X1 U21963 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19896), .B1(
        n19902), .B2(n19756), .ZN(n19727) );
  OAI211_X1 U21964 ( .C1(n19754), .C2(n19899), .A(n19728), .B(n19727), .ZN(
        P2_U3147) );
  AOI22_X1 U21965 ( .A1(n19901), .A2(n19758), .B1(n19900), .B2(n19755), .ZN(
        n19730) );
  AOI22_X1 U21966 ( .A1(n19757), .A2(n19902), .B1(n19903), .B2(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n19729) );
  OAI211_X1 U21967 ( .C1(n19749), .C2(n19906), .A(n19730), .B(n19729), .ZN(
        P2_U3139) );
  AOI22_X1 U21968 ( .A1(n19915), .A2(n19756), .B1(n19755), .B2(n19907), .ZN(
        n19732) );
  AOI22_X1 U21969 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19910), .B1(
        n19758), .B2(n19909), .ZN(n19731) );
  OAI211_X1 U21970 ( .C1(n19754), .C2(n19906), .A(n19732), .B(n19731), .ZN(
        P2_U3131) );
  AOI22_X1 U21971 ( .A1(n19831), .A2(n19756), .B1(n19755), .B2(n19914), .ZN(
        n19734) );
  AOI22_X1 U21972 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19758), .ZN(n19733) );
  OAI211_X1 U21973 ( .C1(n19754), .C2(n19913), .A(n19734), .B(n19733), .ZN(
        P2_U3123) );
  AOI22_X1 U21974 ( .A1(n19928), .A2(n19756), .B1(n19755), .B2(n19920), .ZN(
        n19736) );
  AOI22_X1 U21975 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19758), .ZN(n19735) );
  OAI211_X1 U21976 ( .C1(n19754), .C2(n19925), .A(n19736), .B(n19735), .ZN(
        P2_U3115) );
  AOI22_X1 U21977 ( .A1(n19927), .A2(n19758), .B1(n19926), .B2(n19755), .ZN(
        n19738) );
  AOI22_X1 U21978 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19929), .B1(
        n19834), .B2(n19756), .ZN(n19737) );
  OAI211_X1 U21979 ( .C1(n19754), .C2(n19837), .A(n19738), .B(n19737), .ZN(
        P2_U3107) );
  AOI22_X1 U21980 ( .A1(n19933), .A2(n19758), .B1(n19932), .B2(n19755), .ZN(
        n19740) );
  AOI22_X1 U21981 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19934), .B1(
        n19939), .B2(n19756), .ZN(n19739) );
  OAI211_X1 U21982 ( .C1(n19754), .C2(n19937), .A(n19740), .B(n19739), .ZN(
        P2_U3099) );
  AOI22_X1 U21983 ( .A1(n19946), .A2(n19756), .B1(n19938), .B2(n19755), .ZN(
        n19742) );
  AOI22_X1 U21984 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19941), .B1(
        n19758), .B2(n19940), .ZN(n19741) );
  OAI211_X1 U21985 ( .C1(n19754), .C2(n19743), .A(n19742), .B(n19741), .ZN(
        P2_U3091) );
  INV_X1 U21986 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n19746) );
  AOI22_X1 U21987 ( .A1(n19757), .A2(n19946), .B1(n19945), .B2(n19755), .ZN(
        n19745) );
  AOI22_X1 U21988 ( .A1(n19758), .A2(n19947), .B1(n19953), .B2(n19756), .ZN(
        n19744) );
  OAI211_X1 U21989 ( .C1(n19951), .C2(n19746), .A(n19745), .B(n19744), .ZN(
        P2_U3083) );
  AOI22_X1 U21990 ( .A1(n19757), .A2(n19953), .B1(n19952), .B2(n19755), .ZN(
        n19748) );
  AOI22_X1 U21991 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19955), .B1(
        n19758), .B2(n19954), .ZN(n19747) );
  OAI211_X1 U21992 ( .C1(n19749), .C2(n19965), .A(n19748), .B(n19747), .ZN(
        P2_U3075) );
  AOI22_X1 U21993 ( .A1(n19960), .A2(n19758), .B1(n19755), .B2(n19959), .ZN(
        n19751) );
  AOI22_X1 U21994 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n19756), .ZN(n19750) );
  OAI211_X1 U21995 ( .C1(n19754), .C2(n19965), .A(n19751), .B(n19750), .ZN(
        P2_U3067) );
  AOI22_X1 U21996 ( .A1(n19967), .A2(n19758), .B1(n19755), .B2(n19966), .ZN(
        n19753) );
  AOI22_X1 U21997 ( .A1(n19968), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n19978), .B2(n19756), .ZN(n19752) );
  OAI211_X1 U21998 ( .C1(n19754), .C2(n19971), .A(n19753), .B(n19752), .ZN(
        P2_U3059) );
  AOI22_X1 U21999 ( .A1(n19975), .A2(n19756), .B1(n19974), .B2(n19755), .ZN(
        n19760) );
  AOI22_X1 U22000 ( .A1(n19758), .A2(n19979), .B1(n19978), .B2(n19757), .ZN(
        n19759) );
  OAI211_X1 U22001 ( .C1(n19984), .C2(n19761), .A(n19760), .B(n19759), .ZN(
        P2_U3051) );
  AOI22_X1 U22002 ( .A1(n19763), .A2(n19762), .B1(n19859), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U22003 ( .A1(n19765), .A2(BUF1_REG_18__SCAN_IN), .B1(n19764), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U22004 ( .A1(n19767), .A2(n19862), .B1(n19860), .B2(n19766), .ZN(
        n19768) );
  NAND3_X1 U22005 ( .A1(n19770), .A2(n19769), .A3(n19768), .ZN(P2_U2901) );
  AOI22_X1 U22006 ( .A1(n19874), .A2(n19805), .B1(n19873), .B2(n19802), .ZN(
        n19772) );
  AOI22_X1 U22007 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19877), .B1(
        n19975), .B2(n19804), .ZN(n19771) );
  OAI211_X1 U22008 ( .C1(n19791), .C2(n19886), .A(n19772), .B(n19771), .ZN(
        P2_U3170) );
  AOI22_X1 U22009 ( .A1(n19881), .A2(n19805), .B1(n19880), .B2(n19802), .ZN(
        n19774) );
  AOI22_X1 U22010 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19803), .ZN(n19773) );
  OAI211_X1 U22011 ( .C1(n19801), .C2(n19886), .A(n19774), .B(n19773), .ZN(
        P2_U3162) );
  AOI22_X1 U22012 ( .A1(n19888), .A2(n19805), .B1(n19802), .B2(n19887), .ZN(
        n19776) );
  AOI22_X1 U22013 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19803), .ZN(n19775) );
  OAI211_X1 U22014 ( .C1(n19801), .C2(n19893), .A(n19776), .B(n19775), .ZN(
        P2_U3154) );
  AOI22_X1 U22015 ( .A1(n19895), .A2(n19805), .B1(n19894), .B2(n19802), .ZN(
        n19778) );
  AOI22_X1 U22016 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19896), .B1(
        n19902), .B2(n19803), .ZN(n19777) );
  OAI211_X1 U22017 ( .C1(n19801), .C2(n19899), .A(n19778), .B(n19777), .ZN(
        P2_U3146) );
  AOI22_X1 U22018 ( .A1(n19915), .A2(n19803), .B1(n19802), .B2(n19907), .ZN(
        n19780) );
  AOI22_X1 U22019 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19910), .B1(
        n19805), .B2(n19909), .ZN(n19779) );
  OAI211_X1 U22020 ( .C1(n19801), .C2(n19906), .A(n19780), .B(n19779), .ZN(
        P2_U3130) );
  AOI22_X1 U22021 ( .A1(n19915), .A2(n19804), .B1(n19802), .B2(n19914), .ZN(
        n19782) );
  AOI22_X1 U22022 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19805), .ZN(n19781) );
  OAI211_X1 U22023 ( .C1(n19791), .C2(n19925), .A(n19782), .B(n19781), .ZN(
        P2_U3122) );
  AOI22_X1 U22024 ( .A1(n19831), .A2(n19804), .B1(n19802), .B2(n19920), .ZN(
        n19784) );
  AOI22_X1 U22025 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19805), .ZN(n19783) );
  OAI211_X1 U22026 ( .C1(n19791), .C2(n19837), .A(n19784), .B(n19783), .ZN(
        P2_U3114) );
  AOI22_X1 U22027 ( .A1(n19927), .A2(n19805), .B1(n19926), .B2(n19802), .ZN(
        n19786) );
  AOI22_X1 U22028 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19929), .B1(
        n19928), .B2(n19804), .ZN(n19785) );
  OAI211_X1 U22029 ( .C1(n19791), .C2(n19937), .A(n19786), .B(n19785), .ZN(
        P2_U3106) );
  AOI22_X1 U22030 ( .A1(n19933), .A2(n19805), .B1(n19932), .B2(n19802), .ZN(
        n19788) );
  AOI22_X1 U22031 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19934), .B1(
        n19939), .B2(n19803), .ZN(n19787) );
  OAI211_X1 U22032 ( .C1(n19801), .C2(n19937), .A(n19788), .B(n19787), .ZN(
        P2_U3098) );
  AOI22_X1 U22033 ( .A1(n19804), .A2(n19939), .B1(n19938), .B2(n19802), .ZN(
        n19790) );
  AOI22_X1 U22034 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19941), .B1(
        n19805), .B2(n19940), .ZN(n19789) );
  OAI211_X1 U22035 ( .C1(n19791), .C2(n19944), .A(n19790), .B(n19789), .ZN(
        P2_U3090) );
  INV_X1 U22036 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19794) );
  AOI22_X1 U22037 ( .A1(n19804), .A2(n19946), .B1(n19945), .B2(n19802), .ZN(
        n19793) );
  AOI22_X1 U22038 ( .A1(n19805), .A2(n19947), .B1(n19953), .B2(n19803), .ZN(
        n19792) );
  OAI211_X1 U22039 ( .C1(n19951), .C2(n19794), .A(n19793), .B(n19792), .ZN(
        P2_U3082) );
  AOI22_X1 U22040 ( .A1(n19846), .A2(n19803), .B1(n19952), .B2(n19802), .ZN(
        n19796) );
  AOI22_X1 U22041 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19955), .B1(
        n19805), .B2(n19954), .ZN(n19795) );
  OAI211_X1 U22042 ( .C1(n19801), .C2(n19849), .A(n19796), .B(n19795), .ZN(
        P2_U3074) );
  AOI22_X1 U22043 ( .A1(n19960), .A2(n19805), .B1(n19802), .B2(n19959), .ZN(
        n19798) );
  AOI22_X1 U22044 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n19803), .ZN(n19797) );
  OAI211_X1 U22045 ( .C1(n19801), .C2(n19965), .A(n19798), .B(n19797), .ZN(
        P2_U3066) );
  AOI22_X1 U22046 ( .A1(n19967), .A2(n19805), .B1(n19802), .B2(n19966), .ZN(
        n19800) );
  AOI22_X1 U22047 ( .A1(n19968), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n19978), .B2(n19803), .ZN(n19799) );
  OAI211_X1 U22048 ( .C1(n19801), .C2(n19971), .A(n19800), .B(n19799), .ZN(
        P2_U3058) );
  AOI22_X1 U22049 ( .A1(n19975), .A2(n19803), .B1(n19974), .B2(n19802), .ZN(
        n19807) );
  AOI22_X1 U22050 ( .A1(n19805), .A2(n19979), .B1(n19978), .B2(n19804), .ZN(
        n19806) );
  OAI211_X1 U22051 ( .C1(n19984), .C2(n19808), .A(n19807), .B(n19806), .ZN(
        P2_U3050) );
  AOI22_X1 U22052 ( .A1(n19860), .A2(n19809), .B1(n19859), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19815) );
  AOI21_X1 U22053 ( .B1(n19811), .B2(n19861), .A(n19810), .ZN(n19813) );
  OR2_X1 U22054 ( .A1(n19813), .A2(n19812), .ZN(n19814) );
  OAI211_X1 U22055 ( .C1(n19816), .C2(n19868), .A(n19815), .B(n19814), .ZN(
        P2_U2918) );
  AOI22_X1 U22056 ( .A1(n19874), .A2(n17376), .B1(n19873), .B2(n19853), .ZN(
        n19818) );
  INV_X1 U22057 ( .A(n19852), .ZN(n19855) );
  AOI22_X1 U22058 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19877), .B1(
        n19975), .B2(n19855), .ZN(n19817) );
  OAI211_X1 U22059 ( .C1(n19842), .C2(n19886), .A(n19818), .B(n19817), .ZN(
        P2_U3169) );
  AOI22_X1 U22060 ( .A1(n19881), .A2(n17376), .B1(n19880), .B2(n19853), .ZN(
        n19820) );
  AOI22_X1 U22061 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19854), .ZN(n19819) );
  OAI211_X1 U22062 ( .C1(n19852), .C2(n19886), .A(n19820), .B(n19819), .ZN(
        P2_U3161) );
  AOI22_X1 U22063 ( .A1(n19888), .A2(n17376), .B1(n19853), .B2(n19887), .ZN(
        n19822) );
  AOI22_X1 U22064 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19890), .B1(
        n19882), .B2(n19855), .ZN(n19821) );
  OAI211_X1 U22065 ( .C1(n19842), .C2(n19899), .A(n19822), .B(n19821), .ZN(
        P2_U3153) );
  AOI22_X1 U22066 ( .A1(n19895), .A2(n17376), .B1(n19894), .B2(n19853), .ZN(
        n19824) );
  AOI22_X1 U22067 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19896), .B1(
        n19902), .B2(n19854), .ZN(n19823) );
  OAI211_X1 U22068 ( .C1(n19852), .C2(n19899), .A(n19824), .B(n19823), .ZN(
        P2_U3145) );
  AOI22_X1 U22069 ( .A1(n19901), .A2(n17376), .B1(n19900), .B2(n19853), .ZN(
        n19826) );
  AOI22_X1 U22070 ( .A1(n19902), .A2(n19855), .B1(n19903), .B2(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n19825) );
  OAI211_X1 U22071 ( .C1(n19842), .C2(n19906), .A(n19826), .B(n19825), .ZN(
        P2_U3137) );
  AOI22_X1 U22072 ( .A1(n19915), .A2(n19854), .B1(n19853), .B2(n19907), .ZN(
        n19828) );
  AOI22_X1 U22073 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19910), .B1(
        n17376), .B2(n19909), .ZN(n19827) );
  OAI211_X1 U22074 ( .C1(n19852), .C2(n19906), .A(n19828), .B(n19827), .ZN(
        P2_U3129) );
  AOI22_X1 U22075 ( .A1(n19915), .A2(n19855), .B1(n19853), .B2(n19914), .ZN(
        n19830) );
  AOI22_X1 U22076 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n17376), .ZN(n19829) );
  OAI211_X1 U22077 ( .C1(n19842), .C2(n19925), .A(n19830), .B(n19829), .ZN(
        P2_U3121) );
  AOI22_X1 U22078 ( .A1(n19831), .A2(n19855), .B1(n19853), .B2(n19920), .ZN(
        n19833) );
  AOI22_X1 U22079 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n17376), .ZN(n19832) );
  OAI211_X1 U22080 ( .C1(n19842), .C2(n19837), .A(n19833), .B(n19832), .ZN(
        P2_U3113) );
  AOI22_X1 U22081 ( .A1(n19927), .A2(n17376), .B1(n19926), .B2(n19853), .ZN(
        n19836) );
  AOI22_X1 U22082 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19929), .B1(
        n19834), .B2(n19854), .ZN(n19835) );
  OAI211_X1 U22083 ( .C1(n19852), .C2(n19837), .A(n19836), .B(n19835), .ZN(
        P2_U3105) );
  AOI22_X1 U22084 ( .A1(n19933), .A2(n17376), .B1(n19932), .B2(n19853), .ZN(
        n19839) );
  AOI22_X1 U22085 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19934), .B1(
        n19939), .B2(n19854), .ZN(n19838) );
  OAI211_X1 U22086 ( .C1(n19852), .C2(n19937), .A(n19839), .B(n19838), .ZN(
        P2_U3097) );
  AOI22_X1 U22087 ( .A1(n19855), .A2(n19939), .B1(n19938), .B2(n19853), .ZN(
        n19841) );
  AOI22_X1 U22088 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19941), .B1(
        n17376), .B2(n19940), .ZN(n19840) );
  OAI211_X1 U22089 ( .C1(n19842), .C2(n19944), .A(n19841), .B(n19840), .ZN(
        P2_U3089) );
  INV_X1 U22090 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n19845) );
  AOI22_X1 U22091 ( .A1(n19855), .A2(n19946), .B1(n19945), .B2(n19853), .ZN(
        n19844) );
  AOI22_X1 U22092 ( .A1(n17376), .A2(n19947), .B1(n19953), .B2(n19854), .ZN(
        n19843) );
  OAI211_X1 U22093 ( .C1(n19951), .C2(n19845), .A(n19844), .B(n19843), .ZN(
        P2_U3081) );
  AOI22_X1 U22094 ( .A1(n19854), .A2(n19846), .B1(n19952), .B2(n19853), .ZN(
        n19848) );
  AOI22_X1 U22095 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19955), .B1(
        n17376), .B2(n19954), .ZN(n19847) );
  OAI211_X1 U22096 ( .C1(n19852), .C2(n19849), .A(n19848), .B(n19847), .ZN(
        P2_U3073) );
  AOI22_X1 U22097 ( .A1(n19967), .A2(n17376), .B1(n19853), .B2(n19966), .ZN(
        n19851) );
  AOI22_X1 U22098 ( .A1(n19968), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n19854), .B2(n19978), .ZN(n19850) );
  OAI211_X1 U22099 ( .C1(n19852), .C2(n19971), .A(n19851), .B(n19850), .ZN(
        P2_U3057) );
  AOI22_X1 U22100 ( .A1(n19975), .A2(n19854), .B1(n19974), .B2(n19853), .ZN(
        n19857) );
  AOI22_X1 U22101 ( .A1(n17376), .A2(n19979), .B1(n19978), .B2(n19855), .ZN(
        n19856) );
  OAI211_X1 U22102 ( .C1(n19984), .C2(n19858), .A(n19857), .B(n19856), .ZN(
        P2_U3049) );
  AOI22_X1 U22103 ( .A1(n19860), .A2(n19864), .B1(n19859), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19867) );
  INV_X1 U22104 ( .A(n19861), .ZN(n19863) );
  OAI211_X1 U22105 ( .C1(n19865), .C2(n19864), .A(n19863), .B(n19862), .ZN(
        n19866) );
  OAI211_X1 U22106 ( .C1(n19870), .C2(n19868), .A(n19867), .B(n19866), .ZN(
        P2_U2919) );
  AOI22_X1 U22107 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19875), .ZN(n19958) );
  NOR2_X2 U22108 ( .A1(n19870), .A2(n19869), .ZN(n19980) );
  NOR2_X2 U22109 ( .A1(n19872), .A2(n19871), .ZN(n19973) );
  AOI22_X1 U22110 ( .A1(n19874), .A2(n19980), .B1(n19873), .B2(n19973), .ZN(
        n19879) );
  AOI22_X1 U22111 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19876), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19875), .ZN(n19972) );
  INV_X1 U22112 ( .A(n19972), .ZN(n19977) );
  AOI22_X1 U22113 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19877), .B1(
        n19975), .B2(n19977), .ZN(n19878) );
  OAI211_X1 U22114 ( .C1(n19958), .C2(n19886), .A(n19879), .B(n19878), .ZN(
        P2_U3168) );
  AOI22_X1 U22115 ( .A1(n19881), .A2(n19980), .B1(n19880), .B2(n19973), .ZN(
        n19885) );
  AOI22_X1 U22116 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19976), .ZN(n19884) );
  OAI211_X1 U22117 ( .C1(n19972), .C2(n19886), .A(n19885), .B(n19884), .ZN(
        P2_U3160) );
  AOI22_X1 U22118 ( .A1(n19888), .A2(n19980), .B1(n19973), .B2(n19887), .ZN(
        n19892) );
  AOI22_X1 U22119 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19890), .B1(
        n19889), .B2(n19976), .ZN(n19891) );
  OAI211_X1 U22120 ( .C1(n19972), .C2(n19893), .A(n19892), .B(n19891), .ZN(
        P2_U3152) );
  AOI22_X1 U22121 ( .A1(n19895), .A2(n19980), .B1(n19894), .B2(n19973), .ZN(
        n19898) );
  AOI22_X1 U22122 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19896), .B1(
        n19902), .B2(n19976), .ZN(n19897) );
  OAI211_X1 U22123 ( .C1(n19972), .C2(n19899), .A(n19898), .B(n19897), .ZN(
        P2_U3144) );
  AOI22_X1 U22124 ( .A1(n19901), .A2(n19980), .B1(n19900), .B2(n19973), .ZN(
        n19905) );
  AOI22_X1 U22125 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19903), .B1(
        n19977), .B2(n19902), .ZN(n19904) );
  OAI211_X1 U22126 ( .C1(n19958), .C2(n19906), .A(n19905), .B(n19904), .ZN(
        P2_U3136) );
  AOI22_X1 U22127 ( .A1(n19908), .A2(n19977), .B1(n19973), .B2(n19907), .ZN(
        n19912) );
  AOI22_X1 U22128 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19910), .B1(
        n19980), .B2(n19909), .ZN(n19911) );
  OAI211_X1 U22129 ( .C1(n19958), .C2(n19913), .A(n19912), .B(n19911), .ZN(
        P2_U3128) );
  AOI22_X1 U22130 ( .A1(n19915), .A2(n19977), .B1(n19973), .B2(n19914), .ZN(
        n19919) );
  AOI22_X1 U22131 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19980), .ZN(n19918) );
  OAI211_X1 U22132 ( .C1(n19958), .C2(n19925), .A(n19919), .B(n19918), .ZN(
        P2_U3120) );
  AOI22_X1 U22133 ( .A1(n19976), .A2(n19928), .B1(n19973), .B2(n19920), .ZN(
        n19924) );
  AOI22_X1 U22134 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19980), .ZN(n19923) );
  OAI211_X1 U22135 ( .C1(n19972), .C2(n19925), .A(n19924), .B(n19923), .ZN(
        P2_U3112) );
  AOI22_X1 U22136 ( .A1(n19927), .A2(n19980), .B1(n19926), .B2(n19973), .ZN(
        n19931) );
  AOI22_X1 U22137 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19929), .B1(
        n19928), .B2(n19977), .ZN(n19930) );
  OAI211_X1 U22138 ( .C1(n19958), .C2(n19937), .A(n19931), .B(n19930), .ZN(
        P2_U3104) );
  AOI22_X1 U22139 ( .A1(n19933), .A2(n19980), .B1(n19932), .B2(n19973), .ZN(
        n19936) );
  AOI22_X1 U22140 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19934), .B1(
        n19939), .B2(n19976), .ZN(n19935) );
  OAI211_X1 U22141 ( .C1(n19972), .C2(n19937), .A(n19936), .B(n19935), .ZN(
        P2_U3096) );
  AOI22_X1 U22142 ( .A1(n19977), .A2(n19939), .B1(n19938), .B2(n19973), .ZN(
        n19943) );
  AOI22_X1 U22143 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19941), .B1(
        n19980), .B2(n19940), .ZN(n19942) );
  OAI211_X1 U22144 ( .C1(n19958), .C2(n19944), .A(n19943), .B(n19942), .ZN(
        P2_U3088) );
  INV_X1 U22145 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19950) );
  AOI22_X1 U22146 ( .A1(n19977), .A2(n19946), .B1(n19945), .B2(n19973), .ZN(
        n19949) );
  AOI22_X1 U22147 ( .A1(n19980), .A2(n19947), .B1(n19953), .B2(n19976), .ZN(
        n19948) );
  OAI211_X1 U22148 ( .C1(n19951), .C2(n19950), .A(n19949), .B(n19948), .ZN(
        P2_U3080) );
  AOI22_X1 U22149 ( .A1(n19977), .A2(n19953), .B1(n19952), .B2(n19973), .ZN(
        n19957) );
  AOI22_X1 U22150 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19955), .B1(
        n19980), .B2(n19954), .ZN(n19956) );
  OAI211_X1 U22151 ( .C1(n19958), .C2(n19965), .A(n19957), .B(n19956), .ZN(
        P2_U3072) );
  AOI22_X1 U22152 ( .A1(n19960), .A2(n19980), .B1(n19973), .B2(n19959), .ZN(
        n19964) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19962), .B1(
        n19961), .B2(n19976), .ZN(n19963) );
  OAI211_X1 U22154 ( .C1(n19972), .C2(n19965), .A(n19964), .B(n19963), .ZN(
        P2_U3064) );
  AOI22_X1 U22155 ( .A1(n19967), .A2(n19980), .B1(n19973), .B2(n19966), .ZN(
        n19970) );
  AOI22_X1 U22156 ( .A1(n19968), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n19976), .B2(n19978), .ZN(n19969) );
  OAI211_X1 U22157 ( .C1(n19972), .C2(n19971), .A(n19970), .B(n19969), .ZN(
        P2_U3056) );
  AOI22_X1 U22158 ( .A1(n19976), .A2(n19975), .B1(n19974), .B2(n19973), .ZN(
        n19982) );
  AOI22_X1 U22159 ( .A1(n19980), .A2(n19979), .B1(n19978), .B2(n19977), .ZN(
        n19981) );
  OAI211_X1 U22160 ( .C1(n19984), .C2(n19983), .A(n19982), .B(n19981), .ZN(
        P2_U3048) );
  INV_X1 U22161 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20307) );
  INV_X1 U22162 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n19985) );
  AOI222_X1 U22163 ( .A1(n20307), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20310), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n19985), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n19986) );
  OAI22_X1 U22164 ( .A1(n20029), .A2(P3_ADDRESS_REG_0__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n20034), .ZN(n19987) );
  INV_X1 U22165 ( .A(n19987), .ZN(U376) );
  OAI22_X1 U22166 ( .A1(n20029), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n20034), .ZN(n19988) );
  INV_X1 U22167 ( .A(n19988), .ZN(U365) );
  OAI22_X1 U22168 ( .A1(n20029), .A2(P3_ADDRESS_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n20034), .ZN(n19989) );
  INV_X1 U22169 ( .A(n19989), .ZN(U354) );
  OAI22_X1 U22170 ( .A1(n20029), .A2(P3_ADDRESS_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n20034), .ZN(n19990) );
  INV_X1 U22171 ( .A(n19990), .ZN(U353) );
  OAI22_X1 U22172 ( .A1(n20029), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n20034), .ZN(n19991) );
  INV_X1 U22173 ( .A(n19991), .ZN(U352) );
  OAI22_X1 U22174 ( .A1(n20029), .A2(P3_ADDRESS_REG_5__SCAN_IN), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(n19986), .ZN(n19992) );
  INV_X1 U22175 ( .A(n19992), .ZN(U351) );
  INV_X2 U22176 ( .A(n20029), .ZN(n20034) );
  OAI22_X1 U22177 ( .A1(n20029), .A2(P3_ADDRESS_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n20034), .ZN(n19993) );
  INV_X1 U22178 ( .A(n19993), .ZN(U350) );
  AOI22_X1 U22179 ( .A1(n20034), .A2(n19995), .B1(n19994), .B2(n20029), .ZN(
        U349) );
  AOI22_X1 U22180 ( .A1(n20034), .A2(n19997), .B1(n19996), .B2(n20029), .ZN(
        U348) );
  AOI22_X1 U22181 ( .A1(n20034), .A2(n19999), .B1(n19998), .B2(n20029), .ZN(
        U347) );
  AOI22_X1 U22182 ( .A1(n20034), .A2(n20001), .B1(n20000), .B2(n20029), .ZN(
        U375) );
  OAI22_X1 U22183 ( .A1(n20029), .A2(P3_ADDRESS_REG_11__SCAN_IN), .B1(
        P2_ADDRESS_REG_11__SCAN_IN), .B2(n20034), .ZN(n20002) );
  INV_X1 U22184 ( .A(n20002), .ZN(U374) );
  OAI22_X1 U22185 ( .A1(n20029), .A2(P3_ADDRESS_REG_12__SCAN_IN), .B1(
        P2_ADDRESS_REG_12__SCAN_IN), .B2(n20034), .ZN(n20003) );
  INV_X1 U22186 ( .A(n20003), .ZN(U373) );
  OAI22_X1 U22187 ( .A1(n20029), .A2(P3_ADDRESS_REG_13__SCAN_IN), .B1(
        P2_ADDRESS_REG_13__SCAN_IN), .B2(n20034), .ZN(n20004) );
  INV_X1 U22188 ( .A(n20004), .ZN(U372) );
  AOI22_X1 U22189 ( .A1(n20034), .A2(n20006), .B1(n20005), .B2(n20029), .ZN(
        U371) );
  AOI22_X1 U22190 ( .A1(n20034), .A2(n20008), .B1(n20007), .B2(n20029), .ZN(
        U370) );
  AOI22_X1 U22191 ( .A1(n20034), .A2(n20010), .B1(n20009), .B2(n20029), .ZN(
        U369) );
  AOI22_X1 U22192 ( .A1(n20034), .A2(n20012), .B1(n20011), .B2(n20029), .ZN(
        U368) );
  OAI22_X1 U22193 ( .A1(n20029), .A2(P3_ADDRESS_REG_18__SCAN_IN), .B1(
        P2_ADDRESS_REG_18__SCAN_IN), .B2(n20034), .ZN(n20013) );
  INV_X1 U22194 ( .A(n20013), .ZN(U367) );
  OAI22_X1 U22195 ( .A1(n20029), .A2(P3_ADDRESS_REG_19__SCAN_IN), .B1(
        P2_ADDRESS_REG_19__SCAN_IN), .B2(n20034), .ZN(n20014) );
  INV_X1 U22196 ( .A(n20014), .ZN(U366) );
  INV_X1 U22197 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U22198 ( .A1(n20034), .A2(n20016), .B1(n20015), .B2(n20029), .ZN(
        U364) );
  OAI22_X1 U22199 ( .A1(n20029), .A2(P3_ADDRESS_REG_21__SCAN_IN), .B1(
        P2_ADDRESS_REG_21__SCAN_IN), .B2(n20034), .ZN(n20017) );
  INV_X1 U22200 ( .A(n20017), .ZN(U363) );
  OAI22_X1 U22201 ( .A1(n20029), .A2(P3_ADDRESS_REG_22__SCAN_IN), .B1(
        P2_ADDRESS_REG_22__SCAN_IN), .B2(n20034), .ZN(n20018) );
  INV_X1 U22202 ( .A(n20018), .ZN(U362) );
  AOI22_X1 U22203 ( .A1(n20034), .A2(n20020), .B1(n20019), .B2(n20029), .ZN(
        U361) );
  AOI22_X1 U22204 ( .A1(n19986), .A2(n20022), .B1(n20021), .B2(n20029), .ZN(
        U360) );
  AOI22_X1 U22205 ( .A1(n20034), .A2(n20024), .B1(n20023), .B2(n20029), .ZN(
        U359) );
  AOI22_X1 U22206 ( .A1(n20034), .A2(n20026), .B1(n20025), .B2(n20029), .ZN(
        U358) );
  AOI22_X1 U22207 ( .A1(n20034), .A2(n20028), .B1(n20027), .B2(n20029), .ZN(
        U357) );
  AOI22_X1 U22208 ( .A1(n19986), .A2(n20031), .B1(n20030), .B2(n20029), .ZN(
        U356) );
  AOI22_X1 U22209 ( .A1(n20034), .A2(n20033), .B1(n20032), .B2(n20029), .ZN(
        U355) );
  AOI22_X1 U22210 ( .A1(n21456), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20036) );
  OAI21_X1 U22211 ( .B1(n20037), .B2(n20066), .A(n20036), .ZN(P1_U2936) );
  AOI22_X1 U22212 ( .A1(n20053), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20038) );
  OAI21_X1 U22213 ( .B1(n20039), .B2(n20066), .A(n20038), .ZN(P1_U2935) );
  AOI22_X1 U22214 ( .A1(n20053), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20040) );
  OAI21_X1 U22215 ( .B1(n20041), .B2(n20066), .A(n20040), .ZN(P1_U2934) );
  AOI22_X1 U22216 ( .A1(n20053), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20042) );
  OAI21_X1 U22217 ( .B1(n20043), .B2(n20066), .A(n20042), .ZN(P1_U2933) );
  AOI22_X1 U22218 ( .A1(n20053), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20044) );
  OAI21_X1 U22219 ( .B1(n20045), .B2(n20066), .A(n20044), .ZN(P1_U2932) );
  AOI22_X1 U22220 ( .A1(n20053), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20046) );
  OAI21_X1 U22221 ( .B1(n13283), .B2(n20066), .A(n20046), .ZN(P1_U2931) );
  AOI22_X1 U22222 ( .A1(n20053), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20047) );
  OAI21_X1 U22223 ( .B1(n13290), .B2(n20066), .A(n20047), .ZN(P1_U2930) );
  AOI22_X1 U22224 ( .A1(n20053), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20048) );
  OAI21_X1 U22225 ( .B1(n13294), .B2(n20066), .A(n20048), .ZN(P1_U2929) );
  AOI22_X1 U22226 ( .A1(n20053), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20049) );
  OAI21_X1 U22227 ( .B1(n20050), .B2(n20066), .A(n20049), .ZN(P1_U2928) );
  AOI22_X1 U22228 ( .A1(n21456), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20051) );
  OAI21_X1 U22229 ( .B1(n20052), .B2(n20066), .A(n20051), .ZN(P1_U2927) );
  AOI22_X1 U22230 ( .A1(n20053), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20054) );
  OAI21_X1 U22231 ( .B1(n20055), .B2(n20066), .A(n20054), .ZN(P1_U2926) );
  AOI22_X1 U22232 ( .A1(n21456), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20056) );
  OAI21_X1 U22233 ( .B1(n20057), .B2(n20066), .A(n20056), .ZN(P1_U2925) );
  AOI22_X1 U22234 ( .A1(n21456), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20058) );
  OAI21_X1 U22235 ( .B1(n20059), .B2(n20066), .A(n20058), .ZN(P1_U2924) );
  AOI22_X1 U22236 ( .A1(n21456), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20061) );
  OAI21_X1 U22237 ( .B1(n20062), .B2(n20066), .A(n20061), .ZN(P1_U2923) );
  AOI22_X1 U22238 ( .A1(n21456), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20063) );
  OAI21_X1 U22239 ( .B1(n20064), .B2(n20066), .A(n20063), .ZN(P1_U2922) );
  AOI22_X1 U22240 ( .A1(n21456), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20060), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20065) );
  OAI21_X1 U22241 ( .B1(n20067), .B2(n20066), .A(n20065), .ZN(P1_U2921) );
  INV_X1 U22242 ( .A(n20104), .ZN(n20090) );
  OAI222_X1 U22243 ( .A1(n20092), .A2(n21673), .B1(n20068), .B2(n22398), .C1(
        n21674), .C2(n20090), .ZN(P1_U3197) );
  INV_X1 U22244 ( .A(n20092), .ZN(n20103) );
  AOI222_X1 U22245 ( .A1(n20103), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n20104), .ZN(n20069) );
  INV_X1 U22246 ( .A(n20069), .ZN(P1_U3198) );
  AOI222_X1 U22247 ( .A1(n20103), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20104), .ZN(n20070) );
  INV_X1 U22248 ( .A(n20070), .ZN(P1_U3199) );
  AOI222_X1 U22249 ( .A1(n20103), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20104), .ZN(n20071) );
  INV_X1 U22250 ( .A(n20071), .ZN(P1_U3200) );
  AOI22_X1 U22251 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20103), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20100), .ZN(n20072) );
  OAI21_X1 U22252 ( .B1(n21696), .B2(n20090), .A(n20072), .ZN(P1_U3201) );
  AOI22_X1 U22253 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20104), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20100), .ZN(n20073) );
  OAI21_X1 U22254 ( .B1(n21717), .B2(n20092), .A(n20073), .ZN(P1_U3202) );
  AOI22_X1 U22255 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20103), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20100), .ZN(n20074) );
  OAI21_X1 U22256 ( .B1(n21717), .B2(n20090), .A(n20074), .ZN(P1_U3203) );
  AOI22_X1 U22257 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20104), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20100), .ZN(n20075) );
  OAI21_X1 U22258 ( .B1(n21743), .B2(n20092), .A(n20075), .ZN(P1_U3204) );
  AOI22_X1 U22259 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20103), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20100), .ZN(n20076) );
  OAI21_X1 U22260 ( .B1(n21743), .B2(n20090), .A(n20076), .ZN(P1_U3205) );
  AOI22_X1 U22261 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20104), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20100), .ZN(n20077) );
  OAI21_X1 U22262 ( .B1(n20078), .B2(n20092), .A(n20077), .ZN(P1_U3206) );
  AOI222_X1 U22263 ( .A1(n20103), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20104), .ZN(n20079) );
  INV_X1 U22264 ( .A(n20079), .ZN(P1_U3207) );
  AOI222_X1 U22265 ( .A1(n20103), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20104), .ZN(n20080) );
  INV_X1 U22266 ( .A(n20080), .ZN(P1_U3208) );
  AOI22_X1 U22267 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n20103), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20100), .ZN(n20081) );
  OAI21_X1 U22268 ( .B1(n20082), .B2(n20090), .A(n20081), .ZN(P1_U3209) );
  INV_X1 U22269 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20084) );
  AOI22_X1 U22270 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n20103), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20100), .ZN(n20083) );
  OAI21_X1 U22271 ( .B1(n20084), .B2(n20090), .A(n20083), .ZN(P1_U3210) );
  AOI22_X1 U22272 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n20104), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n22395), .ZN(n20085) );
  OAI21_X1 U22273 ( .B1(n21745), .B2(n20092), .A(n20085), .ZN(P1_U3211) );
  AOI22_X1 U22274 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n20103), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n22395), .ZN(n20086) );
  OAI21_X1 U22275 ( .B1(n21745), .B2(n20090), .A(n20086), .ZN(P1_U3212) );
  AOI22_X1 U22276 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n20104), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n22395), .ZN(n20087) );
  OAI21_X1 U22277 ( .B1(n21757), .B2(n20092), .A(n20087), .ZN(P1_U3213) );
  AOI222_X1 U22278 ( .A1(n20104), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20103), .ZN(n20088) );
  INV_X1 U22279 ( .A(n20088), .ZN(P1_U3214) );
  AOI22_X1 U22280 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n20103), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n22395), .ZN(n20089) );
  OAI21_X1 U22281 ( .B1(n21775), .B2(n20090), .A(n20089), .ZN(P1_U3215) );
  AOI22_X1 U22282 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n20104), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n22395), .ZN(n20091) );
  OAI21_X1 U22283 ( .B1(n21807), .B2(n20092), .A(n20091), .ZN(P1_U3216) );
  AOI222_X1 U22284 ( .A1(n20103), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20104), .ZN(n20093) );
  INV_X1 U22285 ( .A(n20093), .ZN(P1_U3217) );
  AOI222_X1 U22286 ( .A1(n20104), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20103), .ZN(n20094) );
  INV_X1 U22287 ( .A(n20094), .ZN(P1_U3218) );
  AOI222_X1 U22288 ( .A1(n20104), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20103), .ZN(n20095) );
  INV_X1 U22289 ( .A(n20095), .ZN(P1_U3219) );
  AOI222_X1 U22290 ( .A1(n20103), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20104), .ZN(n20096) );
  INV_X1 U22291 ( .A(n20096), .ZN(P1_U3220) );
  AOI222_X1 U22292 ( .A1(n20103), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20104), .ZN(n20097) );
  INV_X1 U22293 ( .A(n20097), .ZN(P1_U3221) );
  AOI222_X1 U22294 ( .A1(n20103), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20104), .ZN(n20098) );
  INV_X1 U22295 ( .A(n20098), .ZN(P1_U3222) );
  AOI222_X1 U22296 ( .A1(n20103), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20104), .ZN(n20099) );
  INV_X1 U22297 ( .A(n20099), .ZN(P1_U3223) );
  AOI222_X1 U22298 ( .A1(n20103), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20100), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20104), .ZN(n20101) );
  INV_X1 U22299 ( .A(n20101), .ZN(P1_U3224) );
  AOI222_X1 U22300 ( .A1(n20104), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n22395), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20103), .ZN(n20102) );
  INV_X1 U22301 ( .A(n20102), .ZN(P1_U3225) );
  AOI222_X1 U22302 ( .A1(n20104), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n22395), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20103), .ZN(n20105) );
  INV_X1 U22303 ( .A(n20105), .ZN(P1_U3226) );
  OAI22_X1 U22304 ( .A1(n22395), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22398), .ZN(n20106) );
  INV_X1 U22305 ( .A(n20106), .ZN(P1_U3458) );
  AOI221_X1 U22306 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20117) );
  NOR4_X1 U22307 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20110) );
  NOR4_X1 U22308 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20109) );
  NOR4_X1 U22309 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20108) );
  NOR4_X1 U22310 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20107) );
  NAND4_X1 U22311 ( .A1(n20110), .A2(n20109), .A3(n20108), .A4(n20107), .ZN(
        n20116) );
  NOR4_X1 U22312 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20114) );
  AOI211_X1 U22313 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20113) );
  NOR4_X1 U22314 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20112) );
  NOR4_X1 U22315 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20111) );
  NAND4_X1 U22316 ( .A1(n20114), .A2(n20113), .A3(n20112), .A4(n20111), .ZN(
        n20115) );
  NOR2_X1 U22317 ( .A1(n20116), .A2(n20115), .ZN(n20129) );
  MUX2_X1 U22318 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n20117), .S(n20129), 
        .Z(P1_U2808) );
  OAI22_X1 U22319 ( .A1(n22395), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22398), .ZN(n20118) );
  INV_X1 U22320 ( .A(n20118), .ZN(P1_U3459) );
  AOI21_X1 U22321 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20119) );
  OAI221_X1 U22322 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20119), .C1(n21674), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20129), .ZN(n20120) );
  OAI21_X1 U22323 ( .B1(n20129), .B2(n20121), .A(n20120), .ZN(P1_U3481) );
  OAI22_X1 U22324 ( .A1(n22395), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22398), .ZN(n20122) );
  INV_X1 U22325 ( .A(n20122), .ZN(P1_U3460) );
  NOR3_X1 U22326 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20123) );
  OAI21_X1 U22327 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20123), .A(n20129), .ZN(
        n20124) );
  OAI21_X1 U22328 ( .B1(n20129), .B2(n20125), .A(n20124), .ZN(P1_U2807) );
  OAI22_X1 U22329 ( .A1(n22395), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22398), .ZN(n20126) );
  INV_X1 U22330 ( .A(n20126), .ZN(P1_U3461) );
  OAI21_X1 U22331 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20129), .ZN(n20127) );
  OAI21_X1 U22332 ( .B1(n20129), .B2(n20128), .A(n20127), .ZN(P1_U3482) );
  AOI22_X1 U22333 ( .A1(n20133), .A2(n20132), .B1(n20131), .B2(n20130), .ZN(
        n20134) );
  OAI21_X1 U22334 ( .B1(n20136), .B2(n20135), .A(n20134), .ZN(P1_U2859) );
  AOI22_X1 U22335 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20142) );
  INV_X1 U22336 ( .A(n20137), .ZN(n21652) );
  OAI21_X1 U22337 ( .B1(n11018), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11017), .ZN(n21636) );
  INV_X1 U22338 ( .A(n21636), .ZN(n20140) );
  AOI22_X1 U22339 ( .A1(n21652), .A2(n20236), .B1(n20237), .B2(n20140), .ZN(
        n20141) );
  OAI211_X1 U22340 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20240), .A(
        n20142), .B(n20141), .ZN(P1_U2998) );
  AOI22_X1 U22341 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n20149) );
  OAI21_X1 U22342 ( .B1(n20145), .B2(n20144), .A(n20143), .ZN(n20146) );
  INV_X1 U22343 ( .A(n20146), .ZN(n21476) );
  AOI22_X1 U22344 ( .A1(n20147), .A2(n20236), .B1(n20237), .B2(n21476), .ZN(
        n20148) );
  OAI211_X1 U22345 ( .C1(n20240), .C2(n20150), .A(n20149), .B(n20148), .ZN(
        P1_U2997) );
  AOI22_X1 U22346 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n20157) );
  OAI21_X1 U22347 ( .B1(n11022), .B2(n20152), .A(n11021), .ZN(n20154) );
  INV_X1 U22348 ( .A(n20154), .ZN(n21493) );
  INV_X1 U22349 ( .A(n20155), .ZN(n21665) );
  AOI22_X1 U22350 ( .A1(n21493), .A2(n20237), .B1(n20236), .B2(n21665), .ZN(
        n20156) );
  OAI211_X1 U22351 ( .C1(n20240), .C2(n21667), .A(n20157), .B(n20156), .ZN(
        P1_U2996) );
  AOI22_X1 U22352 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20163) );
  OAI21_X1 U22353 ( .B1(n11019), .B2(n20159), .A(n20158), .ZN(n20161) );
  INV_X1 U22354 ( .A(n20161), .ZN(n21490) );
  AOI22_X1 U22355 ( .A1(n21490), .A2(n20237), .B1(n20236), .B2(n21680), .ZN(
        n20162) );
  OAI211_X1 U22356 ( .C1(n20240), .C2(n21676), .A(n20163), .B(n20162), .ZN(
        P1_U2995) );
  AOI22_X1 U22357 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n20170) );
  OAI21_X1 U22358 ( .B1(n20164), .B2(n20166), .A(n20165), .ZN(n20167) );
  INV_X1 U22359 ( .A(n20167), .ZN(n21507) );
  AOI22_X1 U22360 ( .A1(n21507), .A2(n20237), .B1(n20236), .B2(n20168), .ZN(
        n20169) );
  OAI211_X1 U22361 ( .C1(n20240), .C2(n21689), .A(n20170), .B(n20169), .ZN(
        P1_U2994) );
  AOI22_X1 U22362 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n20176) );
  NAND2_X1 U22363 ( .A1(n20172), .A2(n20171), .ZN(n20173) );
  NAND2_X1 U22364 ( .A1(n20174), .A2(n20173), .ZN(n21498) );
  AOI22_X1 U22365 ( .A1(n21498), .A2(n20237), .B1(n20236), .B2(n21704), .ZN(
        n20175) );
  OAI211_X1 U22366 ( .C1(n20240), .C2(n21702), .A(n20176), .B(n20175), .ZN(
        P1_U2993) );
  AOI22_X1 U22367 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n20182) );
  AOI21_X1 U22368 ( .B1(n20179), .B2(n20178), .A(n11206), .ZN(n21517) );
  AOI22_X1 U22369 ( .A1(n21517), .A2(n20237), .B1(n20236), .B2(n20180), .ZN(
        n20181) );
  OAI211_X1 U22370 ( .C1(n20240), .C2(n21712), .A(n20182), .B(n20181), .ZN(
        P1_U2992) );
  MUX2_X1 U22371 ( .A(n20184), .B(n20183), .S(n20231), .Z(n20185) );
  NAND2_X1 U22372 ( .A1(n20185), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n20190) );
  OAI21_X1 U22373 ( .B1(n20185), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n20190), .ZN(n21541) );
  AOI22_X1 U22374 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n20189) );
  AOI22_X1 U22375 ( .A1(n20187), .A2(n20236), .B1(n20222), .B2(n20186), .ZN(
        n20188) );
  OAI211_X1 U22376 ( .C1(n21822), .C2(n21541), .A(n20189), .B(n20188), .ZN(
        P1_U2989) );
  NOR2_X1 U22377 ( .A1(n11483), .A2(n12179), .ZN(n20191) );
  MUX2_X1 U22378 ( .A(n20231), .B(n20191), .S(n20190), .Z(n20192) );
  XOR2_X1 U22379 ( .A(n12191), .B(n20192), .Z(n21570) );
  AOI22_X1 U22380 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n20197) );
  INV_X1 U22381 ( .A(n20193), .ZN(n20194) );
  AOI22_X1 U22382 ( .A1(n20195), .A2(n20236), .B1(n20222), .B2(n20194), .ZN(
        n20196) );
  OAI211_X1 U22383 ( .C1(n21570), .C2(n21822), .A(n20197), .B(n20196), .ZN(
        P1_U2988) );
  OAI21_X1 U22384 ( .B1(n20200), .B2(n20199), .A(n20198), .ZN(n20201) );
  INV_X1 U22385 ( .A(n20201), .ZN(n21558) );
  AOI22_X1 U22386 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n20206) );
  NOR2_X1 U22387 ( .A1(n20240), .A2(n20202), .ZN(n20203) );
  AOI21_X1 U22388 ( .B1(n20204), .B2(n20236), .A(n20203), .ZN(n20205) );
  OAI211_X1 U22389 ( .C1(n21558), .C2(n21822), .A(n20206), .B(n20205), .ZN(
        P1_U2987) );
  XNOR2_X1 U22390 ( .A(n12179), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n20207) );
  XNOR2_X1 U22391 ( .A(n20208), .B(n20207), .ZN(n21580) );
  AOI22_X1 U22392 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n20213) );
  INV_X1 U22393 ( .A(n20209), .ZN(n20211) );
  AOI22_X1 U22394 ( .A1(n20211), .A2(n20236), .B1(n20222), .B2(n20210), .ZN(
        n20212) );
  OAI211_X1 U22395 ( .C1(n21822), .C2(n21580), .A(n20213), .B(n20212), .ZN(
        P1_U2984) );
  OAI21_X1 U22396 ( .B1(n20216), .B2(n20215), .A(n20214), .ZN(n20219) );
  NOR2_X1 U22397 ( .A1(n11209), .A2(n21589), .ZN(n20218) );
  OAI21_X1 U22398 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n12179), .A(
        n20219), .ZN(n20217) );
  OAI21_X1 U22399 ( .B1(n20219), .B2(n20218), .A(n20217), .ZN(n20220) );
  XOR2_X1 U22400 ( .A(n20220), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .Z(
        n21595) );
  AOI22_X1 U22401 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n20225) );
  AOI22_X1 U22402 ( .A1(n20223), .A2(n20236), .B1(n20222), .B2(n20221), .ZN(
        n20224) );
  OAI211_X1 U22403 ( .C1(n21595), .C2(n21822), .A(n20225), .B(n20224), .ZN(
        P1_U2982) );
  AOI22_X1 U22404 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n20229) );
  MUX2_X1 U22405 ( .A(n12197), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .S(
        n20231), .Z(n20226) );
  XNOR2_X1 U22406 ( .A(n20227), .B(n20226), .ZN(n21618) );
  AOI22_X1 U22407 ( .A1(n21618), .A2(n20237), .B1(n21772), .B2(n20236), .ZN(
        n20228) );
  OAI211_X1 U22408 ( .C1(n20240), .C2(n21767), .A(n20229), .B(n20228), .ZN(
        P1_U2980) );
  AOI22_X1 U22409 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n20230), .B1(
        n21639), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n20239) );
  OAI22_X1 U22410 ( .A1(n20231), .A2(n12355), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n12197), .ZN(n20232) );
  NOR2_X1 U22411 ( .A1(n20233), .A2(n20232), .ZN(n20234) );
  XNOR2_X1 U22412 ( .A(n20234), .B(n21629), .ZN(n21623) );
  AOI22_X1 U22413 ( .A1(n21623), .A2(n20237), .B1(n20236), .B2(n20235), .ZN(
        n20238) );
  OAI211_X1 U22414 ( .C1(n20240), .C2(n21796), .A(n20239), .B(n20238), .ZN(
        P1_U2978) );
  OAI222_X1 U22415 ( .A1(n22398), .A2(n20242), .B1(n22398), .B2(n20241), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(n22395), .ZN(P1_U2804) );
  INV_X1 U22416 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20245) );
  AOI22_X1 U22417 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n10994), .ZN(n20244) );
  OAI21_X1 U22418 ( .B1(n20245), .B2(n20309), .A(n20244), .ZN(U247) );
  INV_X1 U22419 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20247) );
  AOI22_X1 U22420 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n10994), .ZN(n20246) );
  OAI21_X1 U22421 ( .B1(n20247), .B2(n20309), .A(n20246), .ZN(U246) );
  INV_X1 U22422 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20249) );
  AOI22_X1 U22423 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n10994), .ZN(n20248) );
  OAI21_X1 U22424 ( .B1(n20249), .B2(n20309), .A(n20248), .ZN(U245) );
  INV_X1 U22425 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20251) );
  AOI22_X1 U22426 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n10994), .ZN(n20250) );
  OAI21_X1 U22427 ( .B1(n20251), .B2(n20309), .A(n20250), .ZN(U244) );
  AOI22_X1 U22428 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n10994), .ZN(n20252) );
  OAI21_X1 U22429 ( .B1(n20253), .B2(n20309), .A(n20252), .ZN(U243) );
  INV_X1 U22430 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20255) );
  AOI22_X1 U22431 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10994), .ZN(n20254) );
  OAI21_X1 U22432 ( .B1(n20255), .B2(n20309), .A(n20254), .ZN(U242) );
  AOI22_X1 U22433 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10994), .ZN(n20256) );
  OAI21_X1 U22434 ( .B1(n20257), .B2(n20309), .A(n20256), .ZN(U241) );
  INV_X1 U22435 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20259) );
  AOI22_X1 U22436 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10994), .ZN(n20258) );
  OAI21_X1 U22437 ( .B1(n20259), .B2(n20309), .A(n20258), .ZN(U240) );
  AOI22_X1 U22438 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10994), .ZN(n20260) );
  OAI21_X1 U22439 ( .B1(n20261), .B2(n20309), .A(n20260), .ZN(U239) );
  AOI22_X1 U22440 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10994), .ZN(n20262) );
  OAI21_X1 U22441 ( .B1(n20263), .B2(n20309), .A(n20262), .ZN(U238) );
  AOI22_X1 U22442 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10994), .ZN(n20264) );
  OAI21_X1 U22443 ( .B1(n20265), .B2(n20309), .A(n20264), .ZN(U237) );
  INV_X1 U22444 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20267) );
  AOI22_X1 U22445 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10994), .ZN(n20266) );
  OAI21_X1 U22446 ( .B1(n20267), .B2(n20309), .A(n20266), .ZN(U236) );
  INV_X1 U22447 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20269) );
  AOI22_X1 U22448 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10994), .ZN(n20268) );
  OAI21_X1 U22449 ( .B1(n20269), .B2(n20309), .A(n20268), .ZN(U235) );
  INV_X1 U22450 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20271) );
  AOI22_X1 U22451 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10994), .ZN(n20270) );
  OAI21_X1 U22452 ( .B1(n20271), .B2(n20309), .A(n20270), .ZN(U234) );
  INV_X1 U22453 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20273) );
  AOI22_X1 U22454 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10994), .ZN(n20272) );
  OAI21_X1 U22455 ( .B1(n20273), .B2(n20309), .A(n20272), .ZN(U233) );
  INV_X1 U22456 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20275) );
  AOI22_X1 U22457 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10994), .ZN(n20274) );
  OAI21_X1 U22458 ( .B1(n20275), .B2(n20309), .A(n20274), .ZN(U232) );
  AOI22_X1 U22459 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10994), .ZN(n20276) );
  OAI21_X1 U22460 ( .B1(n20277), .B2(n20309), .A(n20276), .ZN(U231) );
  AOI22_X1 U22461 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10994), .ZN(n20278) );
  OAI21_X1 U22462 ( .B1(n20279), .B2(n20309), .A(n20278), .ZN(U230) );
  AOI22_X1 U22463 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10994), .ZN(n20280) );
  OAI21_X1 U22464 ( .B1(n20281), .B2(n20309), .A(n20280), .ZN(U229) );
  AOI22_X1 U22465 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n10994), .ZN(n20282) );
  OAI21_X1 U22466 ( .B1(n20283), .B2(n20309), .A(n20282), .ZN(U228) );
  AOI22_X1 U22467 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n10994), .ZN(n20284) );
  OAI21_X1 U22468 ( .B1(n20285), .B2(n20309), .A(n20284), .ZN(U227) );
  AOI22_X1 U22469 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n10994), .ZN(n20286) );
  OAI21_X1 U22470 ( .B1(n20287), .B2(n20309), .A(n20286), .ZN(U226) );
  AOI22_X1 U22471 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10994), .ZN(n20288) );
  OAI21_X1 U22472 ( .B1(n20289), .B2(n20309), .A(n20288), .ZN(U225) );
  AOI22_X1 U22473 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n10994), .ZN(n20290) );
  OAI21_X1 U22474 ( .B1(n20291), .B2(n20309), .A(n20290), .ZN(U224) );
  AOI22_X1 U22475 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10994), .ZN(n20292) );
  OAI21_X1 U22476 ( .B1(n20293), .B2(n20309), .A(n20292), .ZN(U223) );
  AOI22_X1 U22477 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10994), .ZN(n20294) );
  OAI21_X1 U22478 ( .B1(n20295), .B2(n20309), .A(n20294), .ZN(U222) );
  AOI22_X1 U22479 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10994), .ZN(n20297) );
  OAI21_X1 U22480 ( .B1(n20298), .B2(n20309), .A(n20297), .ZN(U221) );
  AOI22_X1 U22481 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10994), .ZN(n20299) );
  OAI21_X1 U22482 ( .B1(n20300), .B2(n20309), .A(n20299), .ZN(U220) );
  AOI22_X1 U22483 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10994), .ZN(n20301) );
  OAI21_X1 U22484 ( .B1(n20302), .B2(n20309), .A(n20301), .ZN(U219) );
  AOI22_X1 U22485 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10994), .ZN(n20303) );
  OAI21_X1 U22486 ( .B1(n20304), .B2(n20309), .A(n20303), .ZN(U218) );
  AOI22_X1 U22487 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20296), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10994), .ZN(n20305) );
  OAI21_X1 U22488 ( .B1(n20306), .B2(n20309), .A(n20305), .ZN(U217) );
  OAI222_X1 U22489 ( .A1(U212), .A2(n20310), .B1(n20309), .B2(n20308), .C1(
        U214), .C2(n20307), .ZN(U216) );
  INV_X1 U22490 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20311) );
  AOI22_X1 U22491 ( .A1(n22398), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20311), 
        .B2(n22395), .ZN(P1_U3483) );
  OAI21_X1 U22492 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20779), .A(n20312), 
        .ZN(n20313) );
  AOI211_X1 U22493 ( .C1(n20314), .C2(n20313), .A(n21900), .B(n21417), .ZN(
        n20315) );
  OAI21_X1 U22494 ( .B1(n20315), .B2(n21438), .A(n21430), .ZN(n20321) );
  OAI21_X1 U22495 ( .B1(n21900), .B2(n20317), .A(n20316), .ZN(n20318) );
  AOI21_X1 U22496 ( .B1(n20319), .B2(n21414), .A(n20318), .ZN(n20320) );
  MUX2_X1 U22497 ( .A(n20321), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n20320), 
        .Z(P3_U3296) );
  AND2_X2 U22498 ( .A1(n20323), .A2(n20782), .ZN(n20364) );
  AOI22_X1 U22499 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20363), .ZN(n20325) );
  OAI21_X1 U22500 ( .B1(n20941), .B2(n20366), .A(n20325), .ZN(P3_U2768) );
  AOI22_X1 U22501 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20363), .ZN(n20326) );
  OAI21_X1 U22502 ( .B1(n20878), .B2(n20366), .A(n20326), .ZN(P3_U2769) );
  AOI22_X1 U22503 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20363), .ZN(n20327) );
  OAI21_X1 U22504 ( .B1(n20859), .B2(n20366), .A(n20327), .ZN(P3_U2770) );
  AOI22_X1 U22505 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20363), .ZN(n20328) );
  OAI21_X1 U22506 ( .B1(n20861), .B2(n20366), .A(n20328), .ZN(P3_U2771) );
  AOI22_X1 U22507 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20363), .ZN(n20329) );
  OAI21_X1 U22508 ( .B1(n20860), .B2(n20366), .A(n20329), .ZN(P3_U2772) );
  AOI22_X1 U22509 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20357), .ZN(n20330) );
  OAI21_X1 U22510 ( .B1(n20858), .B2(n20366), .A(n20330), .ZN(P3_U2773) );
  AOI22_X1 U22511 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20357), .ZN(n20331) );
  OAI21_X1 U22512 ( .B1(n20862), .B2(n20366), .A(n20331), .ZN(P3_U2774) );
  AOI22_X1 U22513 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20357), .ZN(n20332) );
  OAI21_X1 U22514 ( .B1(n20930), .B2(n20366), .A(n20332), .ZN(P3_U2775) );
  AOI22_X1 U22515 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20357), .ZN(n20333) );
  OAI21_X1 U22516 ( .B1(n20922), .B2(n20366), .A(n20333), .ZN(P3_U2776) );
  AOI22_X1 U22517 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20357), .ZN(n20334) );
  OAI21_X1 U22518 ( .B1(n20885), .B2(n20366), .A(n20334), .ZN(P3_U2777) );
  AOI22_X1 U22519 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20357), .ZN(n20335) );
  OAI21_X1 U22520 ( .B1(n20336), .B2(n20366), .A(n20335), .ZN(P3_U2778) );
  AOI22_X1 U22521 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20357), .ZN(n20337) );
  OAI21_X1 U22522 ( .B1(n20915), .B2(n20366), .A(n20337), .ZN(P3_U2779) );
  AOI22_X1 U22523 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20363), .ZN(n20338) );
  OAI21_X1 U22524 ( .B1(n20339), .B2(n20366), .A(n20338), .ZN(P3_U2780) );
  AOI22_X1 U22525 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20363), .ZN(n20340) );
  OAI21_X1 U22526 ( .B1(n20341), .B2(n20366), .A(n20340), .ZN(P3_U2781) );
  AOI22_X1 U22527 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20364), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20363), .ZN(n20342) );
  OAI21_X1 U22528 ( .B1(n20903), .B2(n20366), .A(n20342), .ZN(P3_U2782) );
  AOI22_X1 U22529 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20363), .ZN(n20343) );
  OAI21_X1 U22530 ( .B1(n20976), .B2(n20366), .A(n20343), .ZN(P3_U2783) );
  AOI22_X1 U22531 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20363), .ZN(n20344) );
  OAI21_X1 U22532 ( .B1(n20345), .B2(n20366), .A(n20344), .ZN(P3_U2784) );
  AOI22_X1 U22533 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20363), .ZN(n20346) );
  OAI21_X1 U22534 ( .B1(n20774), .B2(n20366), .A(n20346), .ZN(P3_U2785) );
  AOI22_X1 U22535 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20363), .ZN(n20347) );
  OAI21_X1 U22536 ( .B1(n20775), .B2(n20366), .A(n20347), .ZN(P3_U2786) );
  AOI22_X1 U22537 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20363), .ZN(n20348) );
  OAI21_X1 U22538 ( .B1(n20824), .B2(n20366), .A(n20348), .ZN(P3_U2787) );
  AOI22_X1 U22539 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20363), .ZN(n20349) );
  OAI21_X1 U22540 ( .B1(n20772), .B2(n20366), .A(n20349), .ZN(P3_U2788) );
  AOI22_X1 U22541 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20363), .ZN(n20350) );
  OAI21_X1 U22542 ( .B1(n20811), .B2(n20366), .A(n20350), .ZN(P3_U2789) );
  AOI22_X1 U22543 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20363), .ZN(n20351) );
  OAI21_X1 U22544 ( .B1(n20773), .B2(n20366), .A(n20351), .ZN(P3_U2790) );
  AOI22_X1 U22545 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20363), .ZN(n20352) );
  OAI21_X1 U22546 ( .B1(n20963), .B2(n20366), .A(n20352), .ZN(P3_U2791) );
  AOI22_X1 U22547 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20357), .ZN(n20353) );
  OAI21_X1 U22548 ( .B1(n20783), .B2(n20366), .A(n20353), .ZN(P3_U2792) );
  AOI22_X1 U22549 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20357), .ZN(n20354) );
  OAI21_X1 U22550 ( .B1(n20802), .B2(n20366), .A(n20354), .ZN(P3_U2793) );
  AOI22_X1 U22551 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20357), .ZN(n20355) );
  OAI21_X1 U22552 ( .B1(n20356), .B2(n20366), .A(n20355), .ZN(P3_U2794) );
  AOI22_X1 U22553 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20357), .ZN(n20358) );
  OAI21_X1 U22554 ( .B1(n20359), .B2(n20366), .A(n20358), .ZN(P3_U2795) );
  AOI22_X1 U22555 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20363), .ZN(n20360) );
  OAI21_X1 U22556 ( .B1(n20361), .B2(n20366), .A(n20360), .ZN(P3_U2796) );
  AOI22_X1 U22557 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20363), .ZN(n20362) );
  OAI21_X1 U22558 ( .B1(n20947), .B2(n20366), .A(n20362), .ZN(P3_U2797) );
  AOI22_X1 U22559 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20364), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20363), .ZN(n20365) );
  OAI21_X1 U22560 ( .B1(n20367), .B2(n20366), .A(n20365), .ZN(P3_U2798) );
  NAND2_X1 U22561 ( .A1(n20368), .A2(n20379), .ZN(n20981) );
  INV_X1 U22562 ( .A(n20981), .ZN(n20985) );
  NAND2_X1 U22563 ( .A1(n20370), .A2(n20369), .ZN(n20771) );
  INV_X1 U22564 ( .A(n20771), .ZN(n20397) );
  AOI22_X1 U22565 ( .A1(n20727), .A2(n20371), .B1(n20985), .B2(n20397), .ZN(
        n20377) );
  INV_X1 U22566 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20536) );
  NAND2_X1 U22567 ( .A1(n20741), .A2(n20580), .ZN(n20755) );
  OAI21_X1 U22568 ( .B1(n20536), .B2(n20755), .A(n20762), .ZN(n20375) );
  AOI21_X1 U22569 ( .B1(n20580), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21422), .ZN(n20438) );
  OAI22_X1 U22570 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20492), .B1(n20765), 
        .B2(n20372), .ZN(n20373) );
  AOI221_X1 U22571 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20375), .C1(
        n20374), .C2(n20438), .A(n20373), .ZN(n20376) );
  OAI211_X1 U22572 ( .C1(n20385), .C2(n20768), .A(n20377), .B(n20376), .ZN(
        P3_U2670) );
  OAI22_X1 U22573 ( .A1(n20378), .A2(n20762), .B1(n20765), .B2(n20388), .ZN(
        n20382) );
  INV_X1 U22574 ( .A(n20379), .ZN(n21006) );
  NOR2_X1 U22575 ( .A1(n21006), .A2(n21394), .ZN(n21000) );
  NOR2_X1 U22576 ( .A1(n20380), .A2(n21000), .ZN(n20994) );
  NOR2_X1 U22577 ( .A1(n21422), .A2(n20580), .ZN(n20504) );
  INV_X1 U22578 ( .A(n20504), .ZN(n20544) );
  OAI22_X1 U22579 ( .A1(n20994), .A2(n20771), .B1(n20544), .B2(n20383), .ZN(
        n20381) );
  AOI211_X1 U22580 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n20430), .A(n20382), .B(
        n20381), .ZN(n20393) );
  AOI21_X1 U22581 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20384), .A(
        n20523), .ZN(n20395) );
  OAI211_X1 U22582 ( .C1(n20384), .C2(n20383), .A(n20741), .B(n20395), .ZN(
        n20392) );
  NOR2_X1 U22583 ( .A1(n20386), .A2(n20385), .ZN(n20398) );
  INV_X1 U22584 ( .A(n20398), .ZN(n20387) );
  OAI211_X1 U22585 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20456), .B(n20387), .ZN(n20391) );
  OAI211_X1 U22586 ( .C1(n20389), .C2(n20388), .A(n20727), .B(n20396), .ZN(
        n20390) );
  NAND4_X1 U22587 ( .A1(n20393), .A2(n20392), .A3(n20391), .A4(n20390), .ZN(
        P3_U2669) );
  XNOR2_X1 U22588 ( .A(n20395), .B(n20394), .ZN(n20405) );
  AOI211_X1 U22589 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n20396), .A(n20421), .B(
        n20764), .ZN(n20403) );
  AOI21_X1 U22590 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21013), .A(
        n21029), .ZN(n21015) );
  OR2_X1 U22591 ( .A1(n21015), .A2(n11661), .ZN(n21025) );
  AOI22_X1 U22592 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n20430), .B1(n20397), 
        .B2(n21025), .ZN(n20400) );
  OAI211_X1 U22593 ( .C1(P3_REIP_REG_3__SCAN_IN), .C2(n20398), .A(n20456), .B(
        n20407), .ZN(n20399) );
  OAI211_X1 U22594 ( .C1(n20762), .C2(n20401), .A(n20400), .B(n20399), .ZN(
        n20402) );
  AOI211_X1 U22595 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n20749), .A(n20403), .B(
        n20402), .ZN(n20404) );
  OAI21_X1 U22596 ( .B1(n20405), .B2(n21422), .A(n20404), .ZN(P3_U2668) );
  OAI21_X1 U22597 ( .B1(n20406), .B2(n20521), .A(n20580), .ZN(n20425) );
  NOR3_X1 U22598 ( .A1(n20412), .A2(n21422), .A3(n20425), .ZN(n20419) );
  AOI211_X1 U22599 ( .C1(n20408), .C2(n20407), .A(n20432), .B(n20492), .ZN(
        n20418) );
  AOI21_X1 U22600 ( .B1(n20409), .B2(n21413), .A(n20771), .ZN(n20417) );
  NOR2_X1 U22601 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21422), .ZN(
        n20410) );
  AOI21_X1 U22602 ( .B1(n20411), .B2(n20410), .A(n20504), .ZN(n20415) );
  INV_X1 U22603 ( .A(n20412), .ZN(n20414) );
  AOI22_X1 U22604 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20430), .B1(n20749), 
        .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n20413) );
  OAI211_X1 U22605 ( .C1(n20415), .C2(n20414), .A(n20413), .B(n21329), .ZN(
        n20416) );
  NOR4_X1 U22606 ( .A1(n20419), .A2(n20418), .A3(n20417), .A4(n20416), .ZN(
        n20423) );
  OAI211_X1 U22607 ( .C1(n20421), .C2(n20420), .A(n20727), .B(n20427), .ZN(
        n20422) );
  OAI211_X1 U22608 ( .C1(n20762), .C2(n20424), .A(n20423), .B(n20422), .ZN(
        P3_U2667) );
  XNOR2_X1 U22609 ( .A(n20426), .B(n20425), .ZN(n20437) );
  AOI211_X1 U22610 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n20427), .A(n20447), .B(
        n20764), .ZN(n20428) );
  AOI21_X1 U22611 ( .B1(n20718), .B2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20428), .ZN(n20436) );
  INV_X1 U22612 ( .A(n20429), .ZN(n20445) );
  NOR2_X1 U22613 ( .A1(n20492), .A2(n20445), .ZN(n20431) );
  NOR2_X1 U22614 ( .A1(n20430), .A2(n20431), .ZN(n20442) );
  INV_X1 U22615 ( .A(n20442), .ZN(n20460) );
  AOI22_X1 U22616 ( .A1(n20432), .A2(n20431), .B1(n20749), .B2(
        P3_EBX_REG_5__SCAN_IN), .ZN(n20433) );
  INV_X1 U22617 ( .A(n20433), .ZN(n20434) );
  AOI211_X1 U22618 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n20460), .A(n10995), .B(
        n20434), .ZN(n20435) );
  OAI211_X1 U22619 ( .C1(n21422), .C2(n20437), .A(n20436), .B(n20435), .ZN(
        P3_U2666) );
  AOI22_X1 U22620 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n20450) );
  NOR2_X1 U22621 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20492), .ZN(n20461) );
  OAI21_X1 U22622 ( .B1(n20482), .B2(n20521), .A(n20580), .ZN(n20451) );
  NOR3_X1 U22623 ( .A1(n20439), .A2(n21422), .A3(n20451), .ZN(n20444) );
  INV_X1 U22624 ( .A(n20438), .ZN(n20543) );
  OAI21_X1 U22625 ( .B1(n20504), .B2(n20440), .A(n20439), .ZN(n20441) );
  OAI22_X1 U22626 ( .A1(n20442), .A2(n21102), .B1(n20543), .B2(n20441), .ZN(
        n20443) );
  AOI211_X1 U22627 ( .C1(n20461), .C2(n20445), .A(n20444), .B(n20443), .ZN(
        n20449) );
  OAI211_X1 U22628 ( .C1(n20447), .C2(n20446), .A(n20727), .B(n20453), .ZN(
        n20448) );
  NAND4_X1 U22629 ( .A1(n20450), .A2(n20449), .A3(n21329), .A4(n20448), .ZN(
        P3_U2665) );
  XNOR2_X1 U22630 ( .A(n20452), .B(n20451), .ZN(n20464) );
  AOI211_X1 U22631 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n20453), .A(n20468), .B(
        n20764), .ZN(n20454) );
  AOI211_X1 U22632 ( .C1(n20749), .C2(P3_EBX_REG_7__SCAN_IN), .A(n10995), .B(
        n20454), .ZN(n20463) );
  NAND2_X1 U22633 ( .A1(n20456), .A2(n20455), .ZN(n20458) );
  OAI22_X1 U22634 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20458), .B1(n20762), 
        .B2(n20457), .ZN(n20459) );
  AOI221_X1 U22635 ( .B1(n20461), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n20460), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n20459), .ZN(n20462) );
  OAI211_X1 U22636 ( .C1(n21422), .C2(n20464), .A(n20463), .B(n20462), .ZN(
        P3_U2664) );
  NOR2_X1 U22637 ( .A1(n20482), .A2(n20521), .ZN(n20465) );
  AOI21_X1 U22638 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20465), .A(
        n20523), .ZN(n20466) );
  XNOR2_X1 U22639 ( .A(n20467), .B(n20466), .ZN(n20476) );
  AND2_X1 U22640 ( .A1(n20477), .A2(n20727), .ZN(n20480) );
  OAI21_X1 U22641 ( .B1(n20470), .B2(n20468), .A(n20480), .ZN(n20469) );
  OAI21_X1 U22642 ( .B1(n20470), .B2(n20765), .A(n20469), .ZN(n20471) );
  AOI211_X1 U22643 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n20718), .A(
        n10995), .B(n20471), .ZN(n20475) );
  NOR2_X1 U22644 ( .A1(n20492), .A2(n20483), .ZN(n20473) );
  OAI21_X1 U22645 ( .B1(n20472), .B2(n20492), .A(n20768), .ZN(n20499) );
  OAI21_X1 U22646 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n20473), .A(n20499), .ZN(
        n20474) );
  OAI211_X1 U22647 ( .C1(n20476), .C2(n21422), .A(n20475), .B(n20474), .ZN(
        P3_U2663) );
  OAI21_X1 U22648 ( .B1(n20764), .B2(n20477), .A(n20765), .ZN(n20478) );
  AOI22_X1 U22649 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20499), .B1(
        P3_EBX_REG_9__SCAN_IN), .B2(n20478), .ZN(n20490) );
  INV_X1 U22650 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20479) );
  AOI22_X1 U22651 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20718), .B1(
        n20480), .B2(n20479), .ZN(n20489) );
  NOR3_X1 U22652 ( .A1(n20482), .A2(n20481), .A3(n20521), .ZN(n20501) );
  NOR2_X1 U22653 ( .A1(n20501), .A2(n20755), .ZN(n20487) );
  NOR4_X1 U22654 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20492), .A3(n20484), .A4(
        n20483), .ZN(n20500) );
  AOI211_X1 U22655 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n20544), .A(
        n20543), .B(n20486), .ZN(n20485) );
  AOI211_X1 U22656 ( .C1(n20487), .C2(n20486), .A(n20500), .B(n20485), .ZN(
        n20488) );
  NAND4_X1 U22657 ( .A1(n20490), .A2(n20489), .A3(n20488), .A4(n21329), .ZN(
        P3_U2662) );
  NOR3_X1 U22658 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20492), .A3(n20491), 
        .ZN(n20498) );
  OAI211_X1 U22659 ( .C1(n20494), .C2(n20493), .A(n20727), .B(n20509), .ZN(
        n20495) );
  OAI211_X1 U22660 ( .C1(n20496), .C2(n20762), .A(n21329), .B(n20495), .ZN(
        n20497) );
  AOI211_X1 U22661 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20749), .A(n20498), .B(
        n20497), .ZN(n20508) );
  OAI21_X1 U22662 ( .B1(n20500), .B2(n20499), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n20507) );
  OAI21_X1 U22663 ( .B1(n20522), .B2(n20521), .A(n20580), .ZN(n20510) );
  INV_X1 U22664 ( .A(n20510), .ZN(n20512) );
  INV_X1 U22665 ( .A(n20501), .ZN(n20502) );
  AOI21_X1 U22666 ( .B1(n20505), .B2(n20502), .A(n21422), .ZN(n20503) );
  OAI22_X1 U22667 ( .A1(n20505), .A2(n20512), .B1(n20504), .B2(n20503), .ZN(
        n20506) );
  NAND3_X1 U22668 ( .A1(n20508), .A2(n20507), .A3(n20506), .ZN(P3_U2661) );
  NAND2_X1 U22669 ( .A1(n20766), .A2(n20552), .ZN(n20520) );
  AOI211_X1 U22670 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n20509), .A(n20531), .B(
        n20764), .ZN(n20517) );
  INV_X1 U22671 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20515) );
  INV_X1 U22672 ( .A(n20511), .ZN(n20513) );
  OAI221_X1 U22673 ( .B1(n20513), .B2(n20512), .C1(n20511), .C2(n20510), .A(
        n20741), .ZN(n20514) );
  OAI211_X1 U22674 ( .C1(n20765), .C2(n20515), .A(n21329), .B(n20514), .ZN(
        n20516) );
  AOI211_X1 U22675 ( .C1(n20718), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20517), .B(n20516), .ZN(n20518) );
  OAI221_X1 U22676 ( .B1(n20520), .B2(n21146), .C1(n20520), .C2(n20519), .A(
        n20518), .ZN(P3_U2660) );
  AOI22_X1 U22677 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n20534) );
  INV_X1 U22678 ( .A(n20520), .ZN(n20547) );
  NOR2_X1 U22679 ( .A1(n20522), .A2(n20521), .ZN(n20524) );
  AOI21_X1 U22680 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n20524), .A(
        n20523), .ZN(n20526) );
  OAI21_X1 U22681 ( .B1(n20527), .B2(n20526), .A(n20741), .ZN(n20525) );
  AOI21_X1 U22682 ( .B1(n20527), .B2(n20526), .A(n20525), .ZN(n20528) );
  AOI221_X1 U22683 ( .B1(n20547), .B2(P3_REIP_REG_12__SCAN_IN), .C1(n20576), 
        .C2(n20529), .A(n20528), .ZN(n20533) );
  OAI211_X1 U22684 ( .C1(n20531), .C2(n20530), .A(n20727), .B(n20539), .ZN(
        n20532) );
  NAND4_X1 U22685 ( .A1(n20534), .A2(n20533), .A3(n21329), .A4(n20532), .ZN(
        P3_U2659) );
  INV_X1 U22686 ( .A(n20542), .ZN(n20535) );
  AOI211_X1 U22687 ( .C1(n20537), .C2(n20536), .A(n20535), .B(n20755), .ZN(
        n20538) );
  AOI211_X1 U22688 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n20718), .A(
        n10995), .B(n20538), .ZN(n20551) );
  AOI211_X1 U22689 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n20539), .A(n20563), .B(
        n20764), .ZN(n20540) );
  AOI21_X1 U22690 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n20749), .A(n20540), .ZN(
        n20550) );
  INV_X1 U22691 ( .A(n20541), .ZN(n20545) );
  AOI211_X1 U22692 ( .C1(n20545), .C2(n20544), .A(n20543), .B(n20542), .ZN(
        n20546) );
  AOI21_X1 U22693 ( .B1(n20547), .B2(P3_REIP_REG_13__SCAN_IN), .A(n20546), 
        .ZN(n20549) );
  OAI211_X1 U22694 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(P3_REIP_REG_12__SCAN_IN), .A(n20576), .B(n20554), .ZN(n20548) );
  NAND4_X1 U22695 ( .A1(n20551), .A2(n20550), .A3(n20549), .A4(n20548), .ZN(
        P3_U2658) );
  INV_X1 U22696 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20566) );
  INV_X1 U22697 ( .A(n20577), .ZN(n20553) );
  OAI21_X1 U22698 ( .B1(n20553), .B2(n20552), .A(n20766), .ZN(n20585) );
  INV_X1 U22699 ( .A(n20554), .ZN(n20555) );
  AOI21_X1 U22700 ( .B1(n20555), .B2(n20576), .A(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n20560) );
  OAI21_X1 U22701 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20556), .A(
        n20580), .ZN(n20557) );
  XNOR2_X1 U22702 ( .A(n20558), .B(n20557), .ZN(n20559) );
  OAI22_X1 U22703 ( .A1(n20585), .A2(n20560), .B1(n21422), .B2(n20559), .ZN(
        n20561) );
  AOI211_X1 U22704 ( .C1(n20749), .C2(P3_EBX_REG_14__SCAN_IN), .A(n10995), .B(
        n20561), .ZN(n20565) );
  OAI211_X1 U22705 ( .C1(n20563), .C2(n20562), .A(n20727), .B(n20571), .ZN(
        n20564) );
  OAI211_X1 U22706 ( .C1(n20762), .C2(n20566), .A(n20565), .B(n20564), .ZN(
        P3_U2657) );
  OAI21_X1 U22707 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20567), .A(
        n20580), .ZN(n20569) );
  OAI21_X1 U22708 ( .B1(n20570), .B2(n20569), .A(n20741), .ZN(n20568) );
  AOI21_X1 U22709 ( .B1(n20570), .B2(n20569), .A(n20568), .ZN(n20575) );
  AOI211_X1 U22710 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n20571), .A(n20593), .B(
        n20764), .ZN(n20574) );
  AOI22_X1 U22711 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n20572) );
  INV_X1 U22712 ( .A(n20572), .ZN(n20573) );
  NOR4_X1 U22713 ( .A1(n10995), .A2(n20575), .A3(n20574), .A4(n20573), .ZN(
        n20578) );
  NAND3_X1 U22714 ( .A1(n20577), .A2(n20576), .A3(n20579), .ZN(n20584) );
  OAI211_X1 U22715 ( .C1(n20585), .C2(n20579), .A(n20578), .B(n20584), .ZN(
        P3_U2656) );
  AOI22_X1 U22716 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n20596) );
  OAI21_X1 U22717 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20581), .A(
        n20580), .ZN(n20582) );
  XNOR2_X1 U22718 ( .A(n20583), .B(n20582), .ZN(n20590) );
  AOI21_X1 U22719 ( .B1(n20585), .B2(n20584), .A(n21342), .ZN(n20589) );
  NOR3_X1 U22720 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20587), .A3(n20586), 
        .ZN(n20588) );
  AOI211_X1 U22721 ( .C1(n20590), .C2(n20741), .A(n20589), .B(n20588), .ZN(
        n20595) );
  OAI211_X1 U22722 ( .C1(n20593), .C2(n20592), .A(n20727), .B(n20591), .ZN(
        n20594) );
  NAND4_X1 U22723 ( .A1(n20596), .A2(n20595), .A3(n21329), .A4(n20594), .ZN(
        P3_U2655) );
  NOR2_X1 U22724 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n20623), .ZN(n20613) );
  OAI211_X1 U22725 ( .C1(n20597), .C2(n20599), .A(n20727), .B(n20607), .ZN(
        n20598) );
  OAI211_X1 U22726 ( .C1(n20765), .C2(n20599), .A(n21329), .B(n20598), .ZN(
        n20600) );
  AOI211_X1 U22727 ( .C1(n20718), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20613), .B(n20600), .ZN(n20605) );
  OAI211_X1 U22728 ( .C1(n20603), .C2(n20602), .A(n20741), .B(n20601), .ZN(
        n20604) );
  OAI211_X1 U22729 ( .C1(n20606), .C2(n21326), .A(n20605), .B(n20604), .ZN(
        P3_U2653) );
  NOR3_X1 U22730 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n21326), .A3(n20623), 
        .ZN(n20612) );
  AOI211_X1 U22731 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n20607), .A(n20629), .B(
        n20764), .ZN(n20611) );
  OAI22_X1 U22732 ( .A1(n20609), .A2(n20762), .B1(n20765), .B2(n20608), .ZN(
        n20610) );
  NOR4_X1 U22733 ( .A1(n10995), .A2(n20612), .A3(n20611), .A4(n20610), .ZN(
        n20620) );
  OAI21_X1 U22734 ( .B1(n20614), .B2(n20613), .A(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n20619) );
  OAI211_X1 U22735 ( .C1(n20617), .C2(n20616), .A(n20741), .B(n20615), .ZN(
        n20618) );
  NAND3_X1 U22736 ( .A1(n20620), .A2(n20619), .A3(n20618), .ZN(P3_U2652) );
  AOI22_X1 U22737 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n20633) );
  AND2_X1 U22738 ( .A1(n20766), .A2(n20621), .ZN(n20648) );
  NOR4_X1 U22739 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20623), .A3(n21326), 
        .A4(n20622), .ZN(n20624) );
  AOI21_X1 U22740 ( .B1(n20648), .B2(P3_REIP_REG_20__SCAN_IN), .A(n20624), 
        .ZN(n20632) );
  OAI211_X1 U22741 ( .C1(n20627), .C2(n20626), .A(n20741), .B(n20625), .ZN(
        n20631) );
  OAI211_X1 U22742 ( .C1(n20629), .C2(n20628), .A(n20727), .B(n20634), .ZN(
        n20630) );
  NAND4_X1 U22743 ( .A1(n20633), .A2(n20632), .A3(n20631), .A4(n20630), .ZN(
        P3_U2651) );
  INV_X1 U22744 ( .A(n20658), .ZN(n20644) );
  AOI211_X1 U22745 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n20634), .A(n20653), .B(
        n20764), .ZN(n20638) );
  OAI22_X1 U22746 ( .A1(n20636), .A2(n20762), .B1(n20765), .B2(n20635), .ZN(
        n20637) );
  AOI211_X1 U22747 ( .C1(n20648), .C2(P3_REIP_REG_21__SCAN_IN), .A(n20638), 
        .B(n20637), .ZN(n20643) );
  OAI211_X1 U22748 ( .C1(n20641), .C2(n20640), .A(n20741), .B(n20639), .ZN(
        n20642) );
  OAI211_X1 U22749 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n20644), .A(n20643), 
        .B(n20642), .ZN(P3_U2650) );
  AOI22_X1 U22750 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n20657) );
  AOI22_X1 U22751 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .B1(n20646), .B2(n20645), .ZN(n20647) );
  AOI22_X1 U22752 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20648), .B1(n20658), 
        .B2(n20647), .ZN(n20656) );
  OAI211_X1 U22753 ( .C1(n20651), .C2(n20650), .A(n20741), .B(n20649), .ZN(
        n20655) );
  OAI211_X1 U22754 ( .C1(n20653), .C2(n20652), .A(n20727), .B(n20660), .ZN(
        n20654) );
  NAND4_X1 U22755 ( .A1(n20657), .A2(n20656), .A3(n20655), .A4(n20654), .ZN(
        P3_U2649) );
  NAND3_X1 U22756 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n20658), .ZN(n20669) );
  NOR2_X1 U22757 ( .A1(n20719), .A2(n20659), .ZN(n20673) );
  AOI211_X1 U22758 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n20660), .A(n20678), .B(
        n20764), .ZN(n20663) );
  AOI22_X1 U22759 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n20661) );
  INV_X1 U22760 ( .A(n20661), .ZN(n20662) );
  AOI211_X1 U22761 ( .C1(n20673), .C2(P3_REIP_REG_23__SCAN_IN), .A(n20663), 
        .B(n20662), .ZN(n20668) );
  OAI211_X1 U22762 ( .C1(n20666), .C2(n20665), .A(n20741), .B(n20664), .ZN(
        n20667) );
  OAI211_X1 U22763 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n20669), .A(n20668), 
        .B(n20667), .ZN(P3_U2648) );
  AOI22_X1 U22764 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n20682) );
  INV_X1 U22765 ( .A(n20670), .ZN(n20672) );
  AOI22_X1 U22766 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20673), .B1(n20672), 
        .B2(n20671), .ZN(n20681) );
  OAI211_X1 U22767 ( .C1(n20676), .C2(n20675), .A(n20741), .B(n20674), .ZN(
        n20680) );
  OAI211_X1 U22768 ( .C1(n20678), .C2(n20677), .A(n20727), .B(n20684), .ZN(
        n20679) );
  NAND4_X1 U22769 ( .A1(n20682), .A2(n20681), .A3(n20680), .A4(n20679), .ZN(
        P3_U2647) );
  NAND2_X1 U22770 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20683), .ZN(n20695) );
  AOI211_X1 U22771 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n20684), .A(n20702), .B(
        n20764), .ZN(n20688) );
  OAI22_X1 U22772 ( .A1(n20686), .A2(n20762), .B1(n20765), .B2(n20685), .ZN(
        n20687) );
  AOI211_X1 U22773 ( .C1(n20697), .C2(n20689), .A(n20688), .B(n20687), .ZN(
        n20694) );
  OAI211_X1 U22774 ( .C1(n20692), .C2(n20691), .A(n20741), .B(n20690), .ZN(
        n20693) );
  OAI211_X1 U22775 ( .C1(n20719), .C2(n20695), .A(n20694), .B(n20693), .ZN(
        P3_U2646) );
  AOI22_X1 U22776 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n20706) );
  NOR2_X1 U22777 ( .A1(n20719), .A2(n20696), .ZN(n20711) );
  OAI221_X1 U22778 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(P3_REIP_REG_25__SCAN_IN), .C1(P3_REIP_REG_26__SCAN_IN), .C2(n20697), .A(n20711), .ZN(n20705) );
  OAI211_X1 U22779 ( .C1(n20700), .C2(n20699), .A(n20741), .B(n20698), .ZN(
        n20704) );
  OAI211_X1 U22780 ( .C1(n20702), .C2(n20701), .A(n20727), .B(n20707), .ZN(
        n20703) );
  NAND4_X1 U22781 ( .A1(n20706), .A2(n20705), .A3(n20704), .A4(n20703), .ZN(
        P3_U2645) );
  AOI211_X1 U22782 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n20707), .A(n20729), .B(
        n20764), .ZN(n20710) );
  OAI22_X1 U22783 ( .A1(n11261), .A2(n20762), .B1(n20765), .B2(n20708), .ZN(
        n20709) );
  AOI211_X1 U22784 ( .C1(n20711), .C2(P3_REIP_REG_27__SCAN_IN), .A(n20710), 
        .B(n20709), .ZN(n20716) );
  OAI211_X1 U22785 ( .C1(n20714), .C2(n20713), .A(n20741), .B(n20712), .ZN(
        n20715) );
  OAI211_X1 U22786 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n20717), .A(n20716), 
        .B(n20715), .ZN(P3_U2644) );
  AOI22_X1 U22787 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20718), .B1(
        n20749), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n20733) );
  NOR2_X1 U22788 ( .A1(n20719), .A2(n20720), .ZN(n20723) );
  AOI22_X1 U22789 ( .A1(n20723), .A2(n20722), .B1(n20721), .B2(n20720), .ZN(
        n20732) );
  OAI211_X1 U22790 ( .C1(n20726), .C2(n20725), .A(n20741), .B(n20724), .ZN(
        n20731) );
  OAI211_X1 U22791 ( .C1(n20729), .C2(n20728), .A(n20727), .B(n20736), .ZN(
        n20730) );
  NAND4_X1 U22792 ( .A1(n20733), .A2(n20732), .A3(n20731), .A4(n20730), .ZN(
        P3_U2643) );
  INV_X1 U22793 ( .A(n20734), .ZN(n20735) );
  AOI21_X1 U22794 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n20736), .A(n20735), .ZN(
        n20740) );
  OAI22_X1 U22795 ( .A1(n20738), .A2(n20762), .B1(n20765), .B2(n20737), .ZN(
        n20739) );
  AOI211_X1 U22796 ( .C1(n20751), .C2(P3_REIP_REG_29__SCAN_IN), .A(n20740), 
        .B(n20739), .ZN(n20745) );
  OAI211_X1 U22797 ( .C1(n20743), .C2(n20742), .A(n20741), .B(n20756), .ZN(
        n20744) );
  OAI211_X1 U22798 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n20746), .A(n20745), 
        .B(n20744), .ZN(P3_U2642) );
  AOI22_X1 U22799 ( .A1(n20749), .A2(P3_EBX_REG_31__SCAN_IN), .B1(n20748), 
        .B2(n20747), .ZN(n20761) );
  NOR2_X1 U22800 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20750), .ZN(n20759) );
  INV_X1 U22801 ( .A(n20751), .ZN(n20753) );
  AOI21_X1 U22802 ( .B1(n20754), .B2(n20753), .A(n20752), .ZN(n20758) );
  NAND2_X1 U22803 ( .A1(n20765), .A2(n20764), .ZN(n20767) );
  AOI22_X1 U22804 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n20767), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n20766), .ZN(n20770) );
  NAND3_X1 U22805 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20768), .A3(
        n20996), .ZN(n20769) );
  OAI211_X1 U22806 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20771), .A(
        n20770), .B(n20769), .ZN(P3_U2671) );
  NAND2_X1 U22807 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n20785) );
  NOR2_X1 U22808 ( .A1(n20824), .A2(n20772), .ZN(n20810) );
  NOR4_X1 U22809 ( .A1(n20775), .A2(n20774), .A3(n20773), .A4(n20811), .ZN(
        n20776) );
  NAND4_X1 U22810 ( .A1(n20810), .A2(P3_EAX_REG_0__SCAN_IN), .A3(
        P3_EAX_REG_1__SCAN_IN), .A4(n20776), .ZN(n20958) );
  NOR2_X1 U22811 ( .A1(n20809), .A2(n20966), .ZN(n20790) );
  INV_X1 U22812 ( .A(n20790), .ZN(n20975) );
  INV_X1 U22813 ( .A(n20807), .ZN(n20801) );
  NAND2_X1 U22814 ( .A1(n20809), .A2(n20843), .ZN(n20968) );
  AOI22_X1 U22815 ( .A1(n20798), .A2(P3_EAX_REG_12__SCAN_IN), .B1(
        P3_EAX_REG_13__SCAN_IN), .B2(n20968), .ZN(n20791) );
  NAND4_X1 U22816 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_13__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n20784)
         );
  NOR3_X1 U22817 ( .A1(n20958), .A2(n20785), .A3(n20784), .ZN(n20844) );
  NAND2_X1 U22818 ( .A1(n20786), .A2(n20843), .ZN(n20839) );
  NOR2_X2 U22819 ( .A1(n20787), .A2(n20966), .ZN(n20972) );
  AOI22_X1 U22820 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20973), .B1(n20972), .B2(
        n20788), .ZN(n20789) );
  OAI221_X1 U22821 ( .B1(n20791), .B2(n20844), .C1(n20791), .C2(n20790), .A(
        n20789), .ZN(P3_U2722) );
  INV_X1 U22822 ( .A(n20798), .ZN(n20795) );
  NAND2_X1 U22823 ( .A1(n20795), .A2(P3_EAX_REG_12__SCAN_IN), .ZN(n20794) );
  AOI22_X1 U22824 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20973), .B1(n20972), .B2(
        n20792), .ZN(n20793) );
  OAI221_X1 U22825 ( .B1(n20795), .B2(P3_EAX_REG_12__SCAN_IN), .C1(n20794), 
        .C2(n20946), .A(n20793), .ZN(P3_U2723) );
  INV_X1 U22826 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n20799) );
  AOI22_X1 U22827 ( .A1(n20807), .A2(P3_EAX_REG_10__SCAN_IN), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n20968), .ZN(n20797) );
  OAI222_X1 U22828 ( .A1(n20839), .A2(n20799), .B1(n20798), .B2(n20797), .C1(
        n20956), .C2(n20796), .ZN(P3_U2724) );
  AOI22_X1 U22829 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20973), .B1(n20972), .B2(
        n20800), .ZN(n20804) );
  OAI221_X1 U22830 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n20807), .C1(n20802), 
        .C2(n20801), .A(n20968), .ZN(n20803) );
  NAND2_X1 U22831 ( .A1(n20804), .A2(n20803), .ZN(P3_U2725) );
  INV_X1 U22832 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n20808) );
  AOI22_X1 U22833 ( .A1(n20814), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n20968), .ZN(n20806) );
  OAI222_X1 U22834 ( .A1(n20839), .A2(n20808), .B1(n20807), .B2(n20806), .C1(
        n20956), .C2(n20805), .ZN(P3_U2726) );
  NAND3_X1 U22835 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(n20843), .ZN(n20967) );
  NOR2_X1 U22836 ( .A1(n20809), .A2(n20967), .ZN(n20834) );
  NAND2_X1 U22837 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n20838), .ZN(n20823) );
  NAND2_X1 U22838 ( .A1(n20810), .A2(n20832), .ZN(n20815) );
  NOR2_X1 U22839 ( .A1(n20811), .A2(n20815), .ZN(n20819) );
  AOI21_X1 U22840 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n20968), .A(n20819), .ZN(
        n20813) );
  OAI222_X1 U22841 ( .A1(n20934), .A2(n20839), .B1(n20814), .B2(n20813), .C1(
        n20956), .C2(n20812), .ZN(P3_U2728) );
  INV_X1 U22842 ( .A(n20815), .ZN(n20822) );
  AOI21_X1 U22843 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20968), .A(n20822), .ZN(
        n20818) );
  INV_X1 U22844 ( .A(n20816), .ZN(n20817) );
  OAI222_X1 U22845 ( .A1(n20865), .A2(n20839), .B1(n20819), .B2(n20818), .C1(
        n20956), .C2(n20817), .ZN(P3_U2729) );
  AOI22_X1 U22846 ( .A1(n20832), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n20968), .ZN(n20821) );
  OAI222_X1 U22847 ( .A1(n20848), .A2(n20839), .B1(n20822), .B2(n20821), .C1(
        n20956), .C2(n20820), .ZN(P3_U2730) );
  NOR2_X1 U22848 ( .A1(n20824), .A2(n20823), .ZN(n20828) );
  AOI21_X1 U22849 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20968), .A(n20832), .ZN(
        n20827) );
  INV_X1 U22850 ( .A(n20825), .ZN(n20826) );
  OAI222_X1 U22851 ( .A1(n20829), .A2(n20839), .B1(n20828), .B2(n20827), .C1(
        n20956), .C2(n20826), .ZN(P3_U2731) );
  AOI21_X1 U22852 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20968), .A(n20838), .ZN(
        n20831) );
  OAI222_X1 U22853 ( .A1(n20833), .A2(n20839), .B1(n20832), .B2(n20831), .C1(
        n20956), .C2(n20830), .ZN(P3_U2732) );
  AOI21_X1 U22854 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n20968), .A(n20834), .ZN(
        n20837) );
  INV_X1 U22855 ( .A(n20835), .ZN(n20836) );
  OAI222_X1 U22856 ( .A1(n20876), .A2(n20839), .B1(n20838), .B2(n20837), .C1(
        n20956), .C2(n20836), .ZN(P3_U2733) );
  NAND2_X1 U22857 ( .A1(n20840), .A2(n20946), .ZN(n20933) );
  AOI22_X1 U22858 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n20938), .B1(n20972), .B2(
        n20842), .ZN(n20847) );
  NAND2_X1 U22859 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .ZN(n20845) );
  NAND2_X1 U22860 ( .A1(n20844), .A2(n20843), .ZN(n20948) );
  NAND2_X1 U22861 ( .A1(n20959), .A2(n20940), .ZN(n20877) );
  INV_X1 U22862 ( .A(n20867), .ZN(n20872) );
  NOR2_X1 U22863 ( .A1(n20845), .A2(n20872), .ZN(n20852) );
  NOR2_X1 U22864 ( .A1(n20946), .A2(n20852), .ZN(n20857) );
  AND2_X1 U22865 ( .A1(n20858), .A2(n20852), .ZN(n20856) );
  AOI21_X1 U22866 ( .B1(n20857), .B2(P3_EAX_REG_21__SCAN_IN), .A(n20856), .ZN(
        n20846) );
  OAI211_X1 U22867 ( .C1(n20848), .C2(n20933), .A(n20847), .B(n20846), .ZN(
        P3_U2714) );
  NAND2_X1 U22868 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n20867), .ZN(n20866) );
  AOI22_X1 U22869 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20939), .B1(n20972), .B2(
        n20849), .ZN(n20851) );
  AOI22_X1 U22870 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n20938), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n20857), .ZN(n20850) );
  OAI211_X1 U22871 ( .C1(n20852), .C2(n20866), .A(n20851), .B(n20850), .ZN(
        P3_U2715) );
  INV_X1 U22872 ( .A(n20938), .ZN(n20928) );
  OAI22_X1 U22873 ( .A1(n20854), .A2(n20956), .B1(n20853), .B2(n20928), .ZN(
        n20855) );
  AOI221_X1 U22874 ( .B1(n20857), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n20856), 
        .C2(P3_EAX_REG_22__SCAN_IN), .A(n20855), .ZN(n20864) );
  NOR4_X1 U22875 ( .A1(n20861), .A2(n20860), .A3(n20859), .A4(n20858), .ZN(
        n20884) );
  NAND3_X1 U22876 ( .A1(n20884), .A2(n20873), .A3(n20862), .ZN(n20863) );
  OAI211_X1 U22877 ( .C1(n20933), .C2(n20865), .A(n20864), .B(n20863), .ZN(
        P3_U2713) );
  AOI22_X1 U22878 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20939), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20938), .ZN(n20869) );
  OAI211_X1 U22879 ( .C1(n20867), .C2(P3_EAX_REG_19__SCAN_IN), .A(n20968), .B(
        n20866), .ZN(n20868) );
  OAI211_X1 U22880 ( .C1(n20870), .C2(n20956), .A(n20869), .B(n20868), .ZN(
        P3_U2716) );
  AOI22_X1 U22881 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n20938), .B1(n20972), .B2(
        n20871), .ZN(n20875) );
  OAI211_X1 U22882 ( .C1(n20873), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20968), .B(
        n20872), .ZN(n20874) );
  OAI211_X1 U22883 ( .C1(n20933), .C2(n20876), .A(n20875), .B(n20874), .ZN(
        P3_U2717) );
  AOI22_X1 U22884 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20939), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20938), .ZN(n20882) );
  OAI21_X1 U22885 ( .B1(n20878), .B2(n20946), .A(n20877), .ZN(n20880) );
  NAND2_X1 U22886 ( .A1(n20880), .A2(n20879), .ZN(n20881) );
  OAI211_X1 U22887 ( .C1(n20883), .C2(n20956), .A(n20882), .B(n20881), .ZN(
        P3_U2718) );
  AOI22_X1 U22888 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20939), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20938), .ZN(n20888) );
  NAND4_X1 U22889 ( .A1(n20940), .A2(n20884), .A3(P3_EAX_REG_17__SCAN_IN), 
        .A4(P3_EAX_REG_22__SCAN_IN), .ZN(n20931) );
  NAND2_X1 U22890 ( .A1(n20959), .A2(n20929), .ZN(n20921) );
  AOI211_X1 U22891 ( .C1(n20885), .C2(n20923), .A(n20891), .B(n20946), .ZN(
        n20886) );
  INV_X1 U22892 ( .A(n20886), .ZN(n20887) );
  OAI211_X1 U22893 ( .C1(n20889), .C2(n20956), .A(n20888), .B(n20887), .ZN(
        P3_U2710) );
  INV_X1 U22894 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n20894) );
  AOI22_X1 U22895 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n20938), .B1(n20972), .B2(
        n20890), .ZN(n20893) );
  OAI211_X1 U22896 ( .C1(n20891), .C2(P3_EAX_REG_26__SCAN_IN), .A(n20968), .B(
        n20914), .ZN(n20892) );
  OAI211_X1 U22897 ( .C1(n20933), .C2(n20894), .A(n20893), .B(n20892), .ZN(
        P3_U2709) );
  NAND2_X1 U22898 ( .A1(n20913), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n20910) );
  NAND2_X1 U22899 ( .A1(n20905), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n20904) );
  NOR2_X1 U22900 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n20904), .ZN(n20896) );
  NAND2_X1 U22901 ( .A1(n20968), .A2(n20904), .ZN(n20902) );
  OAI21_X1 U22902 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n20975), .A(n20902), .ZN(
        n20895) );
  AOI22_X1 U22903 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n20896), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n20895), .ZN(n20897) );
  OAI21_X1 U22904 ( .B1(n20898), .B2(n20928), .A(n20897), .ZN(P3_U2704) );
  OAI22_X1 U22905 ( .A1(n20899), .A2(n20956), .B1(n15699), .B2(n20928), .ZN(
        n20900) );
  AOI21_X1 U22906 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n20939), .A(n20900), .ZN(
        n20901) );
  OAI221_X1 U22907 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n20904), .C1(n20903), 
        .C2(n20902), .A(n20901), .ZN(P3_U2705) );
  AOI22_X1 U22908 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20939), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20938), .ZN(n20907) );
  OAI211_X1 U22909 ( .C1(n20905), .C2(P3_EAX_REG_29__SCAN_IN), .A(n20968), .B(
        n20904), .ZN(n20906) );
  OAI211_X1 U22910 ( .C1(n20908), .C2(n20956), .A(n20907), .B(n20906), .ZN(
        P3_U2706) );
  AOI22_X1 U22911 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20939), .B1(n20972), .B2(
        n20909), .ZN(n20912) );
  OAI211_X1 U22912 ( .C1(n20913), .C2(P3_EAX_REG_28__SCAN_IN), .A(n20968), .B(
        n20910), .ZN(n20911) );
  OAI211_X1 U22913 ( .C1(n20928), .C2(n16486), .A(n20912), .B(n20911), .ZN(
        P3_U2707) );
  AOI22_X1 U22914 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20939), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20938), .ZN(n20918) );
  AOI211_X1 U22915 ( .C1(n20915), .C2(n20914), .A(n20913), .B(n20946), .ZN(
        n20916) );
  INV_X1 U22916 ( .A(n20916), .ZN(n20917) );
  OAI211_X1 U22917 ( .C1(n20919), .C2(n20956), .A(n20918), .B(n20917), .ZN(
        P3_U2708) );
  INV_X1 U22918 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n20927) );
  AOI22_X1 U22919 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20939), .B1(n20972), .B2(
        n20920), .ZN(n20926) );
  OAI21_X1 U22920 ( .B1(n20922), .B2(n20946), .A(n20921), .ZN(n20924) );
  NAND2_X1 U22921 ( .A1(n20924), .A2(n20923), .ZN(n20925) );
  OAI211_X1 U22922 ( .C1(n20928), .C2(n20927), .A(n20926), .B(n20925), .ZN(
        P3_U2711) );
  AOI211_X1 U22923 ( .C1(n20931), .C2(n20930), .A(n20946), .B(n20929), .ZN(
        n20936) );
  OAI22_X1 U22924 ( .A1(n20934), .A2(n20933), .B1(n20956), .B2(n20932), .ZN(
        n20935) );
  AOI211_X1 U22925 ( .C1(n20938), .C2(BUF2_REG_23__SCAN_IN), .A(n20936), .B(
        n20935), .ZN(n20937) );
  INV_X1 U22926 ( .A(n20937), .ZN(P3_U2712) );
  AOI22_X1 U22927 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20939), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20938), .ZN(n20944) );
  AOI211_X1 U22928 ( .C1(n20952), .C2(n20941), .A(n20946), .B(n20940), .ZN(
        n20942) );
  INV_X1 U22929 ( .A(n20942), .ZN(n20943) );
  OAI211_X1 U22930 ( .C1(n20945), .C2(n20956), .A(n20944), .B(n20943), .ZN(
        P3_U2719) );
  AOI211_X1 U22931 ( .C1(n20948), .C2(n20947), .A(n20946), .B(n20953), .ZN(
        n20949) );
  AOI21_X1 U22932 ( .B1(n20973), .B2(BUF2_REG_14__SCAN_IN), .A(n20949), .ZN(
        n20950) );
  OAI21_X1 U22933 ( .B1(n20951), .B2(n20956), .A(n20950), .ZN(P3_U2721) );
  OAI211_X1 U22934 ( .C1(n20953), .C2(P3_EAX_REG_15__SCAN_IN), .A(n20968), .B(
        n20952), .ZN(n20955) );
  NAND2_X1 U22935 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20973), .ZN(n20954) );
  OAI211_X1 U22936 ( .C1(n20957), .C2(n20956), .A(n20955), .B(n20954), .ZN(
        P3_U2720) );
  AOI21_X1 U22937 ( .B1(n20959), .B2(n20958), .A(n20966), .ZN(n20962) );
  AOI22_X1 U22938 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20973), .B1(n20972), .B2(
        n20960), .ZN(n20961) );
  OAI221_X1 U22939 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n20964), .C1(n20963), 
        .C2(n20962), .A(n20961), .ZN(P3_U2727) );
  AOI22_X1 U22940 ( .A1(n20973), .A2(BUF2_REG_1__SCAN_IN), .B1(n20972), .B2(
        n20965), .ZN(n20970) );
  NOR2_X1 U22941 ( .A1(n20966), .A2(n20976), .ZN(n20977) );
  OAI211_X1 U22942 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n20977), .A(n20968), .B(
        n20967), .ZN(n20969) );
  NAND2_X1 U22943 ( .A1(n20970), .A2(n20969), .ZN(P3_U2734) );
  AOI22_X1 U22944 ( .A1(n20973), .A2(BUF2_REG_0__SCAN_IN), .B1(n20972), .B2(
        n20971), .ZN(n20974) );
  OAI221_X1 U22945 ( .B1(n20977), .B2(n20976), .C1(n20977), .C2(n20975), .A(
        n20974), .ZN(P3_U2735) );
  NOR2_X1 U22946 ( .A1(n21075), .A2(n20978), .ZN(n20980) );
  OAI22_X1 U22947 ( .A1(n21003), .A2(n21162), .B1(n20980), .B2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21389) );
  INV_X1 U22948 ( .A(n20996), .ZN(n21024) );
  AOI222_X1 U22949 ( .A1(n21137), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21389), 
        .B2(n21024), .C1(n21003), .C2(n21026), .ZN(n20979) );
  AOI22_X1 U22950 ( .A1(n21030), .A2(n21003), .B1(n20979), .B2(n21027), .ZN(
        P3_U3290) );
  AOI21_X1 U22951 ( .B1(n21075), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n21367), .ZN(n20990) );
  OAI22_X1 U22952 ( .A1(n20981), .A2(n20980), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20990), .ZN(n21390) );
  AOI22_X1 U22953 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20983), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n20982), .ZN(n20997) );
  NAND2_X1 U22954 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20998) );
  INV_X1 U22955 ( .A(n20998), .ZN(n20984) );
  AOI222_X1 U22956 ( .A1(n21390), .A2(n21024), .B1(n20985), .B2(n21026), .C1(
        n20997), .C2(n20984), .ZN(n20986) );
  AOI22_X1 U22957 ( .A1(n21030), .A2(n20991), .B1(n20986), .B2(n21027), .ZN(
        P3_U3289) );
  AOI22_X1 U22958 ( .A1(n20989), .A2(n11040), .B1(n20988), .B2(n20987), .ZN(
        n21017) );
  AOI211_X1 U22959 ( .C1(n21010), .C2(n21017), .A(n21006), .B(n21394), .ZN(
        n20993) );
  AOI211_X1 U22960 ( .C1(n21394), .C2(n20991), .A(n20990), .B(n21013), .ZN(
        n20992) );
  AOI211_X1 U22961 ( .C1(n21386), .C2(n20994), .A(n20993), .B(n20992), .ZN(
        n21395) );
  OAI222_X1 U22962 ( .A1(n20998), .A2(n20997), .B1(n20996), .B2(n21395), .C1(
        n20995), .C2(n21429), .ZN(n20999) );
  AOI22_X1 U22963 ( .A1(n21026), .A2(n21000), .B1(n21027), .B2(n20999), .ZN(
        n21001) );
  OAI21_X1 U22964 ( .B1(n21394), .B2(n21027), .A(n21001), .ZN(P3_U3288) );
  AOI21_X1 U22965 ( .B1(n21002), .B2(n21003), .A(n21012), .ZN(n21022) );
  NAND2_X1 U22966 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21003), .ZN(
        n21009) );
  OAI211_X1 U22967 ( .C1(n21006), .C2(n21005), .A(n21386), .B(n21004), .ZN(
        n21007) );
  OAI22_X1 U22968 ( .A1(n21010), .A2(n21009), .B1(n21008), .B2(n21007), .ZN(
        n21021) );
  OAI22_X1 U22969 ( .A1(n21029), .A2(n21013), .B1(n21012), .B2(n21011), .ZN(
        n21014) );
  INV_X1 U22970 ( .A(n21014), .ZN(n21018) );
  INV_X1 U22971 ( .A(n21015), .ZN(n21016) );
  OAI22_X1 U22972 ( .A1(n21019), .A2(n21018), .B1(n21017), .B2(n21016), .ZN(
        n21020) );
  NOR3_X1 U22973 ( .A1(n21022), .A2(n21021), .A3(n21020), .ZN(n21402) );
  INV_X1 U22974 ( .A(n21402), .ZN(n21023) );
  AOI22_X1 U22975 ( .A1(n21026), .A2(n21025), .B1(n21024), .B2(n21023), .ZN(
        n21028) );
  AOI22_X1 U22976 ( .A1(n21030), .A2(n21029), .B1(n21028), .B2(n21027), .ZN(
        P3_U3285) );
  NOR2_X1 U22977 ( .A1(n21031), .A2(n21263), .ZN(n21281) );
  AOI22_X1 U22978 ( .A1(n21373), .A2(n21033), .B1(n21032), .B2(n21281), .ZN(
        n21046) );
  NOR2_X1 U22979 ( .A1(n21386), .A2(n21367), .ZN(n21356) );
  NAND2_X1 U22980 ( .A1(n21035), .A2(n21034), .ZN(n21036) );
  AOI22_X1 U22981 ( .A1(n21386), .A2(n21037), .B1(n21367), .B2(n21036), .ZN(
        n21296) );
  AOI22_X1 U22982 ( .A1(n21293), .A2(n21039), .B1(n21384), .B2(n21038), .ZN(
        n21040) );
  OAI211_X1 U22983 ( .C1(n21042), .C2(n21356), .A(n21296), .B(n21040), .ZN(
        n21198) );
  AOI21_X1 U22984 ( .B1(n21075), .B2(n21041), .A(n21263), .ZN(n21294) );
  OAI21_X1 U22985 ( .B1(n21363), .B2(n21042), .A(n21294), .ZN(n21043) );
  OAI211_X1 U22986 ( .C1(n21198), .C2(n21043), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n21329), .ZN(n21044) );
  NAND3_X1 U22987 ( .A1(n21046), .A2(n21045), .A3(n21044), .ZN(P3_U2841) );
  NOR2_X1 U22988 ( .A1(n21263), .A2(n21268), .ZN(n21172) );
  NOR2_X1 U22989 ( .A1(n21386), .A2(n21075), .ZN(n21303) );
  AOI221_X1 U22990 ( .B1(n21303), .B2(n21137), .C1(n21162), .C2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n21263), .ZN(n21047) );
  AOI221_X1 U22991 ( .B1(n21172), .B2(n21049), .C1(n21110), .C2(n21048), .A(
        n21047), .ZN(n21051) );
  NAND2_X1 U22992 ( .A1(n10995), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n21050) );
  OAI211_X1 U22993 ( .C1(n21275), .C2(n21137), .A(n21051), .B(n21050), .ZN(
        P3_U2862) );
  AOI22_X1 U22994 ( .A1(n10995), .A2(P3_REIP_REG_1__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21238), .ZN(n21058) );
  NOR2_X1 U22995 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21367), .ZN(
        n21052) );
  NOR2_X1 U22996 ( .A1(n21285), .A2(n21052), .ZN(n21054) );
  NOR2_X1 U22997 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21303), .ZN(
        n21053) );
  MUX2_X1 U22998 ( .A(n21054), .B(n21053), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n21056) );
  AOI22_X1 U22999 ( .A1(n21369), .A2(n21056), .B1(n21110), .B2(n21055), .ZN(
        n21057) );
  OAI211_X1 U23000 ( .C1(n21059), .C2(n21246), .A(n21058), .B(n21057), .ZN(
        P3_U2861) );
  INV_X1 U23001 ( .A(n21117), .ZN(n21060) );
  AOI211_X1 U23002 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n21060), .A(
        n21362), .B(n11701), .ZN(n21062) );
  NAND2_X1 U23003 ( .A1(n21072), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21074) );
  AOI21_X1 U23004 ( .B1(n21071), .B2(n21074), .A(n21312), .ZN(n21061) );
  AOI211_X1 U23005 ( .C1(n21063), .C2(n21084), .A(n21062), .B(n21061), .ZN(
        n21065) );
  AOI21_X1 U23006 ( .B1(n21162), .B2(n21137), .A(n21362), .ZN(n21070) );
  NAND3_X1 U23007 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21070), .A3(
        n11701), .ZN(n21064) );
  OAI211_X1 U23008 ( .C1(n21066), .C2(n21268), .A(n21065), .B(n21064), .ZN(
        n21068) );
  AOI21_X1 U23009 ( .B1(n21369), .B2(n21068), .A(n21067), .ZN(n21069) );
  OAI21_X1 U23010 ( .B1(n11701), .B2(n21275), .A(n21069), .ZN(P3_U2860) );
  AOI22_X1 U23011 ( .A1(n10995), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21238), .ZN(n21079) );
  AOI22_X1 U23012 ( .A1(n21072), .A2(n21070), .B1(n21386), .B2(n21071), .ZN(
        n21096) );
  OAI22_X1 U23013 ( .A1(n21162), .A2(n21072), .B1(n21071), .B2(n21312), .ZN(
        n21073) );
  AOI211_X1 U23014 ( .C1(n21075), .C2(n21074), .A(n11704), .B(n21073), .ZN(
        n21081) );
  AOI211_X1 U23015 ( .C1(n21096), .C2(n11704), .A(n21081), .B(n21263), .ZN(
        n21076) );
  AOI21_X1 U23016 ( .B1(n21077), .B2(n21110), .A(n21076), .ZN(n21078) );
  OAI211_X1 U23017 ( .C1(n21246), .C2(n21080), .A(n21079), .B(n21078), .ZN(
        P3_U2859) );
  NOR3_X1 U23018 ( .A1(n21285), .A2(n21081), .A3(n21095), .ZN(n21083) );
  NOR3_X1 U23019 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21096), .A3(
        n11704), .ZN(n21082) );
  AOI211_X1 U23020 ( .C1(n21085), .C2(n21084), .A(n21083), .B(n21082), .ZN(
        n21090) );
  OAI22_X1 U23021 ( .A1(n21095), .A2(n21275), .B1(n21246), .B2(n21086), .ZN(
        n21088) );
  NOR2_X1 U23022 ( .A1(n21088), .A2(n21087), .ZN(n21089) );
  OAI21_X1 U23023 ( .B1(n21090), .B2(n21263), .A(n21089), .ZN(P3_U2858) );
  INV_X1 U23024 ( .A(n21091), .ZN(n21092) );
  NOR2_X1 U23025 ( .A1(n21117), .A2(n21263), .ZN(n21318) );
  OAI21_X1 U23026 ( .B1(n21092), .B2(n21312), .A(n21318), .ZN(n21094) );
  OAI221_X1 U23027 ( .B1(n21094), .B2(n21093), .C1(n21094), .C2(n21321), .A(
        n21329), .ZN(n21101) );
  NOR3_X1 U23028 ( .A1(n21096), .A2(n21095), .A3(n11704), .ZN(n21100) );
  OAI221_X1 U23029 ( .B1(n21097), .B2(n21100), .C1(n21097), .C2(n11283), .A(
        n21369), .ZN(n21099) );
  OAI211_X1 U23030 ( .C1(n11283), .C2(n21101), .A(n21099), .B(n21098), .ZN(
        P3_U2857) );
  NAND2_X1 U23031 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21100), .ZN(
        n21111) );
  NOR3_X1 U23032 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21263), .A3(
        n21111), .ZN(n21104) );
  OAI22_X1 U23033 ( .A1(n21329), .A2(n21102), .B1(n21112), .B2(n21101), .ZN(
        n21103) );
  AOI211_X1 U23034 ( .C1(n21105), .C2(n21110), .A(n21104), .B(n21103), .ZN(
        n21106) );
  OAI21_X1 U23035 ( .B1(n21246), .B2(n21107), .A(n21106), .ZN(P3_U2856) );
  AOI22_X1 U23036 ( .A1(n10995), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21238), .ZN(n21120) );
  AOI22_X1 U23037 ( .A1(n21110), .A2(n21109), .B1(n21172), .B2(n21108), .ZN(
        n21119) );
  OAI22_X1 U23038 ( .A1(n21114), .A2(n21362), .B1(n21113), .B2(n21312), .ZN(
        n21115) );
  OR3_X1 U23039 ( .A1(n21117), .A2(n21116), .A3(n21115), .ZN(n21121) );
  OAI211_X1 U23040 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n21140), .A(
        n21369), .B(n21121), .ZN(n21118) );
  NAND3_X1 U23041 ( .A1(n21120), .A2(n21119), .A3(n21118), .ZN(P3_U2855) );
  AOI22_X1 U23042 ( .A1(n10995), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21238), .ZN(n21128) );
  NAND3_X1 U23043 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21336), .A3(
        n21121), .ZN(n21124) );
  NAND3_X1 U23044 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21140), .A3(
        n21122), .ZN(n21123) );
  OAI211_X1 U23045 ( .C1(n21125), .C2(n21219), .A(n21124), .B(n21123), .ZN(
        n21126) );
  AOI22_X1 U23046 ( .A1(n21369), .A2(n21126), .B1(n21373), .B2(n21125), .ZN(
        n21127) );
  OAI211_X1 U23047 ( .C1(n21246), .C2(n21129), .A(n21128), .B(n21127), .ZN(
        P3_U2854) );
  AOI21_X1 U23048 ( .B1(n21136), .B2(n21130), .A(n21162), .ZN(n21133) );
  NAND2_X1 U23049 ( .A1(n21386), .A2(n21131), .ZN(n21181) );
  OAI21_X1 U23050 ( .B1(n21132), .B2(n21268), .A(n21181), .ZN(n21364) );
  AOI211_X1 U23051 ( .C1(n21386), .C2(n21134), .A(n21133), .B(n21364), .ZN(
        n21151) );
  NAND2_X1 U23052 ( .A1(n21219), .A2(n21268), .ZN(n21148) );
  NOR2_X1 U23053 ( .A1(n21135), .A2(n21219), .ZN(n21365) );
  INV_X1 U23054 ( .A(n21136), .ZN(n21353) );
  NOR2_X1 U23055 ( .A1(n21353), .A2(n21137), .ZN(n21361) );
  OAI221_X1 U23056 ( .B1(n21363), .B2(n21361), .C1(n21363), .C2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n21369), .ZN(n21138) );
  AOI211_X1 U23057 ( .C1(n21142), .C2(n21148), .A(n21365), .B(n21138), .ZN(
        n21354) );
  OAI211_X1 U23058 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n21363), .A(
        n21151), .B(n21354), .ZN(n21139) );
  NAND2_X1 U23059 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21139), .ZN(
        n21147) );
  NAND3_X1 U23060 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21140), .ZN(n21185) );
  NAND2_X1 U23061 ( .A1(n21141), .A2(n21185), .ZN(n21153) );
  NAND2_X1 U23062 ( .A1(n21369), .A2(n21153), .ZN(n21377) );
  NOR3_X1 U23063 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21142), .A3(
        n21377), .ZN(n21143) );
  AOI21_X1 U23064 ( .B1(n21373), .B2(n21144), .A(n21143), .ZN(n21145) );
  OAI221_X1 U23065 ( .B1(n10995), .B2(n21147), .C1(n21329), .C2(n21146), .A(
        n21145), .ZN(P3_U2851) );
  AOI21_X1 U23066 ( .B1(n21152), .B2(n21361), .A(n21363), .ZN(n21161) );
  INV_X1 U23067 ( .A(n21148), .ZN(n21320) );
  NAND2_X1 U23068 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21149) );
  AOI21_X1 U23069 ( .B1(n21367), .B2(n21149), .A(n21365), .ZN(n21150) );
  OAI211_X1 U23070 ( .C1(n21152), .C2(n21320), .A(n21151), .B(n21150), .ZN(
        n21347) );
  NOR3_X1 U23071 ( .A1(n21161), .A2(n21347), .A3(n11751), .ZN(n21159) );
  OAI221_X1 U23072 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21154), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n21153), .A(n21369), .ZN(
        n21158) );
  AOI22_X1 U23073 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21238), .B1(
        n21373), .B2(n21155), .ZN(n21157) );
  OAI211_X1 U23074 ( .C1(n21159), .C2(n21158), .A(n21157), .B(n21156), .ZN(
        P3_U2850) );
  NOR2_X1 U23075 ( .A1(n21160), .A2(n21185), .ZN(n21168) );
  INV_X1 U23076 ( .A(n21181), .ZN(n21165) );
  AOI21_X1 U23077 ( .B1(n21386), .B2(n11751), .A(n21161), .ZN(n21345) );
  OAI221_X1 U23078 ( .B1(n21163), .B2(n21162), .C1(n21163), .C2(n21303), .A(
        n21345), .ZN(n21164) );
  AOI211_X1 U23079 ( .C1(n21367), .C2(n21353), .A(n21165), .B(n21164), .ZN(
        n21166) );
  INV_X1 U23080 ( .A(n21166), .ZN(n21167) );
  MUX2_X1 U23081 ( .A(n21168), .B(n21167), .S(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n21169) );
  AOI21_X1 U23082 ( .B1(n21293), .B2(n21170), .A(n21169), .ZN(n21176) );
  AOI22_X1 U23083 ( .A1(n10995), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21238), .ZN(n21175) );
  AOI22_X1 U23084 ( .A1(n21373), .A2(n21173), .B1(n21172), .B2(n21171), .ZN(
        n21174) );
  OAI211_X1 U23085 ( .C1(n21176), .C2(n21263), .A(n21175), .B(n21174), .ZN(
        P3_U2848) );
  NOR2_X1 U23086 ( .A1(n21177), .A2(n21219), .ZN(n21190) );
  AOI21_X1 U23087 ( .B1(n21363), .B2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n21178), .ZN(n21179) );
  AOI21_X1 U23088 ( .B1(n21367), .B2(n21180), .A(n21179), .ZN(n21182) );
  OAI211_X1 U23089 ( .C1(n21183), .C2(n21312), .A(n21182), .B(n21181), .ZN(
        n21335) );
  NAND2_X1 U23090 ( .A1(n21183), .A2(n21335), .ZN(n21184) );
  OAI22_X1 U23091 ( .A1(n21268), .A2(n21186), .B1(n21185), .B2(n21184), .ZN(
        n21187) );
  AOI21_X1 U23092 ( .B1(n21188), .B2(n21190), .A(n21187), .ZN(n21195) );
  AOI22_X1 U23093 ( .A1(n10995), .A2(P3_REIP_REG_15__SCAN_IN), .B1(n21373), 
        .B2(n21189), .ZN(n21194) );
  INV_X1 U23094 ( .A(n21190), .ZN(n21191) );
  OAI211_X1 U23095 ( .C1(n21192), .C2(n21268), .A(n21369), .B(n21191), .ZN(
        n21337) );
  OAI211_X1 U23096 ( .C1(n21335), .C2(n21337), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n21329), .ZN(n21193) );
  OAI211_X1 U23097 ( .C1(n21195), .C2(n21263), .A(n21194), .B(n21193), .ZN(
        P3_U2847) );
  INV_X1 U23098 ( .A(n21276), .ZN(n21200) );
  OAI22_X1 U23099 ( .A1(n21363), .A2(n21196), .B1(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n21356), .ZN(n21197) );
  NOR2_X1 U23100 ( .A1(n21198), .A2(n21197), .ZN(n21199) );
  MUX2_X1 U23101 ( .A(n21200), .B(n21199), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n21204) );
  AOI22_X1 U23102 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21238), .B1(
        n21373), .B2(n21201), .ZN(n21203) );
  NAND2_X1 U23103 ( .A1(n10995), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21202) );
  OAI211_X1 U23104 ( .C1(n21263), .C2(n21204), .A(n21203), .B(n21202), .ZN(
        P3_U2840) );
  OAI21_X1 U23105 ( .B1(n21207), .B2(n21206), .A(n21205), .ZN(n21213) );
  NAND2_X1 U23106 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21208) );
  NOR3_X1 U23107 ( .A1(n21208), .A2(n21267), .A3(n21271), .ZN(n21209) );
  OAI21_X1 U23108 ( .B1(n21285), .B2(n21209), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21222) );
  INV_X1 U23109 ( .A(n21210), .ZN(n21212) );
  AOI222_X1 U23110 ( .A1(n21213), .A2(n21222), .B1(n21384), .B2(n21212), .C1(
        n21293), .C2(n21211), .ZN(n21217) );
  AOI22_X1 U23111 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21238), .B1(
        n21373), .B2(n21214), .ZN(n21216) );
  NAND2_X1 U23112 ( .A1(n10995), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21215) );
  OAI211_X1 U23113 ( .C1(n21217), .C2(n21263), .A(n21216), .B(n21215), .ZN(
        P3_U2837) );
  NAND2_X1 U23114 ( .A1(n21218), .A2(n21229), .ZN(n21225) );
  NOR2_X1 U23115 ( .A1(n21220), .A2(n21219), .ZN(n21221) );
  AOI211_X1 U23116 ( .C1(n21336), .C2(n21222), .A(n21221), .B(n21229), .ZN(
        n21223) );
  OAI22_X1 U23117 ( .A1(n21236), .A2(n21246), .B1(n21223), .B2(n21263), .ZN(
        n21224) );
  AOI22_X1 U23118 ( .A1(n21373), .A2(n21226), .B1(n21225), .B2(n21224), .ZN(
        n21228) );
  OAI211_X1 U23119 ( .C1(n21275), .C2(n21229), .A(n21228), .B(n21227), .ZN(
        P3_U2836) );
  INV_X1 U23120 ( .A(n21230), .ZN(n21242) );
  INV_X1 U23121 ( .A(n21231), .ZN(n21232) );
  AOI211_X1 U23122 ( .C1(n21293), .C2(n21234), .A(n21233), .B(n21232), .ZN(
        n21235) );
  OAI22_X1 U23123 ( .A1(n21236), .A2(n21246), .B1(n21235), .B2(n21263), .ZN(
        n21239) );
  AOI222_X1 U23124 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21239), 
        .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21238), .C1(n21239), 
        .C2(n21237), .ZN(n21241) );
  OAI211_X1 U23125 ( .C1(n21242), .C2(n21333), .A(n21241), .B(n21240), .ZN(
        P3_U2835) );
  AOI21_X1 U23126 ( .B1(n21244), .B2(n21293), .A(n21243), .ZN(n21248) );
  INV_X1 U23127 ( .A(n21245), .ZN(n21247) );
  OAI22_X1 U23128 ( .A1(n21248), .A2(n21263), .B1(n21247), .B2(n21246), .ZN(
        n21261) );
  AOI21_X1 U23129 ( .B1(n21250), .B2(n21261), .A(n21249), .ZN(n21256) );
  OAI211_X1 U23130 ( .C1(n21263), .C2(n21254), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n21329), .ZN(n21255) );
  OAI211_X1 U23131 ( .C1(n21257), .C2(n21333), .A(n21256), .B(n21255), .ZN(
        P3_U2833) );
  AOI22_X1 U23132 ( .A1(n10995), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n21373), 
        .B2(n21258), .ZN(n21266) );
  INV_X1 U23133 ( .A(n21259), .ZN(n21260) );
  NAND3_X1 U23134 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21261), .A3(
        n21262), .ZN(n21265) );
  OAI211_X1 U23135 ( .C1(n21263), .C2(n21262), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n21329), .ZN(n21264) );
  NAND3_X1 U23136 ( .A1(n21266), .A2(n21265), .A3(n21264), .ZN(P3_U2832) );
  NAND2_X1 U23137 ( .A1(n21386), .A2(n21267), .ZN(n21273) );
  OAI21_X1 U23138 ( .B1(n21269), .B2(n21268), .A(n21275), .ZN(n21270) );
  AOI211_X1 U23139 ( .C1(n21293), .C2(n21272), .A(n21271), .B(n21270), .ZN(
        n21284) );
  NAND3_X1 U23140 ( .A1(n21273), .A2(n10990), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21274) );
  NAND2_X1 U23141 ( .A1(n21274), .A2(n21329), .ZN(n21282) );
  NAND3_X1 U23142 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21276), .A3(
        n21275), .ZN(n21279) );
  AOI22_X1 U23143 ( .A1(n10995), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n21373), 
        .B2(n21277), .ZN(n21278) );
  OAI221_X1 U23144 ( .B1(n21282), .B2(n21280), .C1(n21282), .C2(n21279), .A(
        n21278), .ZN(P3_U2839) );
  INV_X1 U23145 ( .A(n21281), .ZN(n21308) );
  AOI211_X1 U23146 ( .C1(n21285), .C2(n10990), .A(n21283), .B(n21282), .ZN(
        n21286) );
  AOI211_X1 U23147 ( .C1(n21373), .C2(n21288), .A(n21287), .B(n21286), .ZN(
        n21289) );
  OAI21_X1 U23148 ( .B1(n21308), .B2(n21290), .A(n21289), .ZN(P3_U2838) );
  AOI22_X1 U23149 ( .A1(n21293), .A2(n21292), .B1(n21384), .B2(n21291), .ZN(
        n21295) );
  NAND3_X1 U23150 ( .A1(n21296), .A2(n21295), .A3(n21294), .ZN(n21297) );
  NAND2_X1 U23151 ( .A1(n21297), .A2(n21329), .ZN(n21301) );
  AOI22_X1 U23152 ( .A1(n10995), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n21373), 
        .B2(n21298), .ZN(n21299) );
  OAI221_X1 U23153 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21308), 
        .C1(n21300), .C2(n21301), .A(n21299), .ZN(P3_U2843) );
  NAND2_X1 U23154 ( .A1(n21300), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21302) );
  OAI21_X1 U23155 ( .B1(n21303), .B2(n21302), .A(n21301), .ZN(n21305) );
  AOI22_X1 U23156 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21305), .B1(
        n21373), .B2(n21304), .ZN(n21307) );
  OAI211_X1 U23157 ( .C1(n21309), .C2(n21308), .A(n21307), .B(n21306), .ZN(
        P3_U2842) );
  NOR3_X1 U23158 ( .A1(n21365), .A2(n21311), .A3(n21310), .ZN(n21319) );
  AOI21_X1 U23159 ( .B1(n21314), .B2(n21313), .A(n21312), .ZN(n21315) );
  AOI221_X1 U23160 ( .B1(n21316), .B2(n21321), .C1(n21338), .C2(n21321), .A(
        n21315), .ZN(n21317) );
  OAI211_X1 U23161 ( .C1(n21320), .C2(n21319), .A(n21318), .B(n21317), .ZN(
        n21328) );
  OAI221_X1 U23162 ( .B1(n21328), .B2(n21321), .C1(n21328), .C2(n21330), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21327) );
  NOR2_X1 U23163 ( .A1(n21322), .A2(n21377), .ZN(n21339) );
  AOI22_X1 U23164 ( .A1(n21373), .A2(n21324), .B1(n21339), .B2(n21323), .ZN(
        n21325) );
  OAI221_X1 U23165 ( .B1(n10995), .B2(n21327), .C1(n21329), .C2(n21326), .A(
        n21325), .ZN(P3_U2844) );
  OAI221_X1 U23166 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n21329), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n10995), .A(n21328), .ZN(
        n21332) );
  NAND3_X1 U23167 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21339), .A3(
        n21330), .ZN(n21331) );
  OAI211_X1 U23168 ( .C1(n21334), .C2(n21333), .A(n21332), .B(n21331), .ZN(
        P3_U2845) );
  OAI221_X1 U23169 ( .B1(n21337), .B2(n21336), .C1(n21337), .C2(n21335), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21343) );
  AOI22_X1 U23170 ( .A1(n21340), .A2(n21373), .B1(n21339), .B2(n21338), .ZN(
        n21341) );
  OAI221_X1 U23171 ( .B1(n10995), .B2(n21343), .C1(n21329), .C2(n21342), .A(
        n21341), .ZN(P3_U2846) );
  AOI22_X1 U23172 ( .A1(n10995), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21373), 
        .B2(n21344), .ZN(n21349) );
  NAND2_X1 U23173 ( .A1(n21369), .A2(n21345), .ZN(n21346) );
  OAI211_X1 U23174 ( .C1(n21347), .C2(n21346), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n21329), .ZN(n21348) );
  OAI211_X1 U23175 ( .C1(n21350), .C2(n21377), .A(n21349), .B(n21348), .ZN(
        P3_U2849) );
  NAND2_X1 U23176 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21351), .ZN(
        n21360) );
  AOI22_X1 U23177 ( .A1(n10995), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21373), 
        .B2(n21352), .ZN(n21359) );
  NAND2_X1 U23178 ( .A1(n21367), .A2(n21353), .ZN(n21355) );
  OAI211_X1 U23179 ( .C1(n21356), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n21355), .B(n21354), .ZN(n21357) );
  OAI211_X1 U23180 ( .C1(n21364), .C2(n21357), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21329), .ZN(n21358) );
  OAI211_X1 U23181 ( .C1(n21360), .C2(n21377), .A(n21359), .B(n21358), .ZN(
        P3_U2852) );
  AOI211_X1 U23182 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n21363), .A(
        n21362), .B(n21361), .ZN(n21371) );
  AOI211_X1 U23183 ( .C1(n21367), .C2(n21366), .A(n21365), .B(n21364), .ZN(
        n21368) );
  NAND2_X1 U23184 ( .A1(n21369), .A2(n21368), .ZN(n21370) );
  OAI21_X1 U23185 ( .B1(n21371), .B2(n21370), .A(n21329), .ZN(n21375) );
  AOI22_X1 U23186 ( .A1(n10995), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n21373), 
        .B2(n21372), .ZN(n21374) );
  OAI221_X1 U23187 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21377), .C1(
        n21376), .C2(n21375), .A(n21374), .ZN(P3_U2853) );
  NAND2_X1 U23188 ( .A1(n21900), .A2(n18415), .ZN(n21428) );
  INV_X1 U23189 ( .A(n21378), .ZN(n21421) );
  INV_X1 U23190 ( .A(n21379), .ZN(n21415) );
  OAI22_X1 U23191 ( .A1(n21382), .A2(n21381), .B1(n21405), .B2(n21380), .ZN(
        n21383) );
  AOI221_X1 U23192 ( .B1(n21386), .B2(n21385), .C1(n21384), .C2(n21385), .A(
        n21383), .ZN(n21442) );
  NOR2_X1 U23193 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21411) );
  OAI222_X1 U23194 ( .A1(n21390), .A2(n21389), .B1(n21390), .B2(n21388), .C1(
        n21389), .C2(n21387), .ZN(n21392) );
  OAI21_X1 U23195 ( .B1(n21392), .B2(n21393), .A(n21391), .ZN(n21397) );
  MUX2_X1 U23196 ( .A(n21395), .B(n21394), .S(n21393), .Z(n21399) );
  INV_X1 U23197 ( .A(n21399), .ZN(n21396) );
  OAI222_X1 U23198 ( .A1(n21398), .A2(n21397), .B1(n21398), .B2(n21396), .C1(
        n21397), .C2(n21396), .ZN(n21400) );
  INV_X1 U23199 ( .A(n21400), .ZN(n21410) );
  OAI221_X1 U23200 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n21400), .A(n21399), .ZN(
        n21401) );
  NOR2_X1 U23201 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(P3_MORE_REG_SCAN_IN), .ZN(
        n21408) );
  NAND3_X1 U23202 ( .A1(n21405), .A2(n21404), .A3(n11138), .ZN(n21439) );
  OAI211_X1 U23203 ( .C1(n21408), .C2(n21439), .A(n21407), .B(n21406), .ZN(
        n21409) );
  AOI211_X1 U23204 ( .C1(n21416), .C2(n21415), .A(n21414), .B(n21434), .ZN(
        n21423) );
  AOI21_X1 U23205 ( .B1(n21900), .B2(n21417), .A(n21423), .ZN(n21437) );
  NAND3_X1 U23206 ( .A1(n21419), .A2(n21437), .A3(n21418), .ZN(n21420) );
  NAND4_X1 U23207 ( .A1(n21422), .A2(n21428), .A3(n21421), .A4(n21420), .ZN(
        P3_U2997) );
  NOR2_X1 U23208 ( .A1(n21423), .A2(n21438), .ZN(n21427) );
  INV_X1 U23209 ( .A(n21424), .ZN(n21425) );
  OAI21_X1 U23210 ( .B1(n21427), .B2(n21426), .A(n21425), .ZN(P3_U3282) );
  OAI211_X1 U23211 ( .C1(n21430), .C2(n21429), .A(n21438), .B(n21428), .ZN(
        n21431) );
  INV_X1 U23212 ( .A(n21431), .ZN(n21432) );
  AOI211_X1 U23213 ( .C1(n21440), .C2(n21434), .A(n21433), .B(n21432), .ZN(
        n21435) );
  OAI221_X1 U23214 ( .B1(n21438), .B2(n21437), .C1(n21438), .C2(n21436), .A(
        n21435), .ZN(P3_U2996) );
  NAND2_X1 U23215 ( .A1(n21440), .A2(n21439), .ZN(n21444) );
  NAND2_X1 U23216 ( .A1(n21444), .A2(P3_MORE_REG_SCAN_IN), .ZN(n21441) );
  OAI21_X1 U23217 ( .B1(n21444), .B2(n21442), .A(n21441), .ZN(P3_U3295) );
  AOI21_X1 U23218 ( .B1(n21444), .B2(P3_FLUSH_REG_SCAN_IN), .A(n21443), .ZN(
        n21445) );
  INV_X1 U23219 ( .A(n21445), .ZN(P3_U2637) );
  AOI21_X1 U23220 ( .B1(n21447), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21446), 
        .ZN(n21450) );
  NOR2_X1 U23221 ( .A1(n21448), .A2(n21447), .ZN(n21449) );
  NOR4_X1 U23222 ( .A1(n21450), .A2(n21449), .A3(n21866), .A4(n13234), .ZN(
        n21452) );
  OAI21_X1 U23223 ( .B1(n21452), .B2(n21832), .A(n21451), .ZN(n21458) );
  AOI211_X1 U23224 ( .C1(n21456), .C2(n21455), .A(n21454), .B(n21453), .ZN(
        n21457) );
  MUX2_X1 U23225 ( .A(n21458), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21457), 
        .Z(P1_U3485) );
  AOI22_X1 U23226 ( .A1(n21625), .A2(n21460), .B1(n21624), .B2(n21459), .ZN(
        n21471) );
  NAND2_X1 U23227 ( .A1(n21639), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n21470) );
  INV_X1 U23228 ( .A(n21461), .ZN(n21502) );
  NAND2_X1 U23229 ( .A1(n21502), .A2(n21573), .ZN(n21499) );
  NOR2_X1 U23230 ( .A1(n21462), .A2(n21499), .ZN(n21555) );
  NOR2_X1 U23231 ( .A1(n21549), .A2(n21463), .ZN(n21566) );
  NAND3_X1 U23232 ( .A1(n21465), .A2(n21566), .A3(n21464), .ZN(n21469) );
  OAI21_X1 U23233 ( .B1(n21467), .B2(n21466), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21468) );
  NAND4_X1 U23234 ( .A1(n21471), .A2(n21470), .A3(n21469), .A4(n21468), .ZN(
        P1_U3017) );
  NAND2_X1 U23235 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21573), .ZN(
        n21480) );
  NOR3_X1 U23236 ( .A1(n21472), .A2(n21632), .A3(n21501), .ZN(n21473) );
  AOI211_X1 U23237 ( .C1(n21632), .C2(n21551), .A(n21473), .B(n21481), .ZN(
        n21478) );
  OAI22_X1 U23238 ( .A1(n21642), .A2(n21474), .B1(n21673), .B2(n21596), .ZN(
        n21475) );
  NOR2_X1 U23239 ( .A1(n21501), .A2(n21485), .ZN(n21482) );
  AOI211_X1 U23240 ( .C1(n21476), .C2(n21624), .A(n21475), .B(n21482), .ZN(
        n21477) );
  OAI221_X1 U23241 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21480), .C1(
        n21479), .C2(n21478), .A(n21477), .ZN(P1_U3029) );
  INV_X1 U23242 ( .A(n21484), .ZN(n21483) );
  AOI211_X1 U23243 ( .C1(n21551), .C2(n21483), .A(n21482), .B(n21481), .ZN(
        n21495) );
  AOI22_X1 U23244 ( .A1(n21575), .A2(n21485), .B1(n21484), .B2(n21573), .ZN(
        n21497) );
  AOI211_X1 U23245 ( .C1(n21492), .C2(n21496), .A(n21497), .B(n21486), .ZN(
        n21489) );
  INV_X1 U23246 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21487) );
  OAI22_X1 U23247 ( .A1(n21642), .A2(n21668), .B1(n21487), .B2(n21596), .ZN(
        n21488) );
  AOI211_X1 U23248 ( .C1(n21490), .C2(n21624), .A(n21489), .B(n21488), .ZN(
        n21491) );
  OAI21_X1 U23249 ( .B1(n21495), .B2(n21492), .A(n21491), .ZN(P1_U3027) );
  AOI222_X1 U23250 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n21639), .B1(n21625), 
        .B2(n21661), .C1(n21624), .C2(n21493), .ZN(n21494) );
  OAI221_X1 U23251 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21497), .C1(
        n21496), .C2(n21495), .A(n21494), .ZN(P1_U3028) );
  AOI22_X1 U23252 ( .A1(n21498), .A2(n21624), .B1(n21639), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n21505) );
  INV_X1 U23253 ( .A(n21549), .ZN(n21518) );
  NOR2_X1 U23254 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21499), .ZN(
        n21511) );
  OR2_X1 U23255 ( .A1(n21501), .A2(n21500), .ZN(n21508) );
  OAI211_X1 U23256 ( .C1(n21503), .C2(n21502), .A(n21508), .B(n21554), .ZN(
        n21506) );
  NOR2_X1 U23257 ( .A1(n21511), .A2(n21506), .ZN(n21532) );
  NAND2_X1 U23258 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21532), .ZN(
        n21514) );
  OAI21_X1 U23259 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21518), .A(
        n21514), .ZN(n21504) );
  OAI211_X1 U23260 ( .C1(n21699), .C2(n21642), .A(n21505), .B(n21504), .ZN(
        P1_U3025) );
  AOI22_X1 U23261 ( .A1(n21507), .A2(n21624), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n21506), .ZN(n21513) );
  OAI22_X1 U23262 ( .A1(n21596), .A2(n21696), .B1(n21509), .B2(n21508), .ZN(
        n21510) );
  AOI211_X1 U23263 ( .C1(n21625), .C2(n21685), .A(n21511), .B(n21510), .ZN(
        n21512) );
  NAND2_X1 U23264 ( .A1(n21513), .A2(n21512), .ZN(P1_U3026) );
  NAND2_X1 U23265 ( .A1(n21515), .A2(n21514), .ZN(n21524) );
  OAI22_X1 U23266 ( .A1(n21711), .A2(n21642), .B1(n21717), .B2(n21596), .ZN(
        n21516) );
  AOI21_X1 U23267 ( .B1(n21517), .B2(n21624), .A(n21516), .ZN(n21519) );
  NAND3_X1 U23268 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21522), .A3(
        n21518), .ZN(n21525) );
  OAI211_X1 U23269 ( .C1(n21522), .C2(n21524), .A(n21519), .B(n21525), .ZN(
        P1_U3024) );
  INV_X1 U23270 ( .A(n21520), .ZN(n21528) );
  NOR4_X1 U23271 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21549), .A3(
        n21522), .A4(n21521), .ZN(n21527) );
  AOI21_X1 U23272 ( .B1(n21525), .B2(n21524), .A(n21523), .ZN(n21526) );
  AOI211_X1 U23273 ( .C1(n21528), .C2(n21624), .A(n21527), .B(n21526), .ZN(
        n21530) );
  NAND2_X1 U23274 ( .A1(n21639), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n21529) );
  OAI211_X1 U23275 ( .C1(n21642), .C2(n21722), .A(n21530), .B(n21529), .ZN(
        P1_U3023) );
  INV_X1 U23276 ( .A(n21531), .ZN(n21535) );
  OAI21_X1 U23277 ( .B1(n21534), .B2(n21533), .A(n21532), .ZN(n21544) );
  AOI22_X1 U23278 ( .A1(n21535), .A2(n21624), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21544), .ZN(n21539) );
  NOR2_X1 U23279 ( .A1(n21596), .A2(n21743), .ZN(n21537) );
  NOR3_X1 U23280 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21549), .A3(
        n21536), .ZN(n21545) );
  AOI211_X1 U23281 ( .C1(n21625), .C2(n21736), .A(n21537), .B(n21545), .ZN(
        n21538) );
  NAND2_X1 U23282 ( .A1(n21539), .A2(n21538), .ZN(P1_U3022) );
  NAND2_X1 U23283 ( .A1(n21540), .A2(n12323), .ZN(n21542) );
  OAI22_X1 U23284 ( .A1(n21549), .A2(n21542), .B1(n21635), .B2(n21541), .ZN(
        n21543) );
  AOI221_X1 U23285 ( .B1(n21545), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n21544), .C2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n21543), .ZN(
        n21547) );
  NAND2_X1 U23286 ( .A1(n21639), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n21546) );
  OAI211_X1 U23287 ( .C1(n21642), .C2(n21548), .A(n21547), .B(n21546), .ZN(
        P1_U3021) );
  NOR2_X1 U23288 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21549), .ZN(
        n21561) );
  AOI22_X1 U23289 ( .A1(n21575), .A2(n21552), .B1(n21551), .B2(n21550), .ZN(
        n21553) );
  NAND2_X1 U23290 ( .A1(n21554), .A2(n21553), .ZN(n21567) );
  AOI21_X1 U23291 ( .B1(n21555), .B2(n12191), .A(n21567), .ZN(n21557) );
  OAI22_X1 U23292 ( .A1(n21558), .A2(n21635), .B1(n21557), .B2(n21556), .ZN(
        n21559) );
  AOI21_X1 U23293 ( .B1(n21561), .B2(n21560), .A(n21559), .ZN(n21563) );
  NAND2_X1 U23294 ( .A1(n21639), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n21562) );
  OAI211_X1 U23295 ( .C1(n21642), .C2(n21564), .A(n21563), .B(n21562), .ZN(
        P1_U3019) );
  AOI22_X1 U23296 ( .A1(n21639), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n21625), 
        .B2(n21565), .ZN(n21569) );
  AOI22_X1 U23297 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21567), .B1(
        n21566), .B2(n12191), .ZN(n21568) );
  OAI211_X1 U23298 ( .C1(n21570), .C2(n21635), .A(n21569), .B(n21568), .ZN(
        P1_U3020) );
  INV_X1 U23299 ( .A(n21571), .ZN(n21572) );
  AOI22_X1 U23300 ( .A1(n21575), .A2(n21574), .B1(n21573), .B2(n21572), .ZN(
        n21598) );
  NOR2_X1 U23301 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21598), .ZN(
        n21603) );
  AOI21_X1 U23302 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n21639), .A(n21603), 
        .ZN(n21579) );
  INV_X1 U23303 ( .A(n21576), .ZN(n21602) );
  AOI22_X1 U23304 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21602), .B1(
        n21625), .B2(n21577), .ZN(n21578) );
  OAI211_X1 U23305 ( .C1(n21635), .C2(n21580), .A(n21579), .B(n21578), .ZN(
        P1_U3016) );
  INV_X1 U23306 ( .A(n21581), .ZN(n21582) );
  OAI22_X1 U23307 ( .A1(n21582), .A2(n21635), .B1(n21642), .B2(n21764), .ZN(
        n21583) );
  AOI21_X1 U23308 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n21591), .A(
        n21583), .ZN(n21587) );
  INV_X1 U23309 ( .A(n21598), .ZN(n21584) );
  NAND3_X1 U23310 ( .A1(n21585), .A2(n12349), .A3(n21584), .ZN(n21586) );
  OAI211_X1 U23311 ( .C1(n21757), .C2(n21596), .A(n21587), .B(n21586), .ZN(
        P1_U3013) );
  OAI21_X1 U23312 ( .B1(n21598), .B2(n21589), .A(n21588), .ZN(n21590) );
  AOI22_X1 U23313 ( .A1(n21625), .A2(n21592), .B1(n21591), .B2(n21590), .ZN(
        n21594) );
  NAND2_X1 U23314 ( .A1(n21639), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n21593) );
  OAI211_X1 U23315 ( .C1(n21595), .C2(n21635), .A(n21594), .B(n21593), .ZN(
        P1_U3014) );
  NOR2_X1 U23316 ( .A1(n21596), .A2(n21745), .ZN(n21600) );
  NOR3_X1 U23317 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21598), .A3(
        n21597), .ZN(n21599) );
  AOI211_X1 U23318 ( .C1(n21624), .C2(n21601), .A(n21600), .B(n21599), .ZN(
        n21605) );
  OAI21_X1 U23319 ( .B1(n21603), .B2(n21602), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21604) );
  OAI211_X1 U23320 ( .C1(n21642), .C2(n21748), .A(n21605), .B(n21604), .ZN(
        P1_U3015) );
  NOR2_X1 U23321 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12197), .ZN(
        n21607) );
  AOI22_X1 U23322 ( .A1(n21639), .A2(P1_REIP_REG_20__SCAN_IN), .B1(n21607), 
        .B2(n21606), .ZN(n21613) );
  NAND2_X1 U23323 ( .A1(n21608), .A2(n21615), .ZN(n21609) );
  NAND2_X1 U23324 ( .A1(n12197), .A2(n21609), .ZN(n21614) );
  AOI21_X1 U23325 ( .B1(n21621), .B2(n21614), .A(n12355), .ZN(n21610) );
  AOI21_X1 U23326 ( .B1(n21611), .B2(n21624), .A(n21610), .ZN(n21612) );
  OAI211_X1 U23327 ( .C1(n21642), .C2(n21783), .A(n21613), .B(n21612), .ZN(
        P1_U3011) );
  AOI21_X1 U23328 ( .B1(n21616), .B2(n21615), .A(n21614), .ZN(n21617) );
  AOI21_X1 U23329 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n21639), .A(n21617), 
        .ZN(n21620) );
  AOI22_X1 U23330 ( .A1(n21625), .A2(n21770), .B1(n21624), .B2(n21618), .ZN(
        n21619) );
  OAI211_X1 U23331 ( .C1(n21621), .C2(n12197), .A(n21620), .B(n21619), .ZN(
        P1_U3012) );
  AOI21_X1 U23332 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n21639), .A(n21622), 
        .ZN(n21627) );
  AOI22_X1 U23333 ( .A1(n21625), .A2(n21800), .B1(n21624), .B2(n21623), .ZN(
        n21626) );
  OAI211_X1 U23334 ( .C1(n21629), .C2(n21628), .A(n21627), .B(n21626), .ZN(
        P1_U3010) );
  INV_X1 U23335 ( .A(n21630), .ZN(n21638) );
  NAND3_X1 U23336 ( .A1(n21633), .A2(n21632), .A3(n21631), .ZN(n21634) );
  OAI21_X1 U23337 ( .B1(n21636), .B2(n21635), .A(n21634), .ZN(n21637) );
  AOI21_X1 U23338 ( .B1(n21638), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n21637), .ZN(n21641) );
  NAND2_X1 U23339 ( .A1(n21639), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21640) );
  OAI211_X1 U23340 ( .C1(n21643), .C2(n21642), .A(n21641), .B(n21640), .ZN(
        P1_U3030) );
  INV_X1 U23341 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21645) );
  AOI22_X1 U23342 ( .A1(n21720), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n21721), 
        .B2(n21674), .ZN(n21644) );
  OAI21_X1 U23343 ( .B1(n21820), .B2(n21645), .A(n21644), .ZN(n21646) );
  AOI21_X1 U23344 ( .B1(n22053), .B2(n21647), .A(n21646), .ZN(n21654) );
  INV_X1 U23345 ( .A(n21648), .ZN(n21650) );
  OAI22_X1 U23346 ( .A1(n21650), .A2(n21812), .B1(n21649), .B2(n21765), .ZN(
        n21651) );
  AOI21_X1 U23347 ( .B1(n21652), .B2(n21679), .A(n21651), .ZN(n21653) );
  OAI211_X1 U23348 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n21795), .A(
        n21654), .B(n21653), .ZN(P1_U2839) );
  INV_X1 U23349 ( .A(n14694), .ZN(n21663) );
  INV_X1 U23350 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21672) );
  AOI221_X1 U23351 ( .B1(n21674), .B2(n21721), .C1(n21673), .C2(n21721), .A(
        n21720), .ZN(n21655) );
  NAND2_X1 U23352 ( .A1(n21672), .A2(n21655), .ZN(n21659) );
  NAND2_X1 U23353 ( .A1(n21792), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n21658) );
  INV_X1 U23354 ( .A(n21655), .ZN(n21656) );
  AOI22_X1 U23355 ( .A1(n21810), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n21656), .ZN(n21657) );
  OAI211_X1 U23356 ( .C1(n21659), .C2(n21732), .A(n21658), .B(n21657), .ZN(
        n21660) );
  AOI21_X1 U23357 ( .B1(n21801), .B2(n21661), .A(n21660), .ZN(n21662) );
  OAI21_X1 U23358 ( .B1(n21663), .B2(n21669), .A(n21662), .ZN(n21664) );
  AOI21_X1 U23359 ( .B1(n21665), .B2(n21679), .A(n21664), .ZN(n21666) );
  OAI21_X1 U23360 ( .B1(n21667), .B2(n21795), .A(n21666), .ZN(P1_U2837) );
  OAI22_X1 U23361 ( .A1(n21670), .A2(n21669), .B1(n21812), .B2(n21668), .ZN(
        n21671) );
  AOI211_X1 U23362 ( .C1(n21792), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21769), .B(n21671), .ZN(n21682) );
  AOI21_X1 U23363 ( .B1(n21721), .B2(n21684), .A(n21720), .ZN(n21697) );
  NOR3_X1 U23364 ( .A1(n21674), .A2(n21673), .A3(n21672), .ZN(n21675) );
  AOI21_X1 U23365 ( .B1(n21675), .B2(n21721), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n21677) );
  OAI22_X1 U23366 ( .A1(n21697), .A2(n21677), .B1(n21676), .B2(n21795), .ZN(
        n21678) );
  AOI21_X1 U23367 ( .B1(n21680), .B2(n21679), .A(n21678), .ZN(n21681) );
  OAI211_X1 U23368 ( .C1(n21683), .C2(n21765), .A(n21682), .B(n21681), .ZN(
        P1_U2836) );
  NOR3_X1 U23369 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21684), .A3(n21732), .ZN(
        n21694) );
  AOI22_X1 U23370 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n21810), .B1(n21801), .B2(
        n21685), .ZN(n21687) );
  OAI211_X1 U23371 ( .C1(n21820), .C2(n21688), .A(n21687), .B(n21686), .ZN(
        n21693) );
  OAI22_X1 U23372 ( .A1(n21691), .A2(n21690), .B1(n21689), .B2(n21795), .ZN(
        n21692) );
  NOR3_X1 U23373 ( .A1(n21694), .A2(n21693), .A3(n21692), .ZN(n21695) );
  OAI21_X1 U23374 ( .B1(n21697), .B2(n21696), .A(n21695), .ZN(P1_U2835) );
  AOI21_X1 U23375 ( .B1(n21721), .B2(n21708), .A(n21720), .ZN(n21718) );
  AOI21_X1 U23376 ( .B1(n21698), .B2(n21721), .A(P1_REIP_REG_6__SCAN_IN), .ZN(
        n21707) );
  OAI22_X1 U23377 ( .A1(n21700), .A2(n21765), .B1(n21812), .B2(n21699), .ZN(
        n21701) );
  AOI211_X1 U23378 ( .C1(n21792), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n21769), .B(n21701), .ZN(n21706) );
  NOR2_X1 U23379 ( .A1(n21795), .A2(n21702), .ZN(n21703) );
  AOI21_X1 U23380 ( .B1(n21704), .B2(n21771), .A(n21703), .ZN(n21705) );
  OAI211_X1 U23381 ( .C1(n21718), .C2(n21707), .A(n21706), .B(n21705), .ZN(
        P1_U2834) );
  NOR3_X1 U23382 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n21708), .A3(n21732), .ZN(
        n21709) );
  AOI211_X1 U23383 ( .C1(n21792), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n21769), .B(n21709), .ZN(n21710) );
  OAI21_X1 U23384 ( .B1(n21812), .B2(n21711), .A(n21710), .ZN(n21715) );
  OAI22_X1 U23385 ( .A1(n21713), .A2(n21813), .B1(n21712), .B2(n21795), .ZN(
        n21714) );
  AOI211_X1 U23386 ( .C1(P1_EBX_REG_7__SCAN_IN), .C2(n21810), .A(n21715), .B(
        n21714), .ZN(n21716) );
  OAI21_X1 U23387 ( .B1(n21718), .B2(n21717), .A(n21716), .ZN(P1_U2833) );
  AOI21_X1 U23388 ( .B1(n21719), .B2(n21721), .A(P1_REIP_REG_8__SCAN_IN), .ZN(
        n21729) );
  AOI21_X1 U23389 ( .B1(n21721), .B2(n21733), .A(n21720), .ZN(n21742) );
  OAI22_X1 U23390 ( .A1(n21723), .A2(n21765), .B1(n21812), .B2(n21722), .ZN(
        n21724) );
  AOI211_X1 U23391 ( .C1(n21792), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n21769), .B(n21724), .ZN(n21728) );
  AOI22_X1 U23392 ( .A1(n21726), .A2(n21771), .B1(n21816), .B2(n21725), .ZN(
        n21727) );
  OAI211_X1 U23393 ( .C1(n21729), .C2(n21742), .A(n21728), .B(n21727), .ZN(
        P1_U2832) );
  AOI21_X1 U23394 ( .B1(n21810), .B2(P1_EBX_REG_9__SCAN_IN), .A(n21769), .ZN(
        n21730) );
  OAI21_X1 U23395 ( .B1(n21820), .B2(n21731), .A(n21730), .ZN(n21735) );
  NOR3_X1 U23396 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n21733), .A3(n21732), .ZN(
        n21734) );
  AOI211_X1 U23397 ( .C1(n21801), .C2(n21736), .A(n21735), .B(n21734), .ZN(
        n21737) );
  OAI21_X1 U23398 ( .B1(n21738), .B2(n21813), .A(n21737), .ZN(n21739) );
  AOI21_X1 U23399 ( .B1(n21740), .B2(n21816), .A(n21739), .ZN(n21741) );
  OAI21_X1 U23400 ( .B1(n21743), .B2(n21742), .A(n21741), .ZN(P1_U2831) );
  AOI211_X1 U23401 ( .C1(n21746), .C2(n21745), .A(n21804), .B(n21744), .ZN(
        n21747) );
  AOI211_X1 U23402 ( .C1(n21792), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n21769), .B(n21747), .ZN(n21753) );
  OAI22_X1 U23403 ( .A1(n21749), .A2(n21813), .B1(n21812), .B2(n21748), .ZN(
        n21750) );
  AOI21_X1 U23404 ( .B1(n21751), .B2(n21816), .A(n21750), .ZN(n21752) );
  OAI211_X1 U23405 ( .C1(n21754), .C2(n21765), .A(n21753), .B(n21752), .ZN(
        P1_U2824) );
  AOI21_X1 U23406 ( .B1(n21810), .B2(P1_EBX_REG_18__SCAN_IN), .A(n21769), .ZN(
        n21755) );
  OAI21_X1 U23407 ( .B1(n21820), .B2(n21756), .A(n21755), .ZN(n21758) );
  AND2_X1 U23408 ( .A1(n21757), .A2(n21776), .ZN(n21773) );
  AOI211_X1 U23409 ( .C1(n21774), .C2(P1_REIP_REG_18__SCAN_IN), .A(n21758), 
        .B(n21773), .ZN(n21759) );
  OAI21_X1 U23410 ( .B1(n21760), .B2(n21813), .A(n21759), .ZN(n21761) );
  AOI21_X1 U23411 ( .B1(n21762), .B2(n21816), .A(n21761), .ZN(n21763) );
  OAI21_X1 U23412 ( .B1(n21812), .B2(n21764), .A(n21763), .ZN(P1_U2822) );
  INV_X1 U23413 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21766) );
  OAI22_X1 U23414 ( .A1(n21767), .A2(n21795), .B1(n21766), .B2(n21765), .ZN(
        n21768) );
  AOI211_X1 U23415 ( .C1(n21792), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n21769), .B(n21768), .ZN(n21780) );
  AOI22_X1 U23416 ( .A1(n21772), .A2(n21771), .B1(n21801), .B2(n21770), .ZN(
        n21779) );
  OAI21_X1 U23417 ( .B1(n21774), .B2(n21773), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n21778) );
  NAND3_X1 U23418 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n21776), .A3(n21775), 
        .ZN(n21777) );
  NAND4_X1 U23419 ( .A1(n21780), .A2(n21779), .A3(n21778), .A4(n21777), .ZN(
        P1_U2821) );
  AOI21_X1 U23420 ( .B1(n21791), .B2(n21790), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n21789) );
  NAND2_X1 U23421 ( .A1(n21782), .A2(n21781), .ZN(n21794) );
  AOI22_X1 U23422 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n21792), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(n21810), .ZN(n21788) );
  OAI22_X1 U23423 ( .A1(n21784), .A2(n21813), .B1(n21812), .B2(n21783), .ZN(
        n21785) );
  AOI21_X1 U23424 ( .B1(n21786), .B2(n21816), .A(n21785), .ZN(n21787) );
  OAI211_X1 U23425 ( .C1(n21789), .C2(n21794), .A(n21788), .B(n21787), .ZN(
        P1_U2820) );
  NAND3_X1 U23426 ( .A1(n21791), .A2(P1_REIP_REG_20__SCAN_IN), .A3(n21790), 
        .ZN(n21806) );
  AOI22_X1 U23427 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n21792), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(n21810), .ZN(n21793) );
  OAI221_X1 U23428 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n21806), .C1(n21807), 
        .C2(n21794), .A(n21793), .ZN(n21799) );
  OAI22_X1 U23429 ( .A1(n21797), .A2(n21813), .B1(n21796), .B2(n21795), .ZN(
        n21798) );
  AOI211_X1 U23430 ( .C1(n21801), .C2(n21800), .A(n21799), .B(n21798), .ZN(
        n21802) );
  INV_X1 U23431 ( .A(n21802), .ZN(P1_U2819) );
  NOR3_X1 U23432 ( .A1(n21805), .A2(n21804), .A3(n21803), .ZN(n21809) );
  NOR3_X1 U23433 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n21807), .A3(n21806), 
        .ZN(n21808) );
  AOI211_X1 U23434 ( .C1(n21810), .C2(P1_EBX_REG_22__SCAN_IN), .A(n21809), .B(
        n21808), .ZN(n21819) );
  OAI22_X1 U23435 ( .A1(n21814), .A2(n21813), .B1(n21812), .B2(n21811), .ZN(
        n21815) );
  AOI21_X1 U23436 ( .B1(n21817), .B2(n21816), .A(n21815), .ZN(n21818) );
  OAI211_X1 U23437 ( .C1(n21821), .C2(n21820), .A(n21819), .B(n21818), .ZN(
        P1_U2818) );
  OAI21_X1 U23438 ( .B1(n21824), .B2(n21823), .A(n21822), .ZN(P1_U2806) );
  OAI22_X1 U23439 ( .A1(n21828), .A2(n21827), .B1(n21826), .B2(n21825), .ZN(
        n21830) );
  MUX2_X1 U23440 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21830), .S(
        n21829), .Z(P1_U3469) );
  INV_X1 U23441 ( .A(n21831), .ZN(n21837) );
  NOR2_X1 U23442 ( .A1(n21837), .A2(n21832), .ZN(n21836) );
  AOI22_X1 U23443 ( .A1(n21836), .A2(n21834), .B1(n21833), .B2(n13234), .ZN(
        P1_U3163) );
  OAI21_X1 U23444 ( .B1(n21836), .B2(n22021), .A(n21835), .ZN(P1_U3466) );
  AOI21_X1 U23445 ( .B1(n21839), .B2(n21838), .A(n21837), .ZN(n21840) );
  OAI22_X1 U23446 ( .A1(n21842), .A2(n21841), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21840), .ZN(n21843) );
  OAI21_X1 U23447 ( .B1(n21845), .B2(n21844), .A(n21843), .ZN(P1_U3161) );
  AOI21_X1 U23448 ( .B1(n21848), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21847), 
        .ZN(n21846) );
  INV_X1 U23449 ( .A(n21846), .ZN(P1_U2805) );
  AOI21_X1 U23450 ( .B1(n21848), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21847), 
        .ZN(n21849) );
  INV_X1 U23451 ( .A(n21849), .ZN(P1_U3465) );
  INV_X1 U23452 ( .A(n21850), .ZN(n21851) );
  OAI21_X1 U23453 ( .B1(n21853), .B2(n14662), .A(n21851), .ZN(P2_U2818) );
  OAI21_X1 U23454 ( .B1(n21853), .B2(n21852), .A(n21851), .ZN(P2_U3592) );
  INV_X1 U23455 ( .A(n21854), .ZN(n21856) );
  OAI21_X1 U23456 ( .B1(n21858), .B2(n21855), .A(n21856), .ZN(P3_U2636) );
  OAI21_X1 U23457 ( .B1(n21858), .B2(n21857), .A(n21856), .ZN(P3_U3281) );
  INV_X1 U23458 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21859) );
  AOI21_X1 U23459 ( .B1(HOLD), .B2(n21860), .A(n21859), .ZN(n21863) );
  AOI21_X1 U23460 ( .B1(n21900), .B2(P3_STATE_REG_1__SCAN_IN), .A(n21861), 
        .ZN(n21916) );
  AOI21_X1 U23461 ( .B1(n21862), .B2(NA), .A(n21909), .ZN(n21914) );
  OAI22_X1 U23462 ( .A1(n21864), .A2(n21863), .B1(n21916), .B2(n21914), .ZN(
        P3_U3029) );
  NAND2_X1 U23463 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21866), .ZN(n21877) );
  AOI22_X1 U23464 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21877), .B1(NA), .B2(
        n21872), .ZN(n21870) );
  INV_X1 U23465 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21868) );
  AOI21_X1 U23466 ( .B1(n21866), .B2(n21911), .A(n21865), .ZN(n21867) );
  OAI21_X1 U23467 ( .B1(n21873), .B2(n21908), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21878) );
  INV_X1 U23468 ( .A(n21878), .ZN(n21874) );
  OAI33_X1 U23469 ( .A1(n21877), .A2(NA), .A3(n21868), .B1(n21908), .B2(n21867), .B3(n21874), .ZN(n21869) );
  AOI22_X1 U23470 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21870), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(n21869), .ZN(n21871) );
  INV_X1 U23471 ( .A(n21871), .ZN(P1_U3196) );
  NOR2_X1 U23472 ( .A1(n21872), .A2(n21908), .ZN(n21879) );
  AOI22_X1 U23473 ( .A1(n21874), .A2(P1_STATE_REG_0__SCAN_IN), .B1(n21879), 
        .B2(n21873), .ZN(n21876) );
  NAND3_X1 U23474 ( .A1(n21876), .A2(n21875), .A3(n21877), .ZN(P1_U3195) );
  AND2_X1 U23475 ( .A1(n21877), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n21881) );
  AOI211_X1 U23476 ( .C1(NA), .C2(n12216), .A(n21879), .B(n21878), .ZN(n21880)
         );
  OAI22_X1 U23477 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21881), .B1(n22398), 
        .B2(n21880), .ZN(P1_U3194) );
  NOR2_X1 U23478 ( .A1(n21882), .A2(n21908), .ZN(n21886) );
  NAND2_X1 U23479 ( .A1(n21883), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21895) );
  NAND2_X1 U23480 ( .A1(n21895), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n21894) );
  OAI21_X1 U23481 ( .B1(n21884), .B2(n21911), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n21899) );
  AOI22_X1 U23482 ( .A1(n21886), .A2(n21885), .B1(n21894), .B2(n21899), .ZN(
        n21887) );
  OAI21_X1 U23483 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n21888), .A(n21887), .ZN(P2_U3209) );
  NAND2_X1 U23484 ( .A1(n21889), .A2(HOLD), .ZN(n21892) );
  OAI211_X1 U23485 ( .C1(n21890), .C2(n21908), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21891) );
  NAND4_X1 U23486 ( .A1(n21893), .A2(n21892), .A3(n21895), .A4(n21891), .ZN(
        P2_U3210) );
  INV_X1 U23487 ( .A(n21894), .ZN(n21898) );
  OAI22_X1 U23488 ( .A1(NA), .A2(n21895), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21896) );
  OAI211_X1 U23489 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n21896), .ZN(n21897) );
  OAI221_X1 U23490 ( .B1(n21899), .B2(n21898), .C1(n21899), .C2(n21908), .A(
        n21897), .ZN(P2_U3211) );
  NOR2_X1 U23491 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21918)
         );
  OAI21_X1 U23492 ( .B1(n21909), .B2(n21908), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21901) );
  NAND2_X1 U23493 ( .A1(n21900), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n21910) );
  OAI21_X1 U23494 ( .B1(n21918), .B2(n21901), .A(n21910), .ZN(n21904) );
  OAI211_X1 U23495 ( .C1(n21909), .C2(n21908), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21902) );
  AOI21_X1 U23496 ( .B1(n21902), .B2(n21905), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21903) );
  AOI21_X1 U23497 ( .B1(n21905), .B2(n21904), .A(n21903), .ZN(n21906) );
  OAI221_X1 U23498 ( .B1(n11798), .B2(P3_STATE_REG_2__SCAN_IN), .C1(n11798), 
        .C2(n21907), .A(n21906), .ZN(P3_U3030) );
  OAI22_X1 U23499 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n21909), .B2(n21908), .ZN(n21913)
         );
  INV_X1 U23500 ( .A(n21910), .ZN(n21912) );
  OAI221_X1 U23501 ( .B1(n21913), .B2(n21912), .C1(n21913), .C2(n21911), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n21917) );
  INV_X1 U23502 ( .A(n21914), .ZN(n21915) );
  OAI22_X1 U23503 ( .A1(n21918), .A2(n21917), .B1(n21916), .B2(n21915), .ZN(
        P3_U3031) );
  INV_X1 U23504 ( .A(n22389), .ZN(n21920) );
  NAND3_X1 U23505 ( .A1(n21920), .A2(n22077), .A3(n21930), .ZN(n21922) );
  NOR2_X1 U23506 ( .A1(n22043), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22013) );
  INV_X1 U23507 ( .A(n22013), .ZN(n21921) );
  NAND2_X1 U23508 ( .A1(n21922), .A2(n21921), .ZN(n21928) );
  INV_X1 U23509 ( .A(n14536), .ZN(n21923) );
  OR2_X1 U23510 ( .A1(n14694), .A2(n21923), .ZN(n21954) );
  NOR2_X1 U23511 ( .A1(n21954), .A2(n22053), .ZN(n21925) );
  NOR3_X1 U23512 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21938) );
  INV_X1 U23513 ( .A(n21938), .ZN(n21935) );
  NOR2_X1 U23514 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21935), .ZN(
        n22305) );
  AOI22_X1 U23515 ( .A1(n22389), .A2(n22059), .B1(n22049), .B2(n22305), .ZN(
        n21932) );
  INV_X1 U23516 ( .A(n21925), .ZN(n21927) );
  INV_X1 U23517 ( .A(n22305), .ZN(n21926) );
  AOI22_X1 U23518 ( .A1(n21928), .A2(n21927), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21926), .ZN(n21929) );
  OAI211_X1 U23519 ( .C1(n11469), .C2(n13234), .A(n22002), .B(n21929), .ZN(
        n22306) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22306), .B1(
        n22312), .B2(n22078), .ZN(n21931) );
  OAI211_X1 U23521 ( .C1(n22309), .C2(n22069), .A(n21932), .B(n21931), .ZN(
        P1_U3033) );
  INV_X1 U23522 ( .A(n21954), .ZN(n21934) );
  INV_X1 U23523 ( .A(n21933), .ZN(n22030) );
  NOR2_X1 U23524 ( .A1(n22029), .A2(n21935), .ZN(n22310) );
  AOI21_X1 U23525 ( .B1(n21934), .B2(n22030), .A(n22310), .ZN(n21936) );
  OAI22_X1 U23526 ( .A1(n21936), .A2(n22043), .B1(n21935), .B2(n13234), .ZN(
        n22311) );
  AOI22_X1 U23527 ( .A1(n22311), .A2(n22048), .B1(n22049), .B2(n22310), .ZN(
        n21940) );
  OAI211_X1 U23528 ( .C1(n21953), .C2(n22050), .A(n22077), .B(n21936), .ZN(
        n21937) );
  OAI211_X1 U23529 ( .C1(n22077), .C2(n21938), .A(n22035), .B(n21937), .ZN(
        n22313) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22059), .ZN(n21939) );
  OAI211_X1 U23531 ( .C1(n22062), .C2(n22316), .A(n21940), .B(n21939), .ZN(
        P1_U3041) );
  NOR3_X1 U23532 ( .A1(n22320), .A2(n22328), .A3(n22043), .ZN(n21942) );
  NOR2_X1 U23533 ( .A1(n21942), .A2(n22013), .ZN(n21948) );
  INV_X1 U23534 ( .A(n21948), .ZN(n21943) );
  NOR2_X1 U23535 ( .A1(n21954), .A2(n14582), .ZN(n21947) );
  NOR2_X1 U23536 ( .A1(n21979), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21967) );
  NOR3_X1 U23537 ( .A1(n21944), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21951) );
  NAND2_X1 U23538 ( .A1(n22029), .A2(n21951), .ZN(n22317) );
  OAI22_X1 U23539 ( .A1(n22318), .A2(n22062), .B1(n22070), .B2(n22317), .ZN(
        n21945) );
  INV_X1 U23540 ( .A(n21945), .ZN(n21950) );
  NOR2_X1 U23541 ( .A1(n21967), .A2(n13234), .ZN(n21971) );
  AOI21_X1 U23542 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22317), .A(n21971), 
        .ZN(n21946) );
  OAI211_X1 U23543 ( .C1(n21948), .C2(n21947), .A(n22002), .B(n21946), .ZN(
        n22321) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22321), .B1(
        n22320), .B2(n22059), .ZN(n21949) );
  OAI211_X1 U23545 ( .C1(n22324), .C2(n22069), .A(n21950), .B(n21949), .ZN(
        P1_U3049) );
  INV_X1 U23546 ( .A(n21951), .ZN(n21959) );
  OAI21_X1 U23547 ( .B1(n21953), .B2(n21952), .A(n22077), .ZN(n21962) );
  OR2_X1 U23548 ( .A1(n21954), .A2(n22064), .ZN(n21955) );
  OR2_X1 U23549 ( .A1(n22029), .A2(n21959), .ZN(n22325) );
  AND2_X1 U23550 ( .A1(n21955), .A2(n22325), .ZN(n21958) );
  OAI22_X1 U23551 ( .A1(n13234), .A2(n21959), .B1(n21962), .B2(n21958), .ZN(
        n21956) );
  OAI22_X1 U23552 ( .A1(n22326), .A2(n22062), .B1(n22070), .B2(n22325), .ZN(
        n21957) );
  INV_X1 U23553 ( .A(n21957), .ZN(n21964) );
  INV_X1 U23554 ( .A(n21958), .ZN(n21961) );
  AOI21_X1 U23555 ( .B1(n22043), .B2(n21959), .A(n22072), .ZN(n21960) );
  OAI21_X1 U23556 ( .B1(n21962), .B2(n21961), .A(n21960), .ZN(n22329) );
  AOI22_X1 U23557 ( .A1(n22329), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n22059), .B2(n22328), .ZN(n21963) );
  OAI211_X1 U23558 ( .C1(n22332), .C2(n22069), .A(n21964), .B(n21963), .ZN(
        P1_U3057) );
  NOR2_X1 U23559 ( .A1(n22336), .A2(n22043), .ZN(n21965) );
  AOI21_X1 U23560 ( .B1(n21965), .B2(n22334), .A(n22013), .ZN(n21974) );
  INV_X1 U23561 ( .A(n21974), .ZN(n21968) );
  AND2_X1 U23562 ( .A1(n21966), .A2(n22053), .ZN(n21973) );
  INV_X1 U23563 ( .A(n22059), .ZN(n22081) );
  OR3_X1 U23564 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n22067), .ZN(n22333) );
  OAI22_X1 U23565 ( .A1(n22334), .A2(n22081), .B1(n22070), .B2(n22333), .ZN(
        n21969) );
  INV_X1 U23566 ( .A(n21969), .ZN(n21976) );
  INV_X1 U23567 ( .A(n22057), .ZN(n21970) );
  AOI211_X1 U23568 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22333), .A(n21971), 
        .B(n21970), .ZN(n21972) );
  OAI21_X1 U23569 ( .B1(n21974), .B2(n21973), .A(n21972), .ZN(n22337) );
  AOI22_X1 U23570 ( .A1(n22337), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n22078), .B2(n22336), .ZN(n21975) );
  OAI211_X1 U23571 ( .C1(n22340), .C2(n22069), .A(n21976), .B(n21975), .ZN(
        P1_U3081) );
  INV_X1 U23572 ( .A(n21997), .ZN(n21988) );
  NOR3_X1 U23573 ( .A1(n12225), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21992) );
  INV_X1 U23574 ( .A(n21992), .ZN(n21989) );
  NOR2_X1 U23575 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21989), .ZN(
        n22341) );
  AOI21_X1 U23576 ( .B1(n21988), .B2(n14582), .A(n22341), .ZN(n21983) );
  NAND2_X1 U23577 ( .A1(n21980), .A2(n21979), .ZN(n22023) );
  INV_X1 U23578 ( .A(n21999), .ZN(n21981) );
  OAI22_X1 U23579 ( .A1(n21983), .A2(n22043), .B1(n22023), .B2(n21981), .ZN(
        n22342) );
  AOI22_X1 U23580 ( .A1(n22342), .A2(n22048), .B1(n22049), .B2(n22341), .ZN(
        n21987) );
  INV_X1 U23581 ( .A(n22352), .ZN(n21982) );
  OAI21_X1 U23582 ( .B1(n21982), .B2(n22343), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21984) );
  NAND2_X1 U23583 ( .A1(n21984), .A2(n21983), .ZN(n21985) );
  AOI22_X1 U23584 ( .A1(n22344), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n22059), .B2(n22343), .ZN(n21986) );
  OAI211_X1 U23585 ( .C1(n22062), .C2(n22352), .A(n21987), .B(n21986), .ZN(
        P1_U3097) );
  NOR2_X1 U23586 ( .A1(n22029), .A2(n21989), .ZN(n22347) );
  AOI21_X1 U23587 ( .B1(n21988), .B2(n22030), .A(n22347), .ZN(n21990) );
  OAI22_X1 U23588 ( .A1(n21990), .A2(n22043), .B1(n21989), .B2(n13234), .ZN(
        n22348) );
  AOI22_X1 U23589 ( .A1(n22348), .A2(n22048), .B1(n22049), .B2(n22347), .ZN(
        n21995) );
  OAI21_X1 U23590 ( .B1(n21993), .B2(n22050), .A(n21990), .ZN(n21991) );
  OAI221_X1 U23591 ( .B1(n22077), .B2(n21992), .C1(n22043), .C2(n21991), .A(
        n22035), .ZN(n22349) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22349), .B1(
        n22355), .B2(n22078), .ZN(n21994) );
  OAI211_X1 U23593 ( .C1(n22081), .C2(n22352), .A(n21995), .B(n21994), .ZN(
        P1_U3105) );
  NOR3_X1 U23594 ( .A1(n22355), .A2(n22354), .A3(n22043), .ZN(n21996) );
  NOR2_X1 U23595 ( .A1(n21996), .A2(n22013), .ZN(n22009) );
  INV_X1 U23596 ( .A(n22009), .ZN(n22000) );
  NOR2_X1 U23597 ( .A1(n21997), .A2(n14582), .ZN(n22008) );
  NAND2_X1 U23598 ( .A1(n21998), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22003) );
  INV_X1 U23599 ( .A(n22003), .ZN(n22045) );
  NAND2_X1 U23600 ( .A1(n22029), .A2(n22001), .ZN(n22006) );
  INV_X1 U23601 ( .A(n22006), .ZN(n22353) );
  AOI22_X1 U23602 ( .A1(n22355), .A2(n22059), .B1(n22049), .B2(n22353), .ZN(
        n22011) );
  INV_X1 U23603 ( .A(n22002), .ZN(n22005) );
  NAND2_X1 U23604 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22003), .ZN(n22056) );
  INV_X1 U23605 ( .A(n22056), .ZN(n22004) );
  AOI211_X1 U23606 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22006), .A(n22005), 
        .B(n22004), .ZN(n22007) );
  AOI22_X1 U23607 ( .A1(n22356), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n22078), .B2(n22354), .ZN(n22010) );
  OAI211_X1 U23608 ( .C1(n22359), .C2(n22069), .A(n22011), .B(n22010), .ZN(
        P1_U3113) );
  NOR2_X1 U23609 ( .A1(n22362), .A2(n22043), .ZN(n22014) );
  AOI21_X1 U23610 ( .B1(n22014), .B2(n22372), .A(n22013), .ZN(n22026) );
  INV_X1 U23611 ( .A(n22026), .ZN(n22017) );
  OR2_X1 U23612 ( .A1(n14536), .A2(n22015), .ZN(n22065) );
  NOR2_X1 U23613 ( .A1(n22065), .A2(n22053), .ZN(n22025) );
  INV_X1 U23614 ( .A(n22023), .ZN(n22016) );
  NOR3_X1 U23615 ( .A1(n22018), .A2(n12225), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22036) );
  INV_X1 U23616 ( .A(n22036), .ZN(n22031) );
  NOR2_X1 U23617 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22031), .ZN(
        n22020) );
  INV_X1 U23618 ( .A(n22020), .ZN(n22360) );
  OAI22_X1 U23619 ( .A1(n22372), .A2(n22062), .B1(n22070), .B2(n22360), .ZN(
        n22019) );
  INV_X1 U23620 ( .A(n22019), .ZN(n22028) );
  OAI21_X1 U23621 ( .B1(n22021), .B2(n22020), .A(n22057), .ZN(n22022) );
  AOI21_X1 U23622 ( .B1(n22023), .B2(P1_STATE2_REG_2__SCAN_IN), .A(n22022), 
        .ZN(n22024) );
  OAI21_X1 U23623 ( .B1(n22026), .B2(n22025), .A(n22024), .ZN(n22363) );
  AOI22_X1 U23624 ( .A1(n22363), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n22059), .B2(n22362), .ZN(n22027) );
  OAI211_X1 U23625 ( .C1(n22366), .C2(n22069), .A(n22028), .B(n22027), .ZN(
        P1_U3129) );
  NOR2_X1 U23626 ( .A1(n22029), .A2(n22031), .ZN(n22368) );
  INV_X1 U23627 ( .A(n22065), .ZN(n22054) );
  AOI21_X1 U23628 ( .B1(n22054), .B2(n22030), .A(n22368), .ZN(n22032) );
  OAI22_X1 U23629 ( .A1(n22032), .A2(n22043), .B1(n22031), .B2(n13234), .ZN(
        n22367) );
  AOI22_X1 U23630 ( .A1(n22049), .A2(n22368), .B1(n22367), .B2(n22048), .ZN(
        n22040) );
  INV_X1 U23631 ( .A(n22042), .ZN(n22033) );
  OAI211_X1 U23632 ( .C1(n22033), .C2(n22050), .A(n22077), .B(n22032), .ZN(
        n22034) );
  OAI211_X1 U23633 ( .C1(n22077), .C2(n22036), .A(n22035), .B(n22034), .ZN(
        n22369) );
  INV_X1 U23634 ( .A(n22037), .ZN(n22038) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22369), .B1(
        n22378), .B2(n22078), .ZN(n22039) );
  OAI211_X1 U23636 ( .C1(n22081), .C2(n22372), .A(n22040), .B(n22039), .ZN(
        P1_U3137) );
  NOR3_X2 U23637 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12225), .A3(
        n22067), .ZN(n22375) );
  OR2_X1 U23638 ( .A1(n14582), .A2(n22043), .ZN(n22047) );
  NAND2_X1 U23639 ( .A1(n22045), .A2(n22044), .ZN(n22046) );
  OAI21_X1 U23640 ( .B1(n22065), .B2(n22047), .A(n22046), .ZN(n22373) );
  AOI22_X1 U23641 ( .A1(n22049), .A2(n22375), .B1(n22048), .B2(n22373), .ZN(
        n22061) );
  INV_X1 U23642 ( .A(n22378), .ZN(n22051) );
  AOI21_X1 U23643 ( .B1(n22051), .B2(n22393), .A(n22050), .ZN(n22052) );
  AOI21_X1 U23644 ( .B1(n22054), .B2(n22053), .A(n22052), .ZN(n22055) );
  NOR2_X1 U23645 ( .A1(n22055), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22058) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22059), .ZN(n22060) );
  OAI211_X1 U23647 ( .C1(n22062), .C2(n22393), .A(n22061), .B(n22060), .ZN(
        P1_U3145) );
  NAND2_X1 U23648 ( .A1(n22063), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22385) );
  OAI21_X1 U23649 ( .B1(n22065), .B2(n22064), .A(n22385), .ZN(n22066) );
  NAND2_X1 U23650 ( .A1(n22066), .A2(n22077), .ZN(n22073) );
  NOR2_X1 U23651 ( .A1(n12225), .A2(n22067), .ZN(n22076) );
  NAND2_X1 U23652 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22076), .ZN(n22068) );
  AND2_X1 U23653 ( .A1(n22073), .A2(n22068), .ZN(n22384) );
  OAI22_X1 U23654 ( .A1(n22070), .A2(n22385), .B1(n22384), .B2(n22069), .ZN(
        n22071) );
  INV_X1 U23655 ( .A(n22071), .ZN(n22080) );
  AOI21_X1 U23656 ( .B1(n22074), .B2(n22073), .A(n22072), .ZN(n22075) );
  OAI21_X1 U23657 ( .B1(n22077), .B2(n22076), .A(n22075), .ZN(n22390) );
  AOI22_X1 U23658 ( .A1(n22390), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n22078), .B2(n22389), .ZN(n22079) );
  OAI211_X1 U23659 ( .C1(n22081), .C2(n22393), .A(n22080), .B(n22079), .ZN(
        P1_U3153) );
  AOI22_X1 U23660 ( .A1(n22389), .A2(n22108), .B1(n22107), .B2(n22305), .ZN(
        n22083) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22306), .B1(
        n22312), .B2(n22115), .ZN(n22082) );
  OAI211_X1 U23662 ( .C1(n22309), .C2(n22112), .A(n22083), .B(n22082), .ZN(
        P1_U3034) );
  AOI22_X1 U23663 ( .A1(n22311), .A2(n22106), .B1(n22107), .B2(n22310), .ZN(
        n22085) );
  AOI22_X1 U23664 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22108), .ZN(n22084) );
  OAI211_X1 U23665 ( .C1(n22111), .C2(n22316), .A(n22085), .B(n22084), .ZN(
        P1_U3042) );
  OAI22_X1 U23666 ( .A1(n22316), .A2(n22118), .B1(n22113), .B2(n22317), .ZN(
        n22086) );
  INV_X1 U23667 ( .A(n22086), .ZN(n22088) );
  AOI22_X1 U23668 ( .A1(n22321), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n22115), .B2(n22328), .ZN(n22087) );
  OAI211_X1 U23669 ( .C1(n22324), .C2(n22112), .A(n22088), .B(n22087), .ZN(
        P1_U3050) );
  OAI22_X1 U23670 ( .A1(n22326), .A2(n22111), .B1(n22113), .B2(n22325), .ZN(
        n22089) );
  INV_X1 U23671 ( .A(n22089), .ZN(n22091) );
  AOI22_X1 U23672 ( .A1(n22329), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n22108), .B2(n22328), .ZN(n22090) );
  OAI211_X1 U23673 ( .C1(n22332), .C2(n22112), .A(n22091), .B(n22090), .ZN(
        P1_U3058) );
  OAI22_X1 U23674 ( .A1(n22334), .A2(n22118), .B1(n22113), .B2(n22333), .ZN(
        n22092) );
  INV_X1 U23675 ( .A(n22092), .ZN(n22094) );
  AOI22_X1 U23676 ( .A1(n22337), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n22115), .B2(n22336), .ZN(n22093) );
  OAI211_X1 U23677 ( .C1(n22340), .C2(n22112), .A(n22094), .B(n22093), .ZN(
        P1_U3082) );
  AOI22_X1 U23678 ( .A1(n22342), .A2(n22106), .B1(n22107), .B2(n22341), .ZN(
        n22096) );
  AOI22_X1 U23679 ( .A1(n22344), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n22108), .B2(n22343), .ZN(n22095) );
  OAI211_X1 U23680 ( .C1(n22111), .C2(n22352), .A(n22096), .B(n22095), .ZN(
        P1_U3098) );
  AOI22_X1 U23681 ( .A1(n22348), .A2(n22106), .B1(n22107), .B2(n22347), .ZN(
        n22098) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22349), .B1(
        n22355), .B2(n22115), .ZN(n22097) );
  OAI211_X1 U23683 ( .C1(n22118), .C2(n22352), .A(n22098), .B(n22097), .ZN(
        P1_U3106) );
  AOI22_X1 U23684 ( .A1(n22354), .A2(n22115), .B1(n22107), .B2(n22353), .ZN(
        n22100) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22356), .B1(
        n22355), .B2(n22108), .ZN(n22099) );
  OAI211_X1 U23686 ( .C1(n22359), .C2(n22112), .A(n22100), .B(n22099), .ZN(
        P1_U3114) );
  OAI22_X1 U23687 ( .A1(n22372), .A2(n22111), .B1(n22113), .B2(n22360), .ZN(
        n22101) );
  INV_X1 U23688 ( .A(n22101), .ZN(n22103) );
  AOI22_X1 U23689 ( .A1(n22363), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n22108), .B2(n22362), .ZN(n22102) );
  OAI211_X1 U23690 ( .C1(n22366), .C2(n22112), .A(n22103), .B(n22102), .ZN(
        P1_U3130) );
  AOI22_X1 U23691 ( .A1(n22107), .A2(n22368), .B1(n22367), .B2(n22106), .ZN(
        n22105) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22369), .B1(
        n22378), .B2(n22115), .ZN(n22104) );
  OAI211_X1 U23693 ( .C1(n22118), .C2(n22372), .A(n22105), .B(n22104), .ZN(
        P1_U3138) );
  AOI22_X1 U23694 ( .A1(n22107), .A2(n22375), .B1(n22106), .B2(n22373), .ZN(
        n22110) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22108), .ZN(n22109) );
  OAI211_X1 U23696 ( .C1(n22111), .C2(n22393), .A(n22110), .B(n22109), .ZN(
        P1_U3146) );
  OAI22_X1 U23697 ( .A1(n22113), .A2(n22385), .B1(n22384), .B2(n22112), .ZN(
        n22114) );
  INV_X1 U23698 ( .A(n22114), .ZN(n22117) );
  AOI22_X1 U23699 ( .A1(n22390), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n22389), .B2(n22115), .ZN(n22116) );
  OAI211_X1 U23700 ( .C1(n22118), .C2(n22393), .A(n22117), .B(n22116), .ZN(
        P1_U3154) );
  AOI22_X1 U23701 ( .A1(n22389), .A2(n22145), .B1(n22144), .B2(n22305), .ZN(
        n22120) );
  AOI22_X1 U23702 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22306), .B1(
        n22312), .B2(n22152), .ZN(n22119) );
  OAI211_X1 U23703 ( .C1(n22309), .C2(n22149), .A(n22120), .B(n22119), .ZN(
        P1_U3035) );
  AOI22_X1 U23704 ( .A1(n22311), .A2(n22143), .B1(n22144), .B2(n22310), .ZN(
        n22122) );
  AOI22_X1 U23705 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22145), .ZN(n22121) );
  OAI211_X1 U23706 ( .C1(n22148), .C2(n22316), .A(n22122), .B(n22121), .ZN(
        P1_U3043) );
  OAI22_X1 U23707 ( .A1(n22316), .A2(n22155), .B1(n22150), .B2(n22317), .ZN(
        n22123) );
  INV_X1 U23708 ( .A(n22123), .ZN(n22125) );
  AOI22_X1 U23709 ( .A1(n22321), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n22152), .B2(n22328), .ZN(n22124) );
  OAI211_X1 U23710 ( .C1(n22324), .C2(n22149), .A(n22125), .B(n22124), .ZN(
        P1_U3051) );
  OAI22_X1 U23711 ( .A1(n22318), .A2(n22155), .B1(n22150), .B2(n22325), .ZN(
        n22126) );
  INV_X1 U23712 ( .A(n22126), .ZN(n22128) );
  AOI22_X1 U23713 ( .A1(n22329), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n22152), .B2(n22201), .ZN(n22127) );
  OAI211_X1 U23714 ( .C1(n22332), .C2(n22149), .A(n22128), .B(n22127), .ZN(
        P1_U3059) );
  OAI22_X1 U23715 ( .A1(n22334), .A2(n22155), .B1(n22150), .B2(n22333), .ZN(
        n22129) );
  INV_X1 U23716 ( .A(n22129), .ZN(n22131) );
  AOI22_X1 U23717 ( .A1(n22337), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22152), .B2(n22336), .ZN(n22130) );
  OAI211_X1 U23718 ( .C1(n22340), .C2(n22149), .A(n22131), .B(n22130), .ZN(
        P1_U3083) );
  AOI22_X1 U23719 ( .A1(n22342), .A2(n22143), .B1(n22144), .B2(n22341), .ZN(
        n22133) );
  AOI22_X1 U23720 ( .A1(n22344), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n22145), .B2(n22343), .ZN(n22132) );
  OAI211_X1 U23721 ( .C1(n22148), .C2(n22352), .A(n22133), .B(n22132), .ZN(
        P1_U3099) );
  AOI22_X1 U23722 ( .A1(n22348), .A2(n22143), .B1(n22144), .B2(n22347), .ZN(
        n22135) );
  AOI22_X1 U23723 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22349), .B1(
        n22355), .B2(n22152), .ZN(n22134) );
  OAI211_X1 U23724 ( .C1(n22155), .C2(n22352), .A(n22135), .B(n22134), .ZN(
        P1_U3107) );
  AOI22_X1 U23725 ( .A1(n22355), .A2(n22145), .B1(n22144), .B2(n22353), .ZN(
        n22137) );
  AOI22_X1 U23726 ( .A1(n22356), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n22152), .B2(n22354), .ZN(n22136) );
  OAI211_X1 U23727 ( .C1(n22359), .C2(n22149), .A(n22137), .B(n22136), .ZN(
        P1_U3115) );
  OAI22_X1 U23728 ( .A1(n22372), .A2(n22148), .B1(n22150), .B2(n22360), .ZN(
        n22138) );
  INV_X1 U23729 ( .A(n22138), .ZN(n22140) );
  AOI22_X1 U23730 ( .A1(n22363), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22145), .B2(n22362), .ZN(n22139) );
  OAI211_X1 U23731 ( .C1(n22366), .C2(n22149), .A(n22140), .B(n22139), .ZN(
        P1_U3131) );
  AOI22_X1 U23732 ( .A1(n22144), .A2(n22368), .B1(n22367), .B2(n22143), .ZN(
        n22142) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22369), .B1(
        n22378), .B2(n22152), .ZN(n22141) );
  OAI211_X1 U23734 ( .C1(n22155), .C2(n22372), .A(n22142), .B(n22141), .ZN(
        P1_U3139) );
  AOI22_X1 U23735 ( .A1(n22144), .A2(n22375), .B1(n22143), .B2(n22373), .ZN(
        n22147) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22145), .ZN(n22146) );
  OAI211_X1 U23737 ( .C1(n22148), .C2(n22393), .A(n22147), .B(n22146), .ZN(
        P1_U3147) );
  OAI22_X1 U23738 ( .A1(n22150), .A2(n22385), .B1(n22384), .B2(n22149), .ZN(
        n22151) );
  INV_X1 U23739 ( .A(n22151), .ZN(n22154) );
  AOI22_X1 U23740 ( .A1(n22390), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n22389), .B2(n22152), .ZN(n22153) );
  OAI211_X1 U23741 ( .C1(n22155), .C2(n22393), .A(n22154), .B(n22153), .ZN(
        P1_U3155) );
  AOI22_X1 U23742 ( .A1(n22389), .A2(n22182), .B1(n22181), .B2(n22305), .ZN(
        n22157) );
  AOI22_X1 U23743 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22306), .B1(
        n22312), .B2(n22189), .ZN(n22156) );
  OAI211_X1 U23744 ( .C1(n22309), .C2(n22186), .A(n22157), .B(n22156), .ZN(
        P1_U3036) );
  AOI22_X1 U23745 ( .A1(n22311), .A2(n22180), .B1(n22181), .B2(n22310), .ZN(
        n22159) );
  AOI22_X1 U23746 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22182), .ZN(n22158) );
  OAI211_X1 U23747 ( .C1(n22185), .C2(n22316), .A(n22159), .B(n22158), .ZN(
        P1_U3044) );
  OAI22_X1 U23748 ( .A1(n22318), .A2(n22185), .B1(n22187), .B2(n22317), .ZN(
        n22160) );
  INV_X1 U23749 ( .A(n22160), .ZN(n22162) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22321), .B1(
        n22320), .B2(n22182), .ZN(n22161) );
  OAI211_X1 U23751 ( .C1(n22324), .C2(n22186), .A(n22162), .B(n22161), .ZN(
        P1_U3052) );
  OAI22_X1 U23752 ( .A1(n22326), .A2(n22185), .B1(n22187), .B2(n22325), .ZN(
        n22163) );
  INV_X1 U23753 ( .A(n22163), .ZN(n22165) );
  AOI22_X1 U23754 ( .A1(n22329), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22182), .B2(n22328), .ZN(n22164) );
  OAI211_X1 U23755 ( .C1(n22332), .C2(n22186), .A(n22165), .B(n22164), .ZN(
        P1_U3060) );
  OAI22_X1 U23756 ( .A1(n22334), .A2(n22192), .B1(n22187), .B2(n22333), .ZN(
        n22166) );
  INV_X1 U23757 ( .A(n22166), .ZN(n22168) );
  AOI22_X1 U23758 ( .A1(n22337), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22189), .B2(n22336), .ZN(n22167) );
  OAI211_X1 U23759 ( .C1(n22340), .C2(n22186), .A(n22168), .B(n22167), .ZN(
        P1_U3084) );
  AOI22_X1 U23760 ( .A1(n22342), .A2(n22180), .B1(n22181), .B2(n22341), .ZN(
        n22170) );
  AOI22_X1 U23761 ( .A1(n22344), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n22182), .B2(n22343), .ZN(n22169) );
  OAI211_X1 U23762 ( .C1(n22185), .C2(n22352), .A(n22170), .B(n22169), .ZN(
        P1_U3100) );
  AOI22_X1 U23763 ( .A1(n22348), .A2(n22180), .B1(n22181), .B2(n22347), .ZN(
        n22172) );
  AOI22_X1 U23764 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22349), .B1(
        n22355), .B2(n22189), .ZN(n22171) );
  OAI211_X1 U23765 ( .C1(n22192), .C2(n22352), .A(n22172), .B(n22171), .ZN(
        P1_U3108) );
  AOI22_X1 U23766 ( .A1(n22354), .A2(n22189), .B1(n22181), .B2(n22353), .ZN(
        n22174) );
  AOI22_X1 U23767 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22356), .B1(
        n22355), .B2(n22182), .ZN(n22173) );
  OAI211_X1 U23768 ( .C1(n22359), .C2(n22186), .A(n22174), .B(n22173), .ZN(
        P1_U3116) );
  OAI22_X1 U23769 ( .A1(n22372), .A2(n22185), .B1(n22187), .B2(n22360), .ZN(
        n22175) );
  INV_X1 U23770 ( .A(n22175), .ZN(n22177) );
  AOI22_X1 U23771 ( .A1(n22363), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22182), .B2(n22362), .ZN(n22176) );
  OAI211_X1 U23772 ( .C1(n22366), .C2(n22186), .A(n22177), .B(n22176), .ZN(
        P1_U3132) );
  AOI22_X1 U23773 ( .A1(n22181), .A2(n22368), .B1(n22367), .B2(n22180), .ZN(
        n22179) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22369), .B1(
        n22378), .B2(n22189), .ZN(n22178) );
  OAI211_X1 U23775 ( .C1(n22192), .C2(n22372), .A(n22179), .B(n22178), .ZN(
        P1_U3140) );
  AOI22_X1 U23776 ( .A1(n22181), .A2(n22375), .B1(n22180), .B2(n22373), .ZN(
        n22184) );
  AOI22_X1 U23777 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22182), .ZN(n22183) );
  OAI211_X1 U23778 ( .C1(n22185), .C2(n22393), .A(n22184), .B(n22183), .ZN(
        P1_U3148) );
  OAI22_X1 U23779 ( .A1(n22187), .A2(n22385), .B1(n22384), .B2(n22186), .ZN(
        n22188) );
  INV_X1 U23780 ( .A(n22188), .ZN(n22191) );
  AOI22_X1 U23781 ( .A1(n22390), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n22389), .B2(n22189), .ZN(n22190) );
  OAI211_X1 U23782 ( .C1(n22192), .C2(n22393), .A(n22191), .B(n22190), .ZN(
        P1_U3156) );
  AOI22_X1 U23783 ( .A1(n22389), .A2(n22220), .B1(n22219), .B2(n22305), .ZN(
        n22194) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22306), .B1(
        n22312), .B2(n22227), .ZN(n22193) );
  OAI211_X1 U23785 ( .C1(n22309), .C2(n22224), .A(n22194), .B(n22193), .ZN(
        P1_U3037) );
  AOI22_X1 U23786 ( .A1(n22311), .A2(n22218), .B1(n22219), .B2(n22310), .ZN(
        n22196) );
  AOI22_X1 U23787 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22220), .ZN(n22195) );
  OAI211_X1 U23788 ( .C1(n22223), .C2(n22316), .A(n22196), .B(n22195), .ZN(
        P1_U3045) );
  OAI22_X1 U23789 ( .A1(n22318), .A2(n22223), .B1(n22225), .B2(n22317), .ZN(
        n22197) );
  INV_X1 U23790 ( .A(n22197), .ZN(n22199) );
  AOI22_X1 U23791 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22321), .B1(
        n22320), .B2(n22220), .ZN(n22198) );
  OAI211_X1 U23792 ( .C1(n22324), .C2(n22224), .A(n22199), .B(n22198), .ZN(
        P1_U3053) );
  OAI22_X1 U23793 ( .A1(n22318), .A2(n22230), .B1(n22225), .B2(n22325), .ZN(
        n22200) );
  INV_X1 U23794 ( .A(n22200), .ZN(n22203) );
  AOI22_X1 U23795 ( .A1(n22329), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22227), .B2(n22201), .ZN(n22202) );
  OAI211_X1 U23796 ( .C1(n22332), .C2(n22224), .A(n22203), .B(n22202), .ZN(
        P1_U3061) );
  OAI22_X1 U23797 ( .A1(n22334), .A2(n22230), .B1(n22225), .B2(n22333), .ZN(
        n22204) );
  INV_X1 U23798 ( .A(n22204), .ZN(n22206) );
  AOI22_X1 U23799 ( .A1(n22337), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22227), .B2(n22336), .ZN(n22205) );
  OAI211_X1 U23800 ( .C1(n22340), .C2(n22224), .A(n22206), .B(n22205), .ZN(
        P1_U3085) );
  AOI22_X1 U23801 ( .A1(n22342), .A2(n22218), .B1(n22219), .B2(n22341), .ZN(
        n22208) );
  AOI22_X1 U23802 ( .A1(n22344), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n22220), .B2(n22343), .ZN(n22207) );
  OAI211_X1 U23803 ( .C1(n22223), .C2(n22352), .A(n22208), .B(n22207), .ZN(
        P1_U3101) );
  AOI22_X1 U23804 ( .A1(n22348), .A2(n22218), .B1(n22219), .B2(n22347), .ZN(
        n22210) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22349), .B1(
        n22355), .B2(n22227), .ZN(n22209) );
  OAI211_X1 U23806 ( .C1(n22230), .C2(n22352), .A(n22210), .B(n22209), .ZN(
        P1_U3109) );
  AOI22_X1 U23807 ( .A1(n22355), .A2(n22220), .B1(n22219), .B2(n22353), .ZN(
        n22212) );
  AOI22_X1 U23808 ( .A1(n22356), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n22227), .B2(n22354), .ZN(n22211) );
  OAI211_X1 U23809 ( .C1(n22359), .C2(n22224), .A(n22212), .B(n22211), .ZN(
        P1_U3117) );
  OAI22_X1 U23810 ( .A1(n22372), .A2(n22223), .B1(n22225), .B2(n22360), .ZN(
        n22213) );
  INV_X1 U23811 ( .A(n22213), .ZN(n22215) );
  AOI22_X1 U23812 ( .A1(n22363), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n22220), .B2(n22362), .ZN(n22214) );
  OAI211_X1 U23813 ( .C1(n22366), .C2(n22224), .A(n22215), .B(n22214), .ZN(
        P1_U3133) );
  AOI22_X1 U23814 ( .A1(n22219), .A2(n22368), .B1(n22367), .B2(n22218), .ZN(
        n22217) );
  AOI22_X1 U23815 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22369), .B1(
        n22378), .B2(n22227), .ZN(n22216) );
  OAI211_X1 U23816 ( .C1(n22230), .C2(n22372), .A(n22217), .B(n22216), .ZN(
        P1_U3141) );
  AOI22_X1 U23817 ( .A1(n22219), .A2(n22375), .B1(n22218), .B2(n22373), .ZN(
        n22222) );
  AOI22_X1 U23818 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22220), .ZN(n22221) );
  OAI211_X1 U23819 ( .C1(n22223), .C2(n22393), .A(n22222), .B(n22221), .ZN(
        P1_U3149) );
  OAI22_X1 U23820 ( .A1(n22225), .A2(n22385), .B1(n22384), .B2(n22224), .ZN(
        n22226) );
  INV_X1 U23821 ( .A(n22226), .ZN(n22229) );
  AOI22_X1 U23822 ( .A1(n22390), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n22389), .B2(n22227), .ZN(n22228) );
  OAI211_X1 U23823 ( .C1(n22230), .C2(n22393), .A(n22229), .B(n22228), .ZN(
        P1_U3157) );
  AOI22_X1 U23824 ( .A1(n22389), .A2(n22257), .B1(n22256), .B2(n22305), .ZN(
        n22232) );
  AOI22_X1 U23825 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22306), .B1(
        n22312), .B2(n22264), .ZN(n22231) );
  OAI211_X1 U23826 ( .C1(n22309), .C2(n22261), .A(n22232), .B(n22231), .ZN(
        P1_U3038) );
  AOI22_X1 U23827 ( .A1(n22311), .A2(n22255), .B1(n22256), .B2(n22310), .ZN(
        n22234) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22257), .ZN(n22233) );
  OAI211_X1 U23829 ( .C1(n22260), .C2(n22316), .A(n22234), .B(n22233), .ZN(
        P1_U3046) );
  OAI22_X1 U23830 ( .A1(n22318), .A2(n22260), .B1(n22262), .B2(n22317), .ZN(
        n22235) );
  INV_X1 U23831 ( .A(n22235), .ZN(n22237) );
  AOI22_X1 U23832 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22321), .B1(
        n22320), .B2(n22257), .ZN(n22236) );
  OAI211_X1 U23833 ( .C1(n22324), .C2(n22261), .A(n22237), .B(n22236), .ZN(
        P1_U3054) );
  OAI22_X1 U23834 ( .A1(n22326), .A2(n22260), .B1(n22262), .B2(n22325), .ZN(
        n22238) );
  INV_X1 U23835 ( .A(n22238), .ZN(n22240) );
  AOI22_X1 U23836 ( .A1(n22329), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22257), .B2(n22328), .ZN(n22239) );
  OAI211_X1 U23837 ( .C1(n22332), .C2(n22261), .A(n22240), .B(n22239), .ZN(
        P1_U3062) );
  OAI22_X1 U23838 ( .A1(n22334), .A2(n22267), .B1(n22262), .B2(n22333), .ZN(
        n22241) );
  INV_X1 U23839 ( .A(n22241), .ZN(n22243) );
  AOI22_X1 U23840 ( .A1(n22337), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22264), .B2(n22336), .ZN(n22242) );
  OAI211_X1 U23841 ( .C1(n22340), .C2(n22261), .A(n22243), .B(n22242), .ZN(
        P1_U3086) );
  AOI22_X1 U23842 ( .A1(n22342), .A2(n22255), .B1(n22256), .B2(n22341), .ZN(
        n22245) );
  AOI22_X1 U23843 ( .A1(n22344), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n22257), .B2(n22343), .ZN(n22244) );
  OAI211_X1 U23844 ( .C1(n22260), .C2(n22352), .A(n22245), .B(n22244), .ZN(
        P1_U3102) );
  AOI22_X1 U23845 ( .A1(n22348), .A2(n22255), .B1(n22256), .B2(n22347), .ZN(
        n22247) );
  AOI22_X1 U23846 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22349), .B1(
        n22355), .B2(n22264), .ZN(n22246) );
  OAI211_X1 U23847 ( .C1(n22267), .C2(n22352), .A(n22247), .B(n22246), .ZN(
        P1_U3110) );
  AOI22_X1 U23848 ( .A1(n22354), .A2(n22264), .B1(n22256), .B2(n22353), .ZN(
        n22249) );
  AOI22_X1 U23849 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22356), .B1(
        n22355), .B2(n22257), .ZN(n22248) );
  OAI211_X1 U23850 ( .C1(n22359), .C2(n22261), .A(n22249), .B(n22248), .ZN(
        P1_U3118) );
  OAI22_X1 U23851 ( .A1(n22372), .A2(n22260), .B1(n22262), .B2(n22360), .ZN(
        n22250) );
  INV_X1 U23852 ( .A(n22250), .ZN(n22252) );
  AOI22_X1 U23853 ( .A1(n22363), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22257), .B2(n22362), .ZN(n22251) );
  OAI211_X1 U23854 ( .C1(n22366), .C2(n22261), .A(n22252), .B(n22251), .ZN(
        P1_U3134) );
  AOI22_X1 U23855 ( .A1(n22256), .A2(n22368), .B1(n22367), .B2(n22255), .ZN(
        n22254) );
  AOI22_X1 U23856 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22369), .B1(
        n22378), .B2(n22264), .ZN(n22253) );
  OAI211_X1 U23857 ( .C1(n22267), .C2(n22372), .A(n22254), .B(n22253), .ZN(
        P1_U3142) );
  AOI22_X1 U23858 ( .A1(n22256), .A2(n22375), .B1(n22255), .B2(n22373), .ZN(
        n22259) );
  AOI22_X1 U23859 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22257), .ZN(n22258) );
  OAI211_X1 U23860 ( .C1(n22260), .C2(n22393), .A(n22259), .B(n22258), .ZN(
        P1_U3150) );
  OAI22_X1 U23861 ( .A1(n22262), .A2(n22385), .B1(n22384), .B2(n22261), .ZN(
        n22263) );
  INV_X1 U23862 ( .A(n22263), .ZN(n22266) );
  AOI22_X1 U23863 ( .A1(n22390), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n22389), .B2(n22264), .ZN(n22265) );
  OAI211_X1 U23864 ( .C1(n22267), .C2(n22393), .A(n22266), .B(n22265), .ZN(
        P1_U3158) );
  AOI22_X1 U23865 ( .A1(n22389), .A2(n22294), .B1(n22293), .B2(n22305), .ZN(
        n22269) );
  AOI22_X1 U23866 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22306), .B1(
        n22312), .B2(n22301), .ZN(n22268) );
  OAI211_X1 U23867 ( .C1(n22309), .C2(n22298), .A(n22269), .B(n22268), .ZN(
        P1_U3039) );
  AOI22_X1 U23868 ( .A1(n22311), .A2(n22292), .B1(n22293), .B2(n22310), .ZN(
        n22271) );
  AOI22_X1 U23869 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22294), .ZN(n22270) );
  OAI211_X1 U23870 ( .C1(n22297), .C2(n22316), .A(n22271), .B(n22270), .ZN(
        P1_U3047) );
  OAI22_X1 U23871 ( .A1(n22318), .A2(n22297), .B1(n22299), .B2(n22317), .ZN(
        n22272) );
  INV_X1 U23872 ( .A(n22272), .ZN(n22274) );
  AOI22_X1 U23873 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22321), .B1(
        n22320), .B2(n22294), .ZN(n22273) );
  OAI211_X1 U23874 ( .C1(n22324), .C2(n22298), .A(n22274), .B(n22273), .ZN(
        P1_U3055) );
  OAI22_X1 U23875 ( .A1(n22326), .A2(n22297), .B1(n22299), .B2(n22325), .ZN(
        n22275) );
  INV_X1 U23876 ( .A(n22275), .ZN(n22277) );
  AOI22_X1 U23877 ( .A1(n22329), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22294), .B2(n22328), .ZN(n22276) );
  OAI211_X1 U23878 ( .C1(n22332), .C2(n22298), .A(n22277), .B(n22276), .ZN(
        P1_U3063) );
  OAI22_X1 U23879 ( .A1(n22334), .A2(n22304), .B1(n22299), .B2(n22333), .ZN(
        n22278) );
  INV_X1 U23880 ( .A(n22278), .ZN(n22280) );
  AOI22_X1 U23881 ( .A1(n22337), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22301), .B2(n22336), .ZN(n22279) );
  OAI211_X1 U23882 ( .C1(n22340), .C2(n22298), .A(n22280), .B(n22279), .ZN(
        P1_U3087) );
  AOI22_X1 U23883 ( .A1(n22342), .A2(n22292), .B1(n22293), .B2(n22341), .ZN(
        n22282) );
  AOI22_X1 U23884 ( .A1(n22344), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n22294), .B2(n22343), .ZN(n22281) );
  OAI211_X1 U23885 ( .C1(n22297), .C2(n22352), .A(n22282), .B(n22281), .ZN(
        P1_U3103) );
  AOI22_X1 U23886 ( .A1(n22348), .A2(n22292), .B1(n22293), .B2(n22347), .ZN(
        n22284) );
  AOI22_X1 U23887 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22349), .B1(
        n22355), .B2(n22301), .ZN(n22283) );
  OAI211_X1 U23888 ( .C1(n22304), .C2(n22352), .A(n22284), .B(n22283), .ZN(
        P1_U3111) );
  AOI22_X1 U23889 ( .A1(n22354), .A2(n22301), .B1(n22293), .B2(n22353), .ZN(
        n22286) );
  AOI22_X1 U23890 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22356), .B1(
        n22355), .B2(n22294), .ZN(n22285) );
  OAI211_X1 U23891 ( .C1(n22359), .C2(n22298), .A(n22286), .B(n22285), .ZN(
        P1_U3119) );
  OAI22_X1 U23892 ( .A1(n22372), .A2(n22297), .B1(n22299), .B2(n22360), .ZN(
        n22287) );
  INV_X1 U23893 ( .A(n22287), .ZN(n22289) );
  AOI22_X1 U23894 ( .A1(n22363), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22294), .B2(n22362), .ZN(n22288) );
  OAI211_X1 U23895 ( .C1(n22366), .C2(n22298), .A(n22289), .B(n22288), .ZN(
        P1_U3135) );
  AOI22_X1 U23896 ( .A1(n22293), .A2(n22368), .B1(n22367), .B2(n22292), .ZN(
        n22291) );
  AOI22_X1 U23897 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22369), .B1(
        n22378), .B2(n22301), .ZN(n22290) );
  OAI211_X1 U23898 ( .C1(n22304), .C2(n22372), .A(n22291), .B(n22290), .ZN(
        P1_U3143) );
  AOI22_X1 U23899 ( .A1(n22293), .A2(n22375), .B1(n22292), .B2(n22373), .ZN(
        n22296) );
  AOI22_X1 U23900 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22294), .ZN(n22295) );
  OAI211_X1 U23901 ( .C1(n22297), .C2(n22393), .A(n22296), .B(n22295), .ZN(
        P1_U3151) );
  OAI22_X1 U23902 ( .A1(n22299), .A2(n22385), .B1(n22384), .B2(n22298), .ZN(
        n22300) );
  INV_X1 U23903 ( .A(n22300), .ZN(n22303) );
  AOI22_X1 U23904 ( .A1(n22390), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n22389), .B2(n22301), .ZN(n22302) );
  OAI211_X1 U23905 ( .C1(n22304), .C2(n22393), .A(n22303), .B(n22302), .ZN(
        P1_U3159) );
  AOI22_X1 U23906 ( .A1(n22389), .A2(n22377), .B1(n22376), .B2(n22305), .ZN(
        n22308) );
  AOI22_X1 U23907 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22306), .B1(
        n22312), .B2(n22388), .ZN(n22307) );
  OAI211_X1 U23908 ( .C1(n22309), .C2(n22383), .A(n22308), .B(n22307), .ZN(
        P1_U3040) );
  AOI22_X1 U23909 ( .A1(n22311), .A2(n22374), .B1(n22376), .B2(n22310), .ZN(
        n22315) );
  AOI22_X1 U23910 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22377), .ZN(n22314) );
  OAI211_X1 U23911 ( .C1(n22382), .C2(n22316), .A(n22315), .B(n22314), .ZN(
        P1_U3048) );
  OAI22_X1 U23912 ( .A1(n22318), .A2(n22382), .B1(n22386), .B2(n22317), .ZN(
        n22319) );
  INV_X1 U23913 ( .A(n22319), .ZN(n22323) );
  AOI22_X1 U23914 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22321), .B1(
        n22320), .B2(n22377), .ZN(n22322) );
  OAI211_X1 U23915 ( .C1(n22324), .C2(n22383), .A(n22323), .B(n22322), .ZN(
        P1_U3056) );
  OAI22_X1 U23916 ( .A1(n22326), .A2(n22382), .B1(n22386), .B2(n22325), .ZN(
        n22327) );
  INV_X1 U23917 ( .A(n22327), .ZN(n22331) );
  AOI22_X1 U23918 ( .A1(n22329), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n22377), .B2(n22328), .ZN(n22330) );
  OAI211_X1 U23919 ( .C1(n22332), .C2(n22383), .A(n22331), .B(n22330), .ZN(
        P1_U3064) );
  OAI22_X1 U23920 ( .A1(n22334), .A2(n22394), .B1(n22386), .B2(n22333), .ZN(
        n22335) );
  INV_X1 U23921 ( .A(n22335), .ZN(n22339) );
  AOI22_X1 U23922 ( .A1(n22337), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22388), .B2(n22336), .ZN(n22338) );
  OAI211_X1 U23923 ( .C1(n22340), .C2(n22383), .A(n22339), .B(n22338), .ZN(
        P1_U3088) );
  AOI22_X1 U23924 ( .A1(n22342), .A2(n22374), .B1(n22376), .B2(n22341), .ZN(
        n22346) );
  AOI22_X1 U23925 ( .A1(n22344), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n22377), .B2(n22343), .ZN(n22345) );
  OAI211_X1 U23926 ( .C1(n22382), .C2(n22352), .A(n22346), .B(n22345), .ZN(
        P1_U3104) );
  AOI22_X1 U23927 ( .A1(n22348), .A2(n22374), .B1(n22376), .B2(n22347), .ZN(
        n22351) );
  AOI22_X1 U23928 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22349), .B1(
        n22355), .B2(n22388), .ZN(n22350) );
  OAI211_X1 U23929 ( .C1(n22394), .C2(n22352), .A(n22351), .B(n22350), .ZN(
        P1_U3112) );
  AOI22_X1 U23930 ( .A1(n22354), .A2(n22388), .B1(n22376), .B2(n22353), .ZN(
        n22358) );
  AOI22_X1 U23931 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22356), .B1(
        n22355), .B2(n22377), .ZN(n22357) );
  OAI211_X1 U23932 ( .C1(n22359), .C2(n22383), .A(n22358), .B(n22357), .ZN(
        P1_U3120) );
  OAI22_X1 U23933 ( .A1(n22372), .A2(n22382), .B1(n22386), .B2(n22360), .ZN(
        n22361) );
  INV_X1 U23934 ( .A(n22361), .ZN(n22365) );
  AOI22_X1 U23935 ( .A1(n22363), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n22377), .B2(n22362), .ZN(n22364) );
  OAI211_X1 U23936 ( .C1(n22366), .C2(n22383), .A(n22365), .B(n22364), .ZN(
        P1_U3136) );
  AOI22_X1 U23937 ( .A1(n22376), .A2(n22368), .B1(n22367), .B2(n22374), .ZN(
        n22371) );
  AOI22_X1 U23938 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22369), .B1(
        n22378), .B2(n22388), .ZN(n22370) );
  OAI211_X1 U23939 ( .C1(n22394), .C2(n22372), .A(n22371), .B(n22370), .ZN(
        P1_U3144) );
  AOI22_X1 U23940 ( .A1(n22376), .A2(n22375), .B1(n22374), .B2(n22373), .ZN(
        n22381) );
  AOI22_X1 U23941 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22379), .B1(
        n22378), .B2(n22377), .ZN(n22380) );
  OAI211_X1 U23942 ( .C1(n22382), .C2(n22393), .A(n22381), .B(n22380), .ZN(
        P1_U3152) );
  OAI22_X1 U23943 ( .A1(n22386), .A2(n22385), .B1(n22384), .B2(n22383), .ZN(
        n22387) );
  INV_X1 U23944 ( .A(n22387), .ZN(n22392) );
  AOI22_X1 U23945 ( .A1(n22390), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n22389), .B2(n22388), .ZN(n22391) );
  OAI211_X1 U23946 ( .C1(n22394), .C2(n22393), .A(n22392), .B(n22391), .ZN(
        P1_U3160) );
  AOI22_X1 U23947 ( .A1(n22398), .A2(n22397), .B1(n22396), .B2(n22395), .ZN(
        P1_U3486) );
  CLKBUF_X1 U11107 ( .A(n13636), .Z(n11032) );
  CLKBUF_X1 U11124 ( .A(n13636), .Z(n11033) );
  CLKBUF_X2 U11126 ( .A(n11997), .Z(n13659) );
  CLKBUF_X1 U11132 ( .A(n12686), .Z(n14468) );
  CLKBUF_X1 U11133 ( .A(n12144), .Z(n11010) );
  CLKBUF_X1 U11135 ( .A(n12803), .Z(n15513) );
  CLKBUF_X1 U11181 ( .A(n11915), .Z(n10985) );
  CLKBUF_X2 U11220 ( .A(n11931), .Z(n11858) );
  CLKBUF_X1 U11242 ( .A(n13298), .Z(n11011) );
  NAND2_X1 U11247 ( .A1(n12201), .A2(n11209), .ZN(n12204) );
  NAND2_X1 U11266 ( .A1(n16613), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16605) );
  CLKBUF_X1 U11470 ( .A(n16612), .Z(n16627) );
  CLKBUF_X2 U11474 ( .A(n16739), .Z(n17034) );
  NOR2_X2 U11486 ( .A1(n18049), .A2(n17989), .ZN(n17988) );
  OR2_X1 U11489 ( .A1(n11879), .A2(n11878), .ZN(n14683) );
  CLKBUF_X1 U11514 ( .A(n15784), .Z(n15785) );
  CLKBUF_X1 U12270 ( .A(n15815), .Z(n15816) );
  CLKBUF_X1 U13701 ( .A(n17530), .Z(n17538) );
endmodule

