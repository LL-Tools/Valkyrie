

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6597, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794;

  AND2_X1 U7178 ( .A1(n9846), .A2(n9845), .ZN(n14816) );
  OR2_X2 U7179 ( .A1(n9840), .A2(n12816), .ZN(n14991) );
  INV_X2 U7180 ( .A(n7046), .ZN(n10281) );
  CLKBUF_X2 U7181 ( .A(n7987), .Z(n12847) );
  CLKBUF_X2 U7182 ( .A(n9612), .Z(n9912) );
  CLKBUF_X2 U7183 ( .A(n8969), .Z(n9068) );
  OAI211_X1 U7184 ( .C1(n11212), .C2(n8577), .A(n7749), .B(n8560), .ZN(n13106)
         );
  INV_X1 U7185 ( .A(n7040), .ZN(n7904) );
  INV_X2 U7186 ( .A(n8577), .ZN(n9268) );
  NAND2_X1 U7187 ( .A1(n7854), .A2(n7855), .ZN(n15563) );
  CLKBUF_X1 U7189 ( .A(n9527), .Z(n10254) );
  NOR2_X1 U7190 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6659) );
  NOR2_X1 U7191 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6660) );
  NOR2_X1 U7192 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n8181) );
  NOR2_X1 U7193 ( .A1(n7378), .A2(n9903), .ZN(n7375) );
  INV_X1 U7194 ( .A(n9393), .ZN(n9421) );
  NAND2_X1 U7195 ( .A1(n6432), .A2(n9456), .ZN(n9393) );
  INV_X1 U7196 ( .A(n10585), .ZN(n10473) );
  AND2_X1 U7197 ( .A1(n9840), .A2(n9815), .ZN(n14811) );
  NAND2_X1 U7198 ( .A1(n9550), .A2(n9549), .ZN(n11276) );
  OAI21_X1 U7199 ( .B1(n12366), .B2(n12367), .A(n6525), .ZN(n12562) );
  AND2_X1 U7200 ( .A1(n9415), .A2(n9416), .ZN(n13266) );
  AND2_X1 U7201 ( .A1(n8433), .A2(n8453), .ZN(n14323) );
  INV_X1 U7202 ( .A(n10379), .ZN(n8311) );
  NOR2_X1 U7203 ( .A1(n10107), .A2(n14516), .ZN(n12837) );
  INV_X1 U7204 ( .A(n14084), .ZN(n13986) );
  INV_X1 U7205 ( .A(n7087), .ZN(n10034) );
  NAND2_X1 U7206 ( .A1(n9722), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9747) );
  AND2_X1 U7207 ( .A1(n10443), .A2(n10442), .ZN(n11416) );
  AOI21_X1 U7208 ( .B1(n10356), .B2(n10355), .A(n7008), .ZN(n7808) );
  OAI21_X1 U7209 ( .B1(n9731), .B2(n6553), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9866) );
  INV_X1 U7210 ( .A(n8591), .ZN(n9024) );
  AOI211_X1 U7211 ( .C1(n14516), .C2(n10107), .A(n7907), .B(n12837), .ZN(
        n14515) );
  NAND2_X1 U7212 ( .A1(n8202), .A2(n8201), .ZN(n14655) );
  OAI21_X1 U7213 ( .B1(n10618), .B2(n6729), .A(n6535), .ZN(n12815) );
  NAND2_X1 U7214 ( .A1(n9526), .A2(n6846), .ZN(n12148) );
  INV_X1 U7215 ( .A(n13335), .ZN(n13088) );
  INV_X1 U7216 ( .A(n9010), .ZN(n9075) );
  AND3_X1 U7217 ( .A1(n7061), .A2(n7890), .A3(n7060), .ZN(n13774) );
  NAND2_X1 U7218 ( .A1(n8403), .A2(n8402), .ZN(n14086) );
  INV_X1 U7219 ( .A(n14502), .ZN(n14473) );
  NAND2_X1 U7220 ( .A1(n7287), .A2(n6882), .ZN(n14683) );
  INV_X1 U7221 ( .A(n10609), .ZN(n14836) );
  AOI211_X1 U7222 ( .C1(n11244), .C2(n11243), .A(n14854), .B(n11242), .ZN(
        n14856) );
  INV_X1 U7223 ( .A(n12906), .ZN(n12557) );
  AOI21_X2 U7224 ( .B1(n13039), .B2(n12941), .A(n12940), .ZN(n13016) );
  AND2_X1 U7225 ( .A1(n12878), .A2(n6439), .ZN(n6430) );
  NAND2_X2 U7226 ( .A1(n11351), .A2(n10477), .ZN(n11355) );
  AND2_X1 U7227 ( .A1(n11353), .A2(n11354), .ZN(n10477) );
  AOI21_X2 U7228 ( .B1(n11381), .B2(n11382), .A(n7249), .ZN(n11446) );
  OAI22_X2 U7229 ( .A1(n11473), .A2(n11474), .B1(n9208), .B2(n11488), .ZN(
        n11381) );
  NAND2_X2 U7230 ( .A1(n15392), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U7231 ( .A1(n10430), .A2(n10431), .ZN(n11602) );
  INV_X1 U7232 ( .A(n14855), .ZN(n9507) );
  NAND4_X2 U7233 ( .A1(n9489), .A2(n9490), .A3(n9492), .A4(n9491), .ZN(n14855)
         );
  INV_X4 U7234 ( .A(n8561), .ZN(n9279) );
  AOI21_X2 U7235 ( .B1(n14317), .B2(n10085), .A(n10084), .ZN(n14299) );
  INV_X2 U7237 ( .A(n12972), .ZN(n7186) );
  AOI211_X2 U7238 ( .C1(n15175), .C2(n12894), .A(n12893), .B(n12892), .ZN(
        n12895) );
  BUF_X4 U7239 ( .A(n10319), .Z(n6431) );
  INV_X2 U7240 ( .A(n9695), .ZN(n10319) );
  OAI22_X2 U7241 ( .A1(n11222), .A2(n11223), .B1(n9205), .B2(n9204), .ZN(
        n11149) );
  AOI22_X2 U7242 ( .A1(n11134), .A2(n11135), .B1(n11145), .B2(n9203), .ZN(
        n11222) );
  BUF_X2 U7243 ( .A(n9516), .Z(n9779) );
  XNOR2_X1 U7245 ( .A(n7504), .B(P3_IR_REG_21__SCAN_IN), .ZN(n9071) );
  XNOR2_X2 U7246 ( .A(n9337), .B(n13104), .ZN(n12018) );
  XNOR2_X2 U7247 ( .A(n7857), .B(n7856), .ZN(n8505) );
  OAI21_X2 U7248 ( .B1(n7861), .B2(P2_IR_REG_20__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7857) );
  NAND2_X1 U7249 ( .A1(n13644), .A2(n13643), .ZN(n13642) );
  AOI21_X1 U7250 ( .B1(n9922), .B2(n15327), .A(n9921), .ZN(n12891) );
  AND2_X1 U7251 ( .A1(n7373), .A2(n7372), .ZN(n15003) );
  NAND2_X1 U7252 ( .A1(n15057), .A2(n15059), .ZN(n15056) );
  NOR2_X1 U7253 ( .A1(n13203), .A2(n13204), .ZN(n13202) );
  NOR2_X1 U7254 ( .A1(n9837), .A2(n7422), .ZN(n7421) );
  NAND2_X1 U7255 ( .A1(n8451), .A2(n8450), .ZN(n14519) );
  AOI21_X1 U7256 ( .B1(n7571), .B2(n13724), .A(n7570), .ZN(n7569) );
  AND2_X1 U7257 ( .A1(n15004), .A2(n9822), .ZN(n12866) );
  NAND2_X1 U7258 ( .A1(n8396), .A2(n8395), .ZN(n14536) );
  NAND2_X1 U7259 ( .A1(n9801), .A2(n9800), .ZN(n15049) );
  NAND2_X1 U7260 ( .A1(n8257), .A2(n8256), .ZN(n14450) );
  NAND2_X1 U7261 ( .A1(n8139), .A2(n8138), .ZN(n14594) );
  OR2_X1 U7262 ( .A1(n15338), .A2(n14820), .ZN(n15216) );
  INV_X1 U7265 ( .A(n10139), .ZN(n10206) );
  INV_X2 U7266 ( .A(n10439), .ZN(n10643) );
  CLKBUF_X1 U7268 ( .A(n9579), .Z(n14850) );
  CLKBUF_X1 U7269 ( .A(n9965), .Z(n14110) );
  AOI22_X1 U7270 ( .A1(n11209), .A2(n11286), .B1(n9200), .B2(n9199), .ZN(
        n11181) );
  INV_X2 U7271 ( .A(n13818), .ZN(n6433) );
  INV_X2 U7272 ( .A(n10255), .ZN(n9782) );
  INV_X4 U7273 ( .A(n14469), .ZN(n14486) );
  INV_X1 U7274 ( .A(n9880), .ZN(n9877) );
  INV_X1 U7275 ( .A(n7976), .ZN(n6434) );
  CLKBUF_X2 U7276 ( .A(n10018), .Z(n7091) );
  CLKBUF_X2 U7277 ( .A(n7910), .Z(n7040) );
  AND2_X1 U7278 ( .A1(n12014), .A2(n14280), .ZN(n14070) );
  INV_X1 U7279 ( .A(n8505), .ZN(n13756) );
  NAND2_X1 U7280 ( .A1(n8505), .A2(n13757), .ZN(n8504) );
  XNOR2_X1 U7281 ( .A(n7510), .B(n8544), .ZN(n13594) );
  INV_X4 U7282 ( .A(n7944), .ZN(n7007) );
  MUX2_X1 U7283 ( .A(n13509), .B(P3_REG1_REG_28__SCAN_IN), .S(n15637), .Z(
        n13438) );
  MUX2_X1 U7284 ( .A(n13509), .B(P3_REG2_REG_28__SCAN_IN), .S(n15587), .Z(
        n13256) );
  NAND2_X1 U7285 ( .A1(n12815), .A2(n10642), .ZN(n10661) );
  OAI21_X1 U7286 ( .B1(n14292), .B2(n15567), .A(n14295), .ZN(n7109) );
  AOI22_X1 U7287 ( .A1(n6678), .A2(n13731), .B1(n13642), .B2(n7577), .ZN(
        n13742) );
  MUX2_X1 U7288 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n13509), .S(n15631), .Z(
        n13513) );
  AND3_X1 U7289 ( .A1(n14315), .A2(n14314), .A3(n14313), .ZN(n14316) );
  NAND2_X1 U7290 ( .A1(n9442), .A2(n7163), .ZN(n13262) );
  OR2_X1 U7291 ( .A1(n13021), .A2(n6574), .ZN(n6705) );
  NOR2_X1 U7292 ( .A1(n10100), .A2(n7092), .ZN(n14517) );
  NAND2_X1 U7293 ( .A1(n6938), .A2(n6937), .ZN(n8464) );
  AND2_X1 U7294 ( .A1(n13280), .A2(n7081), .ZN(n13445) );
  NOR2_X1 U7295 ( .A1(n7038), .A2(n7037), .ZN(n7036) );
  NAND2_X1 U7296 ( .A1(n13683), .A2(n8407), .ZN(n13644) );
  AOI21_X1 U7297 ( .B1(n7491), .B2(n15482), .A(n7489), .ZN(n12882) );
  OAI21_X1 U7298 ( .B1(n14304), .B2(n6885), .A(n6539), .ZN(n10104) );
  MUX2_X1 U7299 ( .A(n12829), .B(n12828), .S(n14618), .Z(n12830) );
  NAND2_X1 U7300 ( .A1(n7001), .A2(n9415), .ZN(n7159) );
  AOI21_X1 U7301 ( .B1(n14302), .B2(n14481), .A(n14301), .ZN(n14522) );
  OAI211_X1 U7302 ( .C1(n12939), .C2(n12925), .A(n12924), .B(n12923), .ZN(
        n12990) );
  AOI21_X1 U7303 ( .B1(n7089), .B2(n14481), .A(n14320), .ZN(n14529) );
  NAND2_X1 U7304 ( .A1(n7172), .A2(n7171), .ZN(n12939) );
  AND2_X1 U7305 ( .A1(n15017), .A2(n15016), .ZN(n15263) );
  NOR2_X1 U7306 ( .A1(n7137), .A2(n6491), .ZN(n7136) );
  INV_X1 U7307 ( .A(n7723), .ZN(n14284) );
  OAI211_X1 U7308 ( .C1(n12896), .C2(n15353), .A(n12891), .B(n12888), .ZN(
        n10368) );
  XNOR2_X1 U7309 ( .A(n6683), .B(n15235), .ZN(n6720) );
  NAND2_X1 U7310 ( .A1(n9427), .A2(n9426), .ZN(n13250) );
  NAND2_X1 U7311 ( .A1(n15253), .A2(n9861), .ZN(n12896) );
  NAND2_X1 U7312 ( .A1(n13220), .A2(n7526), .ZN(n13187) );
  NAND2_X1 U7313 ( .A1(n12963), .A2(n7174), .ZN(n7172) );
  INV_X1 U7314 ( .A(n6826), .ZN(n13172) );
  OAI22_X1 U7315 ( .A1(n13974), .A2(n7604), .B1(n13973), .B2(n13972), .ZN(
        n13979) );
  OAI211_X1 U7316 ( .C1(n13634), .C2(n8372), .A(n6670), .B(n6669), .ZN(n13613)
         );
  NAND2_X1 U7317 ( .A1(n13634), .A2(n6671), .ZN(n6670) );
  NAND2_X1 U7318 ( .A1(n14333), .A2(n14332), .ZN(n14317) );
  OR2_X1 U7319 ( .A1(n14023), .A2(n14079), .ZN(n14024) );
  NAND2_X1 U7320 ( .A1(n14381), .A2(n10005), .ZN(n14364) );
  NAND2_X1 U7321 ( .A1(n13047), .A2(n13046), .ZN(n13045) );
  NAND2_X1 U7322 ( .A1(n13005), .A2(n12910), .ZN(n13047) );
  NAND2_X1 U7323 ( .A1(n7371), .A2(n7381), .ZN(n15005) );
  NAND2_X1 U7324 ( .A1(n10378), .A2(n10377), .ZN(n14023) );
  AOI21_X1 U7325 ( .B1(n7174), .B2(n7177), .A(n6501), .ZN(n7171) );
  NAND2_X1 U7326 ( .A1(n7423), .A2(n7421), .ZN(n7419) );
  OR3_X1 U7327 ( .A1(n15297), .A2(n15296), .A3(n15295), .ZN(n15371) );
  OAI21_X1 U7328 ( .B1(n10692), .B2(n7539), .A(n7537), .ZN(n9191) );
  INV_X1 U7329 ( .A(n13723), .ZN(n8271) );
  XNOR2_X1 U7330 ( .A(n10317), .B(n10316), .ZN(n14666) );
  OR2_X1 U7331 ( .A1(n14676), .A2(n10374), .ZN(n10376) );
  NOR2_X1 U7332 ( .A1(n13202), .A2(n7263), .ZN(n7262) );
  NAND2_X1 U7333 ( .A1(n10314), .A2(n10268), .ZN(n14676) );
  AND2_X1 U7334 ( .A1(n15074), .A2(n9788), .ZN(n15057) );
  OR2_X1 U7335 ( .A1(n15244), .A2(n15013), .ZN(n9859) );
  NAND2_X1 U7336 ( .A1(n7360), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7359) );
  AND2_X1 U7337 ( .A1(n6920), .A2(n6919), .ZN(n15070) );
  AOI21_X1 U7338 ( .B1(n7780), .B2(n7782), .A(n6532), .ZN(n7778) );
  NAND2_X2 U7339 ( .A1(n6692), .A2(n9852), .ZN(n15244) );
  NOR2_X1 U7340 ( .A1(n13731), .A2(n8421), .ZN(n7577) );
  AOI21_X1 U7341 ( .B1(n7567), .B2(n7572), .A(n7565), .ZN(n7000) );
  NAND2_X1 U7342 ( .A1(n9190), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U7343 ( .A1(n10276), .A2(n10275), .ZN(n15246) );
  NAND2_X1 U7344 ( .A1(n10010), .A2(n10009), .ZN(n14293) );
  NAND2_X1 U7345 ( .A1(n10017), .A2(n10016), .ZN(n14516) );
  INV_X1 U7346 ( .A(n15063), .ZN(n7077) );
  OR2_X1 U7347 ( .A1(n10267), .A2(n10266), .ZN(n10314) );
  AND2_X1 U7348 ( .A1(n7569), .A2(n6616), .ZN(n7567) );
  NAND2_X1 U7349 ( .A1(n9839), .A2(n9838), .ZN(n15258) );
  XNOR2_X1 U7350 ( .A(n13452), .B(n12942), .ZN(n9412) );
  CLKBUF_X1 U7351 ( .A(n15118), .Z(n7051) );
  OR2_X1 U7352 ( .A1(n6568), .A2(n11777), .ZN(n6964) );
  NAND2_X1 U7353 ( .A1(n6925), .A2(n6672), .ZN(n6669) );
  NOR2_X1 U7354 ( .A1(n6672), .A2(n6925), .ZN(n6671) );
  NAND2_X1 U7355 ( .A1(n7475), .A2(n7478), .ZN(n15087) );
  OAI211_X1 U7356 ( .C1(n15118), .C2(n7406), .A(n9776), .B(n7129), .ZN(n15076)
         );
  OR2_X1 U7357 ( .A1(n9189), .A2(n13146), .ZN(n9190) );
  AND2_X1 U7358 ( .A1(n14378), .A2(n10076), .ZN(n7683) );
  NOR2_X1 U7359 ( .A1(n7785), .A2(n14347), .ZN(n7784) );
  XNOR2_X1 U7360 ( .A(n15282), .B(n15072), .ZN(n15059) );
  AND2_X1 U7361 ( .A1(n10077), .A2(n10003), .ZN(n14378) );
  NOR2_X1 U7362 ( .A1(n14541), .A2(n14087), .ZN(n7785) );
  OR2_X1 U7363 ( .A1(n7405), .A2(n7409), .ZN(n7129) );
  NAND2_X1 U7364 ( .A1(n14325), .A2(n7736), .ZN(n7735) );
  XNOR2_X1 U7365 ( .A(n10014), .B(n10013), .ZN(n14678) );
  XNOR2_X1 U7366 ( .A(n9851), .B(n8449), .ZN(n12709) );
  NAND2_X1 U7367 ( .A1(n7323), .A2(n9850), .ZN(n10014) );
  OAI21_X1 U7368 ( .B1(n6481), .B2(n9899), .A(n7483), .ZN(n7479) );
  OR2_X1 U7369 ( .A1(n14634), .A2(n13960), .ZN(n10077) );
  NAND2_X2 U7370 ( .A1(n6679), .A2(n9789), .ZN(n15282) );
  NOR2_X1 U7371 ( .A1(n15107), .A2(n7410), .ZN(n7409) );
  NAND2_X1 U7372 ( .A1(n7616), .A2(n6573), .ZN(n12697) );
  NAND2_X2 U7373 ( .A1(n8352), .A2(n8351), .ZN(n14541) );
  NAND2_X1 U7374 ( .A1(n9812), .A2(n9811), .ZN(n15264) );
  NAND2_X2 U7375 ( .A1(n8346), .A2(n8345), .ZN(n14634) );
  NOR2_X1 U7376 ( .A1(n14706), .A2(n7631), .ZN(n7630) );
  NAND2_X1 U7377 ( .A1(n9153), .A2(n10826), .ZN(n7350) );
  NAND2_X1 U7378 ( .A1(n8444), .A2(n8443), .ZN(n8448) );
  XNOR2_X1 U7379 ( .A(n15115), .B(n15089), .ZN(n15104) );
  XNOR2_X1 U7380 ( .A(n8350), .B(n8385), .ZN(n12398) );
  NAND2_X1 U7381 ( .A1(n12564), .A2(n6649), .ZN(n12951) );
  AND2_X1 U7382 ( .A1(n8290), .A2(n8289), .ZN(n13629) );
  NAND2_X1 U7383 ( .A1(n8446), .A2(SI_26_), .ZN(n8447) );
  NAND2_X1 U7384 ( .A1(n8411), .A2(n8410), .ZN(n14629) );
  OR2_X1 U7385 ( .A1(n12221), .A2(n10374), .ZN(n8346) );
  NAND2_X1 U7386 ( .A1(n15402), .A2(n9779), .ZN(n15370) );
  NAND2_X1 U7387 ( .A1(n9717), .A2(n15183), .ZN(n6856) );
  NAND2_X1 U7388 ( .A1(n8329), .A2(n8328), .ZN(n14638) );
  NAND2_X1 U7389 ( .A1(n8418), .A2(n8417), .ZN(n14085) );
  XNOR2_X1 U7390 ( .A(n9228), .B(n9227), .ZN(n13156) );
  XNOR2_X1 U7391 ( .A(n8445), .B(n8428), .ZN(n12669) );
  NAND2_X1 U7392 ( .A1(n12172), .A2(n7505), .ZN(n6649) );
  AND2_X1 U7393 ( .A1(n6934), .A2(n6932), .ZN(n9899) );
  NAND2_X1 U7394 ( .A1(n8348), .A2(n8347), .ZN(n8350) );
  NAND2_X2 U7395 ( .A1(n9756), .A2(n9755), .ZN(n15115) );
  XNOR2_X1 U7396 ( .A(n9778), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15402) );
  NAND2_X1 U7397 ( .A1(n6687), .A2(n8427), .ZN(n8445) );
  OR2_X1 U7398 ( .A1(n12224), .A2(n10374), .ZN(n8396) );
  NAND2_X2 U7399 ( .A1(n8306), .A2(n8305), .ZN(n14557) );
  OR2_X1 U7400 ( .A1(n12211), .A2(n10374), .ZN(n8329) );
  NAND2_X1 U7401 ( .A1(n6726), .A2(n11526), .ZN(n6725) );
  OR2_X1 U7402 ( .A1(n12224), .A2(n10270), .ZN(n9801) );
  OR2_X1 U7403 ( .A1(n15178), .A2(n15179), .ZN(n9717) );
  NAND2_X1 U7404 ( .A1(n11869), .A2(n11868), .ZN(n12172) );
  NOR2_X1 U7405 ( .A1(n15140), .A2(n7482), .ZN(n7481) );
  NAND2_X1 U7406 ( .A1(n8409), .A2(n8394), .ZN(n12224) );
  AND2_X1 U7407 ( .A1(n8174), .A2(n8151), .ZN(n7589) );
  INV_X1 U7408 ( .A(n15140), .ZN(n15138) );
  NAND2_X1 U7409 ( .A1(n9707), .A2(n9706), .ZN(n15178) );
  NOR2_X1 U7410 ( .A1(n7181), .A2(n6711), .ZN(n6710) );
  OR2_X1 U7411 ( .A1(n12155), .A2(n10374), .ZN(n8306) );
  NAND2_X2 U7412 ( .A1(n7607), .A2(n8275), .ZN(n14433) );
  NAND2_X1 U7413 ( .A1(n11996), .A2(n10059), .ZN(n11999) );
  NAND2_X1 U7414 ( .A1(n13136), .A2(n6604), .ZN(n10695) );
  NAND2_X1 U7415 ( .A1(n8321), .A2(n8304), .ZN(n12155) );
  NAND2_X1 U7416 ( .A1(n8347), .A2(n6749), .ZN(n9777) );
  NAND2_X1 U7417 ( .A1(n6691), .A2(n6690), .ZN(n8409) );
  NOR2_X1 U7418 ( .A1(n7183), .A2(n7182), .ZN(n7181) );
  NAND2_X1 U7419 ( .A1(n6682), .A2(SI_22_), .ZN(n8347) );
  NOR2_X1 U7420 ( .A1(n14060), .A2(n7772), .ZN(n7771) );
  AND2_X1 U7421 ( .A1(n7368), .A2(n6930), .ZN(n6929) );
  NAND2_X1 U7422 ( .A1(n13126), .A2(n13125), .ZN(n13139) );
  AND2_X1 U7423 ( .A1(n15136), .A2(n10221), .ZN(n15164) );
  NAND2_X1 U7424 ( .A1(n9734), .A2(n9733), .ZN(n15149) );
  OR2_X1 U7425 ( .A1(n11745), .A2(n10374), .ZN(n8257) );
  OR2_X1 U7426 ( .A1(n15213), .A2(n14746), .ZN(n10209) );
  NAND2_X1 U7427 ( .A1(n11923), .A2(n6519), .ZN(n11737) );
  AND2_X1 U7428 ( .A1(n12546), .A2(n7369), .ZN(n7368) );
  AND2_X1 U7429 ( .A1(n9787), .A2(n9786), .ZN(n15090) );
  NAND2_X1 U7430 ( .A1(n8186), .A2(n8185), .ZN(n13887) );
  AND2_X2 U7431 ( .A1(n15216), .A2(n10198), .ZN(n12648) );
  OR2_X1 U7432 ( .A1(n15319), .A2(n15193), .ZN(n15136) );
  OR2_X1 U7433 ( .A1(n8390), .A2(SI_24_), .ZN(n8391) );
  NAND2_X1 U7434 ( .A1(n8326), .A2(n8381), .ZN(n8342) );
  NAND2_X1 U7435 ( .A1(n7464), .A2(n7463), .ZN(n11923) );
  OR2_X1 U7436 ( .A1(n8384), .A2(n11524), .ZN(n8319) );
  NAND2_X1 U7437 ( .A1(n9664), .A2(n9663), .ZN(n12552) );
  NAND2_X1 U7438 ( .A1(n13899), .A2(n13893), .ZN(n14651) );
  NOR2_X1 U7439 ( .A1(n12387), .A2(n12386), .ZN(n12385) );
  AND2_X1 U7440 ( .A1(n9647), .A2(n12240), .ZN(n9648) );
  OR2_X1 U7441 ( .A1(n8248), .A2(n8292), .ZN(n8273) );
  OAI21_X1 U7442 ( .B1(n11574), .B2(n6754), .A(n6750), .ZN(n11753) );
  NAND2_X1 U7443 ( .A1(n10037), .A2(n6517), .ZN(n11788) );
  NAND2_X1 U7444 ( .A1(n9711), .A2(n9710), .ZN(n15188) );
  NAND2_X1 U7445 ( .A1(n9721), .A2(n9720), .ZN(n15319) );
  NAND2_X1 U7446 ( .A1(n8163), .A2(n8162), .ZN(n13880) );
  XNOR2_X1 U7447 ( .A(n8180), .B(n8179), .ZN(n11516) );
  AND2_X1 U7448 ( .A1(n8071), .A2(n6940), .ZN(n11837) );
  NAND2_X1 U7449 ( .A1(n8178), .A2(n8177), .ZN(n8180) );
  OR2_X1 U7450 ( .A1(n8297), .A2(n11069), .ZN(n8272) );
  OAI21_X1 U7451 ( .B1(n8297), .B2(n8296), .A(n8295), .ZN(n8301) );
  NAND2_X1 U7452 ( .A1(n9639), .A2(n9638), .ZN(n15349) );
  NAND2_X1 U7453 ( .A1(n8094), .A2(n8093), .ZN(n13860) );
  OAI21_X1 U7454 ( .B1(n8196), .B2(n6482), .A(n8195), .ZN(n8222) );
  OAI21_X2 U7455 ( .B1(n10667), .B2(n10663), .A(n15208), .ZN(n10664) );
  NAND2_X1 U7456 ( .A1(n7340), .A2(n8246), .ZN(n8297) );
  OAI21_X1 U7457 ( .B1(n8187), .B2(n7341), .A(n6684), .ZN(n7340) );
  AND2_X1 U7458 ( .A1(n10051), .A2(n11570), .ZN(n11429) );
  NAND2_X1 U7459 ( .A1(n9598), .A2(n9597), .ZN(n11961) );
  NAND2_X1 U7460 ( .A1(n8060), .A2(n8059), .ZN(n14610) );
  AND3_X1 U7461 ( .A1(n9923), .A2(n11111), .A3(n7454), .ZN(n11949) );
  NAND2_X1 U7462 ( .A1(n8077), .A2(n8076), .ZN(n14604) );
  NAND2_X1 U7463 ( .A1(n8037), .A2(n8036), .ZN(n13840) );
  NAND2_X1 U7464 ( .A1(n7392), .A2(n11113), .ZN(n12120) );
  NAND2_X1 U7465 ( .A1(n9611), .A2(n9610), .ZN(n12217) );
  XNOR2_X1 U7466 ( .A(n8107), .B(n8108), .ZN(n10943) );
  NAND2_X1 U7467 ( .A1(n9628), .A2(n9627), .ZN(n12166) );
  NAND2_X1 U7468 ( .A1(n7100), .A2(n8159), .ZN(n8187) );
  OR2_X1 U7469 ( .A1(n10876), .A2(n10270), .ZN(n9611) );
  AND2_X1 U7470 ( .A1(n10146), .A2(n10147), .ZN(n10335) );
  NAND2_X1 U7471 ( .A1(n9583), .A2(n6945), .ZN(n15503) );
  NOR2_X1 U7472 ( .A1(n9145), .A2(n6820), .ZN(n11153) );
  NAND2_X1 U7473 ( .A1(n7986), .A2(n7985), .ZN(n13813) );
  NAND2_X1 U7474 ( .A1(n8013), .A2(n8012), .ZN(n14614) );
  AND2_X1 U7475 ( .A1(n6823), .A2(n6583), .ZN(n6820) );
  INV_X1 U7476 ( .A(n7403), .ZN(n11203) );
  AND2_X1 U7477 ( .A1(n9319), .A2(n12027), .ZN(n11675) );
  AOI21_X1 U7478 ( .B1(n7599), .B2(n7600), .A(n6685), .ZN(n6684) );
  INV_X1 U7479 ( .A(n9579), .ZN(n11805) );
  INV_X1 U7480 ( .A(n8639), .ZN(n13102) );
  INV_X1 U7481 ( .A(n14849), .ZN(n11938) );
  OAI22_X1 U7482 ( .A1(n11181), .A2(n11182), .B1(n9201), .B2(n6814), .ZN(
        n11134) );
  AND4_X1 U7483 ( .A1(n9619), .A2(n9618), .A3(n9617), .A4(n9616), .ZN(n12162)
         );
  AND4_X1 U7484 ( .A1(n9606), .A2(n9605), .A3(n9604), .A4(n9603), .ZN(n12075)
         );
  AND2_X1 U7485 ( .A1(n7338), .A2(n8057), .ZN(n7071) );
  INV_X2 U7486 ( .A(n13956), .ZN(n13818) );
  NOR2_X2 U7487 ( .A1(n9927), .A2(n9877), .ZN(n10125) );
  NAND2_X1 U7488 ( .A1(n7560), .A2(n6767), .ZN(n7559) );
  NAND4_X1 U7489 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .ZN(n14109)
         );
  AND4_X1 U7490 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n8591)
         );
  OAI21_X1 U7491 ( .B1(n9002), .B2(P3_IR_REG_20__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7504) );
  AND3_X1 U7492 ( .A1(n8559), .A2(n8558), .A3(n6566), .ZN(n9292) );
  NOR2_X1 U7493 ( .A1(n9143), .A2(n6810), .ZN(n11138) );
  NAND4_X1 U7494 ( .A1(n7933), .A2(n7932), .A3(n7931), .A4(n7930), .ZN(n14107)
         );
  XNOR2_X1 U7495 ( .A(n9199), .B(n9173), .ZN(n11209) );
  NAND2_X1 U7496 ( .A1(n6991), .A2(n6990), .ZN(n9002) );
  AND2_X1 U7497 ( .A1(n7265), .A2(n7264), .ZN(n9199) );
  NAND2_X2 U7498 ( .A1(n9486), .A2(n9485), .ZN(n9519) );
  NAND2_X2 U7499 ( .A1(n12885), .A2(n10363), .ZN(n9516) );
  AND2_X1 U7500 ( .A1(n6812), .A2(n6811), .ZN(n9143) );
  CLKBUF_X3 U7501 ( .A(n7929), .Z(n10379) );
  NAND2_X1 U7502 ( .A1(n10122), .A2(n9927), .ZN(n10121) );
  AND2_X1 U7503 ( .A1(n14674), .A2(n7876), .ZN(n7929) );
  INV_X1 U7504 ( .A(n9926), .ZN(n10122) );
  NAND2_X2 U7505 ( .A1(n9168), .A2(n7007), .ZN(n8905) );
  NAND2_X1 U7506 ( .A1(n9934), .A2(n7383), .ZN(n12674) );
  NAND2_X1 U7507 ( .A1(n8547), .A2(n8546), .ZN(n8744) );
  CLKBUF_X1 U7508 ( .A(n9926), .Z(n10324) );
  NAND2_X1 U7509 ( .A1(n13594), .A2(n8547), .ZN(n8969) );
  NAND2_X1 U7510 ( .A1(n9875), .A2(n9876), .ZN(n9927) );
  XNOR2_X1 U7511 ( .A(n9866), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9926) );
  INV_X1 U7512 ( .A(n9485), .ZN(n15401) );
  CLKBUF_X1 U7513 ( .A(n9072), .Z(n12813) );
  MUX2_X1 U7514 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9933), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9934) );
  XNOR2_X1 U7515 ( .A(n9936), .B(n9935), .ZN(n12480) );
  NAND2_X2 U7516 ( .A1(n9072), .A2(n13601), .ZN(n9168) );
  OAI21_X1 U7517 ( .B1(SI_7_), .B2(n7343), .A(n8029), .ZN(n8026) );
  XNOR2_X1 U7518 ( .A(n7858), .B(n7862), .ZN(n12014) );
  XNOR2_X1 U7519 ( .A(n8552), .B(n8551), .ZN(n9072) );
  NAND2_X2 U7520 ( .A1(n8554), .A2(n8553), .ZN(n13601) );
  OAI21_X1 U7521 ( .B1(n9942), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9933) );
  AND2_X1 U7522 ( .A1(n9928), .A2(n9874), .ZN(n9875) );
  OR2_X1 U7523 ( .A1(n9870), .A2(n9863), .ZN(n9864) );
  OAI211_X1 U7524 ( .C1(n7868), .C2(n7867), .A(n8499), .B(n7866), .ZN(n13757)
         );
  XNOR2_X1 U7525 ( .A(n9484), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9485) );
  AND2_X1 U7526 ( .A1(n7853), .A2(n7947), .ZN(n14130) );
  XNOR2_X1 U7527 ( .A(n7874), .B(n7873), .ZN(n7876) );
  NAND2_X1 U7528 ( .A1(n6883), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7722) );
  NOR2_X1 U7529 ( .A1(n7815), .A2(n10784), .ZN(n7895) );
  XNOR2_X1 U7530 ( .A(n8110), .B(SI_11_), .ZN(n8108) );
  NAND2_X1 U7531 ( .A1(n7050), .A2(n7006), .ZN(n8030) );
  NAND2_X1 U7532 ( .A1(n7695), .A2(n6526), .ZN(n8554) );
  NAND2_X1 U7533 ( .A1(n6651), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7510) );
  XNOR2_X1 U7534 ( .A(n8597), .B(P3_IR_REG_4__SCAN_IN), .ZN(n11236) );
  NAND2_X2 U7535 ( .A1(n10801), .A2(P1_U3086), .ZN(n15397) );
  NAND2_X2 U7536 ( .A1(n7007), .A2(P2_U3088), .ZN(n14682) );
  NAND2_X2 U7537 ( .A1(n7007), .A2(P1_U3086), .ZN(n15400) );
  AND3_X1 U7538 ( .A1(n9476), .A2(n9477), .A3(n6451), .ZN(n9931) );
  XNOR2_X1 U7539 ( .A(n8586), .B(P3_IR_REG_3__SCAN_IN), .ZN(n11145) );
  AND2_X1 U7540 ( .A1(n9480), .A2(n7473), .ZN(n7472) );
  XNOR2_X1 U7541 ( .A(n9525), .B(P1_IR_REG_2__SCAN_IN), .ZN(n11247) );
  AND2_X1 U7542 ( .A1(n9493), .A2(n9496), .ZN(n7473) );
  AND4_X1 U7543 ( .A1(n8865), .A2(n8540), .A3(n8539), .A4(n9001), .ZN(n9004)
         );
  NAND4_X1 U7544 ( .A1(n7320), .A2(n15465), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6935) );
  AND3_X1 U7545 ( .A1(n6648), .A2(n6647), .A3(n6646), .ZN(n8761) );
  AND3_X1 U7546 ( .A1(n9479), .A2(n7056), .A3(n9478), .ZN(n6451) );
  AND2_X1 U7547 ( .A1(n9475), .A2(n9929), .ZN(n9476) );
  NAND4_X1 U7548 ( .A1(n8537), .A2(n8649), .A3(n8536), .A4(n8535), .ZN(n8760)
         );
  INV_X1 U7549 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7830) );
  INV_X1 U7550 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7831) );
  INV_X1 U7551 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7832) );
  INV_X1 U7552 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8535) );
  NOR2_X1 U7553 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n8537) );
  INV_X4 U7554 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U7555 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7556 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n14283) );
  INV_X1 U7557 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7320) );
  NOR2_X1 U7558 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n6646) );
  NOR2_X1 U7559 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n6647) );
  INV_X1 U7560 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9623) );
  INV_X1 U7561 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7833) );
  INV_X1 U7562 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7834) );
  INV_X1 U7563 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7835) );
  INV_X1 U7564 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7501) );
  NOR2_X1 U7565 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6661) );
  INV_X1 U7566 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7845) );
  NOR2_X1 U7567 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9470) );
  INV_X1 U7568 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8534) );
  NOR2_X1 U7569 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6637) );
  INV_X1 U7570 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9479) );
  NOR2_X1 U7571 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9676) );
  NOR2_X1 U7572 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n9475) );
  NOR2_X1 U7573 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9675) );
  INV_X1 U7574 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8477) );
  INV_X1 U7575 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8649) );
  INV_X1 U7576 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9551) );
  NOR2_X1 U7577 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n9480) );
  INV_X1 U7578 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9565) );
  INV_X4 U7579 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X2 U7580 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8865) );
  NOR2_X1 U7581 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n6648) );
  NOR2_X1 U7582 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), .ZN(
        n8539) );
  AND2_X4 U7583 ( .A1(n10419), .A2(n10421), .ZN(n6438) );
  NAND2_X2 U7584 ( .A1(n6847), .A2(n9522), .ZN(n14853) );
  INV_X1 U7585 ( .A(n9487), .ZN(n9486) );
  INV_X1 U7586 ( .A(n10585), .ZN(n6436) );
  OR2_X1 U7587 ( .A1(n6734), .A2(n9932), .ZN(n9942) );
  NOR2_X2 U7588 ( .A1(n9712), .A2(n12803), .ZN(n9722) );
  INV_X1 U7589 ( .A(n9516), .ZN(n6437) );
  NAND2_X1 U7590 ( .A1(n7849), .A2(n7007), .ZN(n6668) );
  OAI21_X2 U7591 ( .B1(n13290), .B2(n13289), .A(n9315), .ZN(n13281) );
  XNOR2_X2 U7592 ( .A(n10434), .B(n10449), .ZN(n10445) );
  INV_X4 U7593 ( .A(n6438), .ZN(n10627) );
  NAND2_X2 U7594 ( .A1(n10420), .A2(n14967), .ZN(n12878) );
  INV_X1 U7595 ( .A(n10439), .ZN(n6439) );
  XNOR2_X1 U7596 ( .A(n9864), .B(n9865), .ZN(n9909) );
  XNOR2_X2 U7597 ( .A(n14991), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n12889) );
  NAND2_X1 U7598 ( .A1(n10608), .A2(n10607), .ZN(n14761) );
  OAI21_X1 U7599 ( .B1(n9779), .B2(P1_IR_REG_0__SCAN_IN), .A(n7404), .ZN(n7403) );
  NAND2_X2 U7600 ( .A1(n14688), .A2(n10534), .ZN(n14740) );
  NAND2_X2 U7601 ( .A1(n14775), .A2(n7628), .ZN(n14688) );
  NAND2_X2 U7602 ( .A1(n14777), .A2(n14776), .ZN(n14775) );
  NOR2_X2 U7603 ( .A1(n15158), .A2(n15149), .ZN(n15148) );
  NAND2_X2 U7604 ( .A1(n14756), .A2(n10563), .ZN(n14800) );
  NAND2_X2 U7605 ( .A1(n10560), .A2(n10559), .ZN(n14756) );
  INV_X1 U7606 ( .A(n13956), .ZN(n6440) );
  INV_X1 U7607 ( .A(n13956), .ZN(n6441) );
  AND2_X4 U7608 ( .A1(n14564), .A2(n13756), .ZN(n13761) );
  INV_X4 U7609 ( .A(n13761), .ZN(n13956) );
  NOR2_X2 U7610 ( .A1(n12189), .A2(n13860), .ZN(n7118) );
  NAND2_X2 U7611 ( .A1(n12349), .A2(n7617), .ZN(n7616) );
  NAND2_X2 U7612 ( .A1(n14761), .A2(n14762), .ZN(n10618) );
  NAND2_X2 U7613 ( .A1(n12697), .A2(n10520), .ZN(n14777) );
  NOR3_X2 U7614 ( .A1(n9747), .A2(n14803), .A3(n9746), .ZN(n9757) );
  NAND2_X2 U7615 ( .A1(n12351), .A2(n12350), .ZN(n12349) );
  AND2_X2 U7616 ( .A1(n6725), .A2(n6579), .ZN(n12351) );
  AND2_X4 U7617 ( .A1(n9535), .A2(n9473), .ZN(n9536) );
  OAI222_X1 U7618 ( .A1(P1_U3086), .A2(n10122), .B1(n15400), .B2(n12211), .C1(
        n6700), .C2(n15397), .ZN(P1_U3334) );
  NOR2_X1 U7619 ( .A1(n14365), .A2(n7737), .ZN(n14339) );
  NOR2_X1 U7620 ( .A1(n14365), .A2(n7735), .ZN(n14321) );
  NOR2_X4 U7621 ( .A1(n14365), .A2(n7733), .ZN(n14311) );
  OR2_X2 U7622 ( .A1(n14382), .A2(n14541), .ZN(n14365) );
  INV_X2 U7623 ( .A(n9932), .ZN(n7470) );
  NAND2_X2 U7624 ( .A1(n9502), .A2(n9501), .ZN(n10363) );
  INV_X1 U7625 ( .A(n13791), .ZN(n9970) );
  NAND2_X2 U7626 ( .A1(n7927), .A2(n7928), .ZN(n13791) );
  OAI21_X2 U7627 ( .B1(n14800), .B2(n6732), .A(n6730), .ZN(n14768) );
  NAND2_X1 U7628 ( .A1(n9487), .A2(n15401), .ZN(n9528) );
  XNOR2_X2 U7629 ( .A(n9483), .B(n9482), .ZN(n9487) );
  AOI21_X1 U7630 ( .B1(n7382), .B2(n15004), .A(n15010), .ZN(n7372) );
  NAND2_X1 U7631 ( .A1(n7376), .A2(n6686), .ZN(n7373) );
  AND2_X1 U7632 ( .A1(n7375), .A2(n15004), .ZN(n6686) );
  AOI21_X1 U7633 ( .B1(n7185), .B2(n12584), .A(n7184), .ZN(n7183) );
  INV_X1 U7634 ( .A(n12686), .ZN(n7184) );
  AND2_X1 U7635 ( .A1(n12585), .A2(n13095), .ZN(n7185) );
  NOR2_X1 U7636 ( .A1(n9182), .A2(n11160), .ZN(n9183) );
  OR2_X1 U7637 ( .A1(n10412), .A2(n12975), .ZN(n9443) );
  NAND2_X1 U7638 ( .A1(n10412), .A2(n12975), .ZN(n9444) );
  OR2_X1 U7639 ( .A1(n12934), .A2(n12976), .ZN(n8999) );
  INV_X1 U7640 ( .A(n7876), .ZN(n6770) );
  AND2_X1 U7641 ( .A1(n10012), .A2(n10011), .ZN(n14068) );
  OR2_X1 U7642 ( .A1(n14293), .A2(n14082), .ZN(n10011) );
  INV_X1 U7643 ( .A(n9984), .ZN(n7766) );
  OR2_X1 U7644 ( .A1(n13806), .A2(n13808), .ZN(n10053) );
  INV_X1 U7645 ( .A(n9810), .ZN(n7422) );
  NOR2_X1 U7646 ( .A1(n15059), .A2(n15075), .ZN(n7380) );
  INV_X1 U7647 ( .A(n7479), .ZN(n7478) );
  INV_X1 U7648 ( .A(n9471), .ZN(n7386) );
  INV_X1 U7649 ( .A(n8744), .ZN(n9258) );
  NAND2_X1 U7650 ( .A1(n7559), .A2(n13763), .ZN(n11121) );
  NAND2_X1 U7651 ( .A1(n6770), .A2(n7875), .ZN(n10018) );
  NAND2_X1 U7652 ( .A1(n10002), .A2(n7760), .ZN(n7759) );
  NOR2_X1 U7653 ( .A1(n14394), .A2(n7761), .ZN(n7760) );
  INV_X1 U7654 ( .A(n10001), .ZN(n7761) );
  NAND2_X1 U7655 ( .A1(n11917), .A2(n9593), .ZN(n6862) );
  NAND2_X1 U7656 ( .A1(n6720), .A2(n15327), .ZN(n6719) );
  AOI21_X1 U7657 ( .B1(n13854), .B2(n13853), .A(n7299), .ZN(n7296) );
  NAND2_X1 U7658 ( .A1(n13850), .A2(n13849), .ZN(n7295) );
  INV_X1 U7659 ( .A(n10163), .ZN(n7102) );
  NAND2_X1 U7660 ( .A1(n6455), .A2(n7292), .ZN(n7289) );
  NAND2_X1 U7661 ( .A1(n9363), .A2(n12530), .ZN(n7231) );
  NOR2_X1 U7662 ( .A1(n7606), .A2(n7605), .ZN(n7604) );
  NAND2_X1 U7663 ( .A1(n10237), .A2(n10235), .ZN(n7553) );
  OAI21_X1 U7664 ( .B1(n10232), .B2(n6871), .A(n6461), .ZN(n6874) );
  NAND2_X1 U7665 ( .A1(n7011), .A2(n7010), .ZN(n9413) );
  OAI21_X1 U7666 ( .B1(n9411), .B2(n9412), .A(n9410), .ZN(n7011) );
  NOR2_X1 U7667 ( .A1(n8915), .A2(n8897), .ZN(n8898) );
  INV_X1 U7668 ( .A(n15563), .ZN(n13783) );
  NAND2_X1 U7669 ( .A1(n6694), .A2(n6693), .ZN(n10306) );
  NAND2_X1 U7670 ( .A1(n15013), .A2(n10281), .ZN(n6693) );
  INV_X1 U7671 ( .A(n10219), .ZN(n7480) );
  OR2_X1 U7672 ( .A1(n15115), .A2(n15089), .ZN(n7483) );
  OAI21_X1 U7673 ( .B1(n7944), .B2(n10839), .A(n7019), .ZN(n7974) );
  NAND2_X1 U7674 ( .A1(n7944), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7019) );
  OAI21_X1 U7675 ( .B1(n10774), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n10773), .ZN(
        n10775) );
  OAI21_X1 U7676 ( .B1(n10815), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n10814), .ZN(
        n10816) );
  NAND2_X1 U7677 ( .A1(n15579), .A2(n12825), .ZN(n7169) );
  AND2_X1 U7678 ( .A1(n11307), .A2(n13584), .ZN(n7170) );
  OAI21_X1 U7679 ( .B1(n13228), .B2(n13230), .A(n9273), .ZN(n9452) );
  INV_X1 U7680 ( .A(n13594), .ZN(n8546) );
  OAI21_X1 U7681 ( .B1(n11483), .B2(n11482), .A(n6913), .ZN(n6917) );
  INV_X1 U7682 ( .A(n6914), .ZN(n6913) );
  OAI21_X1 U7683 ( .B1(n11481), .B2(n11482), .A(n6548), .ZN(n6914) );
  AOI21_X1 U7684 ( .B1(n7535), .B2(n7528), .A(n6530), .ZN(n7527) );
  OR2_X1 U7685 ( .A1(n11460), .A2(n9148), .ZN(n9149) );
  NAND2_X1 U7686 ( .A1(n13118), .A2(n6897), .ZN(n9189) );
  NAND2_X1 U7687 ( .A1(n10869), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U7688 ( .A1(n13177), .A2(n9192), .ZN(n9193) );
  NOR2_X1 U7689 ( .A1(n12928), .A2(n6806), .ZN(n6805) );
  INV_X1 U7690 ( .A(n8977), .ZN(n6806) );
  INV_X1 U7691 ( .A(n6988), .ZN(n8950) );
  AND2_X1 U7692 ( .A1(n9045), .A2(n7743), .ZN(n7742) );
  NAND2_X1 U7693 ( .A1(n9044), .A2(n7744), .ZN(n7743) );
  NOR2_X2 U7694 ( .A1(n8728), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7126) );
  AND2_X1 U7695 ( .A1(n9343), .A2(n9334), .ZN(n12134) );
  NAND2_X1 U7696 ( .A1(n13106), .A2(n13500), .ZN(n9322) );
  OR2_X1 U7697 ( .A1(n13553), .A2(n13009), .ZN(n13325) );
  INV_X1 U7698 ( .A(n7703), .ZN(n7702) );
  OAI21_X1 U7699 ( .B1(n7705), .B2(n7704), .A(n9378), .ZN(n7703) );
  AND2_X1 U7700 ( .A1(n7189), .A2(n12331), .ZN(n7193) );
  OR2_X1 U7701 ( .A1(n7752), .A2(n6443), .ZN(n7189) );
  NAND3_X1 U7702 ( .A1(n8542), .A2(n7187), .A3(n7188), .ZN(n8553) );
  AOI21_X1 U7703 ( .B1(n7666), .B2(n7668), .A(n6631), .ZN(n7664) );
  NAND2_X1 U7704 ( .A1(n8754), .A2(n8753), .ZN(n8756) );
  NAND2_X1 U7705 ( .A1(n10856), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8618) );
  INV_X1 U7706 ( .A(n12471), .ZN(n7591) );
  AND2_X1 U7707 ( .A1(n7574), .A2(n13684), .ZN(n6939) );
  INV_X1 U7708 ( .A(n10380), .ZN(n8512) );
  NAND2_X1 U7709 ( .A1(n7673), .A2(n6765), .ZN(n6764) );
  INV_X1 U7710 ( .A(n14038), .ZN(n6765) );
  AND2_X1 U7711 ( .A1(n9994), .A2(n7768), .ZN(n7767) );
  AND2_X1 U7712 ( .A1(n14466), .A2(n9993), .ZN(n9994) );
  INV_X1 U7713 ( .A(n12493), .ZN(n7774) );
  OR2_X1 U7714 ( .A1(n14054), .A2(n7766), .ZN(n7765) );
  AOI21_X1 U7715 ( .B1(n10053), .B2(n10052), .A(n7076), .ZN(n7794) );
  NAND2_X1 U7716 ( .A1(n14107), .A2(n9970), .ZN(n10051) );
  AND2_X1 U7717 ( .A1(n7285), .A2(n7851), .ZN(n7284) );
  INV_X1 U7718 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7285) );
  INV_X1 U7719 ( .A(n12101), .ZN(n7635) );
  NOR2_X1 U7720 ( .A1(n15059), .A2(n7379), .ZN(n7378) );
  NAND2_X1 U7721 ( .A1(n11737), .A2(n6505), .ZN(n12071) );
  INV_X1 U7722 ( .A(n9889), .ZN(n7384) );
  NAND2_X1 U7723 ( .A1(n12071), .A2(n7474), .ZN(n12159) );
  AND2_X1 U7724 ( .A1(n12160), .A2(n9890), .ZN(n7474) );
  CLKBUF_X1 U7725 ( .A(n10121), .Z(n9962) );
  NOR2_X1 U7726 ( .A1(n6470), .A2(n6610), .ZN(n7322) );
  NAND2_X1 U7727 ( .A1(n8409), .A2(n6688), .ZN(n6687) );
  NAND2_X1 U7728 ( .A1(n8390), .A2(SI_24_), .ZN(n8408) );
  NAND2_X1 U7729 ( .A1(n7239), .A2(n10885), .ZN(n10884) );
  OR2_X1 U7730 ( .A1(n10816), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n7239) );
  AOI21_X1 U7731 ( .B1(n6483), .B2(n7183), .A(n7180), .ZN(n7179) );
  NAND2_X1 U7732 ( .A1(n6710), .A2(n12951), .ZN(n6709) );
  INV_X1 U7733 ( .A(n13100), .ZN(n12360) );
  NAND2_X1 U7734 ( .A1(n13495), .A2(n9322), .ZN(n11311) );
  INV_X1 U7735 ( .A(n9292), .ZN(n9017) );
  INV_X1 U7736 ( .A(n13086), .ZN(n12941) );
  NAND2_X1 U7737 ( .A1(n13228), .A2(n13230), .ZN(n9433) );
  INV_X1 U7738 ( .A(n9433), .ZN(n9449) );
  OR2_X1 U7739 ( .A1(n13234), .A2(n12348), .ZN(n9448) );
  NAND2_X1 U7740 ( .A1(n7222), .A2(n9424), .ZN(n7221) );
  NAND2_X1 U7741 ( .A1(n9423), .A2(n9422), .ZN(n7222) );
  INV_X1 U7742 ( .A(n9452), .ZN(n9435) );
  NAND2_X1 U7743 ( .A1(n13594), .A2(n8545), .ZN(n8561) );
  NAND2_X1 U7744 ( .A1(n6910), .A2(n10689), .ZN(n10688) );
  INV_X1 U7745 ( .A(n6911), .ZN(n6910) );
  NOR2_X1 U7746 ( .A1(n7258), .A2(n13160), .ZN(n7257) );
  OR2_X1 U7747 ( .A1(n9193), .A2(n13194), .ZN(n7526) );
  NAND2_X1 U7748 ( .A1(n9193), .A2(n13194), .ZN(n13220) );
  NAND2_X1 U7749 ( .A1(n9162), .A2(n13194), .ZN(n13207) );
  NAND2_X1 U7750 ( .A1(n9427), .A2(n7689), .ZN(n7688) );
  INV_X1 U7751 ( .A(n9441), .ZN(n7689) );
  INV_X1 U7752 ( .A(n13288), .ZN(n9058) );
  INV_X1 U7753 ( .A(n13277), .ZN(n13282) );
  NAND2_X1 U7754 ( .A1(n6988), .A2(n8949), .ZN(n8965) );
  NAND2_X1 U7755 ( .A1(n9310), .A2(n9311), .ZN(n13277) );
  NAND2_X1 U7756 ( .A1(n13315), .A2(n9408), .ZN(n13300) );
  INV_X1 U7757 ( .A(n7205), .ZN(n7204) );
  AOI21_X1 U7758 ( .B1(n7150), .B2(n7152), .A(n7148), .ZN(n7147) );
  INV_X1 U7759 ( .A(n9350), .ZN(n7148) );
  OR2_X1 U7760 ( .A1(n8734), .A2(n7158), .ZN(n7154) );
  INV_X1 U7761 ( .A(n12617), .ZN(n7158) );
  NAND2_X1 U7762 ( .A1(n12522), .A2(n7747), .ZN(n12620) );
  NOR2_X1 U7763 ( .A1(n12617), .A2(n7748), .ZN(n7747) );
  INV_X1 U7764 ( .A(n9034), .ZN(n7748) );
  OR2_X1 U7765 ( .A1(n12615), .A2(n13097), .ZN(n9364) );
  INV_X1 U7766 ( .A(n7718), .ZN(n7717) );
  OAI21_X1 U7767 ( .B1(n6478), .B2(n6449), .A(n9361), .ZN(n7718) );
  INV_X1 U7768 ( .A(n9288), .ZN(n8886) );
  INV_X1 U7769 ( .A(n9168), .ZN(n8885) );
  AND3_X1 U7770 ( .A1(n9130), .A2(n11851), .A3(n9129), .ZN(n11325) );
  NAND2_X1 U7771 ( .A1(n9093), .A2(n9104), .ZN(n10821) );
  NAND2_X1 U7772 ( .A1(n8903), .A2(n8902), .ZN(n6782) );
  NAND2_X1 U7773 ( .A1(n9002), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U7774 ( .A1(n7652), .A2(n7650), .ZN(n8812) );
  NAND2_X1 U7775 ( .A1(n8654), .A2(n8653), .ZN(n8656) );
  NAND2_X1 U7776 ( .A1(n7130), .A2(n8566), .ZN(n8583) );
  AND2_X1 U7777 ( .A1(n8584), .A2(n8567), .ZN(n8582) );
  NAND2_X1 U7778 ( .A1(n13649), .A2(n8220), .ZN(n6923) );
  INV_X1 U7779 ( .A(n11837), .ZN(n7585) );
  NAND2_X1 U7780 ( .A1(n6923), .A2(n6921), .ZN(n13673) );
  NOR2_X1 U7781 ( .A1(n8219), .A2(n6922), .ZN(n6921) );
  INV_X1 U7782 ( .A(n13674), .ZN(n6922) );
  NOR2_X1 U7783 ( .A1(n8524), .A2(n15560), .ZN(n8521) );
  INV_X1 U7784 ( .A(n8525), .ZN(n10899) );
  AND4_X1 U7785 ( .A1(n8069), .A2(n8068), .A3(n8067), .A4(n8066), .ZN(n13837)
         );
  OR2_X1 U7786 ( .A1(n10380), .A2(n11793), .ZN(n7903) );
  AND2_X1 U7787 ( .A1(n7911), .A2(n7914), .ZN(n7560) );
  AND2_X1 U7788 ( .A1(n7913), .A2(n7912), .ZN(n6767) );
  NOR2_X1 U7789 ( .A1(n14223), .A2(n14222), .ZN(n14238) );
  NAND2_X1 U7790 ( .A1(n14254), .A2(n14253), .ZN(n14256) );
  INV_X1 U7791 ( .A(n10098), .ZN(n10025) );
  INV_X1 U7792 ( .A(n10008), .ZN(n6885) );
  NAND2_X1 U7793 ( .A1(n14299), .A2(n14300), .ZN(n7687) );
  NAND2_X1 U7794 ( .A1(n7687), .A2(n7685), .ZN(n10109) );
  NOR2_X1 U7795 ( .A1(n14068), .A2(n7686), .ZN(n7685) );
  INV_X1 U7796 ( .A(n10086), .ZN(n7686) );
  AOI21_X1 U7797 ( .B1(n7784), .B2(n7781), .A(n6536), .ZN(n7780) );
  INV_X1 U7798 ( .A(n6476), .ZN(n7781) );
  XNOR2_X1 U7799 ( .A(n14629), .B(n14085), .ZN(n14332) );
  NAND2_X1 U7800 ( .A1(n14391), .A2(n10075), .ZN(n7684) );
  NAND2_X1 U7801 ( .A1(n7759), .A2(n6524), .ZN(n14381) );
  AOI21_X1 U7802 ( .B1(n7678), .B2(n14493), .A(n6529), .ZN(n7677) );
  NAND2_X1 U7803 ( .A1(n7676), .A2(n12712), .ZN(n7675) );
  NAND2_X1 U7804 ( .A1(n11999), .A2(n6768), .ZN(n12182) );
  NOR2_X1 U7805 ( .A1(n12185), .A2(n6769), .ZN(n6768) );
  INV_X1 U7806 ( .A(n10060), .ZN(n6769) );
  NAND2_X1 U7807 ( .A1(n12002), .A2(n6450), .ZN(n6896) );
  OR2_X1 U7808 ( .A1(n14109), .A2(n11081), .ZN(n9968) );
  NAND2_X1 U7809 ( .A1(n10088), .A2(n10087), .ZN(n14481) );
  OR2_X1 U7810 ( .A1(n10876), .A2(n10374), .ZN(n8060) );
  INV_X1 U7811 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7840) );
  OR2_X1 U7812 ( .A1(n7951), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U7813 ( .A1(n10643), .A2(n12148), .ZN(n10465) );
  INV_X1 U7814 ( .A(n9519), .ZN(n9911) );
  NAND2_X1 U7815 ( .A1(n11824), .A2(n11823), .ZN(n7444) );
  INV_X1 U7816 ( .A(n15029), .ZN(n15032) );
  NOR2_X1 U7817 ( .A1(n7424), .A2(n7486), .ZN(n7485) );
  INV_X1 U7818 ( .A(n12869), .ZN(n7486) );
  NAND2_X1 U7819 ( .A1(n7461), .A2(n15069), .ZN(n6919) );
  NAND2_X1 U7820 ( .A1(n15087), .A2(n15086), .ZN(n6920) );
  OAI21_X1 U7821 ( .B1(n6862), .B2(n6859), .A(n6857), .ZN(n12069) );
  INV_X1 U7822 ( .A(n6858), .ZN(n6857) );
  OAI21_X1 U7823 ( .B1(n6860), .B2(n6859), .A(n12074), .ZN(n6858) );
  INV_X1 U7824 ( .A(n9607), .ZN(n6859) );
  NAND2_X1 U7825 ( .A1(n6862), .A2(n6860), .ZN(n11732) );
  OR2_X1 U7826 ( .A1(n11805), .A2(n11952), .ZN(n9580) );
  NAND2_X1 U7827 ( .A1(n6843), .A2(n10135), .ZN(n6842) );
  INV_X1 U7828 ( .A(n9517), .ZN(n6843) );
  OR2_X1 U7829 ( .A1(n9506), .A2(n14855), .ZN(n9517) );
  INV_X1 U7830 ( .A(n15190), .ZN(n15166) );
  INV_X1 U7831 ( .A(n15192), .ZN(n15168) );
  AND2_X1 U7832 ( .A1(n15147), .A2(n15507), .ZN(n15353) );
  NOR2_X1 U7833 ( .A1(n9472), .A2(n9471), .ZN(n7391) );
  NOR2_X1 U7834 ( .A1(n9937), .A2(n7388), .ZN(n9495) );
  NAND2_X1 U7835 ( .A1(n9479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9940) );
  INV_X1 U7836 ( .A(n9942), .ZN(n7626) );
  NAND2_X1 U7837 ( .A1(n9939), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n9941) );
  NAND2_X1 U7838 ( .A1(n8342), .A2(n8378), .ZN(n6682) );
  OR2_X1 U7839 ( .A1(n7120), .A2(n12451), .ZN(n6963) );
  NAND2_X1 U7840 ( .A1(n7248), .A2(n15410), .ZN(n6969) );
  NOR2_X1 U7841 ( .A1(n7248), .A2(n15410), .ZN(n6970) );
  NAND2_X1 U7842 ( .A1(n6555), .A2(n7194), .ZN(n11331) );
  NOR2_X1 U7843 ( .A1(n7195), .A2(n6510), .ZN(n7194) );
  NOR2_X1 U7844 ( .A1(n10405), .A2(n10404), .ZN(n10406) );
  NOR2_X1 U7845 ( .A1(n10403), .A2(n13048), .ZN(n10404) );
  AOI21_X1 U7846 ( .B1(n11837), .B2(n7584), .A(n7583), .ZN(n7582) );
  INV_X1 U7847 ( .A(n8051), .ZN(n7584) );
  INV_X1 U7848 ( .A(n8071), .ZN(n7583) );
  NAND2_X1 U7849 ( .A1(n11410), .A2(n11409), .ZN(n11582) );
  OR2_X1 U7850 ( .A1(n11585), .A2(n11586), .ZN(n7269) );
  OAI21_X1 U7851 ( .B1(n14278), .B2(n15529), .A(n7282), .ZN(n6771) );
  INV_X1 U7852 ( .A(n15543), .ZN(n7283) );
  INV_X1 U7853 ( .A(n11987), .ZN(n9506) );
  AND2_X1 U7854 ( .A1(n9834), .A2(n9833), .ZN(n15045) );
  INV_X1 U7855 ( .A(n15045), .ZN(n14835) );
  NAND2_X1 U7856 ( .A1(n14983), .A2(n14982), .ZN(n6683) );
  NAND2_X1 U7857 ( .A1(n7419), .A2(n7417), .ZN(n15009) );
  OR2_X1 U7858 ( .A1(n7247), .A2(n11776), .ZN(n7244) );
  NOR2_X1 U7859 ( .A1(n11776), .A2(n15726), .ZN(n7246) );
  NAND2_X1 U7860 ( .A1(n7243), .A2(n7121), .ZN(n7120) );
  NAND2_X1 U7861 ( .A1(n15407), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7243) );
  AND2_X1 U7862 ( .A1(n7247), .A2(n11776), .ZN(n7121) );
  NAND2_X1 U7863 ( .A1(n13809), .A2(n6502), .ZN(n7308) );
  INV_X1 U7864 ( .A(n13841), .ZN(n7319) );
  INV_X1 U7865 ( .A(n13844), .ZN(n7312) );
  INV_X1 U7866 ( .A(n7316), .ZN(n7315) );
  OAI21_X1 U7867 ( .B1(n13843), .B2(n13842), .A(n7317), .ZN(n7316) );
  NAND2_X1 U7868 ( .A1(n6543), .A2(n7319), .ZN(n7317) );
  NAND2_X1 U7869 ( .A1(n13844), .A2(n13832), .ZN(n7314) );
  NOR2_X1 U7870 ( .A1(n7319), .A2(n6543), .ZN(n7318) );
  INV_X1 U7871 ( .A(n13861), .ZN(n7303) );
  NAND2_X1 U7872 ( .A1(n7302), .A2(n7301), .ZN(n7300) );
  INV_X1 U7873 ( .A(n13863), .ZN(n7301) );
  INV_X1 U7874 ( .A(n13862), .ZN(n7302) );
  NAND2_X1 U7875 ( .A1(n7303), .A2(n6475), .ZN(n7298) );
  NAND2_X1 U7876 ( .A1(n10162), .A2(n10163), .ZN(n10161) );
  NAND2_X1 U7877 ( .A1(n13883), .A2(n7291), .ZN(n7290) );
  OAI21_X1 U7878 ( .B1(n12098), .B2(n7610), .A(n7608), .ZN(n13923) );
  INV_X1 U7879 ( .A(n8275), .ZN(n7610) );
  NAND2_X1 U7880 ( .A1(n10169), .A2(n10171), .ZN(n7552) );
  NAND2_X1 U7881 ( .A1(n10172), .A2(n10175), .ZN(n6880) );
  INV_X1 U7882 ( .A(n10172), .ZN(n6881) );
  AND2_X1 U7883 ( .A1(n7225), .A2(n9368), .ZN(n7224) );
  NAND2_X1 U7884 ( .A1(n9384), .A2(n7216), .ZN(n7215) );
  NAND2_X1 U7885 ( .A1(n7218), .A2(n9378), .ZN(n7216) );
  AND2_X1 U7886 ( .A1(n7219), .A2(n9378), .ZN(n7217) );
  NAND2_X1 U7887 ( .A1(n7547), .A2(n7546), .ZN(n10192) );
  NAND2_X1 U7888 ( .A1(n10183), .A2(n10185), .ZN(n7546) );
  NAND2_X1 U7889 ( .A1(n10192), .A2(n10186), .ZN(n6840) );
  NAND2_X1 U7890 ( .A1(n10231), .A2(n6873), .ZN(n6872) );
  INV_X1 U7891 ( .A(n10234), .ZN(n6873) );
  INV_X1 U7892 ( .A(n10235), .ZN(n7554) );
  MUX2_X1 U7893 ( .A(n9406), .B(n9405), .S(n9421), .Z(n9407) );
  NAND2_X1 U7894 ( .A1(n6814), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6813) );
  INV_X1 U7895 ( .A(n11225), .ZN(n6818) );
  NAND2_X1 U7896 ( .A1(n11137), .A2(n11224), .ZN(n6819) );
  INV_X1 U7897 ( .A(n13106), .ZN(n9018) );
  INV_X1 U7898 ( .A(n8824), .ZN(n7649) );
  INV_X1 U7899 ( .A(n13999), .ZN(n6740) );
  INV_X1 U7900 ( .A(n14000), .ZN(n6739) );
  NAND3_X1 U7901 ( .A1(n7305), .A2(n7304), .A3(n6494), .ZN(n6744) );
  AOI21_X1 U7902 ( .B1(n13999), .B2(n14000), .A(n6557), .ZN(n6742) );
  INV_X1 U7903 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6655) );
  AND2_X1 U7904 ( .A1(n7519), .A2(n7517), .ZN(n10272) );
  NOR2_X1 U7905 ( .A1(n6481), .A2(n7477), .ZN(n7476) );
  INV_X1 U7906 ( .A(n7481), .ZN(n7477) );
  NOR2_X1 U7907 ( .A1(n6689), .A2(n8423), .ZN(n6688) );
  INV_X1 U7908 ( .A(n8408), .ZN(n6689) );
  AOI21_X1 U7909 ( .B1(n6558), .B2(n8382), .A(n6465), .ZN(n7328) );
  INV_X1 U7910 ( .A(n8382), .ZN(n7329) );
  NOR2_X1 U7911 ( .A1(n8291), .A2(SI_18_), .ZN(n8296) );
  NOR2_X1 U7912 ( .A1(n8294), .A2(n8293), .ZN(n8295) );
  NAND2_X1 U7913 ( .A1(n6747), .A2(n6477), .ZN(n7341) );
  NAND2_X1 U7914 ( .A1(n7007), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7006) );
  OAI21_X1 U7915 ( .B1(n7944), .B2(n10841), .A(n7073), .ZN(n7945) );
  NAND2_X1 U7916 ( .A1(n7944), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7073) );
  NAND2_X1 U7917 ( .A1(n7945), .A2(SI_5_), .ZN(n7971) );
  NAND2_X1 U7918 ( .A1(n7944), .A2(n10854), .ZN(n6714) );
  NAND2_X1 U7919 ( .A1(n7944), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7074) );
  INV_X1 U7920 ( .A(n11818), .ZN(n9456) );
  NAND2_X1 U7921 ( .A1(n7095), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9174) );
  NOR2_X1 U7922 ( .A1(n11187), .A2(n9178), .ZN(n9179) );
  NOR2_X1 U7923 ( .A1(n11475), .A2(n9146), .ZN(n9147) );
  AND2_X1 U7924 ( .A1(n11488), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U7925 ( .A1(n7365), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U7926 ( .A1(n10800), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7055) );
  INV_X1 U7927 ( .A(n6832), .ZN(n6830) );
  AND2_X1 U7928 ( .A1(n6829), .A2(n6828), .ZN(n6827) );
  NAND2_X1 U7929 ( .A1(n6833), .A2(n13160), .ZN(n6829) );
  NOR2_X1 U7930 ( .A1(n6632), .A2(n13478), .ZN(n6833) );
  NAND2_X1 U7931 ( .A1(n10687), .A2(n7065), .ZN(n9159) );
  AND2_X1 U7932 ( .A1(n13220), .A2(n6473), .ZN(n7521) );
  NAND2_X1 U7933 ( .A1(n13172), .A2(n9161), .ZN(n9162) );
  NOR2_X1 U7934 ( .A1(n8978), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n6989) );
  NOR2_X1 U7935 ( .A1(n8933), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n6988) );
  OR2_X1 U7936 ( .A1(n13520), .A2(n12927), .ZN(n9311) );
  NOR2_X1 U7937 ( .A1(n8873), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n6987) );
  NOR2_X1 U7938 ( .A1(n8889), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7128) );
  NOR2_X1 U7939 ( .A1(n8819), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8833) );
  OR2_X1 U7940 ( .A1(n8713), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U7941 ( .A1(n9328), .A2(n9026), .ZN(n7197) );
  NOR2_X1 U7942 ( .A1(n7201), .A2(n7200), .ZN(n7199) );
  INV_X1 U7943 ( .A(n9026), .ZN(n7201) );
  INV_X1 U7944 ( .A(n9025), .ZN(n7200) );
  NAND2_X1 U7945 ( .A1(n7159), .A2(n7160), .ZN(n9000) );
  AND2_X1 U7946 ( .A1(n9049), .A2(n7740), .ZN(n7739) );
  NAND2_X1 U7947 ( .A1(n7742), .A2(n9043), .ZN(n7740) );
  OR2_X1 U7948 ( .A1(n13546), .A2(n13089), .ZN(n9399) );
  NAND2_X1 U7949 ( .A1(n9010), .A2(n9071), .ZN(n11307) );
  INV_X1 U7950 ( .A(n9377), .ZN(n7704) );
  OR2_X1 U7951 ( .A1(n12632), .A2(n12589), .ZN(n9370) );
  OR2_X1 U7952 ( .A1(n12955), .A2(n13098), .ZN(n9361) );
  INV_X1 U7953 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8551) );
  NOR2_X1 U7954 ( .A1(n8986), .A2(n7661), .ZN(n7660) );
  INV_X1 U7955 ( .A(n8975), .ZN(n7661) );
  INV_X1 U7956 ( .A(n8973), .ZN(n7658) );
  NAND2_X1 U7957 ( .A1(n9004), .A2(n7805), .ZN(n9089) );
  NOR2_X1 U7958 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n8541) );
  INV_X1 U7959 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7503) );
  NOR2_X1 U7960 ( .A1(n8800), .A2(n7651), .ZN(n7650) );
  INV_X1 U7961 ( .A(n8796), .ZN(n7651) );
  INV_X1 U7962 ( .A(n8781), .ZN(n7168) );
  NOR2_X1 U7963 ( .A1(n8760), .A2(n8759), .ZN(n8762) );
  INV_X1 U7964 ( .A(n8659), .ZN(n8658) );
  NAND2_X1 U7965 ( .A1(n10852), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8665) );
  INV_X1 U7966 ( .A(n8584), .ZN(n6799) );
  NAND2_X1 U7967 ( .A1(n10864), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8600) );
  INV_X1 U7968 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8555) );
  OR3_X1 U7969 ( .A1(n8432), .A2(n13736), .A3(n8431), .ZN(n8453) );
  NAND2_X1 U7970 ( .A1(n7141), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8432) );
  INV_X1 U7971 ( .A(n7784), .ZN(n7782) );
  XNOR2_X1 U7972 ( .A(n14536), .B(n14086), .ZN(n14347) );
  NAND2_X1 U7973 ( .A1(n14057), .A2(n6758), .ZN(n6757) );
  INV_X1 U7974 ( .A(n12407), .ZN(n6758) );
  INV_X1 U7975 ( .A(n11749), .ZN(n6752) );
  INV_X1 U7976 ( .A(n10054), .ZN(n6753) );
  NAND2_X1 U7977 ( .A1(n13791), .A2(n9971), .ZN(n11570) );
  NAND2_X1 U7978 ( .A1(n7773), .A2(n7771), .ZN(n14464) );
  OR2_X1 U7979 ( .A1(n8251), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8091) );
  NOR2_X1 U7980 ( .A1(n10304), .A2(n10279), .ZN(n10303) );
  NOR2_X1 U7981 ( .A1(n10246), .A2(n10247), .ZN(n6865) );
  NAND2_X1 U7982 ( .A1(n7105), .A2(n6867), .ZN(n6866) );
  AND2_X1 U7983 ( .A1(n7555), .A2(n6868), .ZN(n6867) );
  NAND2_X1 U7984 ( .A1(n10246), .A2(n10247), .ZN(n6868) );
  NOR2_X1 U7985 ( .A1(n11616), .A2(n7447), .ZN(n7443) );
  NAND2_X1 U7986 ( .A1(n12677), .A2(n6522), .ZN(n12796) );
  NAND2_X1 U7987 ( .A1(n12866), .A2(n9902), .ZN(n7382) );
  NAND2_X1 U7988 ( .A1(n15270), .A2(n15365), .ZN(n6717) );
  NOR2_X1 U7989 ( .A1(n9780), .A2(n14792), .ZN(n7139) );
  NOR2_X1 U7990 ( .A1(n15307), .A2(n15115), .ZN(n7462) );
  NAND2_X1 U7991 ( .A1(n15138), .A2(n15119), .ZN(n6934) );
  AND2_X1 U7992 ( .A1(n15123), .A2(n6933), .ZN(n6932) );
  INV_X1 U7993 ( .A(n15121), .ZN(n6933) );
  NAND2_X1 U7994 ( .A1(n15137), .A2(n9741), .ZN(n9742) );
  INV_X1 U7995 ( .A(n9892), .ZN(n6931) );
  NAND2_X1 U7996 ( .A1(n9892), .A2(n12243), .ZN(n6930) );
  INV_X1 U7997 ( .A(n9893), .ZN(n7370) );
  NOR2_X1 U7998 ( .A1(n15503), .A2(n11424), .ZN(n7456) );
  NAND2_X1 U7999 ( .A1(n14853), .A2(n12148), .ZN(n10135) );
  INV_X1 U8000 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U8001 ( .A1(n9862), .A2(n7056), .ZN(n7639) );
  NOR2_X1 U8002 ( .A1(n7639), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U8003 ( .A1(n8030), .A2(SI_8_), .ZN(n8055) );
  NOR2_X1 U8004 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  NAND3_X1 U8005 ( .A1(n8001), .A2(n8000), .A3(n7999), .ZN(n8008) );
  NAND2_X1 U8006 ( .A1(n8056), .A2(SI_9_), .ZN(n8072) );
  AND2_X1 U8007 ( .A1(n7970), .A2(n7972), .ZN(n7999) );
  OAI21_X1 U8008 ( .B1(n7974), .B2(SI_6_), .A(n8004), .ZN(n8003) );
  NAND2_X1 U8009 ( .A1(n7923), .A2(SI_4_), .ZN(n6918) );
  OAI21_X1 U8010 ( .B1(n7945), .B2(SI_5_), .A(n7971), .ZN(n7969) );
  INV_X1 U8011 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U8012 ( .A1(n10776), .A2(n10814), .ZN(n10815) );
  NAND2_X1 U8013 ( .A1(n10964), .A2(n10963), .ZN(n11097) );
  NAND2_X1 U8014 ( .A1(n12092), .A2(n12093), .ZN(n12455) );
  NAND2_X1 U8015 ( .A1(n13019), .A2(n13018), .ZN(n13020) );
  NAND2_X1 U8016 ( .A1(n6653), .A2(n11549), .ZN(n11561) );
  INV_X1 U8017 ( .A(n11563), .ZN(n6653) );
  NAND2_X1 U8018 ( .A1(n11561), .A2(n6708), .ZN(n11687) );
  AND2_X1 U8019 ( .A1(n11552), .A2(n11551), .ZN(n6708) );
  AND2_X1 U8020 ( .A1(n13029), .A2(n7495), .ZN(n7494) );
  OR2_X1 U8021 ( .A1(n12962), .A2(n7496), .ZN(n7495) );
  INV_X1 U8022 ( .A(n12915), .ZN(n7496) );
  AOI22_X1 U8023 ( .A1(n12583), .A2(n12582), .B1(n12581), .B2(n12580), .ZN(
        n12584) );
  XNOR2_X1 U8024 ( .A(n13532), .B(n7186), .ZN(n12937) );
  INV_X1 U8025 ( .A(n13048), .ZN(n13059) );
  NAND2_X1 U8026 ( .A1(n13602), .A2(n9287), .ZN(n6807) );
  NAND2_X1 U8027 ( .A1(n12899), .A2(n12898), .ZN(n6643) );
  NOR2_X1 U8028 ( .A1(n13505), .A2(n9448), .ZN(n9450) );
  NAND2_X1 U8029 ( .A1(n9259), .A2(n9258), .ZN(n9284) );
  AND4_X1 U8030 ( .A1(n8699), .A2(n8698), .A3(n8697), .A4(n8696), .ZN(n12559)
         );
  AND4_X1 U8031 ( .A1(n8630), .A2(n8629), .A3(n8628), .A4(n8627), .ZN(n8639)
         );
  NAND2_X1 U8032 ( .A1(n8546), .A2(n7508), .ZN(n7507) );
  NOR2_X1 U8033 ( .A1(n7509), .A2(n11334), .ZN(n7508) );
  XNOR2_X1 U8034 ( .A(n8543), .B(n13588), .ZN(n8545) );
  NAND2_X1 U8035 ( .A1(n13587), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8543) );
  NOR2_X1 U8036 ( .A1(n11215), .A2(n15596), .ZN(n11214) );
  OAI21_X1 U8037 ( .B1(n9173), .B2(n9139), .A(n9140), .ZN(n11211) );
  NOR2_X1 U8038 ( .A1(n11211), .A2(n11212), .ZN(n11210) );
  OR2_X1 U8039 ( .A1(n11184), .A2(n11185), .ZN(n6815) );
  AND2_X1 U8040 ( .A1(n9182), .A2(n11160), .ZN(n7107) );
  AOI21_X1 U8041 ( .B1(n11152), .B2(n11476), .A(n11477), .ZN(n11475) );
  INV_X1 U8042 ( .A(n6917), .ZN(n9184) );
  NAND2_X1 U8043 ( .A1(n9147), .A2(n11388), .ZN(n7365) );
  NOR2_X1 U8044 ( .A1(n11455), .A2(n7363), .ZN(n11454) );
  OR2_X1 U8045 ( .A1(n9185), .A2(n11891), .ZN(n9186) );
  OR2_X1 U8046 ( .A1(n11893), .A2(n11892), .ZN(n11895) );
  NAND2_X1 U8047 ( .A1(n7516), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7515) );
  INV_X1 U8048 ( .A(n9153), .ZN(n9154) );
  NOR2_X1 U8049 ( .A1(n10707), .A2(n9218), .ZN(n12387) );
  NAND2_X1 U8050 ( .A1(n9188), .A2(n10826), .ZN(n13115) );
  NAND2_X1 U8051 ( .A1(n9155), .A2(n13110), .ZN(n13109) );
  NAND2_X1 U8052 ( .A1(n12393), .A2(n7350), .ZN(n9155) );
  NAND2_X1 U8053 ( .A1(n7358), .A2(n10684), .ZN(n13131) );
  INV_X1 U8054 ( .A(n7359), .ZN(n7358) );
  NAND2_X1 U8055 ( .A1(n13139), .A2(n6606), .ZN(n13136) );
  NAND2_X1 U8056 ( .A1(n6912), .A2(n9225), .ZN(n10692) );
  NAND2_X1 U8057 ( .A1(n6911), .A2(n10689), .ZN(n6912) );
  INV_X1 U8058 ( .A(n9159), .ZN(n7064) );
  NOR2_X1 U8059 ( .A1(n13156), .A2(n13155), .ZN(n13154) );
  NAND2_X1 U8060 ( .A1(n7250), .A2(n7255), .ZN(n13190) );
  AOI21_X1 U8061 ( .B1(n7257), .B2(n7256), .A(n6625), .ZN(n7255) );
  NAND2_X1 U8062 ( .A1(n7521), .A2(n7526), .ZN(n7523) );
  NAND2_X1 U8063 ( .A1(n7520), .A2(n7525), .ZN(n7522) );
  OR2_X1 U8064 ( .A1(n9393), .A2(n9073), .ZN(n13048) );
  NAND2_X1 U8065 ( .A1(n13281), .A2(n13282), .ZN(n8972) );
  NAND2_X1 U8066 ( .A1(n13520), .A2(n12927), .ZN(n9310) );
  INV_X1 U8067 ( .A(n13279), .ZN(n6783) );
  NAND2_X1 U8068 ( .A1(n7212), .A2(n7211), .ZN(n13276) );
  AOI21_X1 U8069 ( .B1(n13300), .B2(n8941), .A(n7797), .ZN(n13290) );
  NOR2_X1 U8070 ( .A1(n9313), .A2(n13304), .ZN(n7797) );
  OR2_X1 U8071 ( .A1(n13532), .A2(n12941), .ZN(n13299) );
  INV_X1 U8072 ( .A(n9050), .ZN(n7206) );
  INV_X1 U8073 ( .A(n9412), .ZN(n13304) );
  OR2_X1 U8074 ( .A1(n8922), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8933) );
  INV_X1 U8075 ( .A(n6987), .ZN(n8908) );
  NAND2_X1 U8076 ( .A1(n8767), .A2(n8766), .ZN(n8785) );
  INV_X1 U8077 ( .A(n8768), .ZN(n8767) );
  NAND2_X1 U8078 ( .A1(n6986), .A2(n6985), .ZN(n8694) );
  INV_X1 U8079 ( .A(n8675), .ZN(n6986) );
  NAND2_X1 U8080 ( .A1(n8681), .A2(n9354), .ZN(n12271) );
  XNOR2_X1 U8081 ( .A(n13101), .B(n12110), .ZN(n12173) );
  NAND2_X1 U8082 ( .A1(n12132), .A2(n12134), .ZN(n8623) );
  NAND2_X1 U8083 ( .A1(n12028), .A2(n8590), .ZN(n7693) );
  NAND2_X1 U8084 ( .A1(n8602), .A2(n7166), .ZN(n9337) );
  INV_X1 U8085 ( .A(n7167), .ZN(n7166) );
  OAI22_X1 U8086 ( .A1(n9288), .A2(SI_4_), .B1(n9168), .B2(n11236), .ZN(n7167)
         );
  AND2_X1 U8087 ( .A1(n9326), .A2(n9329), .ZN(n12030) );
  INV_X1 U8088 ( .A(n11675), .ZN(n11671) );
  NAND2_X1 U8089 ( .A1(n9000), .A2(n9418), .ZN(n9442) );
  AND2_X1 U8090 ( .A1(n13250), .A2(n10398), .ZN(n7746) );
  NAND2_X1 U8091 ( .A1(n7145), .A2(n7116), .ZN(n13315) );
  AND2_X1 U8092 ( .A1(n7707), .A2(n9406), .ZN(n7116) );
  NAND2_X1 U8093 ( .A1(n13390), .A2(n7708), .ZN(n7145) );
  NAND2_X1 U8094 ( .A1(n7738), .A2(n7739), .ZN(n13336) );
  OR2_X1 U8095 ( .A1(n13543), .A2(n13335), .ZN(n13327) );
  NAND2_X1 U8096 ( .A1(n13390), .A2(n8839), .ZN(n7714) );
  OR2_X1 U8097 ( .A1(n6605), .A2(n7790), .ZN(n7798) );
  NOR2_X1 U8098 ( .A1(n8791), .A2(n7706), .ZN(n7705) );
  NAND2_X1 U8099 ( .A1(n7154), .A2(n6509), .ZN(n8774) );
  INV_X1 U8100 ( .A(n9374), .ZN(n7153) );
  INV_X1 U8101 ( .A(n9369), .ZN(n12749) );
  AOI21_X1 U8102 ( .B1(n12617), .B2(n7157), .A(n7156), .ZN(n7155) );
  INV_X1 U8103 ( .A(n9371), .ZN(n7156) );
  INV_X1 U8104 ( .A(n9364), .ZN(n7157) );
  AOI21_X1 U8105 ( .B1(n7717), .B2(n6449), .A(n12523), .ZN(n7716) );
  NAND2_X1 U8106 ( .A1(n7191), .A2(n7190), .ZN(n12522) );
  AOI21_X1 U8107 ( .B1(n7193), .B2(n7752), .A(n6554), .ZN(n7190) );
  NAND2_X1 U8108 ( .A1(n12044), .A2(n6443), .ZN(n7192) );
  INV_X1 U8109 ( .A(n9354), .ZN(n7721) );
  INV_X1 U8110 ( .A(n15621), .ZN(n15614) );
  NAND2_X1 U8111 ( .A1(n9095), .A2(n9094), .ZN(n11851) );
  OAI21_X1 U8112 ( .B1(n10821), .B2(P3_D_REG_0__SCAN_IN), .A(n9097), .ZN(n9130) );
  NAND2_X1 U8113 ( .A1(n8944), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6809) );
  OR2_X1 U8114 ( .A1(n9007), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n9098) );
  INV_X1 U8115 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n6990) );
  INV_X1 U8116 ( .A(n8868), .ZN(n6991) );
  NAND2_X1 U8117 ( .A1(n8812), .A2(n8811), .ZN(n8815) );
  NAND2_X1 U8118 ( .A1(n8815), .A2(n8814), .ZN(n8825) );
  NAND2_X1 U8119 ( .A1(n8756), .A2(n7653), .ZN(n7652) );
  NOR2_X1 U8120 ( .A1(n8797), .A2(n7654), .ZN(n7653) );
  INV_X1 U8121 ( .A(n8755), .ZN(n7654) );
  NAND2_X1 U8122 ( .A1(n7168), .A2(n9082), .ZN(n9090) );
  NAND2_X1 U8123 ( .A1(n6786), .A2(n6784), .ZN(n8754) );
  AND2_X1 U8124 ( .A1(n6785), .A2(n7641), .ZN(n6784) );
  NAND2_X1 U8125 ( .A1(n8686), .A2(n6787), .ZN(n6786) );
  AOI21_X1 U8126 ( .B1(n7642), .B2(n7644), .A(n6617), .ZN(n7641) );
  AND2_X1 U8127 ( .A1(n8720), .A2(n8702), .ZN(n8703) );
  NAND2_X1 U8128 ( .A1(n8701), .A2(n8700), .ZN(n8704) );
  NAND2_X1 U8129 ( .A1(n8704), .A2(n8703), .ZN(n8721) );
  INV_X1 U8130 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n6645) );
  INV_X1 U8131 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n6644) );
  OR2_X1 U8132 ( .A1(n8706), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U8133 ( .A1(n8635), .A2(n8634), .ZN(n8654) );
  NAND2_X1 U8134 ( .A1(n10854), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8584) );
  OR3_X1 U8135 ( .A1(n12671), .A2(n12481), .A3(n12225), .ZN(n10682) );
  INV_X1 U8136 ( .A(n7140), .ZN(n8165) );
  NAND2_X1 U8137 ( .A1(n6564), .A2(n7574), .ZN(n6937) );
  NAND2_X1 U8138 ( .A1(n13685), .A2(n6939), .ZN(n6938) );
  INV_X1 U8139 ( .A(n7998), .ZN(n7562) );
  AOI21_X1 U8140 ( .B1(n13634), .B2(n8341), .A(n6925), .ZN(n13614) );
  INV_X1 U8141 ( .A(n8290), .ZN(n7570) );
  NAND2_X1 U8142 ( .A1(n6976), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8363) );
  INV_X1 U8143 ( .A(n11979), .ZN(n7580) );
  NAND2_X1 U8144 ( .A1(n6676), .A2(n8050), .ZN(n11721) );
  INV_X1 U8145 ( .A(n14108), .ZN(n11434) );
  INV_X1 U8146 ( .A(n14073), .ZN(n13732) );
  NAND2_X1 U8147 ( .A1(n7587), .A2(n8175), .ZN(n7586) );
  NOR2_X1 U8148 ( .A1(n7588), .A2(n6675), .ZN(n6674) );
  XNOR2_X1 U8149 ( .A(n7136), .B(n14031), .ZN(n7039) );
  NAND2_X1 U8150 ( .A1(n14036), .A2(n7138), .ZN(n7137) );
  AND2_X1 U8151 ( .A1(n8236), .A2(n8235), .ZN(n13896) );
  AND4_X1 U8152 ( .A1(n8083), .A2(n8082), .A3(n8081), .A4(n8080), .ZN(n13848)
         );
  AND4_X1 U8153 ( .A1(n8022), .A2(n8021), .A3(n8020), .A4(n8019), .ZN(n13820)
         );
  NAND2_X1 U8154 ( .A1(n14213), .A2(n12259), .ZN(n12765) );
  NOR2_X1 U8155 ( .A1(n14238), .A2(n6630), .ZN(n14240) );
  NAND2_X1 U8156 ( .A1(n6780), .A2(n6779), .ZN(n7277) );
  INV_X1 U8157 ( .A(n14239), .ZN(n6779) );
  INV_X1 U8158 ( .A(n14240), .ZN(n6780) );
  NAND2_X1 U8159 ( .A1(n10107), .A2(n14023), .ZN(n7724) );
  INV_X1 U8160 ( .A(n10107), .ZN(n6662) );
  NAND2_X1 U8161 ( .A1(n7734), .A2(n14310), .ZN(n7733) );
  INV_X1 U8162 ( .A(n7735), .ZN(n7734) );
  INV_X1 U8163 ( .A(n14364), .ZN(n7787) );
  INV_X1 U8164 ( .A(n7785), .ZN(n7783) );
  INV_X1 U8165 ( .A(n7782), .ZN(n7777) );
  INV_X1 U8166 ( .A(n14378), .ZN(n10004) );
  NAND2_X1 U8167 ( .A1(n7763), .A2(n13709), .ZN(n7762) );
  NAND2_X1 U8168 ( .A1(n6887), .A2(n6886), .ZN(n10002) );
  AND2_X1 U8169 ( .A1(n6578), .A2(n9999), .ZN(n6886) );
  NAND2_X1 U8170 ( .A1(n6762), .A2(n10074), .ZN(n14391) );
  NAND2_X1 U8171 ( .A1(n6766), .A2(n6763), .ZN(n6762) );
  NAND2_X1 U8172 ( .A1(n9990), .A2(n9989), .ZN(n12498) );
  AND2_X1 U8173 ( .A1(n14055), .A2(n10063), .ZN(n7682) );
  AOI21_X1 U8174 ( .B1(n6450), .B2(n7766), .A(n6492), .ZN(n7764) );
  AND2_X1 U8175 ( .A1(n7758), .A2(n11779), .ZN(n7757) );
  NAND2_X1 U8176 ( .A1(n12002), .A2(n14054), .ZN(n12001) );
  NAND2_X1 U8177 ( .A1(n6891), .A2(n9979), .ZN(n11748) );
  NAND2_X1 U8178 ( .A1(n11534), .A2(n14049), .ZN(n6891) );
  OR2_X1 U8179 ( .A1(n11748), .A2(n14050), .ZN(n11746) );
  NAND2_X1 U8180 ( .A1(n7794), .A2(n7681), .ZN(n7680) );
  NAND2_X1 U8181 ( .A1(n11128), .A2(n13774), .ZN(n11376) );
  NAND2_X1 U8182 ( .A1(n9967), .A2(n9966), .ZN(n11079) );
  AND2_X1 U8183 ( .A1(n10802), .A2(n10801), .ZN(n6893) );
  NAND2_X1 U8184 ( .A1(n10034), .A2(n9965), .ZN(n7070) );
  CLKBUF_X1 U8185 ( .A(n10032), .Z(n14426) );
  NAND2_X1 U8186 ( .A1(n6484), .A2(n10103), .ZN(n10105) );
  XNOR2_X1 U8187 ( .A(n7872), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U8188 ( .A1(n14667), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7872) );
  OR2_X1 U8189 ( .A1(n8010), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8033) );
  AND2_X1 U8190 ( .A1(n7952), .A2(n7977), .ZN(n14159) );
  XNOR2_X1 U8191 ( .A(n6773), .B(P2_IR_REG_4__SCAN_IN), .ZN(n14144) );
  NAND2_X1 U8192 ( .A1(n7947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6773) );
  MUX2_X1 U8193 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7852), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7853) );
  NAND2_X1 U8194 ( .A1(n7134), .A2(n7850), .ZN(n7898) );
  AND2_X1 U8195 ( .A1(n7624), .A2(n14809), .ZN(n7623) );
  OR2_X1 U8196 ( .A1(n14732), .A2(n7625), .ZN(n7624) );
  INV_X1 U8197 ( .A(n10626), .ZN(n7625) );
  NAND2_X1 U8198 ( .A1(n7623), .A2(n6728), .ZN(n6727) );
  INV_X1 U8199 ( .A(n10617), .ZN(n6728) );
  NAND2_X1 U8200 ( .A1(n14800), .A2(n14799), .ZN(n7632) );
  INV_X1 U8201 ( .A(n9722), .ZN(n9723) );
  INV_X1 U8202 ( .A(n7636), .ZN(n7634) );
  AND2_X1 U8203 ( .A1(n7635), .A2(n7638), .ZN(n6726) );
  INV_X1 U8204 ( .A(n10570), .ZN(n7631) );
  AND2_X1 U8205 ( .A1(n6495), .A2(n10583), .ZN(n7615) );
  OR2_X1 U8206 ( .A1(n9528), .A2(n9509), .ZN(n9510) );
  NOR2_X1 U8207 ( .A1(n9496), .A2(n9863), .ZN(n9497) );
  OR2_X1 U8208 ( .A1(n10722), .A2(n7431), .ZN(n7430) );
  NAND2_X1 U8209 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n7431) );
  NOR2_X1 U8210 ( .A1(n10949), .A2(n10948), .ZN(n10947) );
  OR2_X1 U8211 ( .A1(n14866), .A2(n14865), .ZN(n7433) );
  AND2_X1 U8212 ( .A1(n7433), .A2(n7432), .ZN(n14874) );
  NAND2_X1 U8213 ( .A1(n14868), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7432) );
  NAND2_X1 U8214 ( .A1(n14874), .A2(n14873), .ZN(n14872) );
  AOI21_X1 U8215 ( .B1(n14898), .B2(n11268), .A(n11267), .ZN(n14915) );
  NAND2_X1 U8216 ( .A1(n12675), .A2(n7448), .ZN(n12790) );
  OR2_X1 U8217 ( .A1(n12676), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7448) );
  NAND2_X1 U8218 ( .A1(n14931), .A2(n14930), .ZN(n14946) );
  OR2_X1 U8219 ( .A1(n14938), .A2(n7426), .ZN(n7425) );
  OR2_X1 U8220 ( .A1(n14956), .A2(n7428), .ZN(n7426) );
  AND3_X1 U8221 ( .A1(n7425), .A2(n7427), .A3(P1_REG1_REG_18__SCAN_IN), .ZN(
        n14953) );
  INV_X1 U8222 ( .A(n12871), .ZN(n7487) );
  NAND2_X1 U8223 ( .A1(n9835), .A2(n12873), .ZN(n15029) );
  NAND2_X1 U8224 ( .A1(n15044), .A2(n7424), .ZN(n6948) );
  NAND2_X1 U8225 ( .A1(n7376), .A2(n7374), .ZN(n15058) );
  INV_X1 U8226 ( .A(n7378), .ZN(n7374) );
  NAND2_X1 U8227 ( .A1(n15078), .A2(n15090), .ZN(n7379) );
  AND2_X1 U8228 ( .A1(n9764), .A2(n9763), .ZN(n15089) );
  INV_X1 U8229 ( .A(n7051), .ZN(n7413) );
  INV_X1 U8230 ( .A(n9754), .ZN(n7410) );
  NAND2_X1 U8231 ( .A1(n7484), .A2(n9899), .ZN(n15122) );
  NAND2_X1 U8232 ( .A1(n15184), .A2(n7481), .ZN(n7484) );
  NAND2_X1 U8233 ( .A1(n12230), .A2(n10342), .ZN(n6928) );
  INV_X1 U8234 ( .A(n9646), .ZN(n7397) );
  NAND2_X1 U8235 ( .A1(n12158), .A2(n9646), .ZN(n12241) );
  CLKBUF_X1 U8236 ( .A(n12156), .Z(n12158) );
  AOI21_X1 U8237 ( .B1(n7465), .B2(n7468), .A(n11920), .ZN(n7463) );
  INV_X1 U8238 ( .A(n9884), .ZN(n7468) );
  NOR2_X1 U8239 ( .A1(n12148), .A2(n11276), .ZN(n7454) );
  NAND2_X1 U8240 ( .A1(n11167), .A2(n11164), .ZN(n7393) );
  INV_X1 U8241 ( .A(n9920), .ZN(n9921) );
  AOI22_X1 U8242 ( .A1(n14833), .A2(n15190), .B1(n15192), .B2(n15242), .ZN(
        n9920) );
  NAND2_X1 U8243 ( .A1(n10314), .A2(n10313), .ZN(n10317) );
  INV_X1 U8244 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U8245 ( .A1(n8445), .A2(n13604), .ZN(n8444) );
  NAND2_X1 U8246 ( .A1(n8409), .A2(n8408), .ZN(n8424) );
  NAND2_X1 U8247 ( .A1(n8342), .A2(n6511), .ZN(n6749) );
  NAND3_X1 U8248 ( .A1(n8007), .A2(n8008), .A3(n7337), .ZN(n7339) );
  AND2_X1 U8249 ( .A1(n8029), .A2(n8055), .ZN(n7337) );
  AND2_X1 U8250 ( .A1(n8072), .A2(n7018), .ZN(n8057) );
  OR2_X1 U8251 ( .A1(n8056), .A2(SI_9_), .ZN(n7018) );
  INV_X1 U8252 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9473) );
  NOR2_X1 U8253 ( .A1(n9537), .A2(n9536), .ZN(n10931) );
  OAI22_X1 U8254 ( .A1(n6638), .A2(n9535), .B1(P1_IR_REG_31__SCAN_IN), .B2(
        P1_IR_REG_3__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U8255 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6638) );
  NAND2_X1 U8256 ( .A1(n6563), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U8257 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7451) );
  NAND2_X1 U8258 ( .A1(n10883), .A2(n10882), .ZN(n10966) );
  OR2_X1 U8259 ( .A1(n10888), .A2(n15551), .ZN(n6960) );
  OR2_X1 U8260 ( .A1(n10968), .A2(n15551), .ZN(n6958) );
  AND2_X1 U8261 ( .A1(n10888), .A2(n15551), .ZN(n6961) );
  NAND2_X1 U8262 ( .A1(n11095), .A2(n11094), .ZN(n11764) );
  XNOR2_X1 U8263 ( .A(n13016), .B(n13017), .ZN(n13021) );
  AND2_X1 U8264 ( .A1(n8939), .A2(n8938), .ZN(n12942) );
  NAND2_X1 U8265 ( .A1(n12963), .A2(n12962), .ZN(n12961) );
  AND2_X1 U8266 ( .A1(n11310), .A2(n13491), .ZN(n7497) );
  NAND2_X1 U8267 ( .A1(n8948), .A2(n8947), .ZN(n13026) );
  INV_X1 U8268 ( .A(n13543), .ZN(n13334) );
  XNOR2_X1 U8269 ( .A(n12939), .B(n12937), .ZN(n13039) );
  AND3_X1 U8270 ( .A1(n8572), .A2(n8571), .A3(n8570), .ZN(n11345) );
  NOR4_X1 U8271 ( .A1(n10408), .A2(n13250), .A3(n9306), .A4(n9305), .ZN(n9307)
         );
  NOR2_X1 U8272 ( .A1(n6432), .A2(n7079), .ZN(n7078) );
  NAND2_X1 U8273 ( .A1(n9010), .A2(n9436), .ZN(n7079) );
  OAI211_X1 U8274 ( .C1(n7221), .C2(n9425), .A(n7220), .B(n9431), .ZN(n9432)
         );
  NAND2_X1 U8275 ( .A1(n7221), .A2(n6490), .ZN(n7220) );
  INV_X1 U8276 ( .A(n12976), .ZN(n13081) );
  NAND2_X1 U8277 ( .A1(n8985), .A2(n8984), .ZN(n13082) );
  NAND2_X1 U8278 ( .A1(n8957), .A2(n8956), .ZN(n13084) );
  INV_X1 U8279 ( .A(n12942), .ZN(n13085) );
  INV_X1 U8280 ( .A(n12559), .ZN(n13099) );
  NAND2_X1 U8281 ( .A1(n8596), .A2(n6497), .ZN(n13104) );
  XNOR2_X1 U8282 ( .A(n8672), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11460) );
  AND2_X1 U8283 ( .A1(n9210), .A2(n11388), .ZN(n7249) );
  NAND2_X1 U8284 ( .A1(n9157), .A2(n13146), .ZN(n10684) );
  NAND2_X1 U8285 ( .A1(n13109), .A2(n9156), .ZN(n9157) );
  NAND2_X1 U8286 ( .A1(n13109), .A2(n6838), .ZN(n7360) );
  NOR2_X1 U8287 ( .A1(n13146), .A2(n6839), .ZN(n6838) );
  INV_X1 U8288 ( .A(n9156), .ZN(n6839) );
  AND2_X1 U8289 ( .A1(n9190), .A2(n10689), .ZN(n13135) );
  NOR2_X1 U8290 ( .A1(n10695), .A2(n10694), .ZN(n10693) );
  AND2_X1 U8291 ( .A1(n9241), .A2(n9197), .ZN(n13222) );
  INV_X1 U8292 ( .A(n13187), .ZN(n7524) );
  INV_X1 U8293 ( .A(n13216), .ZN(n7016) );
  INV_X1 U8294 ( .A(n13140), .ZN(n13226) );
  AND2_X1 U8295 ( .A1(n13205), .A2(n6627), .ZN(n7021) );
  NAND2_X1 U8296 ( .A1(n7355), .A2(n9239), .ZN(n7352) );
  NAND2_X1 U8297 ( .A1(n13217), .A2(n7354), .ZN(n7353) );
  NAND2_X1 U8298 ( .A1(n7356), .A2(n7355), .ZN(n7354) );
  NAND2_X1 U8299 ( .A1(n9239), .A2(n9165), .ZN(n7356) );
  NAND2_X1 U8300 ( .A1(n8805), .A2(n8804), .ZN(n13477) );
  AND3_X1 U8301 ( .A1(n8589), .A2(n8588), .A3(n8587), .ZN(n12038) );
  INV_X1 U8302 ( .A(n13363), .ZN(n13427) );
  AND2_X1 U8303 ( .A1(n9308), .A2(n9075), .ZN(n15579) );
  NAND2_X1 U8304 ( .A1(n9277), .A2(n9276), .ZN(n10412) );
  AND2_X1 U8305 ( .A1(n13237), .A2(n13486), .ZN(n10410) );
  OAI21_X1 U8306 ( .B1(n12827), .B2(n8905), .A(n8906), .ZN(n13538) );
  NAND2_X1 U8307 ( .A1(n8888), .A2(n8887), .ZN(n13553) );
  NAND2_X1 U8308 ( .A1(n8832), .A2(n8831), .ZN(n13559) );
  NAND2_X1 U8309 ( .A1(n8727), .A2(n8726), .ZN(n12615) );
  OR2_X1 U8310 ( .A1(n11721), .A2(n7585), .ZN(n7581) );
  XNOR2_X1 U8311 ( .A(n7937), .B(n7938), .ZN(n13692) );
  NAND2_X1 U8312 ( .A1(n8464), .A2(n8465), .ZN(n12861) );
  NAND2_X1 U8313 ( .A1(n11044), .A2(n11045), .ZN(n11043) );
  AND2_X1 U8314 ( .A1(n11034), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13700) );
  OR2_X1 U8315 ( .A1(n8070), .A2(n6941), .ZN(n6940) );
  AND2_X1 U8316 ( .A1(n8521), .A2(n8502), .ZN(n13714) );
  INV_X1 U8317 ( .A(n13700), .ZN(n13748) );
  NAND2_X1 U8318 ( .A1(n8507), .A2(n14485), .ZN(n13751) );
  INV_X1 U8319 ( .A(n13714), .ZN(n13753) );
  NAND2_X1 U8320 ( .A1(n8359), .A2(n8358), .ZN(n14087) );
  NAND2_X1 U8321 ( .A1(n14116), .A2(n11007), .ZN(n15532) );
  NAND2_X1 U8322 ( .A1(n14142), .A2(n14143), .ZN(n14141) );
  NAND2_X1 U8323 ( .A1(n14127), .A2(n6774), .ZN(n14142) );
  OR2_X1 U8324 ( .A1(n14124), .A2(n10995), .ZN(n6774) );
  XNOR2_X1 U8325 ( .A(n14144), .B(n10996), .ZN(n14143) );
  NAND2_X1 U8326 ( .A1(n14157), .A2(n14158), .ZN(n14156) );
  NOR2_X1 U8327 ( .A1(n11404), .A2(n7270), .ZN(n14197) );
  NOR2_X1 U8328 ( .A1(n11396), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7270) );
  NAND2_X1 U8329 ( .A1(n14197), .A2(n14196), .ZN(n14195) );
  NAND2_X1 U8330 ( .A1(n11582), .A2(n6612), .ZN(n11585) );
  NAND2_X1 U8331 ( .A1(n7269), .A2(n6781), .ZN(n14207) );
  AND2_X1 U8332 ( .A1(n14208), .A2(n7268), .ZN(n6781) );
  NAND2_X1 U8333 ( .A1(n14246), .A2(n14245), .ZN(n14254) );
  XNOR2_X1 U8334 ( .A(n6772), .B(n14565), .ZN(n14278) );
  NAND2_X1 U8335 ( .A1(n14273), .A2(n14272), .ZN(n6772) );
  AND2_X1 U8336 ( .A1(n10903), .A2(n14074), .ZN(n15546) );
  NOR2_X1 U8337 ( .A1(n15552), .A2(n14283), .ZN(n7280) );
  NAND2_X1 U8338 ( .A1(n10104), .A2(n10012), .ZN(n10026) );
  AND2_X1 U8339 ( .A1(n7687), .A2(n10086), .ZN(n10110) );
  XNOR2_X1 U8340 ( .A(n14319), .B(n7090), .ZN(n7089) );
  INV_X1 U8341 ( .A(n14327), .ZN(n7090) );
  NAND2_X1 U8342 ( .A1(n14502), .A2(n10041), .ZN(n14455) );
  AND2_X1 U8343 ( .A1(n14502), .A2(n14031), .ZN(n14507) );
  NAND2_X1 U8344 ( .A1(n7861), .A2(n7846), .ZN(n7287) );
  NOR2_X1 U8345 ( .A1(n12674), .A2(n12480), .ZN(n7627) );
  AND2_X1 U8346 ( .A1(n14822), .A2(n15190), .ZN(n14812) );
  NAND2_X1 U8347 ( .A1(n14769), .A2(n10583), .ZN(n14724) );
  NAND2_X1 U8348 ( .A1(n14768), .A2(n14770), .ZN(n14769) );
  AND2_X1 U8349 ( .A1(n9798), .A2(n9797), .ZN(n15072) );
  NAND2_X1 U8350 ( .A1(n10448), .A2(n10447), .ZN(n11417) );
  NAND2_X1 U8351 ( .A1(n10446), .A2(n11519), .ZN(n10447) );
  NAND2_X1 U8352 ( .A1(n7622), .A2(n10626), .ZN(n7026) );
  INV_X1 U8353 ( .A(n14809), .ZN(n7025) );
  NAND2_X1 U8354 ( .A1(n10656), .A2(n10655), .ZN(n14826) );
  NAND2_X1 U8355 ( .A1(n9775), .A2(n9774), .ZN(n15069) );
  OR2_X1 U8356 ( .A1(n9528), .A2(n9542), .ZN(n9547) );
  OR2_X1 U8357 ( .A1(n10255), .A2(n11993), .ZN(n9490) );
  NOR2_X1 U8358 ( .A1(n10927), .A2(n10928), .ZN(n10979) );
  AOI21_X1 U8359 ( .B1(n6453), .B2(n7442), .A(n6545), .ZN(n7439) );
  NAND2_X1 U8360 ( .A1(n12433), .A2(n12434), .ZN(n12675) );
  XNOR2_X1 U8361 ( .A(n12790), .B(n12797), .ZN(n12793) );
  XNOR2_X1 U8362 ( .A(n14955), .B(n14952), .ZN(n14948) );
  NAND2_X1 U8363 ( .A1(n14948), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14958) );
  NOR2_X1 U8364 ( .A1(n10391), .A2(n15187), .ZN(n14973) );
  NOR2_X1 U8365 ( .A1(n14998), .A2(n15234), .ZN(n14999) );
  INV_X1 U8366 ( .A(n15008), .ZN(n15017) );
  AOI21_X1 U8367 ( .B1(n15255), .B2(n15015), .A(n15014), .ZN(n15016) );
  INV_X1 U8368 ( .A(n12875), .ZN(n12876) );
  NAND2_X1 U8369 ( .A1(n12874), .A2(n15005), .ZN(n7492) );
  AOI22_X1 U8370 ( .A1(n14833), .A2(n15192), .B1(n15190), .B2(n14835), .ZN(
        n12875) );
  AND2_X1 U8371 ( .A1(n15484), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7490) );
  NAND2_X1 U8372 ( .A1(n12398), .A2(n10318), .ZN(n6679) );
  NAND2_X1 U8373 ( .A1(n11732), .A2(n9607), .ZN(n12070) );
  NAND2_X1 U8374 ( .A1(n15482), .A2(n11909), .ZN(n15196) );
  AND2_X1 U8375 ( .A1(n15482), .A2(n14967), .ZN(n15175) );
  AND2_X1 U8376 ( .A1(n15518), .A2(n15504), .ZN(n12215) );
  INV_X1 U8377 ( .A(n15251), .ZN(n6721) );
  AOI21_X1 U8378 ( .B1(n15253), .B2(n15236), .A(n15250), .ZN(n6722) );
  NAND2_X1 U8379 ( .A1(n14678), .A2(n10318), .ZN(n6692) );
  NAND2_X1 U8380 ( .A1(n10318), .A2(n10802), .ZN(n9505) );
  XNOR2_X1 U8381 ( .A(n10966), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n10889) );
  NOR2_X1 U8382 ( .A1(n6966), .A2(n12457), .ZN(n6962) );
  AOI21_X1 U8383 ( .B1(n12639), .B2(n12638), .A(n6550), .ZN(n15409) );
  NOR2_X1 U8384 ( .A1(n13809), .A2(n6502), .ZN(n7309) );
  AOI21_X1 U8385 ( .B1(n7309), .B2(n7308), .A(n6541), .ZN(n7307) );
  INV_X1 U8386 ( .A(n7385), .ZN(n10142) );
  NOR2_X1 U8387 ( .A1(n7318), .A2(n7314), .ZN(n7313) );
  NOR2_X1 U8388 ( .A1(n7315), .A2(n7312), .ZN(n7311) );
  INV_X1 U8389 ( .A(n10155), .ZN(n7551) );
  OAI21_X1 U8390 ( .B1(n10139), .B2(n11952), .A(n6982), .ZN(n10155) );
  NAND2_X1 U8391 ( .A1(n10139), .A2(n14850), .ZN(n6982) );
  NOR2_X1 U8392 ( .A1(n7303), .A2(n6475), .ZN(n7299) );
  OR2_X1 U8393 ( .A1(n7551), .A2(n10156), .ZN(n7550) );
  AND2_X1 U8394 ( .A1(n7300), .A2(n7298), .ZN(n7297) );
  AND2_X1 U8395 ( .A1(n7609), .A2(n13818), .ZN(n7608) );
  NAND2_X1 U8396 ( .A1(n8275), .A2(n10374), .ZN(n7609) );
  AND2_X1 U8397 ( .A1(n13885), .A2(n7293), .ZN(n7292) );
  INV_X1 U8398 ( .A(n13883), .ZN(n7293) );
  INV_X1 U8399 ( .A(n10167), .ZN(n7032) );
  OAI21_X1 U8400 ( .B1(n13929), .B2(n13928), .A(n13930), .ZN(n13925) );
  NOR2_X1 U8401 ( .A1(n7231), .A2(n7229), .ZN(n7228) );
  NAND2_X1 U8402 ( .A1(n12043), .A2(n9352), .ZN(n7229) );
  INV_X1 U8403 ( .A(n9360), .ZN(n7232) );
  NAND2_X1 U8404 ( .A1(n7227), .A2(n7226), .ZN(n7225) );
  INV_X1 U8405 ( .A(n7230), .ZN(n7227) );
  INV_X1 U8406 ( .A(n7231), .ZN(n7226) );
  AOI21_X1 U8407 ( .B1(n7232), .B2(n6504), .A(n12331), .ZN(n7230) );
  AOI21_X1 U8408 ( .B1(n6446), .B2(n6880), .A(n6878), .ZN(n6877) );
  NAND2_X1 U8409 ( .A1(n13953), .A2(n13958), .ZN(n7601) );
  AOI21_X1 U8410 ( .B1(n14541), .B2(n13956), .A(n6534), .ZN(n13968) );
  NAND2_X1 U8411 ( .A1(n7217), .A2(n13391), .ZN(n7214) );
  NAND2_X1 U8412 ( .A1(n7215), .A2(n13391), .ZN(n7213) );
  INV_X1 U8413 ( .A(n13973), .ZN(n7605) );
  AND2_X1 U8414 ( .A1(n12648), .A2(n12552), .ZN(n10197) );
  INV_X1 U8415 ( .A(n11167), .ZN(n10334) );
  NAND2_X1 U8416 ( .A1(n10230), .A2(n10234), .ZN(n6869) );
  NAND2_X1 U8417 ( .A1(n6872), .A2(n10233), .ZN(n6870) );
  NOR2_X1 U8418 ( .A1(n10234), .A2(n10233), .ZN(n6871) );
  NAND2_X1 U8419 ( .A1(n7236), .A2(n7234), .ZN(n7233) );
  OAI21_X1 U8420 ( .B1(n9402), .B2(n7237), .A(n6546), .ZN(n7236) );
  INV_X1 U8421 ( .A(n9407), .ZN(n7235) );
  NAND2_X1 U8422 ( .A1(n7518), .A2(n9877), .ZN(n7517) );
  NAND3_X1 U8423 ( .A1(n7517), .A2(n10123), .A3(n7519), .ZN(n10259) );
  INV_X1 U8424 ( .A(n8300), .ZN(n7330) );
  INV_X1 U8425 ( .A(n8243), .ZN(n6685) );
  INV_X1 U8426 ( .A(n11145), .ZN(n6811) );
  INV_X1 U8427 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n7529) );
  NOR2_X1 U8428 ( .A1(n6632), .A2(n9227), .ZN(n6832) );
  NAND2_X1 U8429 ( .A1(n6832), .A2(n7066), .ZN(n6828) );
  INV_X1 U8430 ( .A(n12173), .ZN(n9347) );
  INV_X1 U8431 ( .A(n7667), .ZN(n7666) );
  OAI21_X1 U8432 ( .B1(n7669), .B2(n7668), .A(n8942), .ZN(n7667) );
  INV_X1 U8433 ( .A(n8929), .ZN(n7668) );
  INV_X1 U8434 ( .A(n7648), .ZN(n7647) );
  OAI21_X1 U8435 ( .B1(n8814), .B2(n7649), .A(n8841), .ZN(n7648) );
  NOR2_X1 U8436 ( .A1(n8363), .A2(n13622), .ZN(n7141) );
  NAND2_X1 U8437 ( .A1(n7771), .A2(n7770), .ZN(n7768) );
  NOR2_X1 U8438 ( .A1(n9995), .A2(n7774), .ZN(n7770) );
  MUX2_X1 U8439 ( .A(n15237), .B(n14986), .S(n10139), .Z(n10290) );
  INV_X1 U8440 ( .A(n10238), .ZN(n7047) );
  NAND2_X1 U8441 ( .A1(n7556), .A2(n10245), .ZN(n7555) );
  INV_X1 U8442 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n15728) );
  INV_X1 U8443 ( .A(n9850), .ZN(n7324) );
  NAND2_X1 U8444 ( .A1(n6746), .A2(n6444), .ZN(n6745) );
  INV_X1 U8445 ( .A(n8188), .ZN(n8191) );
  INV_X1 U8446 ( .A(n7603), .ZN(n6943) );
  AND2_X1 U8447 ( .A1(n8089), .A2(n8109), .ZN(n7603) );
  INV_X1 U8448 ( .A(n8108), .ZN(n8109) );
  NAND2_X1 U8449 ( .A1(n8111), .A2(n10825), .ZN(n8153) );
  OAI21_X1 U8450 ( .B1(n7007), .B2(n10858), .A(n7002), .ZN(n7343) );
  NAND2_X1 U8451 ( .A1(n7007), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7002) );
  OAI21_X1 U8452 ( .B1(n7944), .B2(n7822), .A(n7821), .ZN(n7823) );
  NAND2_X1 U8453 ( .A1(n7944), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7821) );
  INV_X1 U8454 ( .A(n7817), .ZN(n7598) );
  AOI21_X1 U8455 ( .B1(n11773), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11772), .ZN(
        n11774) );
  AND2_X1 U8456 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  NOR2_X1 U8457 ( .A1(n12584), .A2(n13095), .ZN(n7180) );
  NOR2_X1 U8458 ( .A1(n12562), .A2(n7506), .ZN(n7505) );
  INV_X1 U8459 ( .A(n12171), .ZN(n7506) );
  AOI21_X1 U8460 ( .B1(n9414), .B2(n9413), .A(n13277), .ZN(n9419) );
  INV_X1 U8461 ( .A(n9445), .ZN(n9446) );
  OAI21_X1 U8462 ( .B1(n13508), .B2(n12468), .A(n9444), .ZN(n9445) );
  NAND2_X1 U8463 ( .A1(n6819), .A2(n6818), .ZN(n6823) );
  AND3_X1 U8464 ( .A1(n6900), .A2(n6594), .A3(n6901), .ZN(n9182) );
  NAND2_X1 U8465 ( .A1(n6817), .A2(n6816), .ZN(n9145) );
  NAND2_X1 U8466 ( .A1(n7063), .A2(n6821), .ZN(n6816) );
  NAND2_X1 U8467 ( .A1(n6819), .A2(n6523), .ZN(n6817) );
  NOR2_X1 U8468 ( .A1(n13160), .A2(n7545), .ZN(n7543) );
  OAI22_X1 U8469 ( .A1(n7543), .A2(n12786), .B1(n7544), .B2(n9227), .ZN(n7538)
         );
  NOR2_X1 U8470 ( .A1(n13167), .A2(n13155), .ZN(n7252) );
  INV_X1 U8471 ( .A(n6989), .ZN(n8991) );
  INV_X1 U8472 ( .A(n9344), .ZN(n7152) );
  INV_X1 U8473 ( .A(n7151), .ZN(n7150) );
  OAI21_X1 U8474 ( .B1(n8640), .B2(n7152), .A(n9347), .ZN(n7151) );
  AND2_X1 U8475 ( .A1(n7712), .A2(n9389), .ZN(n7710) );
  INV_X1 U8476 ( .A(n8839), .ZN(n7712) );
  AND2_X1 U8477 ( .A1(n7711), .A2(n8917), .ZN(n7708) );
  OR2_X1 U8478 ( .A1(n13538), .A2(n13031), .ZN(n9406) );
  NAND2_X1 U8479 ( .A1(n7187), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U8480 ( .A1(n7696), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7694) );
  INV_X1 U8481 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7696) );
  NOR2_X1 U8482 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n9083) );
  INV_X1 U8483 ( .A(n8811), .ZN(n6796) );
  AOI21_X1 U8484 ( .B1(n7647), .B2(n7649), .A(n7646), .ZN(n7645) );
  INV_X1 U8485 ( .A(n8843), .ZN(n7646) );
  AND2_X1 U8486 ( .A1(n6795), .A2(n7647), .ZN(n6794) );
  OR2_X1 U8487 ( .A1(n7650), .A2(n6796), .ZN(n6795) );
  INV_X1 U8488 ( .A(n7643), .ZN(n7642) );
  OAI21_X1 U8489 ( .B1(n8703), .B2(n7644), .A(n8735), .ZN(n7643) );
  INV_X1 U8490 ( .A(n8720), .ZN(n7644) );
  AND2_X1 U8491 ( .A1(n7642), .A2(n6788), .ZN(n6787) );
  NAND2_X1 U8492 ( .A1(n6789), .A2(n8700), .ZN(n6788) );
  INV_X1 U8493 ( .A(n8685), .ZN(n6789) );
  NAND2_X1 U8494 ( .A1(n6787), .A2(n6790), .ZN(n6785) );
  INV_X1 U8495 ( .A(n8700), .ZN(n6790) );
  INV_X1 U8496 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8613) );
  XNOR2_X1 U8497 ( .A(n14433), .B(n8412), .ZN(n8285) );
  INV_X1 U8498 ( .A(n7577), .ZN(n7576) );
  AOI21_X1 U8499 ( .B1(n7577), .B2(n7575), .A(n6560), .ZN(n7574) );
  INV_X1 U8500 ( .A(n13643), .ZN(n7575) );
  AND2_X1 U8501 ( .A1(n8461), .A2(n8460), .ZN(n12851) );
  NOR2_X1 U8502 ( .A1(n8230), .A2(n8229), .ZN(n6977) );
  NOR2_X1 U8503 ( .A1(n8277), .A2(n8276), .ZN(n7142) );
  NOR2_X1 U8504 ( .A1(n8330), .A2(n13637), .ZN(n6976) );
  NOR2_X1 U8505 ( .A1(n8141), .A2(n8140), .ZN(n7140) );
  OR3_X1 U8506 ( .A1(n8498), .A2(n15557), .A3(n10114), .ZN(n8524) );
  NAND2_X1 U8507 ( .A1(n7591), .A2(n8175), .ZN(n7588) );
  INV_X1 U8508 ( .A(n8132), .ZN(n6675) );
  NAND2_X1 U8509 ( .A1(n6744), .A2(n6742), .ZN(n6741) );
  NAND2_X1 U8510 ( .A1(n6740), .A2(n6739), .ZN(n6738) );
  NOR2_X1 U8511 ( .A1(n7910), .A2(n14504), .ZN(n7088) );
  OR2_X1 U8512 ( .A1(n7910), .A2(n10908), .ZN(n7911) );
  NOR2_X1 U8513 ( .A1(n7275), .A2(n7274), .ZN(n7273) );
  NOR2_X1 U8514 ( .A1(n12771), .A2(n12772), .ZN(n7274) );
  XNOR2_X1 U8515 ( .A(n14516), .B(n14081), .ZN(n10098) );
  INV_X1 U8516 ( .A(n7737), .ZN(n7736) );
  OR2_X1 U8517 ( .A1(n14629), .A2(n14536), .ZN(n7737) );
  OAI21_X1 U8518 ( .B1(n6479), .B2(n10068), .A(n10071), .ZN(n7674) );
  NOR2_X1 U8519 ( .A1(n6479), .A2(n6761), .ZN(n6760) );
  INV_X1 U8520 ( .A(n10067), .ZN(n6761) );
  INV_X1 U8521 ( .A(n10066), .ZN(n7678) );
  NOR2_X1 U8522 ( .A1(n14655), .A2(n13887), .ZN(n7730) );
  NOR2_X1 U8523 ( .A1(n13880), .A2(n14594), .ZN(n6666) );
  AND2_X1 U8524 ( .A1(n6889), .A2(n9981), .ZN(n6888) );
  OR2_X1 U8525 ( .A1(n6892), .A2(n14049), .ZN(n6889) );
  INV_X1 U8526 ( .A(n9979), .ZN(n6892) );
  INV_X1 U8527 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8038) );
  INV_X1 U8528 ( .A(n14042), .ZN(n11120) );
  INV_X1 U8529 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6657) );
  INV_X1 U8530 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6656) );
  INV_X1 U8531 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8115) );
  OR2_X1 U8532 ( .A1(n8091), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8112) );
  XNOR2_X1 U8533 ( .A(n10456), .B(n10427), .ZN(n10458) );
  NAND2_X1 U8534 ( .A1(n10455), .A2(n10454), .ZN(n10456) );
  INV_X1 U8535 ( .A(n6438), .ZN(n10628) );
  NAND2_X1 U8536 ( .A1(n10320), .A2(n10270), .ZN(n7335) );
  NOR2_X1 U8537 ( .A1(n14832), .A2(n7333), .ZN(n7332) );
  NOR2_X1 U8538 ( .A1(n15244), .A2(n7459), .ZN(n7460) );
  OR2_X1 U8539 ( .A1(n15246), .A2(n15258), .ZN(n7459) );
  INV_X1 U8540 ( .A(n12866), .ZN(n12872) );
  NAND2_X1 U8541 ( .A1(n9813), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9828) );
  INV_X1 U8542 ( .A(n9826), .ZN(n9813) );
  NAND2_X1 U8543 ( .A1(n15056), .A2(n6848), .ZN(n7423) );
  NOR2_X1 U8544 ( .A1(n6849), .A2(n15042), .ZN(n6848) );
  INV_X1 U8545 ( .A(n9799), .ZN(n6849) );
  INV_X1 U8546 ( .A(n9897), .ZN(n7482) );
  NOR2_X1 U8547 ( .A1(n15206), .A2(n15188), .ZN(n9925) );
  NOR2_X1 U8548 ( .A1(n9699), .A2(n12442), .ZN(n7143) );
  NOR2_X1 U8549 ( .A1(n12552), .A2(n12322), .ZN(n7458) );
  NOR2_X1 U8550 ( .A1(n9614), .A2(n9613), .ZN(n7144) );
  NOR2_X1 U8551 ( .A1(n9640), .A2(n15650), .ZN(n7059) );
  AND2_X1 U8552 ( .A1(n12080), .A2(n12357), .ZN(n12163) );
  INV_X1 U8553 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9599) );
  NAND2_X1 U8554 ( .A1(n7467), .A2(n9884), .ZN(n7466) );
  INV_X1 U8555 ( .A(n9883), .ZN(n7467) );
  NOR2_X1 U8556 ( .A1(n9556), .A2(n9555), .ZN(n9570) );
  NAND2_X1 U8557 ( .A1(n11279), .A2(n9883), .ZN(n11940) );
  NAND2_X1 U8558 ( .A1(n7106), .A2(n11364), .ZN(n10147) );
  AND2_X1 U8559 ( .A1(n7077), .A2(n6716), .ZN(n12877) );
  NOR2_X1 U8560 ( .A1(n15264), .A2(n6717), .ZN(n6716) );
  NAND2_X1 U8561 ( .A1(n9476), .A2(n9477), .ZN(n9937) );
  OAI21_X1 U8562 ( .B1(n9938), .B2(n9937), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9939) );
  AOI21_X1 U8563 ( .B1(n7328), .B2(n7329), .A(n7326), .ZN(n7325) );
  INV_X1 U8564 ( .A(n8389), .ZN(n7326) );
  NAND2_X1 U8565 ( .A1(n6699), .A2(n6698), .ZN(n6697) );
  NAND2_X1 U8566 ( .A1(n10801), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6698) );
  OR2_X1 U8567 ( .A1(n10801), .A2(n6700), .ZN(n6699) );
  NAND2_X1 U8568 ( .A1(n6697), .A2(SI_21_), .ZN(n8378) );
  NOR2_X1 U8569 ( .A1(n8325), .A2(n8324), .ZN(n8381) );
  NOR2_X1 U8570 ( .A1(n8323), .A2(SI_20_), .ZN(n8324) );
  INV_X1 U8571 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U8572 ( .A1(n7057), .A2(n7056), .ZN(n9938) );
  INV_X1 U8573 ( .A(n9731), .ZN(n7057) );
  NAND2_X1 U8574 ( .A1(n7470), .A2(n9478), .ZN(n9731) );
  NAND2_X1 U8575 ( .A1(n8272), .A2(n8247), .ZN(n8248) );
  XNOR2_X1 U8576 ( .A(n8245), .B(SI_17_), .ZN(n8243) );
  INV_X1 U8577 ( .A(n7341), .ZN(n7599) );
  NAND2_X1 U8578 ( .A1(n6748), .A2(n8221), .ZN(n7600) );
  NAND2_X1 U8579 ( .A1(n6482), .A2(n8195), .ZN(n6748) );
  INV_X1 U8580 ( .A(n8187), .ZN(n8196) );
  OR2_X1 U8581 ( .A1(n9594), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9678) );
  XNOR2_X1 U8582 ( .A(n8187), .B(SI_14_), .ZN(n8176) );
  XNOR2_X1 U8583 ( .A(n8158), .B(SI_13_), .ZN(n8156) );
  OR2_X1 U8584 ( .A1(n9649), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U8585 ( .A1(n6712), .A2(n8153), .ZN(n8134) );
  NAND2_X1 U8586 ( .A1(n8090), .A2(n7603), .ZN(n6712) );
  OR2_X1 U8587 ( .A1(n9636), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U8588 ( .A1(n8074), .A2(SI_10_), .ZN(n8089) );
  NAND2_X1 U8589 ( .A1(n8088), .A2(n8087), .ZN(n8090) );
  OAI21_X1 U8590 ( .B1(n8074), .B2(SI_10_), .A(n8089), .ZN(n8086) );
  NAND2_X1 U8591 ( .A1(n8073), .A2(n8072), .ZN(n8088) );
  OAI21_X1 U8592 ( .B1(n10801), .B2(n10875), .A(n7049), .ZN(n8056) );
  NAND2_X1 U8593 ( .A1(n10801), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U8594 ( .A1(n8055), .A2(n6997), .ZN(n8052) );
  INV_X1 U8595 ( .A(n8030), .ZN(n6999) );
  INV_X1 U8596 ( .A(n6713), .ZN(n7816) );
  NAND2_X1 U8597 ( .A1(n7944), .A2(n8555), .ZN(n7085) );
  AND2_X1 U8598 ( .A1(n10850), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10745) );
  XNOR2_X1 U8599 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n10746) );
  OR2_X1 U8600 ( .A1(n10765), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U8601 ( .A1(n11099), .A2(n11098), .ZN(n11105) );
  OR2_X1 U8602 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n11097), .ZN(n11098) );
  AND2_X1 U8603 ( .A1(n11767), .A2(n11766), .ZN(n11770) );
  OR2_X1 U8604 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n11774), .ZN(n12091) );
  NAND2_X1 U8605 ( .A1(n12455), .A2(n12454), .ZN(n12460) );
  INV_X1 U8606 ( .A(n15408), .ZN(n7248) );
  OR2_X1 U8607 ( .A1(n15412), .A2(n15411), .ZN(n15415) );
  XNOR2_X1 U8608 ( .A(n12173), .B(n7186), .ZN(n12303) );
  XNOR2_X1 U8609 ( .A(n12934), .B(n7186), .ZN(n12969) );
  XNOR2_X1 U8610 ( .A(n12972), .B(n12309), .ZN(n12359) );
  AOI21_X1 U8611 ( .B1(n7494), .B2(n7496), .A(n6542), .ZN(n7493) );
  AND2_X1 U8612 ( .A1(n7175), .A2(n12984), .ZN(n7174) );
  NAND2_X1 U8613 ( .A1(n7493), .A2(n7176), .ZN(n7175) );
  INV_X1 U8614 ( .A(n7494), .ZN(n7176) );
  INV_X1 U8615 ( .A(n7493), .ZN(n7177) );
  NAND2_X1 U8616 ( .A1(n9292), .A2(n13108), .ZN(n9316) );
  INV_X1 U8617 ( .A(n13108), .ZN(n7692) );
  NAND2_X1 U8618 ( .A1(n12951), .A2(n12567), .ZN(n12586) );
  XNOR2_X1 U8619 ( .A(n13520), .B(n7186), .ZN(n12926) );
  XNOR2_X1 U8620 ( .A(n13270), .B(n7186), .ZN(n12929) );
  AND2_X1 U8621 ( .A1(n11305), .A2(n11304), .ZN(n11544) );
  AND2_X1 U8622 ( .A1(n9454), .A2(n7013), .ZN(n7012) );
  AND2_X1 U8623 ( .A1(n9010), .A2(n6432), .ZN(n7013) );
  AND2_X1 U8624 ( .A1(n8998), .A2(n8997), .ZN(n12976) );
  AND2_X1 U8625 ( .A1(n8896), .A2(n8895), .ZN(n13009) );
  AND3_X1 U8626 ( .A1(n8823), .A2(n8822), .A3(n8821), .ZN(n13008) );
  AND4_X1 U8627 ( .A1(n8751), .A2(n8750), .A3(n8749), .A4(n8748), .ZN(n12589)
         );
  OR2_X1 U8628 ( .A1(n9068), .A2(n15759), .ZN(n8715) );
  AND4_X1 U8629 ( .A1(n8611), .A2(n8610), .A3(n8609), .A4(n8608), .ZN(n11863)
         );
  NAND2_X1 U8630 ( .A1(n9268), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7165) );
  NOR2_X1 U8631 ( .A1(n11214), .A2(n9175), .ZN(n11188) );
  NAND2_X1 U8632 ( .A1(n13601), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U8633 ( .A1(n6994), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7265) );
  INV_X1 U8634 ( .A(n13601), .ZN(n6994) );
  NOR2_X1 U8635 ( .A1(n9180), .A2(n9181), .ZN(n11136) );
  AND2_X1 U8636 ( .A1(n9179), .A2(n11145), .ZN(n9180) );
  NAND2_X1 U8637 ( .A1(n11136), .A2(n6899), .ZN(n6900) );
  AND2_X1 U8638 ( .A1(n6902), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U8639 ( .A1(n11136), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n11232) );
  INV_X1 U8640 ( .A(n6823), .ZN(n11227) );
  NAND2_X1 U8641 ( .A1(n7364), .A2(n7363), .ZN(n7362) );
  OAI21_X1 U8642 ( .B1(n11446), .B2(n11447), .A(n6544), .ZN(n11884) );
  AOI21_X1 U8643 ( .B1(n11883), .B2(n11887), .A(n10708), .ZN(n10707) );
  INV_X1 U8644 ( .A(n10711), .ZN(n6837) );
  NAND2_X1 U8645 ( .A1(n7346), .A2(n11889), .ZN(n6834) );
  NAND3_X1 U8646 ( .A1(n7350), .A2(P3_REG1_REG_11__SCAN_IN), .A3(n7349), .ZN(
        n12393) );
  NAND2_X1 U8647 ( .A1(n6898), .A2(n13116), .ZN(n13118) );
  NAND2_X1 U8648 ( .A1(n7515), .A2(n13115), .ZN(n6898) );
  NAND2_X1 U8649 ( .A1(n10692), .A2(n7543), .ZN(n7542) );
  NAND2_X1 U8650 ( .A1(n10692), .A2(n7544), .ZN(n7536) );
  OR2_X1 U8651 ( .A1(n7541), .A2(n7540), .ZN(n13153) );
  NAND2_X1 U8652 ( .A1(n7542), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7541) );
  INV_X1 U8653 ( .A(n13174), .ZN(n7540) );
  OAI21_X1 U8654 ( .B1(n7064), .B2(n6831), .A(n6824), .ZN(n6826) );
  INV_X1 U8655 ( .A(n6833), .ZN(n6831) );
  INV_X1 U8656 ( .A(n6825), .ZN(n6824) );
  NAND2_X1 U8657 ( .A1(n9159), .A2(n13160), .ZN(n13169) );
  NAND2_X1 U8658 ( .A1(n7361), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13170) );
  INV_X1 U8659 ( .A(n13152), .ZN(n7361) );
  NAND2_X1 U8660 ( .A1(n7521), .A2(n6904), .ZN(n6903) );
  AND2_X1 U8661 ( .A1(n7526), .A2(n9238), .ZN(n6904) );
  NAND2_X1 U8662 ( .A1(n7520), .A2(n6472), .ZN(n6906) );
  AND2_X1 U8663 ( .A1(n13222), .A2(n6909), .ZN(n6908) );
  NOR2_X1 U8664 ( .A1(n9232), .A2(n6993), .ZN(n6992) );
  INV_X1 U8665 ( .A(n9233), .ZN(n6993) );
  AOI21_X1 U8666 ( .B1(n13252), .B2(n9258), .A(n9070), .ZN(n10403) );
  NAND2_X1 U8667 ( .A1(n9443), .A2(n9444), .ZN(n10408) );
  NOR2_X1 U8668 ( .A1(n13229), .A2(n12348), .ZN(n10405) );
  NAND2_X1 U8669 ( .A1(n6989), .A2(n15720), .ZN(n9064) );
  OR2_X1 U8670 ( .A1(n9064), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n13231) );
  INV_X1 U8671 ( .A(n7161), .ZN(n7160) );
  OAI21_X1 U8672 ( .B1(n9310), .B2(n7162), .A(n9416), .ZN(n7161) );
  NAND2_X1 U8673 ( .A1(n8964), .A2(n8963), .ZN(n8978) );
  INV_X1 U8674 ( .A(n8965), .ZN(n8964) );
  NAND2_X1 U8675 ( .A1(n8950), .A2(n8934), .ZN(n13308) );
  NAND2_X1 U8676 ( .A1(n6987), .A2(n8907), .ZN(n8922) );
  NAND2_X1 U8677 ( .A1(n7128), .A2(n8854), .ZN(n8873) );
  INV_X1 U8678 ( .A(n7128), .ZN(n8891) );
  NAND2_X1 U8679 ( .A1(n8833), .A2(n15748), .ZN(n8889) );
  NAND2_X1 U8680 ( .A1(n7127), .A2(n8806), .ZN(n8819) );
  INV_X1 U8681 ( .A(n7127), .ZN(n8807) );
  NAND2_X1 U8682 ( .A1(n7126), .A2(n8745), .ZN(n8768) );
  INV_X1 U8683 ( .A(n7126), .ZN(n8746) );
  NAND2_X1 U8684 ( .A1(n6984), .A2(n8693), .ZN(n8713) );
  INV_X1 U8685 ( .A(n8694), .ZN(n6984) );
  NAND2_X1 U8686 ( .A1(n7123), .A2(n8641), .ZN(n8675) );
  INV_X1 U8687 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8641) );
  INV_X1 U8688 ( .A(n8642), .ZN(n7123) );
  AND2_X1 U8689 ( .A1(n7197), .A2(n9027), .ZN(n7196) );
  NAND2_X1 U8690 ( .A1(n12055), .A2(n8640), .ZN(n7149) );
  NAND2_X1 U8691 ( .A1(n7125), .A2(n7124), .ZN(n8642) );
  INV_X1 U8692 ( .A(n8624), .ZN(n7125) );
  NAND2_X1 U8693 ( .A1(n8604), .A2(n8603), .ZN(n8624) );
  INV_X1 U8694 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8603) );
  INV_X1 U8695 ( .A(n8605), .ZN(n8604) );
  NAND2_X1 U8696 ( .A1(n7164), .A2(n9335), .ZN(n12132) );
  NAND2_X1 U8697 ( .A1(n12037), .A2(n11557), .ZN(n8605) );
  NAND2_X1 U8698 ( .A1(n12034), .A2(n9025), .ZN(n12019) );
  NAND2_X1 U8699 ( .A1(n12019), .A2(n12018), .ZN(n12017) );
  NAND2_X1 U8700 ( .A1(n9020), .A2(n11345), .ZN(n12027) );
  INV_X1 U8701 ( .A(n11331), .ZN(n13500) );
  NAND2_X1 U8702 ( .A1(n11309), .A2(n9322), .ZN(n13496) );
  AND2_X1 U8703 ( .A1(n8860), .A2(n8859), .ZN(n13335) );
  INV_X1 U8704 ( .A(n9291), .ZN(n13338) );
  INV_X1 U8705 ( .A(n7741), .ZN(n13330) );
  AOI21_X1 U8706 ( .B1(n13378), .B2(n9042), .A(n9043), .ZN(n7741) );
  OR2_X1 U8707 ( .A1(n13375), .A2(n13382), .ZN(n13376) );
  NAND2_X1 U8708 ( .A1(n7700), .A2(n7698), .ZN(n13406) );
  AOI21_X1 U8709 ( .B1(n7702), .B2(n7704), .A(n7699), .ZN(n7698) );
  INV_X1 U8710 ( .A(n9385), .ZN(n7699) );
  OR2_X1 U8711 ( .A1(n15627), .A2(n15607), .ZN(n13486) );
  OAI21_X1 U8712 ( .B1(n9286), .B2(n7804), .A(n9252), .ZN(n9275) );
  NAND2_X1 U8713 ( .A1(n8553), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8552) );
  OAI21_X1 U8714 ( .B1(n8974), .B2(n7659), .A(n7657), .ZN(n9247) );
  AOI21_X1 U8715 ( .B1(n7660), .B2(n7658), .A(n6629), .ZN(n7657) );
  INV_X1 U8716 ( .A(n7660), .ZN(n7659) );
  NAND2_X1 U8717 ( .A1(n7188), .A2(n8542), .ZN(n6652) );
  NAND2_X1 U8718 ( .A1(n6809), .A2(n6808), .ZN(n8974) );
  NAND2_X1 U8719 ( .A1(n8946), .A2(n15734), .ZN(n6808) );
  NOR2_X1 U8720 ( .A1(n8930), .A2(n7670), .ZN(n7669) );
  INV_X1 U8721 ( .A(n8918), .ZN(n7670) );
  NAND2_X1 U8722 ( .A1(n8866), .A2(n6460), .ZN(n8868) );
  INV_X1 U8723 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7178) );
  NAND2_X1 U8724 ( .A1(n6793), .A2(n6791), .ZN(n8880) );
  AOI21_X1 U8725 ( .B1(n6794), .B2(n6796), .A(n6792), .ZN(n6791) );
  NAND2_X1 U8726 ( .A1(n7652), .A2(n6794), .ZN(n6793) );
  INV_X1 U8727 ( .A(n7645), .ZN(n6792) );
  NAND2_X1 U8728 ( .A1(n8756), .A2(n8755), .ZN(n8798) );
  INV_X1 U8729 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8739) );
  OR2_X1 U8730 ( .A1(n8671), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8688) );
  NAND2_X1 U8731 ( .A1(n8686), .A2(n8685), .ZN(n8701) );
  OAI21_X1 U8732 ( .B1(n8654), .B2(n7656), .A(n6802), .ZN(n8669) );
  AOI21_X1 U8733 ( .B1(n7655), .B2(n6804), .A(n6803), .ZN(n6802) );
  INV_X1 U8734 ( .A(n8653), .ZN(n6804) );
  INV_X1 U8735 ( .A(n8665), .ZN(n6803) );
  AND2_X1 U8736 ( .A1(n8682), .A2(n8667), .ZN(n8668) );
  NAND2_X1 U8737 ( .A1(n8669), .A2(n8668), .ZN(n8683) );
  AND2_X1 U8738 ( .A1(n8634), .A2(n8620), .ZN(n8632) );
  NAND2_X1 U8739 ( .A1(n6800), .A2(n6797), .ZN(n8617) );
  AOI21_X1 U8740 ( .B1(n8598), .B2(n6799), .A(n6798), .ZN(n6797) );
  INV_X1 U8741 ( .A(n8600), .ZN(n6798) );
  AND2_X1 U8742 ( .A1(n8618), .A2(n8601), .ZN(n8616) );
  OR2_X1 U8743 ( .A1(n8759), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8612) );
  XNOR2_X1 U8744 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8565) );
  NAND2_X1 U8745 ( .A1(n8555), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U8746 ( .A1(n7592), .A2(n7591), .ZN(n7590) );
  XNOR2_X1 U8747 ( .A(n7732), .B(n7987), .ZN(n7937) );
  NAND2_X1 U8748 ( .A1(n6977), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8277) );
  INV_X1 U8749 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11587) );
  OR2_X1 U8750 ( .A1(n8121), .A2(n11587), .ZN(n8141) );
  INV_X1 U8751 ( .A(n6977), .ZN(n8258) );
  INV_X1 U8752 ( .A(n14087), .ZN(n14064) );
  XNOR2_X1 U8753 ( .A(n14610), .B(n8412), .ZN(n6941) );
  NAND2_X1 U8754 ( .A1(n6941), .A2(n8070), .ZN(n8071) );
  NAND2_X1 U8755 ( .A1(n7142), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8330) );
  INV_X1 U8756 ( .A(n7142), .ZN(n8307) );
  INV_X1 U8757 ( .A(n6976), .ZN(n8361) );
  INV_X1 U8758 ( .A(n8341), .ZN(n6672) );
  NAND2_X1 U8759 ( .A1(n6975), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8097) );
  INV_X1 U8760 ( .A(n8078), .ZN(n6975) );
  NAND2_X1 U8761 ( .A1(n6974), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8121) );
  INV_X1 U8762 ( .A(n8097), .ZN(n6974) );
  INV_X1 U8763 ( .A(n13725), .ZN(n13734) );
  NAND2_X1 U8764 ( .A1(n8203), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8230) );
  INV_X1 U8765 ( .A(n8209), .ZN(n8203) );
  NAND2_X1 U8766 ( .A1(n7140), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8209) );
  AND2_X1 U8767 ( .A1(n8459), .A2(n8458), .ZN(n13735) );
  AND2_X1 U8768 ( .A1(n8369), .A2(n8368), .ZN(n13960) );
  AND4_X1 U8769 ( .A1(n7995), .A2(n7994), .A3(n7993), .A4(n7992), .ZN(n13815)
         );
  AND4_X1 U8770 ( .A1(n7962), .A2(n7961), .A3(n7960), .A4(n7959), .ZN(n13808)
         );
  NAND2_X1 U8771 ( .A1(n14169), .A2(n7267), .ZN(n15538) );
  NAND2_X1 U8772 ( .A1(n11016), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7267) );
  NAND2_X1 U8773 ( .A1(n15538), .A2(n15539), .ZN(n15536) );
  NAND2_X1 U8774 ( .A1(n12261), .A2(n12262), .ZN(n7268) );
  XNOR2_X1 U8775 ( .A(n7273), .B(n7272), .ZN(n12773) );
  NOR2_X1 U8776 ( .A1(n12773), .A2(n14590), .ZN(n14221) );
  NAND2_X1 U8777 ( .A1(n12763), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n12767) );
  NOR2_X1 U8778 ( .A1(n14221), .A2(n7271), .ZN(n14223) );
  NOR2_X1 U8779 ( .A1(n7273), .A2(n7272), .ZN(n7271) );
  NAND2_X1 U8780 ( .A1(n7277), .A2(n7276), .ZN(n6778) );
  NAND2_X1 U8781 ( .A1(n14261), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7276) );
  AND2_X1 U8782 ( .A1(n6778), .A2(n14255), .ZN(n14271) );
  INV_X1 U8783 ( .A(n14634), .ZN(n14383) );
  NAND2_X1 U8784 ( .A1(n14397), .A2(n14383), .ZN(n14382) );
  AND2_X1 U8785 ( .A1(n14433), .A2(n13708), .ZN(n14404) );
  NAND2_X1 U8786 ( .A1(n6766), .A2(n7673), .ZN(n14425) );
  OR2_X1 U8787 ( .A1(n14420), .A2(n14445), .ZN(n14446) );
  NAND2_X1 U8788 ( .A1(n12500), .A2(n7730), .ZN(n14488) );
  NAND2_X1 U8789 ( .A1(n12500), .A2(n10039), .ZN(n14487) );
  NAND2_X1 U8790 ( .A1(n7775), .A2(n7774), .ZN(n7773) );
  NAND2_X1 U8791 ( .A1(n12411), .A2(n12412), .ZN(n12499) );
  NAND2_X1 U8792 ( .A1(n12293), .A2(n12407), .ZN(n6755) );
  OR2_X1 U8793 ( .A1(n8039), .A2(n8038), .ZN(n8064) );
  NAND2_X1 U8794 ( .A1(n8062), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8078) );
  INV_X1 U8795 ( .A(n8064), .ZN(n8062) );
  NOR2_X2 U8796 ( .A1(n11788), .A2(n14610), .ZN(n12006) );
  INV_X1 U8797 ( .A(n10055), .ZN(n6754) );
  AND2_X1 U8798 ( .A1(n14050), .A2(n6751), .ZN(n6750) );
  AOI21_X1 U8799 ( .B1(n10055), .B2(n6753), .A(n6752), .ZN(n6751) );
  NAND2_X1 U8800 ( .A1(n11535), .A2(n10055), .ZN(n11750) );
  NAND2_X1 U8801 ( .A1(n8015), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8039) );
  INV_X1 U8802 ( .A(n8017), .ZN(n8015) );
  NAND2_X1 U8803 ( .A1(n7988), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8017) );
  INV_X1 U8804 ( .A(n7990), .ZN(n7988) );
  NAND2_X1 U8805 ( .A1(n11574), .A2(n10054), .ZN(n11535) );
  NAND2_X1 U8806 ( .A1(n11578), .A2(n11663), .ZN(n11579) );
  XNOR2_X1 U8807 ( .A(n13813), .B(n13815), .ZN(n14048) );
  AND3_X1 U8808 ( .A1(n7732), .A2(n10035), .A3(n9970), .ZN(n11641) );
  NAND2_X1 U8809 ( .A1(n7955), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7990) );
  INV_X1 U8810 ( .A(n7957), .ZN(n7955) );
  NAND2_X1 U8811 ( .A1(n10035), .A2(n7732), .ZN(n11437) );
  INV_X1 U8812 ( .A(n11376), .ZN(n10035) );
  NAND2_X1 U8813 ( .A1(n11123), .A2(n10047), .ZN(n11083) );
  NOR2_X1 U8814 ( .A1(n13755), .A2(n7559), .ZN(n11124) );
  AND2_X1 U8815 ( .A1(n14516), .A2(n15564), .ZN(n7094) );
  NAND2_X1 U8816 ( .A1(n7558), .A2(n13755), .ZN(n10973) );
  AND2_X1 U8817 ( .A1(n10682), .A2(n12399), .ZN(n8526) );
  OR2_X1 U8818 ( .A1(n7861), .A2(n7864), .ZN(n8499) );
  INV_X1 U8819 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7862) );
  OR2_X1 U8820 ( .A1(n8183), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8198) );
  OR2_X1 U8821 ( .A1(n8112), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U8822 ( .A1(n8032), .A2(n8034), .ZN(n8251) );
  CLKBUF_X1 U8823 ( .A(n7980), .Z(n7981) );
  NOR2_X1 U8824 ( .A1(n14691), .A2(n7629), .ZN(n7628) );
  INV_X1 U8825 ( .A(n10527), .ZN(n7629) );
  NAND2_X1 U8826 ( .A1(n9767), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9780) );
  INV_X1 U8827 ( .A(n9768), .ZN(n9767) );
  OR2_X1 U8828 ( .A1(n9600), .A2(n9599), .ZN(n9614) );
  INV_X1 U8829 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9613) );
  INV_X1 U8830 ( .A(n7144), .ZN(n9630) );
  NAND2_X1 U8831 ( .A1(n10494), .A2(n10495), .ZN(n7636) );
  NAND2_X1 U8832 ( .A1(n9779), .A2(n15404), .ZN(n7404) );
  AOI21_X1 U8833 ( .B1(n6430), .B2(n10460), .A(n6733), .ZN(n11054) );
  OAI22_X1 U8834 ( .A1(n10628), .A2(n7403), .B1(n11244), .B2(n10421), .ZN(
        n6733) );
  INV_X1 U8835 ( .A(n9757), .ZN(n9758) );
  NAND2_X1 U8836 ( .A1(n11054), .A2(n11053), .ZN(n11052) );
  NAND2_X1 U8837 ( .A1(n10458), .A2(n10457), .ZN(n10464) );
  INV_X1 U8838 ( .A(n11602), .ZN(n10444) );
  NAND2_X1 U8839 ( .A1(n10303), .A2(n10280), .ZN(n10287) );
  AND2_X1 U8840 ( .A1(n10310), .A2(n10312), .ZN(n6696) );
  NAND2_X1 U8841 ( .A1(n10284), .A2(n10283), .ZN(n6980) );
  NAND2_X1 U8842 ( .A1(n6866), .A2(n6864), .ZN(n10284) );
  NOR2_X1 U8843 ( .A1(n6865), .A2(n6547), .ZN(n6864) );
  INV_X1 U8844 ( .A(n10357), .ZN(n7008) );
  AND2_X1 U8845 ( .A1(n9821), .A2(n9820), .ZN(n15012) );
  NAND4_X1 U8846 ( .A1(n9561), .A2(n9560), .A3(n9559), .A4(n9558), .ZN(n9579)
         );
  OR2_X1 U8847 ( .A1(n9519), .A2(n15727), .ZN(n9491) );
  NOR2_X1 U8848 ( .A1(n11253), .A2(n6487), .ZN(n10949) );
  AOI21_X1 U8849 ( .B1(n11252), .B2(n10951), .A(n10950), .ZN(n14859) );
  OR2_X1 U8850 ( .A1(n10982), .A2(n10981), .ZN(n7438) );
  NAND2_X1 U8851 ( .A1(n6636), .A2(n10933), .ZN(n10986) );
  OR2_X1 U8852 ( .A1(n14880), .A2(n10934), .ZN(n6636) );
  AND2_X1 U8853 ( .A1(n7438), .A2(n7437), .ZN(n14891) );
  NAND2_X1 U8854 ( .A1(n11262), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U8855 ( .A1(n14891), .A2(n14890), .ZN(n14889) );
  NAND2_X1 U8856 ( .A1(n14907), .A2(n7443), .ZN(n7445) );
  NOR2_X1 U8857 ( .A1(n7443), .A2(n7442), .ZN(n7441) );
  INV_X1 U8858 ( .A(n7444), .ZN(n7442) );
  OAI21_X1 U8859 ( .B1(n12441), .B2(n12439), .A(n12438), .ZN(n12677) );
  XNOR2_X1 U8860 ( .A(n12796), .B(n12797), .ZN(n12680) );
  NAND2_X1 U8861 ( .A1(n14925), .A2(n6613), .ZN(n14931) );
  NAND3_X1 U8862 ( .A1(n12877), .A2(n15357), .A3(n7460), .ZN(n14977) );
  NAND2_X1 U8863 ( .A1(n15013), .A2(n15244), .ZN(n14982) );
  AOI21_X1 U8864 ( .B1(n7420), .B2(n7416), .A(n7415), .ZN(n9860) );
  OAI21_X1 U8865 ( .B1(n7418), .B2(n7421), .A(n9847), .ZN(n7415) );
  NOR2_X1 U8866 ( .A1(n7418), .A2(n15042), .ZN(n7416) );
  INV_X1 U8867 ( .A(n10349), .ZN(n9906) );
  AND2_X1 U8868 ( .A1(n12877), .A2(n15023), .ZN(n15018) );
  INV_X1 U8869 ( .A(n7382), .ZN(n7381) );
  NAND2_X1 U8870 ( .A1(n7376), .A2(n7375), .ZN(n7371) );
  NAND2_X1 U8871 ( .A1(n7077), .A2(n15365), .ZN(n15047) );
  INV_X1 U8872 ( .A(n6717), .ZN(n6715) );
  NAND2_X1 U8873 ( .A1(n7423), .A2(n9810), .ZN(n12864) );
  NAND2_X1 U8874 ( .A1(n15056), .A2(n9799), .ZN(n15043) );
  AND2_X1 U8875 ( .A1(n9826), .A2(n9804), .ZN(n15050) );
  INV_X1 U8876 ( .A(n7139), .ZN(n9791) );
  NAND2_X1 U8877 ( .A1(n6549), .A2(n7414), .ZN(n7406) );
  NAND2_X1 U8878 ( .A1(n6454), .A2(n15148), .ZN(n15094) );
  NAND2_X1 U8879 ( .A1(n15148), .A2(n7462), .ZN(n15111) );
  OAI211_X1 U8880 ( .C1(n12650), .C2(n6853), .A(n6852), .B(n10221), .ZN(n15137) );
  NAND2_X1 U8881 ( .A1(n6856), .A2(n9718), .ZN(n6852) );
  NAND2_X1 U8882 ( .A1(n15184), .A2(n9897), .ZN(n15172) );
  AND3_X1 U8883 ( .A1(n9716), .A2(n9715), .A3(n9714), .ZN(n15167) );
  NAND2_X1 U8884 ( .A1(n9925), .A2(n6724), .ZN(n15158) );
  INV_X1 U8885 ( .A(n6856), .ZN(n6855) );
  AND3_X1 U8886 ( .A1(n12232), .A2(n7457), .A3(n7458), .ZN(n15207) );
  NAND2_X1 U8887 ( .A1(n15207), .A2(n15386), .ZN(n15206) );
  OR2_X1 U8888 ( .A1(n9666), .A2(n9665), .ZN(n9699) );
  INV_X1 U8889 ( .A(n7143), .ZN(n9701) );
  AOI21_X1 U8890 ( .B1(n7368), .B2(n7370), .A(n6528), .ZN(n7366) );
  NAND2_X1 U8891 ( .A1(n6929), .A2(n6931), .ZN(n6927) );
  NAND2_X1 U8892 ( .A1(n12232), .A2(n7458), .ZN(n12653) );
  NAND2_X1 U8893 ( .A1(n7400), .A2(n7399), .ZN(n12551) );
  INV_X1 U8894 ( .A(n7398), .ZN(n7399) );
  NAND2_X1 U8895 ( .A1(n7144), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9640) );
  INV_X1 U8896 ( .A(n7059), .ZN(n9654) );
  AND3_X1 U8897 ( .A1(n11810), .A2(n6445), .A3(n7455), .ZN(n12080) );
  NAND2_X1 U8898 ( .A1(n11810), .A2(n6445), .ZN(n12081) );
  NAND2_X1 U8899 ( .A1(n9570), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U8900 ( .A1(n6971), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9600) );
  INV_X1 U8901 ( .A(n9585), .ZN(n6971) );
  NAND2_X1 U8902 ( .A1(n11810), .A2(n11922), .ZN(n11930) );
  INV_X1 U8903 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U8904 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9556) );
  NAND2_X1 U8905 ( .A1(n12116), .A2(n9541), .ZN(n11275) );
  NAND2_X1 U8906 ( .A1(n12126), .A2(n9923), .ZN(n12125) );
  NOR2_X1 U8907 ( .A1(n9506), .A2(n11203), .ZN(n11111) );
  NAND2_X1 U8908 ( .A1(n15249), .A2(n15248), .ZN(n15250) );
  AND2_X1 U8909 ( .A1(n12071), .A2(n9890), .ZN(n12161) );
  NAND2_X1 U8910 ( .A1(n10851), .A2(n10318), .ZN(n6945) );
  OR2_X1 U8911 ( .A1(n9962), .A2(n9963), .ZN(n15489) );
  INV_X1 U8912 ( .A(n15489), .ZN(n15504) );
  AND2_X1 U8913 ( .A1(n9869), .A2(n6876), .ZN(n6875) );
  AND2_X1 U8914 ( .A1(n9954), .A2(n9953), .ZN(n10830) );
  NAND2_X1 U8915 ( .A1(n10264), .A2(n10263), .ZN(n10267) );
  XNOR2_X1 U8916 ( .A(n10261), .B(n10260), .ZN(n10274) );
  NAND2_X1 U8917 ( .A1(n8448), .A2(n8447), .ZN(n9851) );
  INV_X1 U8918 ( .A(n9931), .ZN(n6734) );
  INV_X1 U8919 ( .A(n8392), .ZN(n6690) );
  INV_X1 U8920 ( .A(n8393), .ZN(n6691) );
  OAI21_X1 U8921 ( .B1(n8349), .B2(SI_23_), .A(n8389), .ZN(n8385) );
  NAND2_X1 U8922 ( .A1(n6681), .A2(n6680), .ZN(n8348) );
  INV_X1 U8923 ( .A(n8386), .ZN(n6680) );
  INV_X1 U8924 ( .A(n9777), .ZN(n6681) );
  OAI21_X1 U8925 ( .B1(SI_21_), .B2(n6697), .A(n8378), .ZN(n8325) );
  AND2_X1 U8926 ( .A1(n7470), .A2(n6876), .ZN(n9870) );
  XNOR2_X1 U8927 ( .A(n9743), .B(n9862), .ZN(n9880) );
  NAND2_X1 U8928 ( .A1(n9938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9743) );
  XNOR2_X1 U8929 ( .A(n8054), .B(n8052), .ZN(n10870) );
  NAND2_X1 U8930 ( .A1(n7595), .A2(n8029), .ZN(n8054) );
  NAND2_X1 U8931 ( .A1(n8028), .A2(n8027), .ZN(n7595) );
  XNOR2_X1 U8932 ( .A(n8028), .B(n8026), .ZN(n10851) );
  OR2_X1 U8933 ( .A1(n9562), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U8934 ( .A1(n9566), .A2(n9565), .ZN(n9594) );
  INV_X1 U8935 ( .A(n9564), .ZN(n9566) );
  NAND2_X1 U8936 ( .A1(n7973), .A2(n8002), .ZN(n7975) );
  XNOR2_X1 U8937 ( .A(n7946), .B(n7969), .ZN(n10840) );
  AND2_X1 U8938 ( .A1(n10763), .A2(n10752), .ZN(n10761) );
  XNOR2_X1 U8939 ( .A(n10815), .B(n10777), .ZN(n10810) );
  XNOR2_X1 U8940 ( .A(n10884), .B(n14877), .ZN(n10879) );
  OR2_X1 U8941 ( .A1(n10884), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10886) );
  NAND2_X1 U8942 ( .A1(n6953), .A2(n11765), .ZN(n11768) );
  NAND2_X1 U8943 ( .A1(n11761), .A2(n11760), .ZN(n6953) );
  OR2_X1 U8944 ( .A1(n11768), .A2(n7096), .ZN(n7247) );
  INV_X1 U8945 ( .A(n11769), .ZN(n7096) );
  OAI22_X1 U8946 ( .A1(n12460), .A2(n12459), .B1(P1_ADDR_REG_12__SCAN_IN), 
        .B2(n13122), .ZN(n12641) );
  NAND2_X1 U8947 ( .A1(n15429), .A2(n7242), .ZN(n7241) );
  OR2_X1 U8948 ( .A1(n15455), .A2(n15454), .ZN(n15464) );
  NAND2_X1 U8949 ( .A1(n6836), .A2(n6835), .ZN(n9153) );
  NAND2_X1 U8950 ( .A1(n10800), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U8951 ( .A1(n12172), .A2(n12171), .ZN(n12558) );
  AND2_X1 U8952 ( .A1(n7500), .A2(n11310), .ZN(n11315) );
  NAND2_X1 U8953 ( .A1(n7173), .A2(n7493), .ZN(n12985) );
  NAND2_X1 U8954 ( .A1(n7494), .A2(n12963), .ZN(n7173) );
  OAI21_X1 U8955 ( .B1(n12963), .B2(n7177), .A(n7174), .ZN(n12983) );
  NAND2_X1 U8956 ( .A1(n11687), .A2(n11686), .ZN(n11867) );
  NAND2_X1 U8957 ( .A1(n6703), .A2(n13023), .ZN(n6702) );
  INV_X1 U8958 ( .A(n13020), .ZN(n6703) );
  AOI21_X1 U8959 ( .B1(n13020), .B2(n6457), .A(n13066), .ZN(n6704) );
  INV_X1 U8960 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11557) );
  AND2_X1 U8961 ( .A1(n11561), .A2(n11551), .ZN(n11553) );
  OAI21_X1 U8962 ( .B1(n12963), .B2(n7496), .A(n7494), .ZN(n13028) );
  NAND2_X1 U8963 ( .A1(n12961), .A2(n12915), .ZN(n13030) );
  OAI21_X1 U8964 ( .B1(n12586), .B2(n12585), .A(n12584), .ZN(n12688) );
  NAND2_X1 U8965 ( .A1(n11340), .A2(n11341), .ZN(n11548) );
  NAND2_X1 U8966 ( .A1(n11326), .A2(n11325), .ZN(n13071) );
  NAND2_X1 U8967 ( .A1(n11330), .A2(n15578), .ZN(n13063) );
  NAND2_X1 U8968 ( .A1(n6643), .A2(n6515), .ZN(n13069) );
  AND2_X1 U8969 ( .A1(n9284), .A2(n9283), .ZN(n12975) );
  NAND2_X1 U8970 ( .A1(n8928), .A2(n8927), .ZN(n13086) );
  INV_X1 U8971 ( .A(n7750), .ZN(n7749) );
  OAI21_X1 U8972 ( .B1(n8561), .B2(n7751), .A(n7507), .ZN(n7750) );
  AND2_X1 U8973 ( .A1(n9243), .A2(n9242), .ZN(n15575) );
  NAND2_X1 U8974 ( .A1(n13601), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n6996) );
  AOI21_X1 U8975 ( .B1(n11483), .B2(n11481), .A(n11482), .ZN(n11480) );
  INV_X1 U8976 ( .A(n7535), .ZN(n7534) );
  NAND2_X1 U8977 ( .A1(n7364), .A2(n7365), .ZN(n11386) );
  NAND2_X1 U8978 ( .A1(n6915), .A2(n7533), .ZN(n7531) );
  NAND2_X1 U8979 ( .A1(n11884), .A2(n11885), .ZN(n11883) );
  AND2_X1 U8980 ( .A1(n7346), .A2(n7345), .ZN(n7347) );
  NAND2_X1 U8981 ( .A1(n9187), .A2(n10702), .ZN(n10706) );
  INV_X1 U8982 ( .A(n7515), .ZN(n7514) );
  NAND2_X1 U8983 ( .A1(n7516), .A2(n13115), .ZN(n12384) );
  INV_X1 U8984 ( .A(n7349), .ZN(n7348) );
  NOR2_X1 U8985 ( .A1(n12385), .A2(n7259), .ZN(n13126) );
  AND2_X1 U8986 ( .A1(n9220), .A2(n12391), .ZN(n7259) );
  NAND2_X1 U8987 ( .A1(n9160), .A2(n13169), .ZN(n13152) );
  NAND2_X1 U8988 ( .A1(n7064), .A2(n9227), .ZN(n9160) );
  INV_X1 U8989 ( .A(n7257), .ZN(n7253) );
  INV_X1 U8990 ( .A(n13154), .ZN(n7254) );
  INV_X1 U8991 ( .A(n13222), .ZN(n13200) );
  NAND2_X1 U8992 ( .A1(n7523), .A2(n7522), .ZN(n13224) );
  NOR2_X1 U8993 ( .A1(n13202), .A2(n6995), .ZN(n13227) );
  AND2_X1 U8994 ( .A1(n13203), .A2(n13204), .ZN(n6995) );
  NAND2_X1 U8995 ( .A1(n9267), .A2(n9266), .ZN(n13234) );
  XNOR2_X1 U8996 ( .A(n10409), .B(n7691), .ZN(n13237) );
  INV_X1 U8997 ( .A(n10408), .ZN(n7691) );
  OAI21_X1 U8998 ( .B1(n9062), .B2(n7672), .A(n13493), .ZN(n7671) );
  NAND2_X1 U8999 ( .A1(n9310), .A2(n8972), .ZN(n13265) );
  AOI21_X1 U9000 ( .B1(n13443), .B2(n15627), .A(n6783), .ZN(n7081) );
  OAI21_X1 U9001 ( .B1(n7738), .B2(n6474), .A(n7204), .ZN(n13303) );
  NAND2_X1 U9002 ( .A1(n7009), .A2(n8932), .ZN(n13452) );
  NAND2_X1 U9003 ( .A1(n8818), .A2(n8817), .ZN(n13414) );
  NAND2_X1 U9004 ( .A1(n7792), .A2(n6443), .ZN(n12272) );
  AND2_X1 U9005 ( .A1(n7693), .A2(n8592), .ZN(n12016) );
  NAND2_X1 U9006 ( .A1(n9022), .A2(n9021), .ZN(n12031) );
  INV_X1 U9007 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n12037) );
  INV_X1 U9008 ( .A(n13314), .ZN(n15594) );
  INV_X1 U9009 ( .A(n15587), .ZN(n15597) );
  OR2_X1 U9010 ( .A1(n11858), .A2(n11857), .ZN(n13363) );
  NAND2_X1 U9011 ( .A1(n9257), .A2(n9256), .ZN(n13228) );
  INV_X1 U9012 ( .A(n13234), .ZN(n13508) );
  AND2_X1 U9013 ( .A1(n10399), .A2(n10398), .ZN(n13246) );
  NAND2_X1 U9014 ( .A1(n8921), .A2(n8920), .ZN(n13532) );
  NAND2_X1 U9015 ( .A1(n13336), .A2(n9050), .ZN(n13317) );
  NAND2_X1 U9016 ( .A1(n8853), .A2(n8852), .ZN(n13543) );
  NAND2_X1 U9017 ( .A1(n6973), .A2(n9287), .ZN(n8853) );
  INV_X1 U9018 ( .A(n11525), .ZN(n6973) );
  NAND2_X1 U9019 ( .A1(n8871), .A2(n8870), .ZN(n13546) );
  NAND2_X1 U9020 ( .A1(n7701), .A2(n9377), .ZN(n12778) );
  NAND2_X1 U9021 ( .A1(n8774), .A2(n7705), .ZN(n7701) );
  NAND2_X1 U9022 ( .A1(n8784), .A2(n8783), .ZN(n13579) );
  NAND2_X1 U9023 ( .A1(n8774), .A2(n9299), .ZN(n13418) );
  NAND2_X1 U9024 ( .A1(n8765), .A2(n8764), .ZN(n12757) );
  NAND2_X1 U9025 ( .A1(n7154), .A2(n7155), .ZN(n12748) );
  NAND2_X1 U9026 ( .A1(n8743), .A2(n8742), .ZN(n12632) );
  NAND2_X1 U9027 ( .A1(n12522), .A2(n9034), .ZN(n12618) );
  NAND2_X1 U9028 ( .A1(n8734), .A2(n9364), .ZN(n12616) );
  OAI21_X1 U9029 ( .B1(n8681), .B2(n6449), .A(n7717), .ZN(n12529) );
  NAND2_X1 U9030 ( .A1(n8712), .A2(n8711), .ZN(n12955) );
  NAND2_X1 U9031 ( .A1(n7192), .A2(n7753), .ZN(n12330) );
  NAND2_X1 U9032 ( .A1(n7720), .A2(n9358), .ZN(n12329) );
  NAND2_X1 U9033 ( .A1(n8681), .A2(n6478), .ZN(n7720) );
  INV_X1 U9034 ( .A(n9130), .ZN(n13584) );
  INV_X1 U9035 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13588) );
  XNOR2_X1 U9036 ( .A(n9085), .B(n9084), .ZN(n12510) );
  NAND2_X1 U9037 ( .A1(n9100), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9085) );
  NAND2_X1 U9038 ( .A1(n6809), .A2(n8946), .ZN(n8959) );
  NAND2_X1 U9039 ( .A1(n9008), .A2(n9098), .ZN(n11818) );
  INV_X1 U9040 ( .A(n8902), .ZN(n7003) );
  NAND2_X1 U9041 ( .A1(n8865), .A2(n8866), .ZN(n8883) );
  NAND2_X1 U9042 ( .A1(n8825), .A2(n8824), .ZN(n8842) );
  NAND2_X1 U9043 ( .A1(n7652), .A2(n8796), .ZN(n8801) );
  NAND2_X1 U9044 ( .A1(n8721), .A2(n8720), .ZN(n8736) );
  NAND2_X1 U9045 ( .A1(n8656), .A2(n7655), .ZN(n8666) );
  NAND2_X1 U9046 ( .A1(n8656), .A2(n8655), .ZN(n8660) );
  XNOR2_X1 U9047 ( .A(n8631), .B(n8649), .ZN(n11488) );
  NAND2_X1 U9048 ( .A1(n6801), .A2(n8584), .ZN(n8599) );
  NAND2_X1 U9049 ( .A1(n8583), .A2(n8582), .ZN(n6801) );
  NAND2_X1 U9050 ( .A1(n8568), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U9051 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7344) );
  INV_X1 U9052 ( .A(SI_0_), .ZN(n10784) );
  INV_X1 U9053 ( .A(n14519), .ZN(n14310) );
  NAND2_X1 U9054 ( .A1(n7590), .A2(n8151), .ZN(n12735) );
  NAND2_X1 U9055 ( .A1(n7571), .A2(n7573), .ZN(n13628) );
  AND2_X1 U9056 ( .A1(n7573), .A2(n6485), .ZN(n13627) );
  NAND2_X1 U9057 ( .A1(n8271), .A2(n8270), .ZN(n7573) );
  NAND2_X1 U9058 ( .A1(n6677), .A2(n7561), .ZN(n11724) );
  AND2_X1 U9059 ( .A1(n11033), .A2(n7916), .ZN(n11045) );
  INV_X1 U9060 ( .A(n13706), .ZN(n7565) );
  AND2_X1 U9061 ( .A1(n6923), .A2(n6924), .ZN(n13675) );
  OR2_X1 U9062 ( .A1(n13615), .A2(n13619), .ZN(n7796) );
  NAND2_X1 U9063 ( .A1(n13685), .A2(n13684), .ZN(n13683) );
  NAND2_X1 U9064 ( .A1(n11721), .A2(n8051), .ZN(n11836) );
  NAND2_X1 U9065 ( .A1(n11836), .A2(n11837), .ZN(n11835) );
  OR2_X1 U9066 ( .A1(n11121), .A2(n14469), .ZN(n11033) );
  NAND2_X1 U9067 ( .A1(n13714), .A2(n6626), .ZN(n11035) );
  NAND2_X1 U9068 ( .A1(n7568), .A2(n7569), .ZN(n13705) );
  OR2_X1 U9069 ( .A1(n8271), .A2(n7572), .ZN(n7568) );
  NAND2_X1 U9070 ( .A1(n7578), .A2(n7579), .ZN(n12248) );
  NAND2_X1 U9071 ( .A1(n13673), .A2(n8242), .ZN(n13723) );
  NAND2_X1 U9072 ( .A1(n13663), .A2(n7968), .ZN(n11197) );
  NAND2_X1 U9073 ( .A1(n13642), .A2(n8422), .ZN(n6678) );
  AND2_X1 U9074 ( .A1(n12014), .A2(n14031), .ZN(n14072) );
  AND2_X1 U9075 ( .A1(n10899), .A2(n8519), .ZN(n14073) );
  INV_X1 U9076 ( .A(n14078), .ZN(n7594) );
  NAND2_X1 U9077 ( .A1(n8518), .A2(n8517), .ZN(n14082) );
  INV_X1 U9078 ( .A(n13735), .ZN(n14083) );
  NAND2_X1 U9079 ( .A1(n8439), .A2(n8438), .ZN(n14084) );
  OR2_X1 U9080 ( .A1(n14353), .A2(n7091), .ZN(n8403) );
  OR2_X1 U9081 ( .A1(n8146), .A2(n8145), .ZN(n14097) );
  NAND4_X1 U9082 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n7877), .ZN(n14108)
         );
  OR2_X1 U9083 ( .A1(n7910), .A2(n11374), .ZN(n7877) );
  INV_X1 U9084 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7134) );
  NAND2_X1 U9085 ( .A1(n11005), .A2(n11004), .ZN(n14116) );
  NAND2_X1 U9086 ( .A1(n15519), .A2(n6775), .ZN(n14128) );
  OR2_X1 U9087 ( .A1(n15523), .A2(n10994), .ZN(n6775) );
  NAND2_X1 U9088 ( .A1(n14129), .A2(n14128), .ZN(n14127) );
  XNOR2_X1 U9089 ( .A(n14130), .B(n10995), .ZN(n14129) );
  NAND2_X1 U9090 ( .A1(n15531), .A2(n14131), .ZN(n11010) );
  NAND2_X1 U9091 ( .A1(n14141), .A2(n6520), .ZN(n14157) );
  NAND2_X1 U9092 ( .A1(n6641), .A2(n11013), .ZN(n14174) );
  NAND2_X1 U9093 ( .A1(n14161), .A2(n14160), .ZN(n6641) );
  NAND2_X1 U9094 ( .A1(n14170), .A2(n14171), .ZN(n14169) );
  NAND2_X1 U9095 ( .A1(n14156), .A2(n6776), .ZN(n14170) );
  OR2_X1 U9096 ( .A1(n14153), .A2(n10997), .ZN(n6776) );
  NAND2_X1 U9097 ( .A1(n15547), .A2(n15548), .ZN(n15545) );
  NAND2_X1 U9098 ( .A1(n15536), .A2(n7266), .ZN(n14185) );
  OR2_X1 U9099 ( .A1(n15542), .A2(n10999), .ZN(n7266) );
  NAND2_X1 U9100 ( .A1(n14185), .A2(n14186), .ZN(n14184) );
  NOR2_X1 U9101 ( .A1(n11001), .A2(n11002), .ZN(n11404) );
  AND2_X1 U9102 ( .A1(n11398), .A2(n11397), .ZN(n14203) );
  NAND2_X1 U9103 ( .A1(n14203), .A2(n14202), .ZN(n14201) );
  NAND2_X1 U9104 ( .A1(n14195), .A2(n6611), .ZN(n11410) );
  NAND2_X1 U9105 ( .A1(n14215), .A2(n14214), .ZN(n14213) );
  AND2_X1 U9106 ( .A1(n7269), .A2(n7268), .ZN(n14209) );
  NAND2_X1 U9107 ( .A1(n14207), .A2(n6521), .ZN(n12266) );
  NAND2_X1 U9108 ( .A1(n6642), .A2(n14232), .ZN(n14249) );
  INV_X1 U9109 ( .A(n7277), .ZN(n14260) );
  NAND2_X1 U9110 ( .A1(n14274), .A2(n14257), .ZN(n14259) );
  NOR2_X1 U9111 ( .A1(n14271), .A2(n6777), .ZN(n14262) );
  NOR2_X1 U9112 ( .A1(n6778), .A2(n14255), .ZN(n6777) );
  INV_X1 U9113 ( .A(n14282), .ZN(n7279) );
  OAI211_X1 U9114 ( .C1(n7726), .C2(n10107), .A(n7725), .B(n7724), .ZN(n7723)
         );
  NAND2_X1 U9115 ( .A1(n14288), .A2(n7727), .ZN(n7726) );
  AOI21_X1 U9116 ( .B1(n6665), .B2(n14023), .A(n7907), .ZN(n7725) );
  NAND2_X1 U9117 ( .A1(n6664), .A2(n6663), .ZN(n12846) );
  OR2_X1 U9118 ( .A1(n12837), .A2(n12838), .ZN(n6664) );
  NAND2_X1 U9119 ( .A1(n7776), .A2(n7780), .ZN(n14331) );
  NAND2_X1 U9120 ( .A1(n14364), .A2(n7777), .ZN(n7776) );
  NAND2_X1 U9121 ( .A1(n7786), .A2(n7777), .ZN(n14351) );
  NAND2_X1 U9122 ( .A1(n7787), .A2(n6476), .ZN(n7786) );
  NAND2_X1 U9123 ( .A1(n7684), .A2(n10076), .ZN(n14374) );
  NAND2_X1 U9124 ( .A1(n7759), .A2(n7762), .ZN(n14379) );
  NAND2_X1 U9125 ( .A1(n10002), .A2(n10001), .ZN(n14395) );
  AND2_X1 U9126 ( .A1(n6887), .A2(n9999), .ZN(n14414) );
  INV_X1 U9127 ( .A(n10040), .ZN(n14432) );
  NAND2_X1 U9128 ( .A1(n10069), .A2(n10068), .ZN(n14441) );
  NAND2_X1 U9129 ( .A1(n14459), .A2(n10067), .ZN(n10069) );
  AND2_X1 U9130 ( .A1(n12182), .A2(n10063), .ZN(n12294) );
  NAND2_X1 U9131 ( .A1(n6896), .A2(n7764), .ZN(n12292) );
  NAND2_X1 U9132 ( .A1(n11999), .A2(n10060), .ZN(n12184) );
  NAND2_X1 U9133 ( .A1(n12001), .A2(n9984), .ZN(n12181) );
  NAND2_X1 U9134 ( .A1(n11746), .A2(n9981), .ZN(n11780) );
  INV_X1 U9135 ( .A(n14507), .ZN(n14492) );
  INV_X1 U9136 ( .A(n14497), .ZN(n14477) );
  AOI22_X1 U9137 ( .A1(n7976), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n10898), .B2(
        n14130), .ZN(n7854) );
  NAND2_X1 U9138 ( .A1(n10898), .A2(n11008), .ZN(n7060) );
  NAND2_X1 U9139 ( .A1(n7976), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U9140 ( .A1(n6894), .A2(n7900), .ZN(n7087) );
  INV_X1 U9141 ( .A(n14455), .ZN(n14511) );
  AND2_X1 U9142 ( .A1(n14293), .A2(n14584), .ZN(n10118) );
  AND2_X1 U9143 ( .A1(n14618), .A2(n15564), .ZN(n14584) );
  INV_X1 U9144 ( .A(n14293), .ZN(n10415) );
  INV_X1 U9145 ( .A(n7109), .ZN(n7108) );
  NAND2_X1 U9146 ( .A1(n14522), .A2(n7097), .ZN(n14625) );
  NOR2_X1 U9147 ( .A1(n14525), .A2(n6518), .ZN(n7097) );
  NAND2_X1 U9148 ( .A1(n14529), .A2(n7036), .ZN(n14626) );
  NOR2_X1 U9149 ( .A1(n14530), .A2(n15567), .ZN(n7038) );
  INV_X1 U9150 ( .A(n14528), .ZN(n7037) );
  INV_X1 U9151 ( .A(n15554), .ZN(n15555) );
  AND2_X1 U9152 ( .A1(n10114), .A2(n15558), .ZN(n15559) );
  INV_X1 U9153 ( .A(n15558), .ZN(n15560) );
  INV_X1 U9154 ( .A(n7875), .ZN(n14674) );
  NAND2_X1 U9155 ( .A1(n7756), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U9156 ( .A1(n8480), .A2(n8479), .ZN(n12671) );
  INV_X1 U9157 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11743) );
  INV_X1 U9158 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11337) );
  INV_X1 U9159 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11517) );
  INV_X1 U9160 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11349) );
  INV_X1 U9161 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11090) );
  INV_X1 U9162 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11066) );
  INV_X1 U9163 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10874) );
  INV_X1 U9164 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10871) );
  INV_X1 U9165 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10860) );
  INV_X1 U9166 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10862) );
  INV_X1 U9167 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10856) );
  INV_X1 U9168 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10864) );
  INV_X1 U9169 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10854) );
  INV_X1 U9170 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10803) );
  INV_X1 U9171 ( .A(n7623), .ZN(n6729) );
  AOI21_X1 U9172 ( .B1(n7623), .B2(n7625), .A(n6552), .ZN(n7621) );
  NAND2_X1 U9173 ( .A1(n14775), .A2(n10527), .ZN(n14690) );
  NOR2_X1 U9174 ( .A1(n10594), .A2(n6533), .ZN(n7613) );
  NAND2_X1 U9175 ( .A1(n7632), .A2(n10570), .ZN(n14707) );
  NAND2_X1 U9176 ( .A1(n7632), .A2(n7630), .ZN(n14708) );
  AND2_X1 U9177 ( .A1(n7616), .A2(n10511), .ZN(n12699) );
  AND3_X1 U9178 ( .A1(n9690), .A2(n9689), .A3(n9688), .ZN(n14746) );
  NAND2_X1 U9179 ( .A1(n6725), .A2(n7633), .ZN(n12100) );
  AOI21_X1 U9180 ( .B1(n7630), .B2(n6731), .A(n6498), .ZN(n6730) );
  INV_X1 U9181 ( .A(n7630), .ZN(n6732) );
  INV_X1 U9182 ( .A(n14799), .ZN(n6731) );
  AND2_X1 U9183 ( .A1(n7614), .A2(n10593), .ZN(n14788) );
  NAND2_X1 U9184 ( .A1(n10502), .A2(n7620), .ZN(n7619) );
  INV_X1 U9185 ( .A(n10503), .ZN(n7620) );
  CLKBUF_X1 U9186 ( .A(n11351), .Z(n11352) );
  AOI21_X1 U9187 ( .B1(n11417), .B2(n11416), .A(n7024), .ZN(n10483) );
  INV_X1 U9188 ( .A(n14826), .ZN(n14801) );
  NAND2_X1 U9189 ( .A1(n11516), .A2(n10318), .ZN(n9684) );
  NAND2_X1 U9190 ( .A1(n6979), .A2(n6978), .ZN(n10360) );
  INV_X1 U9191 ( .A(n6695), .ZN(n6978) );
  NAND2_X1 U9192 ( .A1(n6980), .A2(n6506), .ZN(n6979) );
  OAI211_X1 U9193 ( .C1(n10287), .C2(n6559), .A(n10311), .B(n6696), .ZN(n6695)
         );
  NAND2_X1 U9194 ( .A1(n7808), .A2(n7513), .ZN(n7512) );
  OR2_X1 U9195 ( .A1(n10359), .A2(n10358), .ZN(n7513) );
  OAI21_X1 U9196 ( .B1(n14991), .B2(n9919), .A(n9918), .ZN(n15242) );
  INV_X1 U9197 ( .A(n15013), .ZN(n15243) );
  INV_X1 U9198 ( .A(n14816), .ZN(n14833) );
  INV_X1 U9199 ( .A(n15072), .ZN(n14837) );
  INV_X1 U9200 ( .A(P1_U4016), .ZN(n14854) );
  INV_X1 U9201 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10850) );
  NOR2_X1 U9202 ( .A1(n9500), .A2(n9499), .ZN(n9501) );
  NOR2_X1 U9203 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n9499) );
  INV_X1 U9204 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10747) );
  INV_X1 U9205 ( .A(n7430), .ZN(n10923) );
  OAI21_X1 U9206 ( .B1(n11247), .B2(P1_REG1_REG_2__SCAN_IN), .A(n7029), .ZN(
        n11254) );
  NAND2_X1 U9207 ( .A1(n11247), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7029) );
  NOR2_X1 U9208 ( .A1(n11254), .A2(n11255), .ZN(n11253) );
  AND2_X1 U9209 ( .A1(n7430), .A2(n7429), .ZN(n11255) );
  NAND2_X1 U9210 ( .A1(n10924), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7429) );
  INV_X1 U9211 ( .A(n7433), .ZN(n14864) );
  NAND2_X1 U9212 ( .A1(n14872), .A2(n6486), .ZN(n10927) );
  INV_X1 U9213 ( .A(n7438), .ZN(n11261) );
  OAI21_X1 U9214 ( .B1(n14900), .B2(n14895), .A(n11265), .ZN(n14898) );
  AND2_X1 U9215 ( .A1(n6635), .A2(n6634), .ZN(n14900) );
  INV_X1 U9216 ( .A(n10984), .ZN(n6634) );
  NAND2_X1 U9217 ( .A1(n10986), .A2(n10985), .ZN(n6635) );
  NAND2_X1 U9218 ( .A1(n14889), .A2(n7434), .ZN(n11613) );
  NAND2_X1 U9219 ( .A1(n7436), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U9220 ( .A1(n14907), .A2(n7446), .ZN(n11615) );
  AND2_X1 U9221 ( .A1(n7445), .A2(n7444), .ZN(n12279) );
  NOR2_X1 U9222 ( .A1(n12285), .A2(n12284), .ZN(n12441) );
  AND2_X1 U9223 ( .A1(n12432), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7449) );
  OAI22_X1 U9224 ( .A1(n12793), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n12792), 
        .B2(n12791), .ZN(n12794) );
  INV_X1 U9225 ( .A(n14972), .ZN(n14945) );
  XNOR2_X1 U9226 ( .A(n7027), .B(n14954), .ZN(n14966) );
  NAND2_X1 U9227 ( .A1(n6538), .A2(n7028), .ZN(n7027) );
  INV_X1 U9228 ( .A(n14953), .ZN(n7028) );
  XNOR2_X1 U9229 ( .A(n6640), .B(n6639), .ZN(n14963) );
  INV_X1 U9230 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U9231 ( .A1(n14958), .A2(n14957), .ZN(n6640) );
  AND2_X1 U9232 ( .A1(n7488), .A2(n7487), .ZN(n15033) );
  NAND2_X1 U9233 ( .A1(n6947), .A2(n6946), .ZN(n15276) );
  INV_X1 U9234 ( .A(n15046), .ZN(n6946) );
  AOI21_X1 U9235 ( .B1(n15070), .B2(n9900), .A(n7377), .ZN(n15060) );
  INV_X1 U9236 ( .A(n7379), .ZN(n7377) );
  NAND2_X1 U9237 ( .A1(n7407), .A2(n9765), .ZN(n15085) );
  OAI21_X1 U9238 ( .B1(n7051), .B2(n15123), .A(n7409), .ZN(n7407) );
  NAND2_X1 U9239 ( .A1(n15122), .A2(n10219), .ZN(n15105) );
  NAND2_X1 U9240 ( .A1(n7411), .A2(n9754), .ZN(n15106) );
  NAND2_X1 U9241 ( .A1(n7413), .A2(n7412), .ZN(n7411) );
  NAND2_X1 U9242 ( .A1(n7135), .A2(n10318), .ZN(n9756) );
  INV_X1 U9243 ( .A(n12155), .ZN(n7135) );
  NAND2_X1 U9244 ( .A1(n12316), .A2(n12317), .ZN(n7367) );
  OAI21_X1 U9245 ( .B1(n12158), .B2(n7402), .A(n7401), .ZN(n12313) );
  NAND2_X1 U9246 ( .A1(n12241), .A2(n9648), .ZN(n12315) );
  INV_X1 U9247 ( .A(n15175), .ZN(n15215) );
  NAND2_X1 U9248 ( .A1(n11737), .A2(n9889), .ZN(n12073) );
  AND2_X1 U9249 ( .A1(n6863), .A2(n6862), .ZN(n11734) );
  NAND2_X1 U9250 ( .A1(n11109), .A2(n11108), .ZN(n11107) );
  NAND2_X1 U9251 ( .A1(n7393), .A2(n9517), .ZN(n11109) );
  INV_X1 U9252 ( .A(n15196), .ZN(n15212) );
  NAND2_X1 U9253 ( .A1(n10318), .A2(n10819), .ZN(n9526) );
  AOI21_X1 U9254 ( .B1(n10319), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n6489), .ZN(
        n6846) );
  AND2_X2 U9255 ( .A1(n10367), .A2(n11902), .ZN(n15518) );
  AND2_X1 U9256 ( .A1(n15231), .A2(n15230), .ZN(n15354) );
  INV_X1 U9257 ( .A(n15259), .ZN(n15260) );
  NOR2_X1 U9258 ( .A1(n7113), .A2(n15276), .ZN(n15362) );
  NAND2_X1 U9259 ( .A1(n7115), .A2(n7114), .ZN(n7113) );
  INV_X1 U9260 ( .A(n15277), .ZN(n7114) );
  NAND2_X1 U9261 ( .A1(n15278), .A2(n15494), .ZN(n7115) );
  INV_X1 U9262 ( .A(n15115), .ZN(n15375) );
  AND2_X1 U9263 ( .A1(n10653), .A2(n10833), .ZN(n15790) );
  NAND2_X1 U9264 ( .A1(n9498), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9494) );
  INV_X1 U9265 ( .A(n9951), .ZN(n12222) );
  OR2_X1 U9266 ( .A1(n9777), .A2(n10801), .ZN(n9778) );
  INV_X1 U9267 ( .A(n9927), .ZN(n15403) );
  INV_X1 U9268 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11510) );
  INV_X1 U9269 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11336) );
  INV_X1 U9270 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n15732) );
  INV_X1 U9271 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n15740) );
  INV_X1 U9272 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n11065) );
  INV_X1 U9273 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10919) );
  NAND2_X1 U9274 ( .A1(n6951), .A2(n6950), .ZN(n6949) );
  INV_X1 U9275 ( .A(n8057), .ZN(n6950) );
  NAND2_X1 U9276 ( .A1(n7339), .A2(n7338), .ZN(n6951) );
  INV_X1 U9277 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10852) );
  INV_X1 U9278 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10796) );
  NAND2_X2 U9279 ( .A1(n7453), .A2(n7450), .ZN(n10929) );
  NAND2_X1 U9280 ( .A1(n7452), .A2(n7451), .ZN(n7450) );
  INV_X1 U9281 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7452) );
  XNOR2_X1 U9282 ( .A(n10810), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n10782) );
  NAND3_X1 U9283 ( .A1(n6959), .A2(n6956), .A3(n6954), .ZN(n10970) );
  NAND2_X1 U9284 ( .A1(n6958), .A2(n6957), .ZN(n6956) );
  NAND2_X1 U9285 ( .A1(n10970), .A2(n10971), .ZN(n11095) );
  XNOR2_X1 U9286 ( .A(n11764), .B(n11762), .ZN(n11761) );
  XNOR2_X1 U9287 ( .A(n11768), .B(n11769), .ZN(n15407) );
  AOI21_X1 U9288 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(n12466), .A(n12465), .ZN(
        n12639) );
  NAND2_X1 U9289 ( .A1(n15421), .A2(n15420), .ZN(n15423) );
  NAND2_X1 U9290 ( .A1(n15423), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n15430) );
  NAND2_X1 U9291 ( .A1(n15418), .A2(n15419), .ZN(n15431) );
  INV_X1 U9292 ( .A(n15421), .ZN(n15418) );
  OAI21_X1 U9293 ( .B1(n15446), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n15445), .ZN(
        n15462) );
  NAND2_X1 U9294 ( .A1(n9434), .A2(n6463), .ZN(n7131) );
  AOI21_X1 U9295 ( .B1(n7080), .B2(n7078), .A(n6464), .ZN(n7132) );
  NAND2_X1 U9296 ( .A1(n7360), .A2(n10684), .ZN(n13133) );
  OR4_X1 U9297 ( .A1(n10701), .A2(n10700), .A3(n10699), .A4(n10698), .ZN(
        P3_U3196) );
  NOR2_X1 U9298 ( .A1(n7021), .A2(n7357), .ZN(n7020) );
  NOR2_X1 U9299 ( .A1(n7053), .A2(n6615), .ZN(n7052) );
  NOR2_X1 U9300 ( .A1(n15639), .A2(n12887), .ZN(n7053) );
  NOR2_X1 U9301 ( .A1(n7045), .A2(n6608), .ZN(n7044) );
  NOR2_X1 U9302 ( .A1(n15631), .A2(n10411), .ZN(n7045) );
  NAND2_X1 U9303 ( .A1(n7581), .A2(n7582), .ZN(n11978) );
  NAND2_X1 U9304 ( .A1(n12861), .A2(n6488), .ZN(n12860) );
  OAI21_X1 U9305 ( .B1(n7558), .B2(n14102), .A(n7557), .ZN(P2_U3531) );
  NAND2_X1 U9306 ( .A1(n14102), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7557) );
  INV_X1 U9307 ( .A(n7269), .ZN(n12260) );
  NOR2_X1 U9308 ( .A1(n7280), .A2(n7279), .ZN(n7278) );
  AOI21_X1 U9309 ( .B1(n14515), .B2(n14507), .A(n10046), .ZN(n10101) );
  NAND2_X1 U9310 ( .A1(n15573), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7068) );
  NAND2_X1 U9311 ( .A1(n15570), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7098) );
  XNOR2_X1 U9312 ( .A(n7026), .B(n7025), .ZN(n14819) );
  INV_X1 U9313 ( .A(n6720), .ZN(n15254) );
  OR2_X1 U9314 ( .A1(n12881), .A2(n7490), .ZN(n7489) );
  NAND2_X1 U9315 ( .A1(n15267), .A2(n12880), .ZN(n7491) );
  MUX2_X1 U9316 ( .A(n15227), .B(n15226), .S(n15518), .Z(n15228) );
  OR2_X1 U9317 ( .A1(n15518), .A2(n9916), .ZN(n7394) );
  NAND2_X1 U9318 ( .A1(n15358), .A2(n15518), .ZN(n7395) );
  NAND2_X1 U9319 ( .A1(n15244), .A2(n12215), .ZN(n9964) );
  AOI21_X1 U9320 ( .B1(n15244), .B2(n10371), .A(n10370), .ZN(n10372) );
  AND2_X1 U9321 ( .A1(n6968), .A2(n7120), .ZN(n12452) );
  INV_X1 U9322 ( .A(n7350), .ZN(n13111) );
  AND2_X1 U9323 ( .A1(n9032), .A2(n9031), .ZN(n6443) );
  NAND2_X2 U9324 ( .A1(n10259), .A2(n10127), .ZN(n10139) );
  INV_X1 U9325 ( .A(n15049), .ZN(n15365) );
  OR2_X1 U9326 ( .A1(n8189), .A2(SI_15_), .ZN(n6444) );
  AND2_X1 U9327 ( .A1(n9924), .A2(n7456), .ZN(n6445) );
  AND2_X1 U9328 ( .A1(n6881), .A2(n10174), .ZN(n6446) );
  AND2_X1 U9329 ( .A1(n13880), .A2(n13882), .ZN(n6447) );
  AOI21_X1 U9330 ( .B1(n13277), .B2(n6458), .A(n6562), .ZN(n7209) );
  INV_X1 U9331 ( .A(n7731), .ZN(n7728) );
  INV_X2 U9332 ( .A(n7849), .ZN(n10898) );
  NAND2_X2 U9333 ( .A1(n10422), .A2(n9878), .ZN(n10449) );
  INV_X4 U9334 ( .A(n7907), .ZN(n14469) );
  AND2_X1 U9335 ( .A1(n7849), .A2(n10801), .ZN(n6448) );
  OR2_X1 U9336 ( .A1(n8719), .A2(n7719), .ZN(n6449) );
  INV_X1 U9337 ( .A(n8372), .ZN(n6925) );
  INV_X1 U9338 ( .A(n10593), .ZN(n10594) );
  AND2_X1 U9339 ( .A1(n9985), .A2(n7765), .ZN(n6450) );
  AND2_X1 U9340 ( .A1(n7582), .A2(n7580), .ZN(n6452) );
  NOR2_X1 U9341 ( .A1(n7441), .A2(n12278), .ZN(n6453) );
  AND2_X1 U9342 ( .A1(n7462), .A2(n7461), .ZN(n6454) );
  AND2_X1 U9343 ( .A1(n6556), .A2(n7290), .ZN(n6455) );
  AND4_X1 U9344 ( .A1(n8773), .A2(n8772), .A3(n8771), .A4(n8770), .ZN(n12687)
         );
  INV_X1 U9345 ( .A(n12687), .ZN(n13095) );
  AND2_X1 U9346 ( .A1(n7771), .A2(n14465), .ZN(n6456) );
  AND2_X1 U9347 ( .A1(n6707), .A2(n13085), .ZN(n6457) );
  AND2_X1 U9348 ( .A1(n9055), .A2(n9056), .ZN(n6458) );
  NOR2_X1 U9349 ( .A1(n14527), .A2(n14084), .ZN(n6459) );
  AND2_X1 U9350 ( .A1(n7178), .A2(n8865), .ZN(n6460) );
  AND3_X1 U9351 ( .A1(n6595), .A2(n6870), .A3(n6869), .ZN(n6461) );
  AND2_X1 U9352 ( .A1(n10158), .A2(n10157), .ZN(n6462) );
  AND2_X1 U9353 ( .A1(n9435), .A2(n6623), .ZN(n6463) );
  NAND2_X1 U9354 ( .A1(n10786), .A2(n7501), .ZN(n8568) );
  AND2_X1 U9355 ( .A1(n9449), .A2(n6623), .ZN(n6464) );
  NAND2_X1 U9356 ( .A1(n8388), .A2(n8387), .ZN(n6465) );
  INV_X1 U9357 ( .A(n12043), .ZN(n7754) );
  AND2_X1 U9358 ( .A1(n7764), .A2(n9986), .ZN(n6466) );
  AND2_X1 U9359 ( .A1(n7730), .A2(n7729), .ZN(n6467) );
  AND2_X1 U9360 ( .A1(n9898), .A2(n10201), .ZN(n15140) );
  NOR2_X1 U9361 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n6468) );
  AND2_X1 U9362 ( .A1(n13983), .A2(n13982), .ZN(n6469) );
  NAND2_X2 U9363 ( .A1(n14989), .A2(n15208), .ZN(n15482) );
  INV_X1 U9364 ( .A(n14057), .ZN(n6759) );
  INV_X1 U9365 ( .A(n14584), .ZN(n7043) );
  AND2_X1 U9366 ( .A1(n7324), .A2(n10013), .ZN(n6470) );
  AND2_X1 U9367 ( .A1(n14291), .A2(n14510), .ZN(n6471) );
  INV_X1 U9368 ( .A(n13840), .ZN(n7119) );
  INV_X1 U9369 ( .A(n10320), .ZN(n7333) );
  AND2_X1 U9370 ( .A1(n7525), .A2(n9238), .ZN(n6472) );
  AND2_X1 U9371 ( .A1(n7525), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6473) );
  INV_X1 U9372 ( .A(n11388), .ZN(n6916) );
  INV_X2 U9373 ( .A(n9516), .ZN(n9534) );
  NAND2_X1 U9374 ( .A1(n8990), .A2(n8989), .ZN(n12934) );
  NAND2_X1 U9375 ( .A1(n9290), .A2(n9289), .ZN(n13253) );
  XNOR2_X1 U9376 ( .A(n13840), .B(n14103), .ZN(n14050) );
  NAND2_X1 U9377 ( .A1(n7536), .A2(n13160), .ZN(n13174) );
  NAND4_X1 U9378 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n13105)
         );
  AND4_X1 U9379 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n9020)
         );
  NAND2_X1 U9380 ( .A1(n8962), .A2(n8961), .ZN(n13520) );
  NAND2_X1 U9381 ( .A1(n6928), .A2(n9892), .ZN(n12316) );
  INV_X1 U9382 ( .A(n8547), .ZN(n7509) );
  NAND2_X2 U9383 ( .A1(n9684), .A2(n9683), .ZN(n15213) );
  INV_X1 U9384 ( .A(n15099), .ZN(n7461) );
  INV_X1 U9385 ( .A(n9900), .ZN(n15075) );
  NAND2_X1 U9386 ( .A1(n6673), .A2(n7586), .ZN(n13649) );
  NAND2_X1 U9387 ( .A1(n6807), .A2(n8977), .ZN(n13270) );
  NAND2_X1 U9388 ( .A1(n9997), .A2(n9996), .ZN(n14420) );
  AOI21_X1 U9389 ( .B1(n13420), .B2(n9041), .A(n7798), .ZN(n13378) );
  INV_X1 U9390 ( .A(n7210), .ZN(n7211) );
  MUX2_X1 U9391 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14687), .S(n7849), .Z(n13763)
         );
  INV_X1 U9392 ( .A(n13763), .ZN(n13755) );
  OR2_X1 U9393 ( .A1(n7206), .A2(n9052), .ZN(n6474) );
  AND2_X1 U9394 ( .A1(n13856), .A2(n13855), .ZN(n6475) );
  INV_X1 U9395 ( .A(n7753), .ZN(n7752) );
  AOI21_X1 U9396 ( .B1(n6443), .B2(n12043), .A(n6531), .ZN(n7753) );
  NAND2_X1 U9397 ( .A1(n14541), .A2(n14087), .ZN(n6476) );
  NAND2_X1 U9398 ( .A1(n8224), .A2(n8223), .ZN(n6477) );
  INV_X1 U9399 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7873) );
  INV_X1 U9400 ( .A(n14622), .ZN(n12838) );
  NAND2_X1 U9401 ( .A1(n10376), .A2(n10375), .ZN(n14622) );
  INV_X1 U9402 ( .A(n12185), .ZN(n10061) );
  NOR2_X1 U9403 ( .A1(n7721), .A2(n9359), .ZN(n6478) );
  AND2_X1 U9404 ( .A1(n14450), .A2(n10070), .ZN(n6479) );
  NAND3_X1 U9405 ( .A1(n12648), .A2(n10187), .A3(n10199), .ZN(n6480) );
  OR2_X1 U9406 ( .A1(n15104), .A2(n7480), .ZN(n6481) );
  INV_X1 U9407 ( .A(n13972), .ZN(n7606) );
  NAND2_X1 U9408 ( .A1(n15070), .A2(n7380), .ZN(n7376) );
  XNOR2_X1 U9409 ( .A(n13026), .B(n8958), .ZN(n13289) );
  INV_X1 U9410 ( .A(n13289), .ZN(n7010) );
  NAND2_X1 U9411 ( .A1(n8190), .A2(n8193), .ZN(n6482) );
  INV_X1 U9412 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U9413 ( .A1(n12584), .A2(n13095), .ZN(n6483) );
  CLKBUF_X1 U9414 ( .A(n10439), .Z(n10588) );
  XNOR2_X1 U9415 ( .A(n15258), .B(n14816), .ZN(n15010) );
  AND2_X1 U9416 ( .A1(n14303), .A2(n10008), .ZN(n6484) );
  XNOR2_X1 U9417 ( .A(n14519), .B(n13735), .ZN(n14305) );
  INV_X1 U9418 ( .A(n14305), .ZN(n14300) );
  INV_X1 U9419 ( .A(n12492), .ZN(n7772) );
  NAND2_X1 U9420 ( .A1(n7876), .A2(n7875), .ZN(n7910) );
  INV_X1 U9421 ( .A(n7572), .ZN(n7571) );
  NAND2_X1 U9422 ( .A1(n13629), .A2(n6485), .ZN(n7572) );
  INV_X1 U9423 ( .A(n15123), .ZN(n7412) );
  NAND2_X1 U9424 ( .A1(n8269), .A2(n8268), .ZN(n6485) );
  NAND2_X1 U9425 ( .A1(n7773), .A2(n12492), .ZN(n12716) );
  NAND2_X1 U9426 ( .A1(n7367), .A2(n9893), .ZN(n12545) );
  NAND2_X1 U9427 ( .A1(n7679), .A2(n10066), .ZN(n14479) );
  OR2_X1 U9428 ( .A1(n14879), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U9429 ( .A1(n9150), .A2(n11891), .ZN(n7346) );
  XNOR2_X1 U9430 ( .A(n8651), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11388) );
  AND2_X1 U9431 ( .A1(n9554), .A2(n9553), .ZN(n11952) );
  AND2_X1 U9432 ( .A1(n11247), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6487) );
  AND2_X1 U9433 ( .A1(n8674), .A2(n8673), .ZN(n13490) );
  INV_X1 U9434 ( .A(n11160), .ZN(n6821) );
  XNOR2_X1 U9435 ( .A(n8615), .B(P3_IR_REG_5__SCAN_IN), .ZN(n11160) );
  INV_X1 U9436 ( .A(n9299), .ZN(n7706) );
  AND3_X1 U9437 ( .A1(n12852), .A2(n12856), .A3(n13714), .ZN(n6488) );
  NAND2_X1 U9438 ( .A1(n12549), .A2(n9673), .ZN(n12650) );
  AND2_X1 U9439 ( .A1(n6437), .A2(n11247), .ZN(n6489) );
  INV_X1 U9440 ( .A(n15042), .ZN(n7424) );
  AND3_X1 U9441 ( .A1(n9443), .A2(n9427), .A3(n9393), .ZN(n6490) );
  OR3_X1 U9442 ( .A1(n14067), .A2(n14068), .A3(n14305), .ZN(n6491) );
  INV_X1 U9443 ( .A(n14853), .ZN(n6844) );
  AND2_X1 U9444 ( .A1(n13860), .A2(n14099), .ZN(n6492) );
  NOR2_X1 U9445 ( .A1(n14938), .A2(n7428), .ZN(n6493) );
  OR2_X1 U9446 ( .A1(n6469), .A2(n13987), .ZN(n6494) );
  NAND2_X1 U9447 ( .A1(n9824), .A2(n9823), .ZN(n15035) );
  NOR2_X1 U9448 ( .A1(n14725), .A2(n10592), .ZN(n6495) );
  OR2_X1 U9449 ( .A1(n14071), .A2(n7788), .ZN(n6496) );
  AND3_X1 U9450 ( .A1(n8595), .A2(n8594), .A3(n7165), .ZN(n6497) );
  AND2_X1 U9451 ( .A1(n10577), .A2(n10576), .ZN(n6498) );
  AND3_X1 U9452 ( .A1(n9373), .A2(n12749), .A3(n9372), .ZN(n6499) );
  AND2_X1 U9453 ( .A1(n8085), .A2(n8084), .ZN(n6500) );
  AND2_X1 U9454 ( .A1(n12918), .A2(n13087), .ZN(n6501) );
  AND2_X1 U9455 ( .A1(n13805), .A2(n13804), .ZN(n6502) );
  AND2_X1 U9456 ( .A1(n7409), .A2(n7411), .ZN(n6503) );
  NAND2_X1 U9457 ( .A1(n9357), .A2(n9356), .ZN(n6504) );
  NOR2_X1 U9458 ( .A1(n12074), .A2(n7384), .ZN(n6505) );
  NOR2_X1 U9459 ( .A1(n10287), .A2(n10282), .ZN(n6506) );
  AND2_X1 U9460 ( .A1(n13174), .A2(n7542), .ZN(n6507) );
  INV_X1 U9461 ( .A(n6723), .ZN(n15077) );
  INV_X1 U9462 ( .A(n15264), .ZN(n12868) );
  NAND2_X1 U9463 ( .A1(n7817), .A2(SI_1_), .ZN(n7884) );
  INV_X1 U9464 ( .A(n9358), .ZN(n7719) );
  INV_X1 U9465 ( .A(n12322), .ZN(n12708) );
  NAND2_X1 U9466 ( .A1(n9652), .A2(n9651), .ZN(n12322) );
  AND3_X1 U9467 ( .A1(n8613), .A2(n6645), .A3(n6644), .ZN(n6508) );
  AND2_X1 U9468 ( .A1(n7153), .A2(n7155), .ZN(n6509) );
  NOR2_X1 U9469 ( .A1(n9168), .A2(n9173), .ZN(n6510) );
  AND2_X1 U9470 ( .A1(n8378), .A2(n8919), .ZN(n6511) );
  INV_X1 U9471 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7822) );
  AND2_X1 U9472 ( .A1(n8153), .A2(n8152), .ZN(n6512) );
  AND2_X1 U9473 ( .A1(n10165), .A2(n10164), .ZN(n6513) );
  AND2_X1 U9474 ( .A1(n7786), .A2(n7783), .ZN(n6514) );
  AND2_X1 U9475 ( .A1(n12902), .A2(n12903), .ZN(n6515) );
  INV_X1 U9476 ( .A(n9042), .ZN(n7744) );
  AND2_X1 U9477 ( .A1(n9083), .A2(n9082), .ZN(n6516) );
  AND2_X1 U9478 ( .A1(n7119), .A2(n10036), .ZN(n6517) );
  INV_X1 U9479 ( .A(n6718), .ZN(n15034) );
  NAND2_X1 U9480 ( .A1(n7077), .A2(n6715), .ZN(n6718) );
  INV_X1 U9481 ( .A(n10244), .ZN(n7556) );
  OR2_X1 U9482 ( .A1(n14521), .A2(n14520), .ZN(n6518) );
  AND2_X1 U9483 ( .A1(n6861), .A2(n9888), .ZN(n6519) );
  OR2_X1 U9484 ( .A1(n14138), .A2(n10996), .ZN(n6520) );
  OR2_X1 U9485 ( .A1(n14211), .A2(n12264), .ZN(n6521) );
  OR2_X1 U9486 ( .A1(n12678), .A2(n12679), .ZN(n6522) );
  INV_X1 U9487 ( .A(n7447), .ZN(n7446) );
  AND2_X1 U9488 ( .A1(n6818), .A2(n6821), .ZN(n6523) );
  INV_X1 U9489 ( .A(n7713), .ZN(n13375) );
  NAND2_X1 U9490 ( .A1(n7714), .A2(n9389), .ZN(n7713) );
  XNOR2_X1 U9491 ( .A(n8224), .B(SI_16_), .ZN(n8221) );
  AND2_X1 U9492 ( .A1(n10004), .A2(n7762), .ZN(n6524) );
  INV_X1 U9493 ( .A(n9415), .ZN(n7162) );
  NAND2_X1 U9494 ( .A1(n6807), .A2(n6805), .ZN(n9415) );
  INV_X1 U9495 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7056) );
  INV_X1 U9496 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8544) );
  INV_X1 U9497 ( .A(n6966), .ZN(n6965) );
  NOR2_X1 U9498 ( .A1(n12450), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6966) );
  AND2_X1 U9499 ( .A1(n12364), .A2(n12365), .ZN(n6525) );
  AND2_X1 U9500 ( .A1(n7697), .A2(n7694), .ZN(n6526) );
  INV_X1 U9501 ( .A(n7418), .ZN(n7417) );
  NAND2_X1 U9502 ( .A1(n15010), .A2(n9836), .ZN(n7418) );
  NAND2_X1 U9503 ( .A1(n10501), .A2(n10500), .ZN(n6527) );
  NOR2_X1 U9504 ( .A1(n12552), .A2(n12701), .ZN(n6528) );
  NOR2_X1 U9505 ( .A1(n14655), .A2(n12713), .ZN(n6529) );
  NOR2_X1 U9506 ( .A1(n11460), .A2(n12050), .ZN(n6530) );
  NOR2_X1 U9507 ( .A1(n12485), .A2(n12559), .ZN(n6531) );
  NOR2_X1 U9508 ( .A1(n14629), .A2(n14085), .ZN(n6532) );
  AND2_X1 U9509 ( .A1(n10598), .A2(n10597), .ZN(n6533) );
  AND2_X1 U9510 ( .A1(n14087), .A2(n13818), .ZN(n6534) );
  AND2_X1 U9511 ( .A1(n7621), .A2(n6727), .ZN(n6535) );
  INV_X1 U9512 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10872) );
  AND2_X1 U9513 ( .A1(n14536), .A2(n14086), .ZN(n6536) );
  INV_X1 U9514 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U9515 ( .A1(n15148), .A2(n15132), .ZN(n15110) );
  AND2_X1 U9516 ( .A1(n8025), .A2(n8024), .ZN(n6537) );
  OR2_X1 U9517 ( .A1(n6493), .A2(n14952), .ZN(n6538) );
  AND2_X1 U9518 ( .A1(n14068), .A2(n6884), .ZN(n6539) );
  INV_X1 U9519 ( .A(n14638), .ZN(n7763) );
  OR2_X1 U9520 ( .A1(n6759), .A2(n6447), .ZN(n6540) );
  AND2_X1 U9521 ( .A1(n13812), .A2(n13811), .ZN(n6541) );
  AND3_X1 U9522 ( .A1(n9540), .A2(n9539), .A3(n9538), .ZN(n10469) );
  INV_X1 U9523 ( .A(n10469), .ZN(n7106) );
  AND2_X1 U9524 ( .A1(n12917), .A2(n13088), .ZN(n6542) );
  AND2_X1 U9525 ( .A1(n13835), .A2(n13834), .ZN(n6543) );
  OAI21_X1 U9526 ( .B1(n14676), .B2(n10270), .A(n10269), .ZN(n10333) );
  OR2_X1 U9527 ( .A1(n9211), .A2(n10788), .ZN(n6544) );
  NOR2_X1 U9528 ( .A1(n12283), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6545) );
  AND2_X1 U9529 ( .A1(n9404), .A2(n13338), .ZN(n6546) );
  INV_X1 U9530 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9865) );
  NOR2_X1 U9531 ( .A1(n10249), .A2(n10248), .ZN(n6547) );
  INV_X1 U9532 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9478) );
  INV_X1 U9533 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10858) );
  INV_X1 U9534 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10839) );
  INV_X1 U9535 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10875) );
  INV_X1 U9536 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10841) );
  NAND2_X1 U9537 ( .A1(n11488), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6548) );
  NOR2_X1 U9538 ( .A1(n15123), .A2(n7408), .ZN(n6549) );
  AND2_X1 U9539 ( .A1(n12637), .A2(n15665), .ZN(n6550) );
  INV_X1 U9540 ( .A(n7656), .ZN(n7655) );
  NAND2_X1 U9541 ( .A1(n8658), .A2(n8655), .ZN(n7656) );
  NAND2_X1 U9542 ( .A1(n6918), .A2(n7971), .ZN(n6551) );
  INV_X1 U9543 ( .A(n9176), .ZN(n6814) );
  AND2_X1 U9544 ( .A1(n10636), .A2(n10635), .ZN(n6552) );
  OR2_X1 U9545 ( .A1(n7639), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U9546 ( .A1(n12523), .A2(n12520), .ZN(n6554) );
  OR2_X1 U9547 ( .A1(n9288), .A2(n10792), .ZN(n6555) );
  AND2_X1 U9548 ( .A1(n13911), .A2(n13902), .ZN(n6556) );
  AND2_X1 U9549 ( .A1(n13987), .A2(n6469), .ZN(n6557) );
  OR2_X1 U9550 ( .A1(n8383), .A2(n7330), .ZN(n6558) );
  INV_X1 U9551 ( .A(n7063), .ZN(n6822) );
  NOR2_X1 U9552 ( .A1(n11236), .A2(n9144), .ZN(n7063) );
  OR2_X1 U9553 ( .A1(n10286), .A2(n10285), .ZN(n6559) );
  INV_X1 U9554 ( .A(n14023), .ZN(n14288) );
  AND2_X1 U9555 ( .A1(n8441), .A2(n8440), .ZN(n6560) );
  OR2_X1 U9556 ( .A1(n14365), .A2(n14536), .ZN(n6561) );
  AND2_X1 U9557 ( .A1(n13520), .A2(n13083), .ZN(n6562) );
  INV_X1 U9558 ( .A(n14527), .ZN(n14325) );
  NAND2_X1 U9559 ( .A1(n8430), .A2(n8429), .ZN(n14527) );
  NAND2_X1 U9560 ( .A1(n14024), .A2(n13997), .ZN(n14036) );
  INV_X1 U9561 ( .A(n9055), .ZN(n9057) );
  OR2_X1 U9562 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6563) );
  OR2_X1 U9563 ( .A1(n7576), .A2(n8406), .ZN(n6564) );
  INV_X1 U9564 ( .A(n11448), .ZN(n7532) );
  AND2_X1 U9565 ( .A1(n14531), .A2(n14589), .ZN(n6565) );
  OR2_X1 U9566 ( .A1(n9168), .A2(n10786), .ZN(n6566) );
  AND2_X1 U9567 ( .A1(n13249), .A2(n8999), .ZN(n9418) );
  AND2_X1 U9568 ( .A1(n7254), .A2(n7253), .ZN(n6567) );
  INV_X1 U9569 ( .A(n9427), .ZN(n9440) );
  OR2_X1 U9570 ( .A1(n13253), .A2(n10403), .ZN(n9427) );
  OR2_X1 U9571 ( .A1(n12451), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6568) );
  NOR2_X1 U9572 ( .A1(n13270), .A2(n13082), .ZN(n6569) );
  NOR2_X1 U9573 ( .A1(n14445), .A2(n9998), .ZN(n6570) );
  AND2_X1 U9574 ( .A1(n9322), .A2(n9316), .ZN(n6571) );
  NOR2_X1 U9575 ( .A1(n14622), .A2(n14516), .ZN(n7727) );
  INV_X1 U9576 ( .A(n7727), .ZN(n6665) );
  AND2_X1 U9577 ( .A1(n8156), .A2(n8157), .ZN(n6572) );
  AND2_X1 U9578 ( .A1(n10511), .A2(n12698), .ZN(n6573) );
  OR2_X1 U9579 ( .A1(n6707), .A2(n13085), .ZN(n6574) );
  NOR2_X1 U9580 ( .A1(n14532), .A2(n6565), .ZN(n6575) );
  AND2_X1 U9581 ( .A1(n8600), .A2(n8585), .ZN(n8598) );
  OR2_X1 U9582 ( .A1(n13969), .A2(n13968), .ZN(n6576) );
  NAND2_X2 U9583 ( .A1(n7170), .A2(n7169), .ZN(n12906) );
  INV_X1 U9584 ( .A(n12906), .ZN(n11312) );
  AND2_X1 U9585 ( .A1(n9023), .A2(n9021), .ZN(n6577) );
  NOR2_X1 U9586 ( .A1(n9179), .A2(n11145), .ZN(n9181) );
  INV_X1 U9587 ( .A(n15258), .ZN(n15023) );
  AND2_X1 U9588 ( .A1(n10000), .A2(n14413), .ZN(n6578) );
  AND2_X1 U9589 ( .A1(n7633), .A2(n6527), .ZN(n6579) );
  NAND2_X1 U9590 ( .A1(n14527), .A2(n14084), .ZN(n6580) );
  AND2_X1 U9591 ( .A1(n7187), .A2(n8551), .ZN(n6581) );
  INV_X1 U9592 ( .A(n13885), .ZN(n7291) );
  NAND2_X1 U9593 ( .A1(n10352), .A2(n10323), .ZN(n6582) );
  AND2_X1 U9594 ( .A1(n6822), .A2(n11160), .ZN(n6583) );
  OR2_X1 U9595 ( .A1(n10171), .A2(n10169), .ZN(n6584) );
  INV_X1 U9596 ( .A(n8029), .ZN(n7597) );
  NAND2_X1 U9597 ( .A1(n7343), .A2(SI_7_), .ZN(n8029) );
  OR2_X1 U9598 ( .A1(n10245), .A2(n7556), .ZN(n6585) );
  AND2_X1 U9599 ( .A1(n13918), .A2(n7289), .ZN(n6586) );
  AND2_X1 U9600 ( .A1(n15032), .A2(n7487), .ZN(n6587) );
  AND2_X1 U9601 ( .A1(n7160), .A2(n9306), .ZN(n6588) );
  AND2_X1 U9602 ( .A1(n13998), .A2(n6738), .ZN(n6589) );
  NAND2_X1 U9603 ( .A1(n13968), .A2(n13969), .ZN(n6590) );
  AND2_X1 U9604 ( .A1(n9082), .A2(n7503), .ZN(n6591) );
  INV_X1 U9605 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7871) );
  AND2_X1 U9606 ( .A1(n6581), .A2(n8544), .ZN(n6592) );
  OR2_X1 U9607 ( .A1(n12322), .A2(n14843), .ZN(n6593) );
  INV_X1 U9608 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9496) );
  OR2_X1 U9609 ( .A1(n11236), .A2(n12022), .ZN(n6594) );
  AND2_X1 U9610 ( .A1(n7564), .A2(n11465), .ZN(n7563) );
  NAND2_X1 U9611 ( .A1(n10236), .A2(n7554), .ZN(n6595) );
  OR2_X1 U9612 ( .A1(n13438), .A2(n13437), .ZN(P3_U3487) );
  INV_X1 U9613 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7187) );
  AND2_X1 U9614 ( .A1(n7472), .A2(n9481), .ZN(n6597) );
  OR2_X1 U9615 ( .A1(n13513), .A2(n13512), .ZN(P3_U3455) );
  OR2_X1 U9616 ( .A1(n13256), .A2(n13255), .ZN(P3_U3205) );
  OR2_X1 U9617 ( .A1(n7848), .A2(n7847), .ZN(n6600) );
  BUF_X1 U9618 ( .A(n10139), .Z(n7046) );
  NAND2_X1 U9619 ( .A1(n12423), .A2(n8132), .ZN(n12470) );
  AND2_X1 U9620 ( .A1(n12411), .A2(n6666), .ZN(n12500) );
  INV_X1 U9621 ( .A(n14228), .ZN(n7272) );
  AND2_X1 U9622 ( .A1(n12163), .A2(n12234), .ZN(n12232) );
  AND2_X1 U9623 ( .A1(n7514), .A2(n13115), .ZN(n6601) );
  NAND2_X1 U9624 ( .A1(n12182), .A2(n7682), .ZN(n12293) );
  NAND2_X1 U9625 ( .A1(n6755), .A2(n14057), .ZN(n12406) );
  AND2_X1 U9626 ( .A1(n12232), .A2(n12708), .ZN(n6602) );
  NAND2_X1 U9627 ( .A1(n12017), .A2(n9026), .ZN(n12056) );
  INV_X1 U9628 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7075) );
  NAND2_X1 U9629 ( .A1(n6709), .A2(n7179), .ZN(n12899) );
  NAND2_X1 U9630 ( .A1(n7149), .A2(n9344), .ZN(n11714) );
  NAND2_X1 U9631 ( .A1(n10209), .A2(n10199), .ZN(n15218) );
  INV_X1 U9632 ( .A(n15218), .ZN(n7084) );
  OR2_X1 U9633 ( .A1(n9849), .A2(n13599), .ZN(n6603) );
  INV_X1 U9634 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7435) );
  INV_X1 U9635 ( .A(n7118), .ZN(n7807) );
  INV_X1 U9636 ( .A(n9925), .ZN(n15157) );
  OR2_X1 U9637 ( .A1(n9223), .A2(n13146), .ZN(n6604) );
  NOR2_X1 U9638 ( .A1(n13477), .A2(n13093), .ZN(n6605) );
  INV_X1 U9639 ( .A(n10179), .ZN(n6878) );
  INV_X1 U9640 ( .A(n14557), .ZN(n7058) );
  NOR2_X1 U9641 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9674) );
  AND2_X1 U9642 ( .A1(n13137), .A2(n13138), .ZN(n6606) );
  AND4_X1 U9643 ( .A1(n6657), .A2(n8115), .A3(n6656), .A4(n6655), .ZN(n6607)
         );
  INV_X1 U9644 ( .A(n13167), .ZN(n7256) );
  AND2_X1 U9645 ( .A1(n10412), .A2(n9136), .ZN(n6608) );
  NAND2_X1 U9646 ( .A1(n12500), .A2(n6467), .ZN(n7731) );
  AND2_X1 U9647 ( .A1(n7637), .A2(n7636), .ZN(n6609) );
  AND2_X1 U9648 ( .A1(n10015), .A2(n15760), .ZN(n6610) );
  INV_X1 U9649 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10820) );
  OR2_X1 U9650 ( .A1(n14198), .A2(n11408), .ZN(n6611) );
  OR2_X1 U9651 ( .A1(n11584), .A2(n11583), .ZN(n6612) );
  OR2_X1 U9652 ( .A1(n14927), .A2(n14926), .ZN(n6613) );
  INV_X1 U9653 ( .A(n9765), .ZN(n7408) );
  OR2_X1 U9654 ( .A1(n11777), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6968) );
  NAND2_X1 U9655 ( .A1(n6834), .A2(n6837), .ZN(n6836) );
  AND2_X1 U9656 ( .A1(n7590), .A2(n7589), .ZN(n6614) );
  INV_X1 U9657 ( .A(n15244), .ZN(n14997) );
  NOR2_X1 U9658 ( .A1(n13240), .A2(n13485), .ZN(n6615) );
  NAND2_X1 U9659 ( .A1(n8315), .A2(n8316), .ZN(n6616) );
  INV_X1 U9660 ( .A(n7502), .ZN(n8866) );
  INV_X1 U9661 ( .A(n6967), .ZN(n12465) );
  AND2_X1 U9662 ( .A1(n10945), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6617) );
  INV_X1 U9663 ( .A(n8322), .ZN(n8323) );
  AND2_X1 U9664 ( .A1(n6603), .A2(n10013), .ZN(n6618) );
  AND2_X1 U9665 ( .A1(n7046), .A2(n7335), .ZN(n6619) );
  AND2_X1 U9666 ( .A1(n7792), .A2(n9031), .ZN(n6620) );
  OR2_X1 U9667 ( .A1(n10185), .A2(n10183), .ZN(n6621) );
  AND2_X1 U9668 ( .A1(n11923), .A2(n9888), .ZN(n6622) );
  INV_X1 U9669 ( .A(n8219), .ZN(n6924) );
  AND2_X2 U9670 ( .A1(n10386), .A2(n10117), .ZN(n14618) );
  INV_X1 U9671 ( .A(n15639), .ZN(n15637) );
  INV_X1 U9672 ( .A(n15338), .ZN(n7457) );
  NOR2_X1 U9673 ( .A1(n11449), .A2(n7533), .ZN(n11383) );
  NAND2_X1 U9674 ( .A1(n8120), .A2(n8119), .ZN(n14599) );
  INV_X1 U9675 ( .A(n14599), .ZN(n7117) );
  AND2_X1 U9676 ( .A1(n11949), .A2(n11952), .ZN(n11810) );
  NOR2_X1 U9677 ( .A1(n11376), .A2(n6667), .ZN(n11578) );
  INV_X1 U9678 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6700) );
  AND2_X1 U9679 ( .A1(n9454), .A2(n9075), .ZN(n6623) );
  INV_X1 U9680 ( .A(n13397), .ZN(n13493) );
  AND2_X1 U9681 ( .A1(n10037), .A2(n10036), .ZN(n6624) );
  NOR2_X1 U9682 ( .A1(n9147), .A2(n11388), .ZN(n11455) );
  INV_X1 U9683 ( .A(n15327), .ZN(n15300) );
  AND2_X2 U9684 ( .A1(n9133), .A2(n11328), .ZN(n15631) );
  INV_X1 U9685 ( .A(n6915), .ZN(n11449) );
  NAND2_X1 U9686 ( .A1(n6917), .A2(n6916), .ZN(n6915) );
  INV_X1 U9687 ( .A(n14651), .ZN(n7729) );
  AND2_X1 U9688 ( .A1(n9231), .A2(n13182), .ZN(n6625) );
  INV_X1 U9689 ( .A(n12217), .ZN(n7455) );
  AND3_X1 U9690 ( .A1(n14486), .A2(n11121), .A3(n7559), .ZN(n6626) );
  NAND2_X1 U9691 ( .A1(n7499), .A2(n7498), .ZN(n7500) );
  NAND2_X1 U9692 ( .A1(n11124), .A2(n14042), .ZN(n11123) );
  AND2_X1 U9693 ( .A1(n13217), .A2(n7352), .ZN(n6627) );
  NAND2_X1 U9694 ( .A1(n14714), .A2(n14716), .ZN(n14715) );
  AND2_X1 U9695 ( .A1(n7531), .A2(n11448), .ZN(n6628) );
  NAND2_X1 U9696 ( .A1(n7611), .A2(n10464), .ZN(n11361) );
  INV_X1 U9697 ( .A(n7545), .ZN(n7544) );
  AND2_X1 U9698 ( .A1(n12670), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6629) );
  INV_X1 U9699 ( .A(n7066), .ZN(n7065) );
  NOR2_X1 U9700 ( .A1(n10696), .A2(n13481), .ZN(n7066) );
  AND2_X1 U9701 ( .A1(n11810), .A2(n7456), .ZN(n11735) );
  AND2_X1 U9702 ( .A1(n14243), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6630) );
  AND2_X1 U9703 ( .A1(n12401), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6631) );
  INV_X1 U9704 ( .A(n13219), .ZN(n7525) );
  INV_X1 U9705 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12220) );
  XNOR2_X1 U9706 ( .A(n7869), .B(P2_IR_REG_19__SCAN_IN), .ZN(n14280) );
  INV_X1 U9707 ( .A(n14280), .ZN(n14031) );
  XOR2_X1 U9708 ( .A(n13182), .B(P3_REG1_REG_16__SCAN_IN), .Z(n6632) );
  INV_X1 U9709 ( .A(n6432), .ZN(n12825) );
  AND2_X1 U9710 ( .A1(n9608), .A2(n9596), .ZN(n14901) );
  INV_X1 U9711 ( .A(n14901), .ZN(n7436) );
  AND2_X1 U9712 ( .A1(n6900), .A2(n6901), .ZN(n6633) );
  INV_X1 U9714 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7124) );
  INV_X1 U9715 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n6985) );
  INV_X1 U9716 ( .A(SI_8_), .ZN(n6998) );
  INV_X1 U9717 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7751) );
  INV_X1 U9718 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7022) );
  INV_X1 U9719 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7242) );
  OR2_X1 U9720 ( .A1(n9195), .A2(n9236), .ZN(n6909) );
  AND2_X1 U9721 ( .A1(n9195), .A2(n9236), .ZN(n6907) );
  AND2_X2 U9722 ( .A1(n6637), .A2(n11244), .ZN(n9535) );
  NAND2_X1 U9723 ( .A1(n15532), .A2(n15533), .ZN(n15531) );
  MUX2_X1 U9724 ( .A(n11648), .B(P2_REG2_REG_2__SCAN_IN), .S(n15523), .Z(
        n15533) );
  NAND2_X1 U9725 ( .A1(n7882), .A2(n7979), .ZN(n15523) );
  OR2_X2 U9726 ( .A1(n14256), .A2(n14255), .ZN(n14274) );
  XNOR2_X2 U9727 ( .A(n12765), .B(n12771), .ZN(n12763) );
  NAND2_X1 U9728 ( .A1(n14174), .A2(n14173), .ZN(n11015) );
  NAND2_X1 U9729 ( .A1(n11012), .A2(n11011), .ZN(n14161) );
  OAI211_X1 U9730 ( .C1(n6642), .C2(n14232), .A(n14249), .B(n15546), .ZN(
        n14233) );
  NAND2_X1 U9731 ( .A1(n14231), .A2(n14230), .ZN(n6642) );
  OR2_X2 U9732 ( .A1(n11026), .A2(n11025), .ZN(n11398) );
  NAND2_X1 U9733 ( .A1(n14191), .A2(n11023), .ZN(n11026) );
  NAND2_X1 U9734 ( .A1(n6643), .A2(n12902), .ZN(n13068) );
  NAND3_X1 U9735 ( .A1(n7497), .A2(n7500), .A3(n6650), .ZN(n11339) );
  NAND2_X1 U9736 ( .A1(n11311), .A2(n12557), .ZN(n6650) );
  AND2_X2 U9737 ( .A1(n7692), .A2(n9017), .ZN(n13495) );
  NAND3_X1 U9738 ( .A1(n7188), .A2(n8542), .A3(n6581), .ZN(n6651) );
  AND2_X1 U9739 ( .A1(n9092), .A2(n6652), .ZN(n9104) );
  NAND2_X1 U9740 ( .A1(n11548), .A2(n11547), .ZN(n11563) );
  NAND2_X2 U9741 ( .A1(n13045), .A2(n12912), .ZN(n12963) );
  NAND3_X1 U9742 ( .A1(n13594), .A2(n8545), .A3(P3_REG0_REG_0__SCAN_IN), .ZN(
        n6654) );
  NAND4_X1 U9743 ( .A1(n8550), .A2(n8548), .A3(n8549), .A4(n6654), .ZN(n13108)
         );
  AND4_X2 U9744 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .ZN(n7133)
         );
  NOR2_X2 U9745 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6658) );
  AOI21_X1 U9746 ( .B1(n7727), .B2(n6662), .A(n7907), .ZN(n6663) );
  NAND2_X1 U9747 ( .A1(n12846), .A2(n12842), .ZN(n14620) );
  AND2_X2 U9748 ( .A1(n14396), .A2(n7763), .ZN(n14397) );
  NAND3_X1 U9749 ( .A1(n11701), .A2(n7732), .A3(n9970), .ZN(n6667) );
  NOR2_X1 U9750 ( .A1(n6434), .A2(n11509), .ZN(n8227) );
  NAND2_X1 U9751 ( .A1(n7976), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U9752 ( .A1(n7976), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U9753 ( .A1(n7976), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8345) );
  NAND2_X1 U9754 ( .A1(n7976), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U9755 ( .A1(n7976), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U9756 ( .A1(n7976), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U9757 ( .A1(n7976), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8429) );
  NAND2_X1 U9758 ( .A1(n7976), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U9759 ( .A1(n7976), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U9760 ( .A1(n7976), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10009) );
  NAND2_X1 U9761 ( .A1(n7976), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10375) );
  NAND2_X1 U9762 ( .A1(n7976), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n10377) );
  INV_X4 U9763 ( .A(n6668), .ZN(n7976) );
  OAI22_X1 U9764 ( .A1(n14237), .A2(n7849), .B1(n11337), .B2(n6434), .ZN(n8200) );
  OAI22_X1 U9765 ( .A1(n12261), .A2(n7849), .B1(n11066), .B2(n6434), .ZN(n8118) );
  NAND2_X1 U9766 ( .A1(n12423), .A2(n6674), .ZN(n6673) );
  NAND3_X1 U9767 ( .A1(n7563), .A2(n13663), .A3(n7968), .ZN(n6677) );
  INV_X1 U9768 ( .A(n11724), .ZN(n6676) );
  NAND3_X1 U9769 ( .A1(n11073), .A2(n13692), .A3(n11057), .ZN(n7941) );
  OAI21_X2 U9770 ( .B1(n15003), .B2(n9904), .A(n10349), .ZN(n14983) );
  NAND2_X1 U9771 ( .A1(n14997), .A2(n10139), .ZN(n6694) );
  NAND4_X1 U9772 ( .A1(n6705), .A2(n6704), .A3(n6702), .A4(n6701), .ZN(n6706)
         );
  NAND3_X1 U9773 ( .A1(n13021), .A2(n6707), .A3(n13020), .ZN(n6701) );
  NAND2_X1 U9774 ( .A1(n6706), .A2(n13027), .ZN(P3_U3169) );
  INV_X1 U9775 ( .A(n13023), .ZN(n6707) );
  AOI21_X2 U9776 ( .B1(n11867), .B2(n11866), .A(n11865), .ZN(n11869) );
  INV_X1 U9777 ( .A(n12567), .ZN(n6711) );
  NAND2_X1 U9778 ( .A1(n8762), .A2(n8761), .ZN(n8781) );
  NAND4_X1 U9779 ( .A1(n8762), .A2(n9004), .A3(n8761), .A4(n6516), .ZN(n9100)
         );
  NAND2_X1 U9780 ( .A1(n6713), .A2(n7814), .ZN(n7887) );
  OAI21_X1 U9781 ( .B1(n7944), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n6714), .ZN(
        n6713) );
  NAND4_X1 U9782 ( .A1(n7795), .A2(n6722), .A3(n6721), .A4(n6719), .ZN(n15358)
         );
  NAND3_X1 U9783 ( .A1(n15370), .A2(n6454), .A3(n15148), .ZN(n6723) );
  INV_X1 U9784 ( .A(n15319), .ZN(n6724) );
  NAND2_X1 U9785 ( .A1(n10618), .A2(n10617), .ZN(n14731) );
  NAND3_X2 U9786 ( .A1(n7387), .A2(n9536), .A3(n7386), .ZN(n9932) );
  NAND2_X1 U9787 ( .A1(n6735), .A2(n7594), .ZN(n7593) );
  NAND3_X1 U9788 ( .A1(n6736), .A2(n14035), .A3(n6496), .ZN(n6735) );
  NAND2_X1 U9789 ( .A1(n6737), .A2(n7039), .ZN(n6736) );
  AOI21_X1 U9790 ( .B1(n14071), .B2(n14070), .A(n13756), .ZN(n6737) );
  NAND3_X1 U9791 ( .A1(n6741), .A2(n14036), .A3(n6589), .ZN(n6743) );
  NAND3_X1 U9792 ( .A1(n6743), .A2(n14018), .A3(n14017), .ZN(n14028) );
  NAND2_X1 U9793 ( .A1(n8221), .A2(n6745), .ZN(n6747) );
  INV_X1 U9794 ( .A(n6745), .ZN(n8195) );
  NAND2_X1 U9795 ( .A1(n8194), .A2(n8193), .ZN(n6746) );
  NAND3_X1 U9796 ( .A1(n7062), .A2(n11569), .A3(n7680), .ZN(n11574) );
  OAI22_X2 U9797 ( .A1(n12293), .A2(n6540), .B1(n6756), .B2(n6447), .ZN(n12712) );
  AND2_X1 U9798 ( .A1(n10065), .A2(n6757), .ZN(n6756) );
  NAND2_X1 U9799 ( .A1(n14459), .A2(n6760), .ZN(n6766) );
  NOR2_X1 U9800 ( .A1(n6764), .A2(n10072), .ZN(n6763) );
  AND2_X1 U9801 ( .A1(n10047), .A2(n7070), .ZN(n14042) );
  NAND2_X2 U9802 ( .A1(n14674), .A2(n6770), .ZN(n10380) );
  NAND2_X1 U9803 ( .A1(n6771), .A2(n14280), .ZN(n7281) );
  NAND2_X1 U9804 ( .A1(n12266), .A2(n12265), .ZN(n12770) );
  NAND2_X1 U9805 ( .A1(n6782), .A2(n7666), .ZN(n7663) );
  NAND2_X1 U9806 ( .A1(n6782), .A2(n8918), .ZN(n8931) );
  NAND2_X1 U9807 ( .A1(n6782), .A2(n7669), .ZN(n7665) );
  NAND2_X1 U9808 ( .A1(n8904), .A2(n6782), .ZN(n12827) );
  XNOR2_X1 U9809 ( .A(n13281), .B(n13282), .ZN(n13443) );
  NAND3_X1 U9810 ( .A1(n8598), .A2(n8582), .A3(n8583), .ZN(n6800) );
  INV_X1 U9811 ( .A(n6815), .ZN(n11183) );
  NOR2_X1 U9812 ( .A1(n6812), .A2(n6811), .ZN(n6810) );
  NAND2_X1 U9813 ( .A1(n6815), .A2(n6813), .ZN(n6812) );
  OAI21_X1 U9814 ( .B1(n10687), .B2(n6830), .A(n6827), .ZN(n6825) );
  NAND3_X1 U9815 ( .A1(n7345), .A2(n7346), .A3(P3_REG1_REG_9__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U9816 ( .A1(n6840), .A2(n10197), .ZN(n10200) );
  INV_X1 U9817 ( .A(n6840), .ZN(n10196) );
  NAND2_X1 U9818 ( .A1(n10125), .A2(n10122), .ZN(n7519) );
  NAND2_X1 U9819 ( .A1(n9507), .A2(n9506), .ZN(n10133) );
  NAND3_X1 U9820 ( .A1(n6842), .A2(n7385), .A3(n6841), .ZN(n12117) );
  NAND3_X1 U9821 ( .A1(n10135), .A2(n11167), .A3(n11164), .ZN(n6841) );
  NAND2_X1 U9822 ( .A1(n10133), .A2(n10132), .ZN(n11167) );
  AND3_X1 U9824 ( .A1(n9524), .A2(n9521), .A3(n9523), .ZN(n6847) );
  NAND2_X1 U9825 ( .A1(n14855), .A2(n11987), .ZN(n10132) );
  AND2_X1 U9826 ( .A1(n7419), .A2(n9836), .ZN(n15011) );
  OAI21_X1 U9827 ( .B1(n12650), .B2(n15178), .A(n6855), .ZN(n15177) );
  NAND3_X1 U9828 ( .A1(n6851), .A2(n9718), .A3(n6850), .ZN(n15156) );
  NAND2_X1 U9829 ( .A1(n6855), .A2(n15178), .ZN(n6850) );
  NAND2_X1 U9830 ( .A1(n12650), .A2(n6855), .ZN(n6851) );
  OR2_X1 U9831 ( .A1(n15178), .A2(n6854), .ZN(n6853) );
  INV_X1 U9832 ( .A(n9718), .ZN(n6854) );
  INV_X1 U9833 ( .A(n11733), .ZN(n6861) );
  NOR2_X1 U9834 ( .A1(n7799), .A2(n6861), .ZN(n6860) );
  INV_X1 U9835 ( .A(n7799), .ZN(n6863) );
  NAND2_X1 U9836 ( .A1(n6874), .A2(n7553), .ZN(n10239) );
  NAND2_X1 U9837 ( .A1(n7470), .A2(n6875), .ZN(n9928) );
  OAI22_X1 U9838 ( .A1(n10159), .A2(n6462), .B1(n10157), .B2(n10158), .ZN(
        n10162) );
  OAI21_X1 U9839 ( .B1(n10173), .B2(n6446), .A(n6880), .ZN(n10178) );
  NAND2_X1 U9840 ( .A1(n6879), .A2(n6877), .ZN(n10177) );
  NAND2_X1 U9841 ( .A1(n10173), .A2(n6880), .ZN(n6879) );
  AND2_X1 U9842 ( .A1(n6600), .A2(n6883), .ZN(n6882) );
  NAND2_X1 U9843 ( .A1(n7844), .A2(n7842), .ZN(n6883) );
  NAND2_X1 U9844 ( .A1(n14300), .A2(n10008), .ZN(n6884) );
  NAND2_X1 U9845 ( .A1(n14304), .A2(n14305), .ZN(n14303) );
  NAND3_X1 U9846 ( .A1(n9997), .A2(n6570), .A3(n9996), .ZN(n6887) );
  OAI21_X1 U9847 ( .B1(n11534), .B2(n6892), .A(n6888), .ZN(n6890) );
  NAND2_X1 U9848 ( .A1(n6890), .A2(n7757), .ZN(n9983) );
  NOR2_X1 U9849 ( .A1(n10801), .A2(n10803), .ZN(n6895) );
  OAI21_X1 U9850 ( .B1(n6893), .B2(n6895), .A(n7849), .ZN(n6894) );
  NAND2_X1 U9851 ( .A1(n6896), .A2(n6466), .ZN(n12290) );
  NAND2_X1 U9852 ( .A1(n9181), .A2(n6902), .ZN(n6901) );
  INV_X1 U9853 ( .A(n11231), .ZN(n6902) );
  NAND4_X1 U9854 ( .A1(n6905), .A2(n6908), .A3(n6906), .A4(n6903), .ZN(n9246)
         );
  NAND3_X1 U9855 ( .A1(n7523), .A2(n6907), .A3(n7522), .ZN(n6905) );
  NAND2_X1 U9856 ( .A1(n11151), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n11483) );
  OAI21_X1 U9857 ( .B1(n7923), .B2(SI_4_), .A(n6918), .ZN(n7925) );
  NAND2_X1 U9858 ( .A1(n7943), .A2(n6918), .ZN(n7946) );
  NAND3_X1 U9859 ( .A1(n6926), .A2(n6927), .A3(n7366), .ZN(n12647) );
  NAND2_X1 U9860 ( .A1(n12230), .A2(n6929), .ZN(n6926) );
  XNOR2_X2 U9861 ( .A(n15307), .B(n14839), .ZN(n15123) );
  NAND2_X2 U9862 ( .A1(n9745), .A2(n9744), .ZN(n15307) );
  INV_X2 U9863 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15465) );
  AND2_X4 U9864 ( .A1(n6936), .A2(n6935), .ZN(n7944) );
  NAND4_X1 U9865 ( .A1(n14283), .A2(n7812), .A3(n7813), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6936) );
  NAND3_X1 U9866 ( .A1(n6944), .A2(n6942), .A3(n6572), .ZN(n7100) );
  NAND2_X1 U9867 ( .A1(n6943), .A2(n6512), .ZN(n6942) );
  NAND3_X1 U9868 ( .A1(n8088), .A2(n6512), .A3(n8087), .ZN(n6944) );
  NAND2_X1 U9869 ( .A1(n8007), .A2(n8008), .ZN(n8028) );
  NAND3_X1 U9870 ( .A1(n6948), .A2(n7488), .A3(n15327), .ZN(n6947) );
  NAND2_X1 U9871 ( .A1(n8073), .A2(n6949), .ZN(n10876) );
  NAND2_X1 U9872 ( .A1(n8273), .A2(n6952), .ZN(n11745) );
  NAND3_X1 U9873 ( .A1(n8273), .A2(n6952), .A3(n10318), .ZN(n9734) );
  NAND2_X1 U9874 ( .A1(n8248), .A2(n8292), .ZN(n6952) );
  INV_X1 U9875 ( .A(n10889), .ZN(n6955) );
  NAND2_X1 U9876 ( .A1(n10968), .A2(n6960), .ZN(n6957) );
  NAND3_X1 U9877 ( .A1(n6955), .A2(n10968), .A3(P2_ADDR_REG_7__SCAN_IN), .ZN(
        n6954) );
  NAND2_X1 U9878 ( .A1(n10889), .A2(n10888), .ZN(n10969) );
  NAND2_X1 U9879 ( .A1(n10889), .A2(n6961), .ZN(n6959) );
  NAND2_X1 U9880 ( .A1(n10969), .A2(n10968), .ZN(n11093) );
  NAND3_X1 U9881 ( .A1(n6964), .A2(n6963), .A3(n6965), .ZN(n12458) );
  NAND3_X1 U9882 ( .A1(n6964), .A2(n6963), .A3(n6962), .ZN(n6967) );
  INV_X1 U9883 ( .A(n7120), .ZN(n12088) );
  OAI21_X1 U9884 ( .B1(n15409), .B2(n6970), .A(n6969), .ZN(n15421) );
  NOR2_X1 U9885 ( .A1(n15442), .A2(n15441), .ZN(n15446) );
  AOI22_X1 U9886 ( .A1(n15462), .A2(n15461), .B1(n15460), .B2(n15459), .ZN(
        n15470) );
  NAND3_X1 U9887 ( .A1(n15430), .A2(n15431), .A3(n15429), .ZN(n15434) );
  NAND2_X1 U9888 ( .A1(n12999), .A2(n12998), .ZN(n12997) );
  INV_X1 U9889 ( .A(n10775), .ZN(n7023) );
  NAND2_X1 U9890 ( .A1(n7023), .A2(n7022), .ZN(n10776) );
  NAND3_X1 U9891 ( .A1(n7342), .A2(n10360), .A3(n10362), .ZN(n7005) );
  XNOR2_X1 U9892 ( .A(n6972), .B(n14967), .ZN(n10356) );
  AND2_X1 U9893 ( .A1(n10353), .A2(n10352), .ZN(n6972) );
  NAND2_X1 U9894 ( .A1(n7059), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9666) );
  OAI22_X2 U9895 ( .A1(n13057), .A2(n13058), .B1(n13082), .B2(n12930), .ZN(
        n12971) );
  NAND2_X1 U9896 ( .A1(n7054), .A2(n12391), .ZN(n7516) );
  NAND3_X1 U9897 ( .A1(n7020), .A2(n7260), .A3(n7351), .ZN(P3_U3201) );
  NAND2_X1 U9898 ( .A1(n8619), .A2(n8618), .ZN(n8633) );
  NAND2_X1 U9899 ( .A1(n8880), .A2(n8879), .ZN(n8882) );
  NAND2_X1 U9900 ( .A1(n8848), .A2(n12013), .ZN(n7640) );
  NAND2_X1 U9901 ( .A1(n9251), .A2(n9250), .ZN(n9286) );
  AOI21_X1 U9902 ( .B1(n7210), .B2(n7209), .A(n6569), .ZN(n7207) );
  NAND2_X1 U9903 ( .A1(n9061), .A2(n9060), .ZN(n10399) );
  AOI21_X1 U9904 ( .B1(n9434), .B2(n9435), .A(n9449), .ZN(n9439) );
  INV_X1 U9905 ( .A(n7780), .ZN(n7779) );
  OAI21_X1 U9906 ( .B1(n10407), .B2(n13397), .A(n10406), .ZN(n13242) );
  INV_X1 U9907 ( .A(n7141), .ZN(n8397) );
  AOI21_X1 U9908 ( .B1(n7110), .B2(n6580), .A(n6459), .ZN(n14304) );
  OAI21_X1 U9909 ( .B1(n12886), .B2(n15629), .A(n7044), .ZN(P3_U3456) );
  OAI21_X1 U9910 ( .B1(n9453), .B2(n9452), .A(n9451), .ZN(n9464) );
  NAND2_X1 U9911 ( .A1(n9464), .A2(n7012), .ZN(n9461) );
  NAND2_X1 U9912 ( .A1(n13664), .A2(n13665), .ZN(n13663) );
  NAND2_X1 U9913 ( .A1(n13636), .A2(n13635), .ZN(n13634) );
  AOI21_X1 U9914 ( .B1(n12248), .B2(n12247), .A(n8106), .ZN(n12422) );
  NAND2_X1 U9915 ( .A1(n7548), .A2(n7550), .ZN(n10159) );
  NOR2_X1 U9916 ( .A1(n13694), .A2(n13691), .ZN(n7940) );
  NAND2_X1 U9917 ( .A1(n7936), .A2(n7942), .ZN(n13694) );
  NAND2_X1 U9918 ( .A1(n6981), .A2(n8533), .ZN(P2_U3186) );
  NAND3_X1 U9919 ( .A1(n8503), .A2(n12861), .A3(n13714), .ZN(n6981) );
  NAND3_X1 U9920 ( .A1(n15434), .A2(n7240), .A3(n7241), .ZN(n15442) );
  NAND2_X2 U9921 ( .A1(n13756), .A2(n12014), .ZN(n14033) );
  NAND2_X1 U9922 ( .A1(n12117), .A2(n12119), .ZN(n12116) );
  NAND2_X1 U9923 ( .A1(n7524), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13221) );
  OR2_X1 U9924 ( .A1(n9915), .A2(n10925), .ZN(n9522) );
  INV_X1 U9925 ( .A(n9188), .ZN(n7054) );
  OAI211_X1 U9926 ( .C1(n13227), .C2(n13226), .A(n13225), .B(n7016), .ZN(n7015) );
  AND4_X2 U9927 ( .A1(n8708), .A2(n8538), .A3(n8709), .A4(n8761), .ZN(n8542)
         );
  INV_X2 U9928 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10786) );
  NAND3_X2 U9929 ( .A1(n7501), .A2(n10786), .A3(n8534), .ZN(n8759) );
  NAND2_X1 U9931 ( .A1(n7362), .A2(n11453), .ZN(n11457) );
  NAND2_X1 U9932 ( .A1(n7168), .A2(n6591), .ZN(n7502) );
  INV_X4 U9933 ( .A(n12557), .ZN(n12972) );
  NAND2_X1 U9934 ( .A1(n8090), .A2(n8089), .ZN(n8107) );
  NAND2_X1 U9935 ( .A1(n7596), .A2(n8055), .ZN(n7338) );
  NAND2_X2 U9936 ( .A1(n11419), .A2(n10487), .ZN(n11528) );
  OR2_X2 U9937 ( .A1(n14259), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14275) );
  INV_X1 U9938 ( .A(n11420), .ZN(n7024) );
  AOI21_X1 U9939 ( .B1(n14279), .B2(n15546), .A(n7283), .ZN(n7282) );
  OAI21_X1 U9940 ( .B1(n9058), .B2(n7210), .A(n7209), .ZN(n13267) );
  NOR2_X1 U9941 ( .A1(n13189), .A2(n6992), .ZN(n9234) );
  AOI22_X1 U9942 ( .A1(n11149), .A2(n11150), .B1(n11160), .B2(n9207), .ZN(
        n11473) );
  NAND2_X1 U9943 ( .A1(n7470), .A2(n7471), .ZN(n15392) );
  INV_X1 U9944 ( .A(n10166), .ZN(n7033) );
  NAND2_X1 U9945 ( .A1(n7033), .A2(n7032), .ZN(n10168) );
  OAI21_X1 U9946 ( .B1(n13601), .B2(n11287), .A(n6996), .ZN(n9198) );
  INV_X1 U9947 ( .A(n8052), .ZN(n8053) );
  NAND2_X1 U9948 ( .A1(n6999), .A2(n6998), .ZN(n6997) );
  NAND2_X1 U9949 ( .A1(n7000), .A2(n7566), .ZN(n13636) );
  NAND2_X1 U9950 ( .A1(n7071), .A2(n7339), .ZN(n8073) );
  AOI21_X1 U9951 ( .B1(n14028), .B2(n14027), .A(n14026), .ZN(n14071) );
  INV_X1 U9952 ( .A(n8972), .ZN(n7001) );
  OAI21_X1 U9953 ( .B1(n8027), .B2(n7597), .A(n8053), .ZN(n7596) );
  NAND2_X1 U9954 ( .A1(n8301), .A2(n8300), .ZN(n8384) );
  NAND2_X1 U9955 ( .A1(n7004), .A2(n7003), .ZN(n8904) );
  INV_X1 U9956 ( .A(n8903), .ZN(n7004) );
  OAI211_X1 U9957 ( .C1(n7511), .C2(n10360), .A(n10365), .B(n7005), .ZN(
        P1_U3242) );
  NAND2_X1 U9958 ( .A1(n12226), .A2(n9287), .ZN(n7009) );
  NAND2_X1 U9959 ( .A1(n7665), .A2(n8929), .ZN(n8943) );
  INV_X1 U9960 ( .A(n13262), .ZN(n9077) );
  NOR2_X1 U9961 ( .A1(n13257), .A2(n9078), .ZN(n9134) );
  NOR2_X1 U9962 ( .A1(n13316), .A2(n7235), .ZN(n7234) );
  NAND2_X1 U9963 ( .A1(n7017), .A2(n7014), .ZN(P3_U3200) );
  INV_X1 U9964 ( .A(n7015), .ZN(n7014) );
  NAND2_X1 U9965 ( .A1(n13218), .A2(n13217), .ZN(n7017) );
  NAND2_X1 U9966 ( .A1(n7095), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U9967 ( .A1(n9152), .A2(n9151), .ZN(n7345) );
  NAND2_X1 U9968 ( .A1(n13188), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13208) );
  NAND2_X1 U9969 ( .A1(n11153), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U9970 ( .A1(n7111), .A2(n14517), .ZN(n14624) );
  NAND2_X1 U9971 ( .A1(n14624), .A2(n14618), .ZN(n7069) );
  OAI21_X1 U9972 ( .B1(n14364), .B2(n7779), .A(n7778), .ZN(n10007) );
  BUF_X4 U9973 ( .A(n7944), .Z(n10801) );
  NAND2_X1 U9974 ( .A1(n7067), .A2(n8323), .ZN(n8321) );
  NAND2_X1 U9975 ( .A1(n8319), .A2(n8302), .ZN(n8303) );
  NAND2_X1 U9976 ( .A1(n7414), .A2(n9765), .ZN(n7405) );
  AOI21_X1 U9977 ( .B1(n14917), .B2(n11622), .A(n11621), .ZN(n11825) );
  XNOR2_X2 U9978 ( .A(n9548), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14868) );
  INV_X1 U9979 ( .A(n8568), .ZN(n7095) );
  NAND2_X1 U9980 ( .A1(n10706), .A2(n7055), .ZN(n9188) );
  NOR2_X1 U9981 ( .A1(n9183), .A2(n7107), .ZN(n11151) );
  NAND2_X1 U9982 ( .A1(n10766), .A2(n10773), .ZN(n10774) );
  NAND2_X1 U9983 ( .A1(n7440), .A2(n7439), .ZN(n12280) );
  NAND2_X2 U9984 ( .A1(n11528), .A2(n11527), .ZN(n11526) );
  AOI22_X2 U9985 ( .A1(n11613), .A2(n11612), .B1(n11619), .B2(n15666), .ZN(
        n14909) );
  INV_X1 U9986 ( .A(n11600), .ZN(n10448) );
  NOR2_X1 U9987 ( .A1(n12431), .A2(n7449), .ZN(n12433) );
  NAND2_X1 U9988 ( .A1(n13695), .A2(n7942), .ZN(n13664) );
  INV_X1 U9989 ( .A(n7030), .ZN(n11044) );
  OAI21_X2 U9990 ( .B1(n14348), .B2(n10081), .A(n10083), .ZN(n14333) );
  OAI21_X1 U9991 ( .B1(n7908), .B2(n7909), .A(n7917), .ZN(n7030) );
  NAND2_X1 U9992 ( .A1(n7031), .A2(n10134), .ZN(n10138) );
  NAND3_X1 U9993 ( .A1(n10334), .A2(n10130), .A3(n10131), .ZN(n7031) );
  OAI21_X1 U9994 ( .B1(n10152), .B2(n10151), .A(n10150), .ZN(n10154) );
  OAI21_X1 U9995 ( .B1(n6513), .B2(n7034), .A(n7552), .ZN(n10173) );
  AOI21_X1 U9996 ( .B1(n10200), .B2(n7791), .A(n7046), .ZN(n10212) );
  OAI21_X1 U9997 ( .B1(n7469), .B2(n9932), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9484) );
  NOR2_X1 U9998 ( .A1(n9450), .A2(n9449), .ZN(n9451) );
  NAND2_X1 U9999 ( .A1(n9461), .A2(n9460), .ZN(n9466) );
  OAI22_X1 U10000 ( .A1(n9275), .A2(n9253), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n12863), .ZN(n9265) );
  NAND2_X1 U10001 ( .A1(n10168), .A2(n6584), .ZN(n7034) );
  NAND2_X1 U10002 ( .A1(n7104), .A2(n7101), .ZN(n10166) );
  NAND3_X1 U10003 ( .A1(n7640), .A2(n12154), .A3(n8899), .ZN(n8900) );
  NAND2_X1 U10004 ( .A1(n7035), .A2(n10145), .ZN(n10149) );
  NAND2_X1 U10005 ( .A1(n10138), .A2(n10137), .ZN(n7035) );
  NAND2_X1 U10006 ( .A1(n7663), .A2(n7664), .ZN(n8945) );
  NAND2_X1 U10007 ( .A1(n7048), .A2(n7047), .ZN(n7806) );
  AND2_X1 U10008 ( .A1(n11416), .A2(n11415), .ZN(n10481) );
  NAND2_X1 U10009 ( .A1(n7614), .A2(n7613), .ZN(n14699) );
  NAND2_X1 U10010 ( .A1(n7470), .A2(n9495), .ZN(n7383) );
  NAND2_X1 U10011 ( .A1(n7383), .A2(n9497), .ZN(n9502) );
  NAND2_X1 U10012 ( .A1(n9742), .A2(n10201), .ZN(n15118) );
  NAND2_X1 U10013 ( .A1(n7327), .A2(n7325), .ZN(n8390) );
  NOR2_X1 U10014 ( .A1(n8003), .A2(n8002), .ZN(n8006) );
  NAND2_X1 U10015 ( .A1(n14376), .A2(n10077), .ZN(n14360) );
  AOI21_X1 U10016 ( .B1(n7905), .B2(P2_REG3_REG_1__SCAN_IN), .A(n7088), .ZN(
        n7906) );
  NAND2_X1 U10017 ( .A1(n11781), .A2(n10058), .ZN(n11996) );
  NAND2_X1 U10018 ( .A1(n8408), .A2(n8391), .ZN(n8393) );
  INV_X1 U10019 ( .A(n14628), .ZN(n7041) );
  OAI21_X1 U10020 ( .B1(n14660), .B2(n14343), .A(n7041), .ZN(P2_U3492) );
  INV_X1 U10021 ( .A(n14534), .ZN(n7042) );
  OAI21_X1 U10022 ( .B1(n7043), .B2(n14343), .A(n7042), .ZN(P2_U3524) );
  NAND2_X2 U10023 ( .A1(n7922), .A2(n7921), .ZN(n8001) );
  NAND2_X1 U10024 ( .A1(n7826), .A2(n7827), .ZN(n7922) );
  NAND3_X1 U10025 ( .A1(n7887), .A2(n7883), .A3(n7895), .ZN(n7820) );
  INV_X1 U10026 ( .A(n12770), .ZN(n7275) );
  OAI211_X1 U10027 ( .C1(n14281), .C2(n14280), .A(n7281), .B(n7278), .ZN(
        P2_U3233) );
  NAND2_X1 U10028 ( .A1(n7690), .A2(n7688), .ZN(n10409) );
  NAND2_X1 U10029 ( .A1(n7662), .A2(n8975), .ZN(n8987) );
  INV_X1 U10030 ( .A(n10239), .ZN(n7048) );
  INV_X1 U10031 ( .A(n8303), .ZN(n7067) );
  NAND3_X1 U10032 ( .A1(n15218), .A2(n15203), .A3(n12648), .ZN(n9707) );
  AND3_X2 U10033 ( .A1(n9505), .A2(n9504), .A3(n9503), .ZN(n11987) );
  NAND2_X1 U10034 ( .A1(n7944), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7050) );
  MUX2_X1 U10035 ( .A(n14969), .B(n14968), .S(n14967), .Z(n14971) );
  OAI21_X1 U10036 ( .B1(n12886), .B2(n15637), .A(n7052), .ZN(P3_U3488) );
  AOI22_X2 U10037 ( .A1(n7976), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10898), 
        .B2(n14144), .ZN(n7927) );
  AND2_X2 U10038 ( .A1(n10040), .A2(n7058), .ZN(n14396) );
  NOR2_X2 U10039 ( .A1(n14431), .A2(n14433), .ZN(n10040) );
  AND2_X2 U10040 ( .A1(n7118), .A2(n7117), .ZN(n12411) );
  NAND2_X1 U10041 ( .A1(n7069), .A2(n7068), .ZN(P2_U3528) );
  INV_X1 U10042 ( .A(n7112), .ZN(n7111) );
  NAND2_X1 U10043 ( .A1(n9802), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9826) );
  NAND2_X1 U10044 ( .A1(n7139), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U10045 ( .A1(n9757), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9768) );
  NAND2_X1 U10046 ( .A1(n7143), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9712) );
  NAND2_X1 U10047 ( .A1(n7233), .A2(n9409), .ZN(n9411) );
  INV_X1 U10048 ( .A(n12817), .ZN(n15020) );
  INV_X1 U10049 ( .A(n13350), .ZN(n7238) );
  NAND2_X1 U10050 ( .A1(n9401), .A2(n7238), .ZN(n7237) );
  NAND3_X1 U10051 ( .A1(n11082), .A2(n10049), .A3(n7794), .ZN(n7062) );
  NAND2_X1 U10052 ( .A1(n7684), .A2(n7683), .ZN(n14376) );
  NAND2_X1 U10053 ( .A1(n10113), .A2(n12855), .ZN(n14290) );
  INV_X1 U10054 ( .A(n11455), .ZN(n7364) );
  NAND2_X1 U10055 ( .A1(n9154), .A2(n12391), .ZN(n7349) );
  NAND2_X1 U10056 ( .A1(n11782), .A2(n14052), .ZN(n11781) );
  XNOR2_X1 U10057 ( .A(n10026), .B(n10025), .ZN(n14518) );
  NAND3_X1 U10059 ( .A1(n7820), .A2(n7819), .A3(n7886), .ZN(n7826) );
  NAND2_X1 U10060 ( .A1(n7598), .A2(n10792), .ZN(n7883) );
  OAI21_X1 U10061 ( .B1(n7944), .B2(n7075), .A(n7074), .ZN(n7817) );
  INV_X1 U10062 ( .A(n11573), .ZN(n7076) );
  NAND3_X1 U10063 ( .A1(n8376), .A2(n7796), .A3(n8375), .ZN(n13685) );
  NAND2_X1 U10064 ( .A1(n11074), .A2(n11075), .ZN(n11073) );
  NAND2_X1 U10065 ( .A1(n15018), .A2(n14997), .ZN(n14985) );
  NAND2_X1 U10066 ( .A1(n7395), .A2(n7394), .ZN(P1_U3557) );
  NAND3_X1 U10067 ( .A1(n7903), .A2(n7906), .A3(n7902), .ZN(n9965) );
  OAI22_X1 U10068 ( .A1(n9265), .A2(n9264), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n12897), .ZN(n9255) );
  XNOR2_X1 U10069 ( .A(n9309), .B(n9308), .ZN(n7080) );
  NAND2_X1 U10070 ( .A1(n9058), .A2(n7209), .ZN(n7208) );
  OAI21_X1 U10071 ( .B1(n7739), .B2(n6474), .A(n9051), .ZN(n7205) );
  NAND2_X1 U10072 ( .A1(n7204), .A2(n6474), .ZN(n7202) );
  NAND2_X1 U10073 ( .A1(n7738), .A2(n7204), .ZN(n7203) );
  NAND3_X1 U10074 ( .A1(n15107), .A2(n7082), .A3(n15086), .ZN(n10346) );
  NOR2_X1 U10075 ( .A1(n10345), .A2(n7083), .ZN(n7082) );
  NAND3_X1 U10076 ( .A1(n15138), .A2(n15123), .A3(n7084), .ZN(n7083) );
  NAND2_X1 U10077 ( .A1(n7808), .A2(n6582), .ZN(n7342) );
  OAI21_X1 U10078 ( .B1(n7944), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n7085), .ZN(
        n7815) );
  NAND3_X1 U10079 ( .A1(n10051), .A2(n10050), .A3(n10053), .ZN(n7681) );
  NAND2_X1 U10080 ( .A1(n7954), .A2(n7953), .ZN(n13806) );
  NAND2_X1 U10081 ( .A1(n8001), .A2(n7970), .ZN(n7943) );
  NAND3_X1 U10082 ( .A1(n7844), .A2(n6468), .A3(n7842), .ZN(n14667) );
  INV_X1 U10083 ( .A(n14290), .ZN(n14289) );
  INV_X1 U10084 ( .A(n14533), .ZN(n7122) );
  NAND2_X1 U10085 ( .A1(n7086), .A2(n14298), .ZN(P2_U3237) );
  OAI21_X1 U10086 ( .B1(n14290), .B2(n6471), .A(n14502), .ZN(n7086) );
  NAND2_X1 U10087 ( .A1(n10109), .A2(n10089), .ZN(n10097) );
  NAND2_X1 U10088 ( .A1(n7122), .A2(n6575), .ZN(n14627) );
  NOR2_X1 U10089 ( .A1(n10109), .A2(n10099), .ZN(n7092) );
  NAND2_X1 U10090 ( .A1(n10097), .A2(n10096), .ZN(n10100) );
  NAND2_X1 U10091 ( .A1(n7087), .A2(n11071), .ZN(n10047) );
  OAI21_X1 U10092 ( .B1(n10213), .B2(n10212), .A(n7809), .ZN(n10232) );
  NAND2_X1 U10093 ( .A1(n7207), .A2(n7208), .ZN(n9061) );
  NAND2_X1 U10094 ( .A1(n10156), .A2(n7551), .ZN(n7549) );
  NAND2_X1 U10095 ( .A1(n8864), .A2(n8847), .ZN(n8849) );
  NAND2_X1 U10096 ( .A1(n11339), .A2(n7500), .ZN(n11340) );
  NAND2_X1 U10097 ( .A1(n7099), .A2(n7098), .ZN(P2_U3496) );
  OAI21_X1 U10098 ( .B1(n14518), .B2(n15567), .A(n7093), .ZN(n7112) );
  NOR2_X1 U10099 ( .A1(n14515), .A2(n7094), .ZN(n7093) );
  OAI211_X1 U10100 ( .C1(n14517), .C2(n14473), .A(n10102), .B(n10101), .ZN(
        P2_U3236) );
  NOR2_X1 U10101 ( .A1(n7532), .A2(n7529), .ZN(n7528) );
  INV_X1 U10102 ( .A(n9472), .ZN(n7387) );
  NAND2_X1 U10103 ( .A1(n13277), .A2(n9056), .ZN(n7210) );
  NAND2_X1 U10104 ( .A1(n11083), .A2(n14043), .ZN(n11082) );
  NAND2_X1 U10105 ( .A1(n14624), .A2(n15572), .ZN(n7099) );
  NAND2_X2 U10106 ( .A1(n10904), .A2(n14683), .ZN(n7849) );
  NAND2_X1 U10107 ( .A1(n7103), .A2(n7102), .ZN(n7101) );
  INV_X1 U10108 ( .A(n10162), .ZN(n7103) );
  NAND2_X1 U10109 ( .A1(n10161), .A2(n10160), .ZN(n7104) );
  NAND3_X1 U10110 ( .A1(n10243), .A2(n7806), .A3(n6585), .ZN(n7105) );
  NAND3_X1 U10111 ( .A1(n7389), .A2(n7391), .A3(n9536), .ZN(n9498) );
  NAND2_X1 U10112 ( .A1(n12156), .A2(n7401), .ZN(n7400) );
  XNOR2_X2 U10113 ( .A(n7344), .B(n7501), .ZN(n9173) );
  NAND2_X1 U10114 ( .A1(n10413), .A2(n15572), .ZN(n10418) );
  NAND2_X1 U10115 ( .A1(n14289), .A2(n7108), .ZN(n10413) );
  NAND2_X1 U10116 ( .A1(n8900), .A2(n8899), .ZN(n8903) );
  NAND2_X1 U10117 ( .A1(n13245), .A2(n10400), .ZN(n7745) );
  INV_X1 U10118 ( .A(n14326), .ZN(n7110) );
  AOI21_X2 U10119 ( .B1(n15217), .B2(n9895), .A(n9894), .ZN(n15182) );
  NAND2_X1 U10120 ( .A1(n11281), .A2(n11280), .ZN(n11279) );
  NAND2_X1 U10121 ( .A1(n12870), .A2(n7485), .ZN(n7488) );
  NAND2_X1 U10122 ( .A1(n8862), .A2(n8861), .ZN(n8864) );
  NAND2_X1 U10123 ( .A1(n8899), .A2(n7640), .ZN(n8850) );
  NAND2_X1 U10124 ( .A1(n10080), .A2(n10079), .ZN(n14348) );
  AND3_X2 U10125 ( .A1(n7133), .A2(n7836), .A3(n7837), .ZN(n7844) );
  XNOR2_X1 U10126 ( .A(n7975), .B(n8003), .ZN(n10838) );
  OAI21_X1 U10127 ( .B1(SI_3_), .B2(n7823), .A(n7921), .ZN(n7825) );
  NOR2_X2 U10128 ( .A1(n8785), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7127) );
  NAND2_X1 U10129 ( .A1(n7746), .A2(n10399), .ZN(n13245) );
  INV_X1 U10130 ( .A(n10335), .ZN(n12119) );
  NAND2_X1 U10131 ( .A1(n8564), .A2(n8565), .ZN(n7130) );
  NAND2_X1 U10132 ( .A1(n8849), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8899) );
  NAND4_X1 U10133 ( .A1(n9467), .A2(n7132), .A3(n9468), .A4(n7131), .ZN(
        P3_U3296) );
  INV_X1 U10134 ( .A(n15086), .ZN(n7414) );
  NOR2_X1 U10135 ( .A1(n15261), .A2(n15260), .ZN(n15262) );
  OAI21_X2 U10136 ( .B1(n12211), .B2(n10270), .A(n9766), .ZN(n15099) );
  NAND2_X1 U10137 ( .A1(n9246), .A2(n9245), .ZN(n7357) );
  NAND3_X1 U10138 ( .A1(n15430), .A2(n7242), .A3(n15431), .ZN(n7240) );
  NAND2_X1 U10139 ( .A1(n7245), .A2(n7244), .ZN(n11777) );
  NAND2_X2 U10140 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7957) );
  NAND2_X1 U10141 ( .A1(n7512), .A2(n10362), .ZN(n7511) );
  OR4_X2 U10142 ( .A1(n14066), .A2(n14327), .A3(n14065), .A4(n14363), .ZN(
        n14067) );
  NOR2_X1 U10143 ( .A1(n14069), .A2(n10025), .ZN(n7138) );
  OAI21_X1 U10144 ( .B1(n15011), .B2(n15010), .A(n15009), .ZN(n15255) );
  NOR2_X1 U10145 ( .A1(n15256), .A2(n15507), .ZN(n15261) );
  NAND2_X1 U10146 ( .A1(n15263), .A2(n15262), .ZN(n15359) );
  NAND2_X1 U10147 ( .A1(n12055), .A2(n7150), .ZN(n7146) );
  NAND2_X1 U10148 ( .A1(n7146), .A2(n7147), .ZN(n12042) );
  NAND2_X1 U10149 ( .A1(n7159), .A2(n6588), .ZN(n7163) );
  NAND3_X1 U10150 ( .A1(n7693), .A2(n8592), .A3(n9328), .ZN(n7164) );
  NAND2_X4 U10151 ( .A1(n9168), .A2(n10801), .ZN(n9288) );
  NOR2_X1 U10152 ( .A1(n12585), .A2(n13095), .ZN(n7182) );
  NAND3_X1 U10153 ( .A1(n7186), .A2(n11313), .A3(n13496), .ZN(n11314) );
  INV_X2 U10154 ( .A(n9089), .ZN(n7188) );
  NAND2_X1 U10155 ( .A1(n12044), .A2(n7193), .ZN(n7191) );
  OAI21_X1 U10156 ( .B1(n12044), .B2(n7752), .A(n7193), .ZN(n12521) );
  NOR2_X1 U10157 ( .A1(n8905), .A2(n10791), .ZN(n7195) );
  NAND2_X1 U10158 ( .A1(n12034), .A2(n7199), .ZN(n7198) );
  NAND2_X1 U10159 ( .A1(n7198), .A2(n7196), .ZN(n9029) );
  NAND3_X1 U10160 ( .A1(n7203), .A2(n9412), .A3(n7202), .ZN(n9054) );
  NAND2_X1 U10161 ( .A1(n9058), .A2(n9057), .ZN(n7212) );
  AND2_X1 U10162 ( .A1(n7212), .A2(n9056), .ZN(n13278) );
  OAI21_X1 U10163 ( .B1(n6499), .B2(n7214), .A(n7213), .ZN(n9388) );
  NOR2_X1 U10164 ( .A1(n9377), .A2(n9393), .ZN(n7218) );
  AND2_X1 U10165 ( .A1(n13421), .A2(n9376), .ZN(n7219) );
  NAND2_X1 U10166 ( .A1(n7223), .A2(n7224), .ZN(n9373) );
  NAND3_X1 U10167 ( .A1(n9353), .A2(n7232), .A3(n7228), .ZN(n7223) );
  AOI21_X1 U10168 ( .B1(n15430), .B2(n15431), .A(n15429), .ZN(n15435) );
  NAND2_X1 U10169 ( .A1(n15407), .A2(n7246), .ZN(n7245) );
  INV_X1 U10170 ( .A(n13156), .ZN(n7251) );
  NAND2_X1 U10171 ( .A1(n7251), .A2(n7252), .ZN(n7250) );
  INV_X1 U10172 ( .A(n9228), .ZN(n7258) );
  NAND2_X1 U10173 ( .A1(n7261), .A2(n13140), .ZN(n7260) );
  XNOR2_X1 U10174 ( .A(n7262), .B(n9240), .ZN(n7261) );
  AND2_X1 U10175 ( .A1(n9234), .A2(n13211), .ZN(n7263) );
  NAND2_X1 U10176 ( .A1(n7286), .A2(n7851), .ZN(n7979) );
  NAND2_X1 U10177 ( .A1(n7286), .A2(n7284), .ZN(n7947) );
  INV_X1 U10178 ( .A(n7898), .ZN(n7286) );
  NAND2_X2 U10179 ( .A1(n7844), .A2(n7845), .ZN(n7861) );
  NAND2_X1 U10180 ( .A1(n13884), .A2(n6455), .ZN(n7288) );
  NAND2_X1 U10181 ( .A1(n7288), .A2(n6586), .ZN(n13927) );
  NAND2_X1 U10182 ( .A1(n7294), .A2(n7297), .ZN(n13865) );
  NAND2_X1 U10183 ( .A1(n7296), .A2(n7295), .ZN(n7294) );
  INV_X1 U10184 ( .A(n13980), .ZN(n7304) );
  INV_X1 U10185 ( .A(n13981), .ZN(n7305) );
  OAI21_X1 U10186 ( .B1(n13810), .B2(n7309), .A(n7308), .ZN(n13823) );
  NAND2_X1 U10187 ( .A1(n7306), .A2(n7307), .ZN(n13817) );
  NAND2_X1 U10188 ( .A1(n13810), .A2(n7308), .ZN(n7306) );
  NAND2_X1 U10189 ( .A1(n7310), .A2(n6576), .ZN(n13974) );
  NAND3_X1 U10190 ( .A1(n13965), .A2(n13964), .A3(n6590), .ZN(n7310) );
  AOI21_X1 U10191 ( .B1(n13833), .B2(n7313), .A(n7311), .ZN(n13851) );
  NAND3_X1 U10192 ( .A1(n8448), .A2(n8447), .A3(n6618), .ZN(n7321) );
  NAND2_X1 U10193 ( .A1(n7321), .A2(n7322), .ZN(n10261) );
  NAND3_X1 U10194 ( .A1(n8448), .A2(n6603), .A3(n8447), .ZN(n7323) );
  NAND2_X1 U10195 ( .A1(n8301), .A2(n7328), .ZN(n7327) );
  NAND2_X1 U10196 ( .A1(n14666), .A2(n10318), .ZN(n7334) );
  NAND2_X1 U10197 ( .A1(n7334), .A2(n7332), .ZN(n7331) );
  NAND2_X1 U10198 ( .A1(n7334), .A2(n10320), .ZN(n10395) );
  NAND2_X1 U10199 ( .A1(n7336), .A2(n7331), .ZN(n10329) );
  OAI21_X1 U10200 ( .B1(n14666), .B2(n7333), .A(n6619), .ZN(n7336) );
  OAI21_X1 U10201 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n7347), .A(n11889), .ZN(
        n11898) );
  NOR2_X1 U10202 ( .A1(n7348), .A2(n13111), .ZN(n12392) );
  OR2_X1 U10203 ( .A1(n13205), .A2(n7353), .ZN(n7351) );
  NAND2_X1 U10204 ( .A1(n9235), .A2(n9166), .ZN(n7355) );
  NAND2_X1 U10205 ( .A1(n7359), .A2(n10684), .ZN(n9158) );
  OR2_X1 U10206 ( .A1(n12317), .A2(n7370), .ZN(n7369) );
  NAND2_X1 U10207 ( .A1(n6451), .A2(n9480), .ZN(n7388) );
  NOR2_X1 U10208 ( .A1(n9937), .A2(n7390), .ZN(n7389) );
  NAND3_X1 U10209 ( .A1(n6451), .A2(n9480), .A3(n9496), .ZN(n7390) );
  INV_X1 U10210 ( .A(n7392), .ZN(n11108) );
  INV_X1 U10211 ( .A(n9648), .ZN(n7402) );
  NOR2_X1 U10212 ( .A1(n7396), .A2(n12317), .ZN(n7401) );
  AND2_X1 U10213 ( .A1(n9648), .A2(n7397), .ZN(n7396) );
  OAI21_X1 U10214 ( .B1(n12317), .B2(n9648), .A(n6593), .ZN(n7398) );
  XNOR2_X1 U10215 ( .A(n11167), .B(n7403), .ZN(n11168) );
  INV_X1 U10216 ( .A(n15043), .ZN(n7420) );
  NAND2_X1 U10217 ( .A1(n7425), .A2(n7427), .ZN(n14941) );
  OAI21_X1 U10218 ( .B1(n14938), .B2(n7428), .A(n14956), .ZN(n7427) );
  AND2_X1 U10219 ( .A1(n14939), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7428) );
  NAND2_X1 U10220 ( .A1(n14907), .A2(n6453), .ZN(n7440) );
  INV_X1 U10221 ( .A(n7445), .ZN(n11822) );
  NOR2_X1 U10222 ( .A1(n14910), .A2(n11614), .ZN(n7447) );
  NAND3_X1 U10223 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .A3(P1_IR_REG_0__SCAN_IN), .ZN(n7453) );
  NAND2_X1 U10224 ( .A1(n11111), .A2(n6845), .ZN(n11110) );
  AND2_X1 U10225 ( .A1(n12877), .A2(n7460), .ZN(n14984) );
  AOI21_X2 U10226 ( .B1(n10897), .B2(n9226), .A(n10693), .ZN(n9228) );
  AOI21_X1 U10227 ( .B1(n10931), .B2(P1_REG1_REG_3__SCAN_IN), .A(n10947), .ZN(
        n14866) );
  AOI21_X1 U10228 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10983), .A(n10979), .ZN(
        n10982) );
  NAND2_X1 U10229 ( .A1(n9860), .A2(n9906), .ZN(n15253) );
  NAND2_X1 U10230 ( .A1(n11275), .A2(n11274), .ZN(n11798) );
  NAND2_X1 U10231 ( .A1(n15076), .A2(n15075), .ZN(n15074) );
  NAND2_X1 U10232 ( .A1(n11279), .A2(n7465), .ZN(n7464) );
  AND2_X1 U10233 ( .A1(n9887), .A2(n7466), .ZN(n7465) );
  NAND2_X1 U10234 ( .A1(n9931), .A2(n7472), .ZN(n7469) );
  AND2_X1 U10235 ( .A1(n9931), .A2(n6597), .ZN(n7471) );
  NAND2_X1 U10236 ( .A1(n15184), .A2(n7476), .ZN(n7475) );
  NAND2_X1 U10237 ( .A1(n7488), .A2(n6587), .ZN(n15031) );
  NAND2_X1 U10238 ( .A1(n12870), .A2(n12869), .ZN(n15044) );
  NAND2_X1 U10239 ( .A1(n11308), .A2(n12906), .ZN(n7498) );
  NAND2_X1 U10240 ( .A1(n11312), .A2(n11309), .ZN(n7499) );
  INV_X1 U10241 ( .A(n10121), .ZN(n7518) );
  INV_X1 U10242 ( .A(n13220), .ZN(n7520) );
  NAND2_X1 U10243 ( .A1(n7535), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U10244 ( .A1(n7530), .A2(n7527), .ZN(n9185) );
  NAND2_X1 U10245 ( .A1(n11449), .A2(n11448), .ZN(n7530) );
  NOR2_X1 U10246 ( .A1(n11449), .A2(n7534), .ZN(n11385) );
  NAND2_X1 U10247 ( .A1(n9184), .A2(n11388), .ZN(n7535) );
  INV_X1 U10248 ( .A(n7538), .ZN(n7537) );
  NOR2_X1 U10249 ( .A1(n13160), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7539) );
  NOR2_X1 U10250 ( .A1(n10696), .A2(n13425), .ZN(n7545) );
  NAND3_X1 U10251 ( .A1(n10182), .A2(n10181), .A3(n6621), .ZN(n7547) );
  NAND3_X1 U10252 ( .A1(n10154), .A2(n10153), .A3(n7549), .ZN(n7548) );
  NAND3_X1 U10253 ( .A1(n7844), .A2(n7842), .A3(n7871), .ZN(n7756) );
  NAND2_X1 U10254 ( .A1(n7559), .A2(n14073), .ZN(n11047) );
  NAND2_X1 U10255 ( .A1(n13755), .A2(n7559), .ZN(n13760) );
  NAND3_X1 U10256 ( .A1(n13764), .A2(n13956), .A3(n7559), .ZN(n13765) );
  INV_X1 U10257 ( .A(n7559), .ZN(n7558) );
  NAND2_X1 U10258 ( .A1(n11196), .A2(n7998), .ZN(n7564) );
  AOI21_X1 U10259 ( .B1(n7563), .B2(n7562), .A(n6537), .ZN(n7561) );
  OAI21_X1 U10260 ( .B1(n11197), .B2(n11196), .A(n7998), .ZN(n11464) );
  NAND2_X1 U10261 ( .A1(n8271), .A2(n7567), .ZN(n7566) );
  NAND2_X1 U10262 ( .A1(n11721), .A2(n6452), .ZN(n7578) );
  AOI21_X1 U10263 ( .B1(n6452), .B2(n7585), .A(n6500), .ZN(n7579) );
  INV_X1 U10264 ( .A(n12470), .ZN(n7592) );
  INV_X1 U10265 ( .A(n7589), .ZN(n7587) );
  NAND2_X1 U10266 ( .A1(n7593), .A2(n14077), .ZN(P2_U3328) );
  OAI21_X1 U10267 ( .B1(n8196), .B2(n7600), .A(n7599), .ZN(n8244) );
  NAND3_X1 U10268 ( .A1(n7602), .A2(n13961), .A3(n7601), .ZN(n13965) );
  NAND3_X1 U10269 ( .A1(n13955), .A2(n13954), .A3(n13958), .ZN(n7602) );
  AOI21_X1 U10270 ( .B1(n13955), .B2(n13954), .A(n13953), .ZN(n13963) );
  NOR2_X1 U10271 ( .A1(n13979), .A2(n13978), .ZN(n13980) );
  NAND2_X1 U10272 ( .A1(n12098), .A2(n7072), .ZN(n7607) );
  XNOR2_X2 U10273 ( .A(n8274), .B(n8294), .ZN(n12098) );
  NAND2_X1 U10274 ( .A1(n7612), .A2(n10459), .ZN(n7611) );
  NAND2_X1 U10275 ( .A1(n10463), .A2(n11052), .ZN(n7612) );
  NAND2_X1 U10276 ( .A1(n10463), .A2(n11052), .ZN(n14716) );
  AND2_X1 U10277 ( .A1(n10459), .A2(n10464), .ZN(n14714) );
  NAND2_X1 U10278 ( .A1(n11361), .A2(n11362), .ZN(n11351) );
  NAND2_X1 U10279 ( .A1(n14769), .A2(n7615), .ZN(n7614) );
  NAND2_X1 U10280 ( .A1(n12349), .A2(n7619), .ZN(n12512) );
  INV_X1 U10281 ( .A(n7616), .ZN(n12511) );
  NOR2_X1 U10282 ( .A1(n12513), .A2(n7618), .ZN(n7617) );
  INV_X1 U10283 ( .A(n7619), .ZN(n7618) );
  NAND2_X1 U10284 ( .A1(n14731), .A2(n14732), .ZN(n7622) );
  INV_X2 U10285 ( .A(n10422), .ZN(n10419) );
  NAND2_X2 U10286 ( .A1(n10421), .A2(n10422), .ZN(n10439) );
  NAND2_X1 U10287 ( .A1(n9926), .A2(n6435), .ZN(n10422) );
  NAND2_X2 U10288 ( .A1(n7627), .A2(n9951), .ZN(n10421) );
  AOI21_X2 U10289 ( .B1(n9941), .B2(n9940), .A(n7626), .ZN(n9951) );
  NAND2_X1 U10290 ( .A1(n11526), .A2(n7638), .ZN(n7637) );
  NAND2_X1 U10291 ( .A1(n7635), .A2(n7634), .ZN(n7633) );
  NAND2_X1 U10292 ( .A1(n11526), .A2(n10493), .ZN(n11708) );
  INV_X1 U10293 ( .A(n7637), .ZN(n11707) );
  NOR2_X1 U10294 ( .A1(n11709), .A2(n10492), .ZN(n7638) );
  NAND2_X1 U10295 ( .A1(n8974), .A2(n8973), .ZN(n7662) );
  NAND3_X1 U10296 ( .A1(n7671), .A2(n12932), .A3(n9074), .ZN(n13257) );
  AND2_X1 U10297 ( .A1(n9063), .A2(n9418), .ZN(n7672) );
  INV_X1 U10298 ( .A(n7674), .ZN(n7673) );
  NAND2_X1 U10299 ( .A1(n12712), .A2(n14060), .ZN(n7679) );
  NAND2_X1 U10300 ( .A1(n7675), .A2(n7677), .ZN(n14459) );
  NOR2_X1 U10301 ( .A1(n14480), .A2(n9991), .ZN(n7676) );
  NAND3_X1 U10302 ( .A1(n9000), .A2(n9427), .A3(n9418), .ZN(n7690) );
  NAND3_X1 U10303 ( .A1(n8542), .A2(n7188), .A3(P3_IR_REG_27__SCAN_IN), .ZN(
        n7695) );
  NAND2_X1 U10304 ( .A1(n8774), .A2(n7702), .ZN(n7700) );
  NAND3_X1 U10305 ( .A1(n7711), .A2(n7709), .A3(n8917), .ZN(n7707) );
  NAND2_X1 U10306 ( .A1(n8898), .A2(n9389), .ZN(n7709) );
  NAND2_X1 U10307 ( .A1(n8898), .A2(n7710), .ZN(n7711) );
  NAND2_X1 U10308 ( .A1(n8681), .A2(n7717), .ZN(n7715) );
  NAND2_X1 U10309 ( .A1(n7715), .A2(n7716), .ZN(n8734) );
  XNOR2_X2 U10310 ( .A(n7722), .B(n7871), .ZN(n10904) );
  NAND2_X1 U10311 ( .A1(n7728), .A2(n14648), .ZN(n14431) );
  INV_X2 U10312 ( .A(n15563), .ZN(n7732) );
  NAND2_X1 U10313 ( .A1(n13378), .A2(n7742), .ZN(n7738) );
  XNOR2_X1 U10314 ( .A(n7745), .B(n10408), .ZN(n10407) );
  NAND2_X2 U10315 ( .A1(n8545), .A2(n8546), .ZN(n8577) );
  INV_X1 U10316 ( .A(n12044), .ZN(n7755) );
  NAND2_X1 U10317 ( .A1(n7755), .A2(n7754), .ZN(n7792) );
  NAND2_X1 U10318 ( .A1(n9022), .A2(n6577), .ZN(n12034) );
  NAND3_X1 U10319 ( .A1(n8542), .A2(n6592), .A3(n7188), .ZN(n13587) );
  NAND2_X1 U10320 ( .A1(n14050), .A2(n9981), .ZN(n7758) );
  INV_X1 U10321 ( .A(n12498), .ZN(n7775) );
  NAND2_X1 U10322 ( .A1(n7769), .A2(n7767), .ZN(n9997) );
  NAND2_X1 U10323 ( .A1(n12498), .A2(n6456), .ZN(n7769) );
  OR2_X1 U10324 ( .A1(n14733), .A2(n9519), .ZN(n9834) );
  AND2_X1 U10325 ( .A1(n11307), .A2(n9125), .ZN(n13397) );
  NAND2_X1 U10326 ( .A1(n10368), .A2(n15512), .ZN(n10373) );
  NAND2_X1 U10327 ( .A1(n10368), .A2(n15518), .ZN(n9961) );
  AND2_X1 U10328 ( .A1(n10904), .A2(n10899), .ZN(n13725) );
  NAND2_X1 U10329 ( .A1(n10261), .A2(n10260), .ZN(n10264) );
  OAI211_X1 U10330 ( .C1(n10110), .C2(n10103), .A(n10109), .B(n14481), .ZN(
        n10113) );
  NAND2_X1 U10331 ( .A1(n7969), .A2(n7971), .ZN(n7972) );
  NOR2_X1 U10332 ( .A1(n12864), .A2(n15032), .ZN(n15027) );
  NAND2_X1 U10333 ( .A1(n6551), .A2(n7972), .ZN(n8002) );
  NAND2_X1 U10334 ( .A1(n9185), .A2(n11891), .ZN(n10703) );
  INV_X4 U10335 ( .A(n9527), .ZN(n9915) );
  NOR2_X1 U10336 ( .A1(n9466), .A2(n9465), .ZN(n9467) );
  NAND2_X1 U10337 ( .A1(n9248), .A2(n7803), .ZN(n9251) );
  AOI21_X1 U10338 ( .B1(n10585), .B2(n14855), .A(n10453), .ZN(n10457) );
  INV_X1 U10339 ( .A(n15187), .ZN(n10420) );
  XNOR2_X1 U10340 ( .A(n9176), .B(n9142), .ZN(n11185) );
  XNOR2_X1 U10341 ( .A(n9176), .B(n9177), .ZN(n11189) );
  MUX2_X2 U10342 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14620), .S(n14618), .Z(
        n12840) );
  MUX2_X2 U10343 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14620), .S(n15572), .Z(
        n14621) );
  AND2_X1 U10344 ( .A1(n13613), .A2(n13715), .ZN(n13721) );
  OR2_X1 U10345 ( .A1(n9695), .A2(n7822), .ZN(n9539) );
  OR2_X1 U10346 ( .A1(n9695), .A2(n7075), .ZN(n9504) );
  INV_X1 U10347 ( .A(n8545), .ZN(n8547) );
  AND2_X1 U10348 ( .A1(n9972), .A2(n11572), .ZN(n9973) );
  OR2_X1 U10349 ( .A1(n14110), .A2(n7087), .ZN(n9966) );
  NAND2_X1 U10350 ( .A1(n9439), .A2(n9438), .ZN(n9468) );
  OR2_X1 U10351 ( .A1(n9288), .A2(n10784), .ZN(n8559) );
  NAND2_X1 U10352 ( .A1(n14678), .A2(n7072), .ZN(n10010) );
  NAND2_X1 U10353 ( .A1(n12709), .A2(n7072), .ZN(n8451) );
  INV_X1 U10354 ( .A(n6448), .ZN(n10374) );
  AND2_X1 U10355 ( .A1(n9241), .A2(n6983), .ZN(n13217) );
  CLKBUF_X1 U10356 ( .A(n14304), .Z(n14306) );
  INV_X1 U10357 ( .A(n12500), .ZN(n12718) );
  OR2_X1 U10358 ( .A1(n12853), .A2(n7091), .ZN(n8518) );
  OR2_X1 U10359 ( .A1(n14308), .A2(n7091), .ZN(n8459) );
  OR2_X1 U10360 ( .A1(n10018), .A2(n11440), .ZN(n7931) );
  OR2_X1 U10361 ( .A1(n10018), .A2(n10912), .ZN(n7913) );
  INV_X1 U10362 ( .A(n11579), .ZN(n10037) );
  AND2_X1 U10363 ( .A1(n10721), .A2(n12885), .ZN(n15192) );
  NAND2_X1 U10364 ( .A1(n12709), .A2(n10318), .ZN(n9839) );
  INV_X1 U10365 ( .A(n10318), .ZN(n10270) );
  INV_X1 U10366 ( .A(n14055), .ZN(n9986) );
  NAND2_X1 U10367 ( .A1(n15631), .A2(n15614), .ZN(n13580) );
  INV_X1 U10368 ( .A(n13580), .ZN(n9136) );
  NAND2_X1 U10369 ( .A1(n15639), .A2(n15614), .ZN(n13485) );
  AND2_X1 U10370 ( .A1(n14030), .A2(n14029), .ZN(n7788) );
  AND2_X1 U10371 ( .A1(n11427), .A2(n11630), .ZN(n7789) );
  NOR2_X1 U10372 ( .A1(n9040), .A2(n12780), .ZN(n7790) );
  AND2_X1 U10373 ( .A1(n10199), .A2(n10198), .ZN(n7791) );
  INV_X1 U10374 ( .A(n11961), .ZN(n9924) );
  INV_X1 U10375 ( .A(n14050), .ZN(n9980) );
  NOR4_X1 U10376 ( .A1(n14059), .A2(n14466), .A3(n14480), .A4(n14058), .ZN(
        n7793) );
  OR2_X1 U10377 ( .A1(n15253), .A2(n7800), .ZN(n7795) );
  NOR2_X1 U10378 ( .A1(n9592), .A2(n11920), .ZN(n7799) );
  OR2_X1 U10379 ( .A1(n15252), .A2(n15353), .ZN(n7800) );
  AND2_X1 U10380 ( .A1(n10657), .A2(n14801), .ZN(n7801) );
  AND2_X1 U10381 ( .A1(n15573), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U10382 ( .A1(n14686), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7803) );
  AND2_X1 U10383 ( .A1(n12883), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7804) );
  AND2_X1 U10384 ( .A1(n15579), .A2(n11818), .ZN(n15607) );
  AND2_X1 U10385 ( .A1(n9083), .A2(n8541), .ZN(n7805) );
  INV_X1 U10386 ( .A(n8003), .ZN(n8000) );
  INV_X1 U10387 ( .A(n14614), .ZN(n10036) );
  INV_X1 U10388 ( .A(n10395), .ZN(n15229) );
  AND2_X1 U10389 ( .A1(n10214), .A2(n10211), .ZN(n7809) );
  NOR3_X1 U10390 ( .A1(n14424), .A2(n14415), .A3(n14061), .ZN(n7810) );
  NAND2_X1 U10391 ( .A1(n15512), .A2(n15504), .ZN(n15389) );
  INV_X1 U10392 ( .A(n15389), .ZN(n10371) );
  INV_X1 U10393 ( .A(n10412), .ZN(n13240) );
  AND2_X1 U10394 ( .A1(n9961), .A2(n9960), .ZN(n7811) );
  OR2_X1 U10395 ( .A1(n13774), .A2(n13761), .ZN(n13773) );
  OR2_X1 U10396 ( .A1(n13778), .A2(n13777), .ZN(n13779) );
  OR2_X1 U10397 ( .A1(n13913), .A2(n13912), .ZN(n13917) );
  INV_X1 U10398 ( .A(n13956), .ZN(n13985) );
  INV_X1 U10399 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9142) );
  AND2_X1 U10400 ( .A1(n11430), .A2(n11370), .ZN(n10049) );
  INV_X1 U10401 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9177) );
  INV_X1 U10402 ( .A(n14060), .ZN(n9991) );
  NOR2_X1 U10403 ( .A1(n9176), .A2(n9177), .ZN(n9178) );
  AND2_X1 U10404 ( .A1(n9291), .A2(n9048), .ZN(n9049) );
  INV_X1 U10405 ( .A(n13887), .ZN(n10039) );
  INV_X1 U10406 ( .A(n14753), .ZN(n10559) );
  NAND2_X1 U10407 ( .A1(n15247), .A2(n15246), .ZN(n15248) );
  INV_X1 U10408 ( .A(n9498), .ZN(n9500) );
  INV_X1 U10409 ( .A(n9357), .ZN(n9032) );
  INV_X1 U10410 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8536) );
  OAI21_X1 U10411 ( .B1(n8373), .B2(n14087), .A(n13715), .ZN(n8370) );
  OR2_X1 U10412 ( .A1(n7935), .A2(n7934), .ZN(n7936) );
  NAND2_X1 U10413 ( .A1(n8452), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8510) );
  AND2_X1 U10414 ( .A1(n8181), .A2(n7829), .ZN(n7837) );
  OR2_X1 U10415 ( .A1(n15049), .A2(n14836), .ZN(n9810) );
  INV_X1 U10416 ( .A(n7106), .ZN(n9923) );
  INV_X1 U10417 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n15650) );
  NAND2_X1 U10418 ( .A1(n8189), .A2(SI_15_), .ZN(n8193) );
  AND2_X1 U10419 ( .A1(n15440), .A2(n15439), .ZN(n15449) );
  INV_X1 U10420 ( .A(n11564), .ZN(n11549) );
  INV_X1 U10421 ( .A(n13016), .ZN(n13019) );
  INV_X1 U10422 ( .A(n13084), .ZN(n8958) );
  INV_X1 U10423 ( .A(n12030), .ZN(n9023) );
  INV_X1 U10424 ( .A(n15607), .ZN(n9076) );
  AND3_X1 U10425 ( .A1(n13582), .A2(n13584), .A3(n9129), .ZN(n11327) );
  NAND2_X1 U10426 ( .A1(n10862), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8634) );
  AND2_X1 U10427 ( .A1(n14519), .A2(n15564), .ZN(n14520) );
  NOR2_X1 U10428 ( .A1(n8474), .A2(n7841), .ZN(n7842) );
  OR2_X1 U10429 ( .A1(n15187), .A2(n14967), .ZN(n10668) );
  INV_X1 U10430 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8693) );
  INV_X1 U10431 ( .A(n13082), .ZN(n12928) );
  INV_X1 U10432 ( .A(n8969), .ZN(n9278) );
  AND2_X1 U10433 ( .A1(n9355), .A2(n9354), .ZN(n12043) );
  NAND2_X1 U10434 ( .A1(n9326), .A2(n9023), .ZN(n8592) );
  AND2_X1 U10435 ( .A1(n9284), .A2(n9263), .ZN(n13230) );
  NOR2_X1 U10436 ( .A1(n9077), .A2(n9076), .ZN(n9078) );
  OR2_X1 U10437 ( .A1(n13579), .A2(n13094), .ZN(n9377) );
  INV_X2 U10438 ( .A(n8905), .ZN(n9287) );
  AND2_X1 U10439 ( .A1(n8700), .A2(n8684), .ZN(n8685) );
  AND2_X1 U10440 ( .A1(n11057), .A2(n7920), .ZN(n11075) );
  OR2_X1 U10441 ( .A1(n8523), .A2(n8522), .ZN(n13726) );
  INV_X1 U10442 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11982) );
  OR2_X1 U10443 ( .A1(n14038), .A2(n14404), .ZN(n14424) );
  NAND2_X1 U10444 ( .A1(n12006), .A2(n10038), .ZN(n12189) );
  OR2_X1 U10445 ( .A1(n8499), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8470) );
  INV_X1 U10446 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7851) );
  INV_X1 U10447 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7850) );
  INV_X1 U10448 ( .A(n10492), .ZN(n10493) );
  AND2_X1 U10449 ( .A1(n10665), .A2(n9943), .ZN(n10670) );
  OR2_X1 U10450 ( .A1(n15064), .A2(n9519), .ZN(n9798) );
  INV_X1 U10451 ( .A(n10939), .ZN(n10983) );
  AND2_X1 U10452 ( .A1(n10337), .A2(n9580), .ZN(n9581) );
  AND2_X1 U10453 ( .A1(n9879), .A2(n10449), .ZN(n11957) );
  OR2_X1 U10454 ( .A1(n15518), .A2(n9855), .ZN(n9960) );
  NAND2_X1 U10455 ( .A1(n11105), .A2(n11104), .ZN(n11767) );
  INV_X1 U10456 ( .A(n13066), .ZN(n13044) );
  NAND2_X1 U10457 ( .A1(n11544), .A2(n12227), .ZN(n13074) );
  INV_X1 U10458 ( .A(n12393), .ZN(n13112) );
  INV_X1 U10459 ( .A(n15575), .ZN(n13215) );
  NOR2_X1 U10460 ( .A1(n13360), .A2(n13366), .ZN(n13359) );
  INV_X1 U10461 ( .A(n13490), .ZN(n12309) );
  INV_X1 U10462 ( .A(n15578), .ZN(n15592) );
  NAND2_X1 U10463 ( .A1(n15614), .A2(n11329), .ZN(n15578) );
  INV_X1 U10464 ( .A(n13485), .ZN(n13471) );
  AND2_X1 U10465 ( .A1(n9370), .A2(n9371), .ZN(n12617) );
  NAND2_X1 U10466 ( .A1(n12825), .A2(n11818), .ZN(n15621) );
  NOR2_X1 U10467 ( .A1(n13583), .A2(n11298), .ZN(n11328) );
  INV_X1 U10468 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9001) );
  INV_X1 U10469 ( .A(n13726), .ZN(n13746) );
  OR2_X1 U10470 ( .A1(n10018), .A2(n15522), .ZN(n7891) );
  INV_X1 U10471 ( .A(n15529), .ZN(n15537) );
  NAND2_X1 U10472 ( .A1(n15558), .A2(n8506), .ZN(n14485) );
  INV_X1 U10473 ( .A(n14660), .ZN(n10388) );
  OAI21_X1 U10474 ( .B1(n10415), .B2(n14660), .A(n10414), .ZN(n10416) );
  AND2_X1 U10475 ( .A1(n10976), .A2(n8522), .ZN(n15564) );
  AND2_X1 U10476 ( .A1(n14426), .A2(n11698), .ZN(n15567) );
  AND2_X1 U10477 ( .A1(n15559), .A2(n10115), .ZN(n10386) );
  AND2_X1 U10478 ( .A1(n8482), .A2(n8481), .ZN(n15553) );
  NOR2_X1 U10479 ( .A1(n10667), .A2(n10666), .ZN(n14822) );
  INV_X1 U10480 ( .A(n15370), .ZN(n15078) );
  INV_X1 U10481 ( .A(n14824), .ZN(n14810) );
  OR2_X1 U10482 ( .A1(n10255), .A2(n9518), .ZN(n9524) );
  INV_X1 U10483 ( .A(n14960), .ZN(n14964) );
  OR2_X1 U10484 ( .A1(n9860), .A2(n9906), .ZN(n9861) );
  AND2_X1 U10485 ( .A1(n10721), .A2(n10844), .ZN(n15190) );
  AND2_X1 U10486 ( .A1(n15482), .A2(n11957), .ZN(n15224) );
  NAND2_X1 U10487 ( .A1(n10662), .A2(n15790), .ZN(n15208) );
  AOI21_X1 U10488 ( .B1(n10830), .B2(n10835), .A(n10832), .ZN(n11902) );
  INV_X1 U10489 ( .A(n15353), .ZN(n15494) );
  NOR2_X1 U10490 ( .A1(n11901), .A2(n9959), .ZN(n10367) );
  INV_X1 U10491 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9929) );
  AND2_X1 U10492 ( .A1(n15464), .A2(n15456), .ZN(n15458) );
  AND3_X1 U10493 ( .A1(n9104), .A2(n9103), .A3(n9102), .ZN(n11298) );
  INV_X1 U10494 ( .A(n13074), .ZN(n13011) );
  INV_X1 U10495 ( .A(n13063), .ZN(n13078) );
  AND2_X1 U10496 ( .A1(n9284), .A2(n9272), .ZN(n12348) );
  OAI211_X1 U10497 ( .C1(n8577), .C2(n13478), .A(n8810), .B(n8809), .ZN(n13093) );
  INV_X1 U10498 ( .A(n13217), .ZN(n13165) );
  OR2_X1 U10499 ( .A1(n15587), .A2(n12015), .ZN(n13431) );
  AND3_X2 U10500 ( .A1(n9121), .A2(n11854), .A3(n9120), .ZN(n15639) );
  NAND2_X1 U10501 ( .A1(n12934), .A2(n9136), .ZN(n9137) );
  INV_X1 U10502 ( .A(n15631), .ZN(n15629) );
  INV_X1 U10503 ( .A(n11851), .ZN(n13582) );
  INV_X1 U10504 ( .A(n13751), .ZN(n13738) );
  INV_X1 U10505 ( .A(n13896), .ZN(n14093) );
  AND2_X1 U10506 ( .A1(n10031), .A2(n14485), .ZN(n14490) );
  NAND2_X1 U10507 ( .A1(n14502), .A2(n10033), .ZN(n14497) );
  NOR2_X1 U10508 ( .A1(n10118), .A2(n7802), .ZN(n10119) );
  INV_X1 U10509 ( .A(n14618), .ZN(n15573) );
  INV_X1 U10510 ( .A(n10416), .ZN(n10417) );
  INV_X1 U10511 ( .A(n14450), .ZN(n14648) );
  INV_X1 U10512 ( .A(n15572), .ZN(n15570) );
  NOR2_X1 U10513 ( .A1(n15560), .A2(n15553), .ZN(n15554) );
  AND2_X1 U10514 ( .A1(n8526), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15558) );
  XNOR2_X1 U10515 ( .A(n8469), .B(n8468), .ZN(n12225) );
  INV_X1 U10516 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11509) );
  INV_X1 U10517 ( .A(n15307), .ZN(n15132) );
  INV_X1 U10518 ( .A(n10664), .ZN(n14808) );
  INV_X1 U10519 ( .A(n15012), .ZN(n14834) );
  OR2_X1 U10520 ( .A1(n10727), .A2(n10844), .ZN(n14959) );
  INV_X1 U10521 ( .A(n14965), .ZN(n14940) );
  INV_X1 U10522 ( .A(n15224), .ZN(n15478) );
  INV_X1 U10523 ( .A(n12215), .ZN(n15346) );
  INV_X1 U10524 ( .A(n15518), .ZN(n15516) );
  INV_X1 U10525 ( .A(n10333), .ZN(n15357) );
  INV_X1 U10526 ( .A(n15213), .ZN(n15386) );
  INV_X1 U10527 ( .A(n15512), .ZN(n15510) );
  AND2_X2 U10528 ( .A1(n10367), .A2(n10366), .ZN(n15512) );
  NAND2_X1 U10529 ( .A1(n10831), .A2(n15790), .ZN(n15487) );
  INV_X1 U10530 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11744) );
  INV_X1 U10531 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11092) );
  AND2_X1 U10532 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10901), .ZN(P2_U3947) );
  NAND2_X1 U10533 ( .A1(n10120), .A2(n10119), .ZN(P2_U3527) );
  NAND2_X1 U10534 ( .A1(n10418), .A2(n10417), .ZN(P2_U3495) );
  AND2_X1 U10535 ( .A1(n10683), .A2(n10833), .ZN(P1_U4016) );
  NAND2_X1 U10536 ( .A1(n7811), .A2(n9964), .ZN(P1_U3556) );
  NAND2_X1 U10537 ( .A1(n10373), .A2(n10372), .ZN(P1_U3524) );
  INV_X1 U10538 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7813) );
  INV_X1 U10539 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7812) );
  INV_X1 U10540 ( .A(SI_2_), .ZN(n7814) );
  INV_X1 U10541 ( .A(SI_1_), .ZN(n10792) );
  INV_X1 U10542 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U10543 ( .A1(n7816), .A2(SI_2_), .ZN(n7886) );
  INV_X1 U10544 ( .A(n7884), .ZN(n7818) );
  NAND2_X1 U10545 ( .A1(n7818), .A2(n7887), .ZN(n7819) );
  INV_X1 U10546 ( .A(n7826), .ZN(n7824) );
  NAND2_X1 U10547 ( .A1(n7823), .A2(SI_3_), .ZN(n7921) );
  NAND2_X1 U10548 ( .A1(n7824), .A2(n7825), .ZN(n7828) );
  INV_X1 U10549 ( .A(n7825), .ZN(n7827) );
  AND2_X1 U10550 ( .A1(n7922), .A2(n7828), .ZN(n10823) );
  NOR2_X1 U10551 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7829) );
  INV_X2 U10552 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7948) );
  NAND4_X1 U10553 ( .A1(n7948), .A2(n7832), .A3(n7831), .A4(n7830), .ZN(n7980)
         );
  NAND3_X1 U10554 ( .A1(n7835), .A2(n7834), .A3(n7833), .ZN(n8250) );
  NOR2_X1 U10555 ( .A1(n7980), .A2(n8250), .ZN(n7836) );
  NOR2_X2 U10556 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n7863) );
  NOR2_X1 U10557 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n7839) );
  NOR2_X1 U10558 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n7838) );
  NAND3_X1 U10559 ( .A1(n7863), .A2(n7839), .A3(n7838), .ZN(n8474) );
  NAND3_X1 U10560 ( .A1(n7840), .A2(n8477), .A3(n7845), .ZN(n7841) );
  NAND2_X1 U10561 ( .A1(n8477), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7843) );
  NOR2_X1 U10562 ( .A1(n8474), .A2(n7843), .ZN(n7848) );
  INV_X1 U10563 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7860) );
  XNOR2_X1 U10564 ( .A(n7860), .B(P2_IR_REG_27__SCAN_IN), .ZN(n7847) );
  AND2_X1 U10565 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n7846) );
  NAND2_X1 U10566 ( .A1(n10823), .A2(n6448), .ZN(n7855) );
  NAND2_X1 U10567 ( .A1(n7979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7852) );
  INV_X1 U10568 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10569 ( .A1(n7861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7858) );
  OAI21_X1 U10570 ( .B1(P2_IR_REG_21__SCAN_IN), .B2(P2_IR_REG_20__SCAN_IN), 
        .A(P2_IR_REG_22__SCAN_IN), .ZN(n7859) );
  AND2_X1 U10571 ( .A1(n7859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7868) );
  AND2_X1 U10572 ( .A1(n7860), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U10573 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  AND2_X1 U10574 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n7865) );
  NAND2_X1 U10575 ( .A1(n7861), .A2(n7865), .ZN(n7866) );
  INV_X1 U10576 ( .A(n13757), .ZN(n14076) );
  XNOR2_X1 U10577 ( .A(n14033), .B(n14076), .ZN(n7870) );
  INV_X1 U10578 ( .A(n7844), .ZN(n8254) );
  NAND2_X1 U10579 ( .A1(n8254), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U10580 ( .A1(n7870), .A2(n14031), .ZN(n10032) );
  NAND2_X1 U10581 ( .A1(n10032), .A2(n14033), .ZN(n7901) );
  INV_X1 U10582 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14668) );
  NAND2_X1 U10583 ( .A1(n7929), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7880) );
  OR2_X1 U10584 ( .A1(n7091), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7879) );
  INV_X1 U10585 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10995) );
  OR2_X1 U10586 ( .A1(n10380), .A2(n10995), .ZN(n7878) );
  INV_X1 U10587 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11374) );
  INV_X1 U10588 ( .A(n12014), .ZN(n14041) );
  OR2_X2 U10589 ( .A1(n8504), .A2(n14041), .ZN(n7907) );
  AND2_X1 U10590 ( .A1(n14108), .A2(n14486), .ZN(n7938) );
  NAND2_X1 U10591 ( .A1(n7898), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7881) );
  MUX2_X1 U10592 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7881), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n7882) );
  INV_X1 U10593 ( .A(n15523), .ZN(n11008) );
  NAND2_X1 U10594 ( .A1(n7884), .A2(n7883), .ZN(n7896) );
  INV_X1 U10595 ( .A(n7895), .ZN(n7885) );
  OAI21_X1 U10596 ( .B1(n7896), .B2(n7885), .A(n7884), .ZN(n7889) );
  NAND2_X1 U10597 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  XNOR2_X1 U10598 ( .A(n7889), .B(n7888), .ZN(n10819) );
  NAND2_X1 U10599 ( .A1(n10819), .A2(n6448), .ZN(n7890) );
  XNOR2_X1 U10600 ( .A(n13774), .B(n7987), .ZN(n7919) );
  NAND2_X1 U10601 ( .A1(n7929), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7894) );
  INV_X1 U10602 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10994) );
  OR2_X1 U10603 ( .A1(n10380), .A2(n10994), .ZN(n7893) );
  INV_X1 U10604 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11648) );
  OR2_X1 U10605 ( .A1(n7910), .A2(n11648), .ZN(n7892) );
  INV_X1 U10606 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n15522) );
  NAND2_X1 U10607 ( .A1(n14109), .A2(n7907), .ZN(n7918) );
  NAND2_X1 U10608 ( .A1(n7919), .A2(n7918), .ZN(n11057) );
  XNOR2_X1 U10609 ( .A(n7895), .B(n7896), .ZN(n10802) );
  NAND2_X1 U10610 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7897) );
  MUX2_X1 U10611 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7897), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7899) );
  NAND2_X1 U10612 ( .A1(n7899), .A2(n7898), .ZN(n14113) );
  OR2_X1 U10613 ( .A1(n7849), .A2(n14113), .ZN(n7900) );
  XNOR2_X1 U10614 ( .A(n7901), .B(n10034), .ZN(n7909) );
  NAND2_X1 U10615 ( .A1(n7929), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7902) );
  INV_X1 U10616 ( .A(n10018), .ZN(n7905) );
  NAND2_X1 U10617 ( .A1(n14110), .A2(n7907), .ZN(n7908) );
  NAND2_X1 U10618 ( .A1(n7909), .A2(n7908), .ZN(n7917) );
  NAND2_X1 U10619 ( .A1(n7929), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7914) );
  INV_X1 U10620 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10912) );
  INV_X1 U10621 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10907) );
  OR2_X1 U10622 ( .A1(n10380), .A2(n10907), .ZN(n7912) );
  INV_X1 U10623 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10908) );
  NAND2_X1 U10624 ( .A1(n10801), .A2(SI_0_), .ZN(n7915) );
  XNOR2_X1 U10625 ( .A(n7915), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14687) );
  OR2_X1 U10626 ( .A1(n7987), .A2(n13763), .ZN(n7916) );
  NAND2_X1 U10627 ( .A1(n11043), .A2(n7917), .ZN(n11074) );
  OR2_X1 U10628 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  INV_X1 U10629 ( .A(n8001), .ZN(n7924) );
  MUX2_X1 U10630 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7944), .Z(n7923) );
  NAND2_X1 U10631 ( .A1(n7924), .A2(n7925), .ZN(n7926) );
  INV_X1 U10632 ( .A(n7925), .ZN(n7970) );
  AND2_X1 U10633 ( .A1(n7926), .A2(n7943), .ZN(n10795) );
  NAND2_X1 U10634 ( .A1(n10795), .A2(n6448), .ZN(n7928) );
  INV_X4 U10635 ( .A(n7987), .ZN(n8412) );
  XNOR2_X1 U10636 ( .A(n13791), .B(n8412), .ZN(n7935) );
  NAND2_X1 U10637 ( .A1(n7929), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7933) );
  INV_X1 U10638 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11436) );
  OR2_X1 U10639 ( .A1(n7910), .A2(n11436), .ZN(n7932) );
  OAI21_X1 U10640 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7957), .ZN(n11440) );
  INV_X1 U10641 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10996) );
  OR2_X1 U10642 ( .A1(n10380), .A2(n10996), .ZN(n7930) );
  NAND2_X1 U10643 ( .A1(n14107), .A2(n14486), .ZN(n7934) );
  NAND2_X1 U10644 ( .A1(n7935), .A2(n7934), .ZN(n7942) );
  INV_X1 U10645 ( .A(n7937), .ZN(n7939) );
  AND2_X1 U10646 ( .A1(n7939), .A2(n7938), .ZN(n13691) );
  NAND2_X1 U10647 ( .A1(n7941), .A2(n7940), .ZN(n13695) );
  NAND2_X1 U10648 ( .A1(n10840), .A2(n6448), .ZN(n7954) );
  INV_X1 U10649 ( .A(n7947), .ZN(n7949) );
  NAND2_X1 U10650 ( .A1(n7949), .A2(n7948), .ZN(n7951) );
  NAND2_X1 U10651 ( .A1(n7951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7950) );
  MUX2_X1 U10652 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7950), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n7952) );
  AOI22_X1 U10653 ( .A1(n7976), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10898), 
        .B2(n14159), .ZN(n7953) );
  XNOR2_X1 U10654 ( .A(n13806), .B(n8412), .ZN(n7963) );
  NAND2_X1 U10655 ( .A1(n10379), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7962) );
  INV_X1 U10656 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11640) );
  OR2_X1 U10657 ( .A1(n7910), .A2(n11640), .ZN(n7961) );
  INV_X1 U10658 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U10659 ( .A1(n7957), .A2(n7956), .ZN(n7958) );
  NAND2_X1 U10660 ( .A1(n7990), .A2(n7958), .ZN(n13667) );
  OR2_X1 U10661 ( .A1(n10018), .A2(n13667), .ZN(n7960) );
  INV_X1 U10662 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10997) );
  OR2_X1 U10663 ( .A1(n10380), .A2(n10997), .ZN(n7959) );
  OR2_X1 U10664 ( .A1(n13808), .A2(n14469), .ZN(n7964) );
  NAND2_X1 U10665 ( .A1(n7963), .A2(n7964), .ZN(n7968) );
  INV_X1 U10666 ( .A(n7963), .ZN(n7966) );
  INV_X1 U10667 ( .A(n7964), .ZN(n7965) );
  NAND2_X1 U10668 ( .A1(n7966), .A2(n7965), .ZN(n7967) );
  AND2_X1 U10669 ( .A1(n7968), .A2(n7967), .ZN(n13665) );
  NAND2_X1 U10670 ( .A1(n8001), .A2(n7999), .ZN(n7973) );
  NAND2_X1 U10671 ( .A1(n7974), .A2(SI_6_), .ZN(n8004) );
  NAND2_X1 U10672 ( .A1(n10838), .A2(n6448), .ZN(n7986) );
  NAND2_X1 U10673 ( .A1(n7977), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7978) );
  MUX2_X1 U10674 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7978), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n7984) );
  INV_X1 U10675 ( .A(n7979), .ZN(n7983) );
  INV_X1 U10676 ( .A(n7981), .ZN(n7982) );
  NAND2_X1 U10677 ( .A1(n7983), .A2(n7982), .ZN(n8010) );
  NAND2_X1 U10678 ( .A1(n7984), .A2(n8010), .ZN(n14172) );
  INV_X1 U10679 ( .A(n14172), .ZN(n11016) );
  AOI22_X1 U10680 ( .A1(n7976), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10898), 
        .B2(n11016), .ZN(n7985) );
  XNOR2_X1 U10681 ( .A(n13813), .B(n12847), .ZN(n7997) );
  NAND2_X1 U10682 ( .A1(n10379), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7995) );
  INV_X1 U10683 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11660) );
  OR2_X1 U10684 ( .A1(n7910), .A2(n11660), .ZN(n7994) );
  INV_X1 U10685 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U10686 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  NAND2_X1 U10687 ( .A1(n8017), .A2(n7991), .ZN(n11662) );
  OR2_X1 U10688 ( .A1(n7091), .A2(n11662), .ZN(n7993) );
  INV_X1 U10689 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10998) );
  OR2_X1 U10690 ( .A1(n10380), .A2(n10998), .ZN(n7992) );
  NOR2_X1 U10691 ( .A1(n13815), .A2(n14469), .ZN(n7996) );
  XNOR2_X1 U10692 ( .A(n7997), .B(n7996), .ZN(n11196) );
  NAND2_X1 U10693 ( .A1(n7997), .A2(n7996), .ZN(n7998) );
  INV_X1 U10694 ( .A(n8004), .ZN(n8005) );
  NAND2_X1 U10695 ( .A1(n10851), .A2(n6448), .ZN(n8013) );
  NAND2_X1 U10696 ( .A1(n8010), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8009) );
  MUX2_X1 U10697 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8009), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n8011) );
  AND2_X1 U10698 ( .A1(n8011), .A2(n8033), .ZN(n11018) );
  AOI22_X1 U10699 ( .A1(n7976), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10898), 
        .B2(n11018), .ZN(n8012) );
  XNOR2_X1 U10700 ( .A(n14614), .B(n8412), .ZN(n8023) );
  NAND2_X1 U10701 ( .A1(n7904), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8022) );
  INV_X1 U10702 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8014) );
  OR2_X1 U10703 ( .A1(n8311), .A2(n8014), .ZN(n8021) );
  INV_X1 U10704 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U10705 ( .A1(n8017), .A2(n8016), .ZN(n8018) );
  NAND2_X1 U10706 ( .A1(n8039), .A2(n8018), .ZN(n11540) );
  OR2_X1 U10707 ( .A1(n7091), .A2(n11540), .ZN(n8020) );
  INV_X1 U10708 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10999) );
  OR2_X1 U10709 ( .A1(n10380), .A2(n10999), .ZN(n8019) );
  NOR2_X1 U10710 ( .A1(n13820), .A2(n14469), .ZN(n8024) );
  XNOR2_X1 U10711 ( .A(n8023), .B(n8024), .ZN(n11465) );
  INV_X1 U10712 ( .A(n8023), .ZN(n8025) );
  INV_X1 U10713 ( .A(n8026), .ZN(n8027) );
  NAND2_X1 U10714 ( .A1(n10870), .A2(n6448), .ZN(n8037) );
  NAND2_X1 U10715 ( .A1(n8033), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8031) );
  MUX2_X1 U10716 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8031), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8035) );
  INV_X1 U10717 ( .A(n8033), .ZN(n8034) );
  NAND2_X1 U10718 ( .A1(n8035), .A2(n8251), .ZN(n14187) );
  INV_X1 U10719 ( .A(n14187), .ZN(n11022) );
  AOI22_X1 U10720 ( .A1(n7976), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10898), 
        .B2(n11022), .ZN(n8036) );
  XNOR2_X1 U10721 ( .A(n13840), .B(n8412), .ZN(n8045) );
  NAND2_X1 U10722 ( .A1(n10379), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8044) );
  INV_X1 U10723 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11000) );
  OR2_X1 U10724 ( .A1(n10380), .A2(n11000), .ZN(n8043) );
  NAND2_X1 U10725 ( .A1(n8039), .A2(n8038), .ZN(n8040) );
  NAND2_X1 U10726 ( .A1(n8064), .A2(n8040), .ZN(n11727) );
  OR2_X1 U10727 ( .A1(n7091), .A2(n11727), .ZN(n8042) );
  INV_X1 U10728 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11019) );
  OR2_X1 U10729 ( .A1(n7910), .A2(n11019), .ZN(n8041) );
  NAND4_X1 U10730 ( .A1(n8044), .A2(n8043), .A3(n8042), .A4(n8041), .ZN(n14103) );
  NAND2_X1 U10731 ( .A1(n14103), .A2(n14486), .ZN(n8046) );
  NAND2_X1 U10732 ( .A1(n8045), .A2(n8046), .ZN(n8051) );
  INV_X1 U10733 ( .A(n8045), .ZN(n8048) );
  INV_X1 U10734 ( .A(n8046), .ZN(n8047) );
  NAND2_X1 U10735 ( .A1(n8048), .A2(n8047), .ZN(n8049) );
  NAND2_X1 U10736 ( .A1(n8051), .A2(n8049), .ZN(n11723) );
  INV_X1 U10737 ( .A(n11723), .ZN(n8050) );
  NAND2_X1 U10738 ( .A1(n8251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8058) );
  XNOR2_X1 U10739 ( .A(n8058), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U10740 ( .A1(n7976), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10898), 
        .B2(n11396), .ZN(n8059) );
  NAND2_X1 U10741 ( .A1(n7904), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8069) );
  INV_X1 U10742 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8061) );
  OR2_X1 U10743 ( .A1(n8311), .A2(n8061), .ZN(n8068) );
  INV_X1 U10744 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U10745 ( .A1(n8064), .A2(n8063), .ZN(n8065) );
  NAND2_X1 U10746 ( .A1(n8078), .A2(n8065), .ZN(n11842) );
  OR2_X1 U10747 ( .A1(n7091), .A2(n11842), .ZN(n8067) );
  INV_X1 U10748 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11405) );
  OR2_X1 U10749 ( .A1(n10380), .A2(n11405), .ZN(n8066) );
  OR2_X1 U10750 ( .A1(n13837), .A2(n14469), .ZN(n8070) );
  MUX2_X1 U10751 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10801), .Z(n8074) );
  XNOR2_X1 U10752 ( .A(n8088), .B(n8086), .ZN(n10916) );
  NAND2_X1 U10753 ( .A1(n10916), .A2(n7072), .ZN(n8077) );
  NAND2_X1 U10754 ( .A1(n8091), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8075) );
  XNOR2_X1 U10755 ( .A(n8075), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U10756 ( .A1(n7976), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n11407), 
        .B2(n10898), .ZN(n8076) );
  XNOR2_X1 U10757 ( .A(n14604), .B(n12847), .ZN(n8085) );
  NAND2_X1 U10758 ( .A1(n8512), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8083) );
  INV_X1 U10759 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11399) );
  OR2_X1 U10760 ( .A1(n7040), .A2(n11399), .ZN(n8082) );
  INV_X1 U10761 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15657) );
  OR2_X1 U10762 ( .A1(n8311), .A2(n15657), .ZN(n8081) );
  NAND2_X1 U10763 ( .A1(n8078), .A2(n11982), .ZN(n8079) );
  NAND2_X1 U10764 ( .A1(n8097), .A2(n8079), .ZN(n12004) );
  OR2_X1 U10765 ( .A1(n7091), .A2(n12004), .ZN(n8080) );
  NOR2_X1 U10766 ( .A1(n13848), .A2(n14469), .ZN(n8084) );
  XNOR2_X1 U10767 ( .A(n8085), .B(n8084), .ZN(n11979) );
  INV_X1 U10768 ( .A(n8086), .ZN(n8087) );
  MUX2_X1 U10769 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10801), .Z(n8110) );
  NAND2_X1 U10770 ( .A1(n10943), .A2(n7072), .ZN(n8094) );
  NAND2_X1 U10771 ( .A1(n8112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8092) );
  XNOR2_X1 U10772 ( .A(n8092), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U10773 ( .A1(n11589), .A2(n10898), .B1(n7976), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8093) );
  XNOR2_X1 U10774 ( .A(n13860), .B(n12847), .ZN(n8105) );
  NAND2_X1 U10775 ( .A1(n7904), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8102) );
  INV_X1 U10776 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8095) );
  OR2_X1 U10777 ( .A1(n8311), .A2(n8095), .ZN(n8101) );
  INV_X1 U10778 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10779 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  NAND2_X1 U10780 ( .A1(n8121), .A2(n8098), .ZN(n12252) );
  OR2_X1 U10781 ( .A1(n7091), .A2(n12252), .ZN(n8100) );
  INV_X1 U10782 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11583) );
  OR2_X1 U10783 ( .A1(n10380), .A2(n11583), .ZN(n8099) );
  NAND4_X1 U10784 ( .A1(n8102), .A2(n8101), .A3(n8100), .A4(n8099), .ZN(n14099) );
  NAND2_X1 U10785 ( .A1(n14099), .A2(n14486), .ZN(n8103) );
  XNOR2_X1 U10786 ( .A(n8105), .B(n8103), .ZN(n12247) );
  INV_X1 U10787 ( .A(n8103), .ZN(n8104) );
  AND2_X1 U10788 ( .A1(n8105), .A2(n8104), .ZN(n8106) );
  INV_X1 U10789 ( .A(n8110), .ZN(n8111) );
  INV_X1 U10790 ( .A(SI_11_), .ZN(n10825) );
  MUX2_X1 U10791 ( .A(n11065), .B(n11066), .S(n10801), .Z(n8154) );
  XNOR2_X1 U10792 ( .A(n8154), .B(SI_12_), .ZN(n8133) );
  XNOR2_X1 U10793 ( .A(n8134), .B(n8133), .ZN(n11064) );
  NAND2_X1 U10794 ( .A1(n11064), .A2(n7072), .ZN(n8120) );
  NAND2_X1 U10795 ( .A1(n8114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8113) );
  MUX2_X1 U10796 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8113), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8117) );
  INV_X1 U10797 ( .A(n8114), .ZN(n8116) );
  NAND2_X1 U10798 ( .A1(n8116), .A2(n8115), .ZN(n8160) );
  NAND2_X1 U10799 ( .A1(n8117), .A2(n8160), .ZN(n12261) );
  INV_X1 U10800 ( .A(n8118), .ZN(n8119) );
  XNOR2_X1 U10801 ( .A(n14599), .B(n8412), .ZN(n8127) );
  NAND2_X1 U10802 ( .A1(n10379), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8126) );
  INV_X1 U10803 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n12262) );
  OR2_X1 U10804 ( .A1(n10380), .A2(n12262), .ZN(n8125) );
  NAND2_X1 U10805 ( .A1(n8121), .A2(n11587), .ZN(n8122) );
  NAND2_X1 U10806 ( .A1(n8141), .A2(n8122), .ZN(n12426) );
  OR2_X1 U10807 ( .A1(n7091), .A2(n12426), .ZN(n8124) );
  INV_X1 U10808 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12298) );
  OR2_X1 U10809 ( .A1(n7040), .A2(n12298), .ZN(n8123) );
  NAND4_X1 U10810 ( .A1(n8126), .A2(n8125), .A3(n8124), .A4(n8123), .ZN(n14098) );
  NAND2_X1 U10811 ( .A1(n14098), .A2(n14486), .ZN(n8128) );
  NAND2_X1 U10812 ( .A1(n8127), .A2(n8128), .ZN(n8132) );
  INV_X1 U10813 ( .A(n8127), .ZN(n8130) );
  INV_X1 U10814 ( .A(n8128), .ZN(n8129) );
  NAND2_X1 U10815 ( .A1(n8130), .A2(n8129), .ZN(n8131) );
  AND2_X1 U10816 ( .A1(n8132), .A2(n8131), .ZN(n12424) );
  NAND2_X1 U10817 ( .A1(n12422), .A2(n12424), .ZN(n12423) );
  NAND2_X1 U10818 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  INV_X1 U10819 ( .A(SI_12_), .ZN(n10868) );
  NAND2_X1 U10820 ( .A1(n8154), .A2(n10868), .ZN(n8152) );
  NAND2_X1 U10821 ( .A1(n8135), .A2(n8152), .ZN(n8136) );
  MUX2_X1 U10822 ( .A(n11092), .B(n11090), .S(n10801), .Z(n8158) );
  XNOR2_X1 U10823 ( .A(n8136), .B(n8156), .ZN(n11089) );
  NAND2_X1 U10824 ( .A1(n11089), .A2(n7072), .ZN(n8139) );
  NAND2_X1 U10825 ( .A1(n8160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8137) );
  XNOR2_X1 U10826 ( .A(n8137), .B(P2_IR_REG_13__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U10827 ( .A1(n12263), .A2(n10898), .B1(n7976), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n8138) );
  XNOR2_X1 U10828 ( .A(n14594), .B(n8412), .ZN(n8147) );
  INV_X1 U10829 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U10830 ( .A1(n8141), .A2(n8140), .ZN(n8142) );
  NAND2_X1 U10831 ( .A1(n8165), .A2(n8142), .ZN(n12472) );
  NAND2_X1 U10832 ( .A1(n8512), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8143) );
  OAI21_X1 U10833 ( .B1(n12472), .B2(n7091), .A(n8143), .ZN(n8146) );
  INV_X1 U10834 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U10835 ( .A1(n7929), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8144) );
  OAI21_X1 U10836 ( .B1(n7040), .B2(n12258), .A(n8144), .ZN(n8145) );
  NAND2_X1 U10837 ( .A1(n14097), .A2(n7907), .ZN(n8148) );
  XNOR2_X1 U10838 ( .A(n8147), .B(n8148), .ZN(n12471) );
  INV_X1 U10839 ( .A(n8147), .ZN(n8150) );
  INV_X1 U10840 ( .A(n8148), .ZN(n8149) );
  NAND2_X1 U10841 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  INV_X1 U10842 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U10843 ( .A1(n8155), .A2(SI_12_), .ZN(n8157) );
  INV_X1 U10844 ( .A(SI_13_), .ZN(n10892) );
  NAND2_X1 U10845 ( .A1(n8158), .A2(n10892), .ZN(n8159) );
  MUX2_X1 U10846 ( .A(n15740), .B(n11349), .S(n10801), .Z(n8188) );
  XNOR2_X1 U10847 ( .A(n8176), .B(n8188), .ZN(n11348) );
  NAND2_X1 U10848 ( .A1(n11348), .A2(n7072), .ZN(n8163) );
  OAI21_X1 U10849 ( .B1(n8160), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8161) );
  XNOR2_X1 U10850 ( .A(n8161), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U10851 ( .A1(n12764), .A2(n10898), .B1(n7976), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n8162) );
  XNOR2_X1 U10852 ( .A(n13880), .B(n8412), .ZN(n8169) );
  INV_X1 U10853 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12772) );
  INV_X1 U10854 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10855 ( .A1(n8165), .A2(n8164), .ZN(n8166) );
  NAND2_X1 U10856 ( .A1(n8209), .A2(n8166), .ZN(n12740) );
  OR2_X1 U10857 ( .A1(n12740), .A2(n7091), .ZN(n8168) );
  AOI22_X1 U10858 ( .A1(n7904), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n10379), 
        .B2(P2_REG0_REG_14__SCAN_IN), .ZN(n8167) );
  OAI211_X1 U10859 ( .C1(n10380), .C2(n12772), .A(n8168), .B(n8167), .ZN(
        n14096) );
  NAND2_X1 U10860 ( .A1(n14096), .A2(n7907), .ZN(n8170) );
  NAND2_X1 U10861 ( .A1(n8169), .A2(n8170), .ZN(n8175) );
  INV_X1 U10862 ( .A(n8169), .ZN(n8172) );
  INV_X1 U10863 ( .A(n8170), .ZN(n8171) );
  NAND2_X1 U10864 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  NAND2_X1 U10865 ( .A1(n8175), .A2(n8173), .ZN(n12736) );
  INV_X1 U10866 ( .A(n12736), .ZN(n8174) );
  NAND2_X1 U10867 ( .A1(n8176), .A2(n8188), .ZN(n8178) );
  INV_X1 U10868 ( .A(SI_14_), .ZN(n10896) );
  NAND2_X1 U10869 ( .A1(n8187), .A2(n10896), .ZN(n8177) );
  MUX2_X1 U10870 ( .A(n15732), .B(n11517), .S(n10801), .Z(n8192) );
  XNOR2_X1 U10871 ( .A(n8192), .B(SI_15_), .ZN(n8179) );
  NAND2_X1 U10872 ( .A1(n11516), .A2(n7072), .ZN(n8186) );
  NAND2_X1 U10873 ( .A1(n6607), .A2(n8181), .ZN(n8249) );
  OR2_X1 U10874 ( .A1(n8251), .A2(n8249), .ZN(n8183) );
  NAND2_X1 U10875 ( .A1(n8183), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8182) );
  MUX2_X1 U10876 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8182), .S(
        P2_IR_REG_15__SCAN_IN), .Z(n8184) );
  AND2_X1 U10877 ( .A1(n8184), .A2(n8198), .ZN(n14228) );
  AOI22_X1 U10878 ( .A1(n7976), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n14228), 
        .B2(n10898), .ZN(n8185) );
  XNOR2_X1 U10879 ( .A(n13887), .B(n8412), .ZN(n13650) );
  NAND2_X1 U10880 ( .A1(n8191), .A2(SI_14_), .ZN(n8190) );
  INV_X1 U10881 ( .A(n8192), .ZN(n8189) );
  NOR2_X1 U10882 ( .A1(n8191), .A2(SI_14_), .ZN(n8194) );
  INV_X1 U10883 ( .A(SI_15_), .ZN(n10894) );
  MUX2_X1 U10884 ( .A(n11336), .B(n11337), .S(n10801), .Z(n8224) );
  XNOR2_X1 U10885 ( .A(n8222), .B(n8221), .ZN(n11335) );
  NAND2_X1 U10886 ( .A1(n11335), .A2(n7072), .ZN(n8202) );
  NAND2_X1 U10887 ( .A1(n8198), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8197) );
  MUX2_X1 U10888 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8197), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8199) );
  OR2_X1 U10889 ( .A1(n8198), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U10890 ( .A1(n8199), .A2(n8225), .ZN(n14237) );
  INV_X1 U10891 ( .A(n8200), .ZN(n8201) );
  XNOR2_X1 U10892 ( .A(n14655), .B(n8412), .ZN(n8214) );
  XNOR2_X1 U10893 ( .A(n8230), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n13656) );
  NAND2_X1 U10894 ( .A1(n13656), .A2(n7905), .ZN(n8208) );
  INV_X1 U10895 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14226) );
  NAND2_X1 U10896 ( .A1(n7929), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8205) );
  NAND2_X1 U10897 ( .A1(n8512), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8204) );
  OAI211_X1 U10898 ( .C1(n7040), .C2(n14226), .A(n8205), .B(n8204), .ZN(n8206)
         );
  INV_X1 U10899 ( .A(n8206), .ZN(n8207) );
  NAND2_X1 U10900 ( .A1(n8208), .A2(n8207), .ZN(n14094) );
  NAND2_X1 U10901 ( .A1(n14094), .A2(n7907), .ZN(n8215) );
  NAND2_X1 U10902 ( .A1(n8214), .A2(n8215), .ZN(n13653) );
  INV_X1 U10903 ( .A(n13653), .ZN(n8213) );
  INV_X1 U10904 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14590) );
  INV_X1 U10905 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12768) );
  NAND2_X1 U10906 ( .A1(n8209), .A2(n12768), .ZN(n8210) );
  NAND2_X1 U10907 ( .A1(n8230), .A2(n8210), .ZN(n13749) );
  OR2_X1 U10908 ( .A1(n13749), .A2(n7091), .ZN(n8212) );
  AOI22_X1 U10909 ( .A1(n7904), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n10379), 
        .B2(P2_REG0_REG_15__SCAN_IN), .ZN(n8211) );
  OAI211_X1 U10910 ( .C1(n10380), .C2(n14590), .A(n8212), .B(n8211), .ZN(
        n14095) );
  AND2_X1 U10911 ( .A1(n14095), .A2(n14486), .ZN(n13743) );
  NAND2_X1 U10912 ( .A1(n13653), .A2(n13743), .ZN(n8218) );
  OAI21_X1 U10913 ( .B1(n13650), .B2(n8213), .A(n8218), .ZN(n8220) );
  INV_X1 U10914 ( .A(n8214), .ZN(n8217) );
  INV_X1 U10915 ( .A(n8215), .ZN(n8216) );
  NAND2_X1 U10916 ( .A1(n8217), .A2(n8216), .ZN(n13652) );
  OAI21_X1 U10917 ( .B1(n13650), .B2(n8218), .A(n13652), .ZN(n8219) );
  INV_X1 U10918 ( .A(SI_16_), .ZN(n8223) );
  MUX2_X1 U10919 ( .A(n11510), .B(n11509), .S(n10801), .Z(n8245) );
  XNOR2_X1 U10920 ( .A(n8244), .B(n8243), .ZN(n11508) );
  NAND2_X1 U10921 ( .A1(n11508), .A2(n7072), .ZN(n13899) );
  NAND2_X1 U10922 ( .A1(n8225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8226) );
  XNOR2_X1 U10923 ( .A(n8226), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14261) );
  AOI21_X1 U10924 ( .B1(n14261), .B2(n10898), .A(n8227), .ZN(n13893) );
  XNOR2_X1 U10925 ( .A(n14651), .B(n8412), .ZN(n8237) );
  INV_X1 U10926 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13658) );
  INV_X1 U10927 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8228) );
  OAI21_X1 U10928 ( .B1(n8230), .B2(n13658), .A(n8228), .ZN(n8231) );
  NAND2_X1 U10929 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n8229) );
  AND2_X1 U10930 ( .A1(n8231), .A2(n8258), .ZN(n14472) );
  NAND2_X1 U10931 ( .A1(n14472), .A2(n7905), .ZN(n8236) );
  INV_X1 U10932 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14244) );
  NAND2_X1 U10933 ( .A1(n8512), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U10934 ( .A1(n10379), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8232) );
  OAI211_X1 U10935 ( .C1(n7040), .C2(n14244), .A(n8233), .B(n8232), .ZN(n8234)
         );
  INV_X1 U10936 ( .A(n8234), .ZN(n8235) );
  NAND2_X1 U10937 ( .A1(n14093), .A2(n7907), .ZN(n8238) );
  NAND2_X1 U10938 ( .A1(n8237), .A2(n8238), .ZN(n8242) );
  INV_X1 U10939 ( .A(n8237), .ZN(n8240) );
  INV_X1 U10940 ( .A(n8238), .ZN(n8239) );
  NAND2_X1 U10941 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  AND2_X1 U10942 ( .A1(n8242), .A2(n8241), .ZN(n13674) );
  INV_X1 U10943 ( .A(SI_17_), .ZN(n11042) );
  NAND2_X1 U10944 ( .A1(n8245), .A2(n11042), .ZN(n8246) );
  INV_X1 U10945 ( .A(SI_18_), .ZN(n11069) );
  NAND2_X1 U10946 ( .A1(n8297), .A2(n11069), .ZN(n8247) );
  MUX2_X1 U10947 ( .A(n11744), .B(n11743), .S(n10801), .Z(n8292) );
  OR3_X1 U10948 ( .A1(n8251), .A2(n8250), .A3(n8249), .ZN(n8252) );
  NAND2_X1 U10949 ( .A1(n8252), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8253) );
  MUX2_X1 U10950 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8253), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n8255) );
  AND2_X1 U10951 ( .A1(n8255), .A2(n8254), .ZN(n14255) );
  AOI22_X1 U10952 ( .A1(n7976), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n14255), 
        .B2(n10898), .ZN(n8256) );
  XNOR2_X1 U10953 ( .A(n14450), .B(n8412), .ZN(n8266) );
  INV_X1 U10954 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n14263) );
  NAND2_X1 U10955 ( .A1(n8258), .A2(n14263), .ZN(n8259) );
  NAND2_X1 U10956 ( .A1(n8277), .A2(n8259), .ZN(n14451) );
  OR2_X1 U10957 ( .A1(n14451), .A2(n7091), .ZN(n8265) );
  INV_X1 U10958 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U10959 ( .A1(n8512), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U10960 ( .A1(n10379), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8260) );
  OAI211_X1 U10961 ( .C1(n7040), .C2(n8262), .A(n8261), .B(n8260), .ZN(n8263)
         );
  INV_X1 U10962 ( .A(n8263), .ZN(n8264) );
  NAND2_X1 U10963 ( .A1(n8265), .A2(n8264), .ZN(n14092) );
  NAND2_X1 U10964 ( .A1(n14092), .A2(n7907), .ZN(n8267) );
  XNOR2_X1 U10965 ( .A(n8266), .B(n8267), .ZN(n13724) );
  INV_X1 U10966 ( .A(n13724), .ZN(n8270) );
  INV_X1 U10967 ( .A(n8266), .ZN(n8269) );
  INV_X1 U10968 ( .A(n8267), .ZN(n8268) );
  NAND2_X1 U10969 ( .A1(n8273), .A2(n8272), .ZN(n8274) );
  MUX2_X1 U10970 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10801), .Z(n8298) );
  XNOR2_X1 U10971 ( .A(n8298), .B(SI_19_), .ZN(n8294) );
  AOI22_X1 U10972 ( .A1(n7976), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10898), 
        .B2(n14280), .ZN(n8275) );
  INV_X1 U10973 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U10974 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  AND2_X1 U10975 ( .A1(n8307), .A2(n8278), .ZN(n14434) );
  NAND2_X1 U10976 ( .A1(n14434), .A2(n7905), .ZN(n8284) );
  INV_X1 U10977 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U10978 ( .A1(n8512), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U10979 ( .A1(n10379), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8279) );
  OAI211_X1 U10980 ( .C1(n7040), .C2(n8281), .A(n8280), .B(n8279), .ZN(n8282)
         );
  INV_X1 U10981 ( .A(n8282), .ZN(n8283) );
  NAND2_X1 U10982 ( .A1(n8284), .A2(n8283), .ZN(n14091) );
  NAND2_X1 U10983 ( .A1(n14091), .A2(n7907), .ZN(n8286) );
  NAND2_X1 U10984 ( .A1(n8285), .A2(n8286), .ZN(n8290) );
  INV_X1 U10985 ( .A(n8285), .ZN(n8288) );
  INV_X1 U10986 ( .A(n8286), .ZN(n8287) );
  NAND2_X1 U10987 ( .A1(n8288), .A2(n8287), .ZN(n8289) );
  INV_X1 U10988 ( .A(n8292), .ZN(n8291) );
  NOR2_X1 U10989 ( .A1(n8292), .A2(n11069), .ZN(n8293) );
  INV_X1 U10990 ( .A(n8298), .ZN(n8299) );
  INV_X1 U10991 ( .A(SI_19_), .ZN(n11177) );
  NAND2_X1 U10992 ( .A1(n8299), .A2(n11177), .ZN(n8300) );
  INV_X1 U10993 ( .A(SI_20_), .ZN(n11524) );
  NAND2_X1 U10994 ( .A1(n8384), .A2(n11524), .ZN(n8302) );
  INV_X1 U10995 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12154) );
  INV_X1 U10996 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12013) );
  MUX2_X1 U10997 ( .A(n12154), .B(n12013), .S(n10801), .Z(n8322) );
  NAND2_X1 U10998 ( .A1(n8303), .A2(n8322), .ZN(n8304) );
  XNOR2_X1 U10999 ( .A(n14557), .B(n8412), .ZN(n8315) );
  INV_X1 U11000 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n15695) );
  NAND2_X1 U11001 ( .A1(n8307), .A2(n15695), .ZN(n8308) );
  NAND2_X1 U11002 ( .A1(n8330), .A2(n8308), .ZN(n14410) );
  OR2_X1 U11003 ( .A1(n14410), .A2(n7091), .ZN(n8314) );
  INV_X1 U11004 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n15641) );
  NAND2_X1 U11005 ( .A1(n7904), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U11006 ( .A1(n8512), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8309) );
  OAI211_X1 U11007 ( .C1(n8311), .C2(n15641), .A(n8310), .B(n8309), .ZN(n8312)
         );
  INV_X1 U11008 ( .A(n8312), .ZN(n8313) );
  NAND2_X1 U11009 ( .A1(n8314), .A2(n8313), .ZN(n14090) );
  NAND2_X1 U11010 ( .A1(n14090), .A2(n7907), .ZN(n8316) );
  INV_X1 U11011 ( .A(n8315), .ZN(n8318) );
  INV_X1 U11012 ( .A(n8316), .ZN(n8317) );
  NAND2_X1 U11013 ( .A1(n8318), .A2(n8317), .ZN(n13706) );
  AND2_X1 U11014 ( .A1(n8319), .A2(n8325), .ZN(n8320) );
  NAND2_X1 U11015 ( .A1(n8321), .A2(n8320), .ZN(n8327) );
  NAND2_X1 U11016 ( .A1(n8323), .A2(SI_20_), .ZN(n8377) );
  NAND2_X1 U11017 ( .A1(n8384), .A2(n8377), .ZN(n8326) );
  NAND2_X1 U11018 ( .A1(n8327), .A2(n8342), .ZN(n12211) );
  INV_X1 U11019 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12210) );
  XNOR2_X1 U11020 ( .A(n14638), .B(n12847), .ZN(n8340) );
  INV_X1 U11021 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13637) );
  NAND2_X1 U11022 ( .A1(n8330), .A2(n13637), .ZN(n8331) );
  AND2_X1 U11023 ( .A1(n8361), .A2(n8331), .ZN(n14399) );
  NAND2_X1 U11024 ( .A1(n14399), .A2(n7905), .ZN(n8337) );
  INV_X1 U11025 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U11026 ( .A1(n10379), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U11027 ( .A1(n8512), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8332) );
  OAI211_X1 U11028 ( .C1(n8334), .C2(n7040), .A(n8333), .B(n8332), .ZN(n8335)
         );
  INV_X1 U11029 ( .A(n8335), .ZN(n8336) );
  NAND2_X1 U11030 ( .A1(n8337), .A2(n8336), .ZN(n14089) );
  NAND2_X1 U11031 ( .A1(n14089), .A2(n7907), .ZN(n8338) );
  XNOR2_X1 U11032 ( .A(n8340), .B(n8338), .ZN(n13635) );
  INV_X1 U11033 ( .A(n8338), .ZN(n8339) );
  NAND2_X1 U11034 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  INV_X1 U11035 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8343) );
  MUX2_X1 U11036 ( .A(n8343), .B(n12220), .S(n10801), .Z(n8386) );
  NAND2_X1 U11037 ( .A1(n9777), .A2(n8386), .ZN(n8344) );
  NAND2_X1 U11038 ( .A1(n8348), .A2(n8344), .ZN(n12221) );
  XNOR2_X1 U11039 ( .A(n14634), .B(n12847), .ZN(n8372) );
  MUX2_X1 U11040 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10801), .Z(n8349) );
  NAND2_X1 U11041 ( .A1(n8349), .A2(SI_23_), .ZN(n8389) );
  NAND2_X1 U11042 ( .A1(n12398), .A2(n7072), .ZN(n8352) );
  INV_X1 U11043 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12401) );
  XNOR2_X1 U11044 ( .A(n14541), .B(n12847), .ZN(n8373) );
  INV_X1 U11045 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13622) );
  NAND2_X1 U11046 ( .A1(n8363), .A2(n13622), .ZN(n8353) );
  AND2_X1 U11047 ( .A1(n8397), .A2(n8353), .ZN(n14367) );
  NAND2_X1 U11048 ( .A1(n14367), .A2(n7905), .ZN(n8359) );
  INV_X1 U11049 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8356) );
  NAND2_X1 U11050 ( .A1(n8512), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U11051 ( .A1(n10379), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8354) );
  OAI211_X1 U11052 ( .C1(n7040), .C2(n8356), .A(n8355), .B(n8354), .ZN(n8357)
         );
  INV_X1 U11053 ( .A(n8357), .ZN(n8358) );
  INV_X1 U11054 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U11055 ( .A1(n8361), .A2(n8360), .ZN(n8362) );
  NAND2_X1 U11056 ( .A1(n8363), .A2(n8362), .ZN(n14384) );
  OR2_X1 U11057 ( .A1(n14384), .A2(n7091), .ZN(n8369) );
  INV_X1 U11058 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U11059 ( .A1(n10379), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U11060 ( .A1(n8512), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8364) );
  OAI211_X1 U11061 ( .C1(n7040), .C2(n8366), .A(n8365), .B(n8364), .ZN(n8367)
         );
  INV_X1 U11062 ( .A(n8367), .ZN(n8368) );
  NOR2_X1 U11063 ( .A1(n13960), .A2(n14469), .ZN(n13715) );
  INV_X1 U11064 ( .A(n8370), .ZN(n8371) );
  NAND2_X1 U11065 ( .A1(n13613), .A2(n8371), .ZN(n8376) );
  AND2_X1 U11066 ( .A1(n14087), .A2(n14486), .ZN(n8374) );
  OAI21_X1 U11067 ( .B1(n8374), .B2(n8373), .A(n13614), .ZN(n8375) );
  INV_X1 U11068 ( .A(n8373), .ZN(n13615) );
  INV_X1 U11069 ( .A(n8374), .ZN(n13619) );
  INV_X1 U11070 ( .A(n8381), .ZN(n8383) );
  INV_X1 U11071 ( .A(n8377), .ZN(n8380) );
  INV_X1 U11072 ( .A(SI_22_), .ZN(n8919) );
  OAI21_X1 U11073 ( .B1(n8386), .B2(n8919), .A(n8378), .ZN(n8379) );
  AOI21_X1 U11074 ( .B1(n8381), .B2(n8380), .A(n8379), .ZN(n8382) );
  INV_X1 U11075 ( .A(n8385), .ZN(n8388) );
  NAND2_X1 U11076 ( .A1(n8386), .A2(n8919), .ZN(n8387) );
  INV_X1 U11077 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15734) );
  INV_X1 U11078 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12223) );
  MUX2_X1 U11079 ( .A(n15734), .B(n12223), .S(n10801), .Z(n8392) );
  NAND2_X1 U11080 ( .A1(n8393), .A2(n8392), .ZN(n8394) );
  XNOR2_X1 U11081 ( .A(n14536), .B(n8412), .ZN(n8405) );
  INV_X1 U11082 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13686) );
  NAND2_X1 U11083 ( .A1(n8397), .A2(n13686), .ZN(n8398) );
  NAND2_X1 U11084 ( .A1(n8432), .A2(n8398), .ZN(n14353) );
  INV_X1 U11085 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14352) );
  NAND2_X1 U11086 ( .A1(n8512), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U11087 ( .A1(n10379), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8399) );
  OAI211_X1 U11088 ( .C1(n7040), .C2(n14352), .A(n8400), .B(n8399), .ZN(n8401)
         );
  INV_X1 U11089 ( .A(n8401), .ZN(n8402) );
  NAND2_X1 U11090 ( .A1(n14086), .A2(n7907), .ZN(n8404) );
  NOR2_X1 U11091 ( .A1(n8405), .A2(n8404), .ZN(n8406) );
  AOI21_X1 U11092 ( .B1(n8405), .B2(n8404), .A(n8406), .ZN(n13684) );
  INV_X1 U11093 ( .A(n8406), .ZN(n8407) );
  MUX2_X1 U11094 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10801), .Z(n8425) );
  XNOR2_X1 U11095 ( .A(n8425), .B(SI_25_), .ZN(n8423) );
  XNOR2_X1 U11096 ( .A(n8424), .B(n8423), .ZN(n12478) );
  NAND2_X1 U11097 ( .A1(n12478), .A2(n7072), .ZN(n8411) );
  INV_X1 U11098 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12483) );
  XNOR2_X1 U11099 ( .A(n14629), .B(n8412), .ZN(n8420) );
  XNOR2_X1 U11100 ( .A(n8432), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14340) );
  NAND2_X1 U11101 ( .A1(n14340), .A2(n7905), .ZN(n8418) );
  INV_X1 U11102 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U11103 ( .A1(n8512), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U11104 ( .A1(n10379), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8413) );
  OAI211_X1 U11105 ( .C1(n7040), .C2(n8415), .A(n8414), .B(n8413), .ZN(n8416)
         );
  INV_X1 U11106 ( .A(n8416), .ZN(n8417) );
  NAND2_X1 U11107 ( .A1(n14085), .A2(n7907), .ZN(n8419) );
  NOR2_X1 U11108 ( .A1(n8420), .A2(n8419), .ZN(n8421) );
  AOI21_X1 U11109 ( .B1(n8420), .B2(n8419), .A(n8421), .ZN(n13643) );
  INV_X1 U11110 ( .A(n8421), .ZN(n8422) );
  INV_X1 U11111 ( .A(n8425), .ZN(n8426) );
  INV_X1 U11112 ( .A(SI_25_), .ZN(n13608) );
  NAND2_X1 U11113 ( .A1(n8426), .A2(n13608), .ZN(n8427) );
  INV_X1 U11114 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12672) );
  INV_X1 U11115 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12670) );
  MUX2_X1 U11116 ( .A(n12672), .B(n12670), .S(n10801), .Z(n8442) );
  XNOR2_X1 U11117 ( .A(n8442), .B(SI_26_), .ZN(n8428) );
  NAND2_X1 U11118 ( .A1(n12669), .A2(n7072), .ZN(n8430) );
  XNOR2_X1 U11119 ( .A(n14325), .B(n12847), .ZN(n8441) );
  INV_X1 U11120 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8431) );
  INV_X1 U11121 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13736) );
  OAI21_X1 U11122 ( .B1(n8432), .B2(n8431), .A(n13736), .ZN(n8433) );
  NAND2_X1 U11123 ( .A1(n14323), .A2(n7905), .ZN(n8439) );
  INV_X1 U11124 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U11125 ( .A1(n8512), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U11126 ( .A1(n10379), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8434) );
  OAI211_X1 U11127 ( .C1(n7040), .C2(n8436), .A(n8435), .B(n8434), .ZN(n8437)
         );
  INV_X1 U11128 ( .A(n8437), .ZN(n8438) );
  NAND2_X1 U11129 ( .A1(n14084), .A2(n14486), .ZN(n8440) );
  XNOR2_X1 U11130 ( .A(n8441), .B(n8440), .ZN(n13731) );
  INV_X1 U11131 ( .A(SI_26_), .ZN(n13604) );
  INV_X1 U11132 ( .A(n8442), .ZN(n8443) );
  INV_X1 U11133 ( .A(n8445), .ZN(n8446) );
  MUX2_X1 U11134 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10801), .Z(n9848) );
  XNOR2_X1 U11135 ( .A(n9848), .B(SI_27_), .ZN(n8449) );
  INV_X1 U11136 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14686) );
  XNOR2_X1 U11137 ( .A(n14519), .B(n12847), .ZN(n8461) );
  INV_X1 U11138 ( .A(n8461), .ZN(n8463) );
  INV_X1 U11139 ( .A(n8453), .ZN(n8452) );
  INV_X1 U11140 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U11141 ( .A1(n8453), .A2(n8529), .ZN(n8454) );
  NAND2_X1 U11142 ( .A1(n8510), .A2(n8454), .ZN(n14308) );
  INV_X1 U11143 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n14307) );
  NAND2_X1 U11144 ( .A1(n8512), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U11145 ( .A1(n10379), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8455) );
  OAI211_X1 U11146 ( .C1(n7040), .C2(n14307), .A(n8456), .B(n8455), .ZN(n8457)
         );
  INV_X1 U11147 ( .A(n8457), .ZN(n8458) );
  NOR2_X1 U11148 ( .A1(n13735), .A2(n14469), .ZN(n8460) );
  INV_X1 U11149 ( .A(n8460), .ZN(n8462) );
  AOI21_X1 U11150 ( .B1(n8463), .B2(n8462), .A(n12851), .ZN(n8465) );
  INV_X1 U11151 ( .A(n8464), .ZN(n8467) );
  INV_X1 U11152 ( .A(n8465), .ZN(n8466) );
  NAND2_X1 U11153 ( .A1(n8467), .A2(n8466), .ZN(n8503) );
  NAND2_X1 U11154 ( .A1(n8470), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8469) );
  INV_X1 U11155 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8468) );
  XNOR2_X1 U11156 ( .A(n12225), .B(P2_B_REG_SCAN_IN), .ZN(n8473) );
  OAI21_X1 U11157 ( .B1(n8470), .B2(P2_IR_REG_24__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8472) );
  INV_X1 U11158 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8471) );
  XNOR2_X1 U11159 ( .A(n8472), .B(n8471), .ZN(n12481) );
  NAND2_X1 U11160 ( .A1(n8473), .A2(n12481), .ZN(n8482) );
  OR2_X1 U11161 ( .A1(n7861), .A2(n8474), .ZN(n8476) );
  NAND2_X1 U11162 ( .A1(n8476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8475) );
  MUX2_X1 U11163 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8475), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8480) );
  INV_X1 U11164 ( .A(n8476), .ZN(n8478) );
  NAND2_X1 U11165 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  INV_X1 U11166 ( .A(n12671), .ZN(n8481) );
  NOR4_X1 U11167 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8486) );
  NOR4_X1 U11168 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8485) );
  NOR4_X1 U11169 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8484) );
  NOR4_X1 U11170 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8483) );
  AND4_X1 U11171 ( .A1(n8486), .A2(n8485), .A3(n8484), .A4(n8483), .ZN(n8492)
         );
  NOR2_X1 U11172 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .ZN(
        n8490) );
  NOR4_X1 U11173 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8489) );
  NOR4_X1 U11174 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n8488) );
  NOR4_X1 U11175 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8487) );
  AND4_X1 U11176 ( .A1(n8490), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(n8491)
         );
  NAND2_X1 U11177 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  NAND2_X1 U11178 ( .A1(n15553), .A2(n8493), .ZN(n10028) );
  INV_X1 U11179 ( .A(n10028), .ZN(n8498) );
  INV_X1 U11180 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15556) );
  NAND2_X1 U11181 ( .A1(n15553), .A2(n15556), .ZN(n8495) );
  NAND2_X1 U11182 ( .A1(n12225), .A2(n12671), .ZN(n8494) );
  NAND2_X1 U11183 ( .A1(n8495), .A2(n8494), .ZN(n15557) );
  INV_X1 U11184 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15561) );
  NAND2_X1 U11185 ( .A1(n15553), .A2(n15561), .ZN(n8497) );
  NAND2_X1 U11186 ( .A1(n12481), .A2(n12671), .ZN(n8496) );
  NAND2_X1 U11187 ( .A1(n8497), .A2(n8496), .ZN(n10114) );
  NAND2_X1 U11188 ( .A1(n8499), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8501) );
  INV_X1 U11189 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8500) );
  XNOR2_X1 U11190 ( .A(n8501), .B(n8500), .ZN(n12399) );
  INV_X1 U11191 ( .A(n8504), .ZN(n10976) );
  INV_X1 U11192 ( .A(n14072), .ZN(n8522) );
  NAND2_X1 U11193 ( .A1(n13756), .A2(n14076), .ZN(n8525) );
  NOR2_X1 U11194 ( .A1(n15564), .A2(n10899), .ZN(n8502) );
  NOR2_X1 U11195 ( .A1(n8504), .A2(n12014), .ZN(n10041) );
  NAND2_X1 U11196 ( .A1(n8521), .A2(n10041), .ZN(n8507) );
  AND2_X2 U11197 ( .A1(n14070), .A2(n13757), .ZN(n14564) );
  NAND2_X1 U11198 ( .A1(n14564), .A2(n8505), .ZN(n10115) );
  INV_X1 U11199 ( .A(n10115), .ZN(n8506) );
  INV_X1 U11200 ( .A(n8510), .ZN(n8508) );
  NAND2_X1 U11201 ( .A1(n8508), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n10042) );
  INV_X1 U11202 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U11203 ( .A1(n8510), .A2(n8509), .ZN(n8511) );
  NAND2_X1 U11204 ( .A1(n10042), .A2(n8511), .ZN(n12853) );
  INV_X1 U11205 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U11206 ( .A1(n10379), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U11207 ( .A1(n8512), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8513) );
  OAI211_X1 U11208 ( .C1(n7040), .C2(n8515), .A(n8514), .B(n8513), .ZN(n8516)
         );
  INV_X1 U11209 ( .A(n8516), .ZN(n8517) );
  INV_X1 U11210 ( .A(n14082), .ZN(n8520) );
  INV_X1 U11211 ( .A(n10904), .ZN(n8519) );
  OAI22_X1 U11212 ( .A1(n8520), .A2(n13734), .B1(n13986), .B2(n13732), .ZN(
        n14301) );
  INV_X1 U11213 ( .A(n8521), .ZN(n8523) );
  NAND2_X1 U11214 ( .A1(n8524), .A2(n10115), .ZN(n8528) );
  OR2_X1 U11215 ( .A1(n8525), .A2(n14072), .ZN(n10027) );
  AND2_X1 U11216 ( .A1(n8526), .A2(n10027), .ZN(n8527) );
  NAND2_X1 U11217 ( .A1(n8528), .A2(n8527), .ZN(n11034) );
  OAI22_X1 U11218 ( .A1(n14308), .A2(n13748), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8529), .ZN(n8530) );
  AOI21_X1 U11219 ( .B1(n14301), .B2(n13746), .A(n8530), .ZN(n8531) );
  OAI21_X1 U11220 ( .B1(n14310), .B2(n13738), .A(n8531), .ZN(n8532) );
  INV_X1 U11221 ( .A(n8532), .ZN(n8533) );
  INV_X1 U11222 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n9122) );
  INV_X1 U11223 ( .A(n8759), .ZN(n8709) );
  INV_X1 U11224 ( .A(n8760), .ZN(n8708) );
  NOR2_X1 U11225 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), 
        .ZN(n8538) );
  NOR2_X1 U11226 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), 
        .ZN(n8540) );
  INV_X1 U11227 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n12834) );
  OR2_X1 U11228 ( .A1(n8577), .A2(n12834), .ZN(n8550) );
  INV_X1 U11229 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11287) );
  OR2_X1 U11230 ( .A1(n8969), .A2(n11287), .ZN(n8549) );
  INV_X1 U11231 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11859) );
  OR2_X1 U11232 ( .A1(n8744), .A2(n11859), .ZN(n8548) );
  NAND2_X1 U11233 ( .A1(n8556), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8557) );
  AND2_X1 U11234 ( .A1(n8563), .A2(n8557), .ZN(n10785) );
  OR2_X1 U11235 ( .A1(n8905), .A2(n10785), .ZN(n8558) );
  INV_X1 U11236 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15596) );
  OR2_X1 U11237 ( .A1(n8969), .A2(n15596), .ZN(n8560) );
  INV_X1 U11238 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11334) );
  INV_X1 U11239 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11212) );
  XNOR2_X1 U11240 ( .A(n8563), .B(n8565), .ZN(n10791) );
  NAND2_X1 U11241 ( .A1(n9018), .A2(n11331), .ZN(n11309) );
  NAND2_X1 U11242 ( .A1(n11311), .A2(n11309), .ZN(n11676) );
  NAND2_X1 U11243 ( .A1(n9268), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8576) );
  INV_X1 U11244 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8562) );
  OR2_X1 U11245 ( .A1(n8561), .A2(n8562), .ZN(n8575) );
  OR2_X1 U11246 ( .A1(n8969), .A2(n9177), .ZN(n8574) );
  INV_X1 U11247 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15577) );
  OR2_X1 U11248 ( .A1(n8744), .A2(n15577), .ZN(n8573) );
  OR2_X1 U11249 ( .A1(n9288), .A2(SI_2_), .ZN(n8572) );
  INV_X1 U11250 ( .A(n8563), .ZN(n8564) );
  NAND2_X1 U11251 ( .A1(n10803), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U11252 ( .A1(n10820), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8567) );
  XNOR2_X1 U11253 ( .A(n8583), .B(n8582), .ZN(n10808) );
  OR2_X1 U11254 ( .A1(n8905), .A2(n10808), .ZN(n8571) );
  XNOR2_X2 U11255 ( .A(n8569), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9176) );
  OR2_X1 U11256 ( .A1(n9168), .A2(n9176), .ZN(n8570) );
  INV_X1 U11257 ( .A(n11345), .ZN(n11679) );
  NAND2_X1 U11258 ( .A1(n13105), .A2(n11679), .ZN(n9319) );
  NAND2_X1 U11259 ( .A1(n11676), .A2(n11675), .ZN(n12028) );
  NAND2_X1 U11260 ( .A1(n9279), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8581) );
  INV_X1 U11261 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15632) );
  OR2_X1 U11262 ( .A1(n8577), .A2(n15632), .ZN(n8580) );
  INV_X1 U11263 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n12036) );
  OR2_X1 U11264 ( .A1(n8969), .A2(n12036), .ZN(n8579) );
  OR2_X1 U11265 ( .A1(n8744), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8578) );
  OR2_X1 U11266 ( .A1(n9288), .A2(SI_3_), .ZN(n8589) );
  NAND2_X1 U11267 ( .A1(n7822), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8585) );
  XNOR2_X1 U11268 ( .A(n8599), .B(n8598), .ZN(n10806) );
  OR2_X1 U11269 ( .A1(n8905), .A2(n10806), .ZN(n8588) );
  NAND2_X1 U11270 ( .A1(n8759), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8586) );
  OR2_X1 U11271 ( .A1(n9168), .A2(n11145), .ZN(n8587) );
  NAND2_X1 U11272 ( .A1(n8591), .A2(n12038), .ZN(n9326) );
  AND2_X1 U11273 ( .A1(n12027), .A2(n9326), .ZN(n8590) );
  INV_X1 U11274 ( .A(n12038), .ZN(n15603) );
  NAND2_X1 U11275 ( .A1(n9024), .A2(n15603), .ZN(n9329) );
  NAND2_X1 U11276 ( .A1(n9279), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U11277 ( .A1(n9278), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U11278 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8593) );
  AND2_X1 U11279 ( .A1(n8605), .A2(n8593), .ZN(n12023) );
  OR2_X1 U11280 ( .A1(n8744), .A2(n12023), .ZN(n8594) );
  NAND2_X1 U11281 ( .A1(n8612), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11282 ( .A1(n10796), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8601) );
  XNOR2_X1 U11283 ( .A(n8617), .B(n8616), .ZN(n10804) );
  OR2_X1 U11284 ( .A1(n8905), .A2(n10804), .ZN(n8602) );
  INV_X1 U11285 ( .A(n12018), .ZN(n9328) );
  INV_X1 U11286 ( .A(n13104), .ZN(n11684) );
  INV_X1 U11287 ( .A(n9337), .ZN(n15613) );
  NAND2_X1 U11288 ( .A1(n11684), .A2(n15613), .ZN(n9335) );
  NAND2_X1 U11289 ( .A1(n9279), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8611) );
  INV_X1 U11290 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15635) );
  OR2_X1 U11291 ( .A1(n8577), .A2(n15635), .ZN(n8610) );
  NAND2_X1 U11292 ( .A1(n8605), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8606) );
  AND2_X1 U11293 ( .A1(n8624), .A2(n8606), .ZN(n12133) );
  OR2_X1 U11294 ( .A1(n8744), .A2(n12133), .ZN(n8609) );
  INV_X1 U11295 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n8607) );
  OR2_X1 U11296 ( .A1(n8969), .A2(n8607), .ZN(n8608) );
  INV_X1 U11297 ( .A(n8612), .ZN(n8614) );
  NAND2_X1 U11298 ( .A1(n8614), .A2(n8613), .ZN(n8706) );
  NAND2_X1 U11299 ( .A1(n8706), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8615) );
  OR2_X1 U11300 ( .A1(n9288), .A2(SI_5_), .ZN(n8622) );
  NAND2_X1 U11301 ( .A1(n8617), .A2(n8616), .ZN(n8619) );
  NAND2_X1 U11302 ( .A1(n10841), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8620) );
  XNOR2_X1 U11303 ( .A(n8633), .B(n8632), .ZN(n10817) );
  OR2_X1 U11304 ( .A1(n8905), .A2(n10817), .ZN(n8621) );
  OAI211_X1 U11305 ( .C1(n11160), .C2(n9168), .A(n8622), .B(n8621), .ZN(n15616) );
  INV_X1 U11306 ( .A(n15616), .ZN(n11682) );
  NAND2_X1 U11307 ( .A1(n11863), .A2(n11682), .ZN(n9343) );
  INV_X1 U11308 ( .A(n11863), .ZN(n13103) );
  NAND2_X1 U11309 ( .A1(n13103), .A2(n15616), .ZN(n9334) );
  NAND2_X1 U11310 ( .A1(n8623), .A2(n9343), .ZN(n12055) );
  NAND2_X1 U11311 ( .A1(n9279), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8630) );
  INV_X1 U11312 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n12063) );
  OR2_X1 U11313 ( .A1(n9068), .A2(n12063), .ZN(n8629) );
  NAND2_X1 U11314 ( .A1(n8624), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8625) );
  AND2_X1 U11315 ( .A1(n8642), .A2(n8625), .ZN(n12064) );
  OR2_X1 U11316 ( .A1(n8744), .A2(n12064), .ZN(n8628) );
  INV_X1 U11317 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n8626) );
  OR2_X1 U11318 ( .A1(n8577), .A2(n8626), .ZN(n8627) );
  NAND2_X1 U11319 ( .A1(n8648), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8631) );
  INV_X1 U11320 ( .A(SI_6_), .ZN(n10836) );
  OR2_X1 U11321 ( .A1(n9288), .A2(n10836), .ZN(n8638) );
  NAND2_X1 U11322 ( .A1(n8633), .A2(n8632), .ZN(n8635) );
  XNOR2_X1 U11323 ( .A(n10860), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8636) );
  XNOR2_X1 U11324 ( .A(n8654), .B(n8636), .ZN(n10837) );
  OR2_X1 U11325 ( .A1(n8905), .A2(n10837), .ZN(n8637) );
  OAI211_X1 U11326 ( .C1(n9168), .C2(n11488), .A(n8638), .B(n8637), .ZN(n12066) );
  NAND2_X1 U11327 ( .A1(n8639), .A2(n12066), .ZN(n9344) );
  INV_X1 U11328 ( .A(n12066), .ZN(n15622) );
  NAND2_X1 U11329 ( .A1(n13102), .A2(n15622), .ZN(n9345) );
  NAND2_X1 U11330 ( .A1(n9344), .A2(n9345), .ZN(n12058) );
  INV_X1 U11331 ( .A(n12058), .ZN(n8640) );
  NAND2_X1 U11332 ( .A1(n9279), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U11333 ( .A1(n9278), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U11334 ( .A1(n8642), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8643) );
  AND2_X1 U11335 ( .A1(n8675), .A2(n8643), .ZN(n12180) );
  OR2_X1 U11336 ( .A1(n8744), .A2(n12180), .ZN(n8645) );
  INV_X1 U11337 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15659) );
  OR2_X1 U11338 ( .A1(n8577), .A2(n15659), .ZN(n8644) );
  NAND4_X1 U11339 ( .A1(n8647), .A2(n8646), .A3(n8645), .A4(n8644), .ZN(n13101) );
  INV_X1 U11340 ( .A(n8648), .ZN(n8650) );
  NAND2_X1 U11341 ( .A1(n8650), .A2(n8649), .ZN(n8671) );
  NAND2_X1 U11342 ( .A1(n8671), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8651) );
  OAI22_X1 U11343 ( .A1(n9288), .A2(SI_7_), .B1(n11388), .B2(n9168), .ZN(n8652) );
  INV_X1 U11344 ( .A(n8652), .ZN(n8663) );
  NAND2_X1 U11345 ( .A1(n10839), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U11346 ( .A1(n10860), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U11347 ( .A1(n10858), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U11348 ( .A1(n8665), .A2(n8657), .ZN(n8659) );
  NAND2_X1 U11349 ( .A1(n8660), .A2(n8659), .ZN(n8661) );
  NAND2_X1 U11350 ( .A1(n8666), .A2(n8661), .ZN(n10789) );
  NAND2_X1 U11351 ( .A1(n10789), .A2(n9287), .ZN(n8662) );
  NAND2_X1 U11352 ( .A1(n8663), .A2(n8662), .ZN(n12110) );
  INV_X1 U11353 ( .A(n13101), .ZN(n8664) );
  INV_X1 U11354 ( .A(n12110), .ZN(n12177) );
  NAND2_X1 U11355 ( .A1(n8664), .A2(n12177), .ZN(n9350) );
  NAND2_X1 U11356 ( .A1(n10872), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U11357 ( .A1(n10871), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8667) );
  OR2_X1 U11358 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  NAND2_X1 U11359 ( .A1(n8683), .A2(n8670), .ZN(n10787) );
  OR2_X1 U11360 ( .A1(n10787), .A2(n8905), .ZN(n8674) );
  NAND2_X1 U11361 ( .A1(n8688), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8672) );
  AOI22_X1 U11362 ( .A1(n8886), .A2(SI_8_), .B1(n11460), .B2(n8885), .ZN(n8673) );
  NAND2_X1 U11363 ( .A1(n9279), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11364 ( .A1(n9268), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U11365 ( .A1(n9278), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U11366 ( .A1(n8675), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8676) );
  AND2_X1 U11367 ( .A1(n8694), .A2(n8676), .ZN(n12312) );
  OR2_X1 U11368 ( .A1(n8744), .A2(n12312), .ZN(n8677) );
  NAND4_X1 U11369 ( .A1(n8680), .A2(n8679), .A3(n8678), .A4(n8677), .ZN(n13100) );
  NAND2_X1 U11370 ( .A1(n13490), .A2(n13100), .ZN(n9355) );
  NAND2_X1 U11371 ( .A1(n12360), .A2(n12309), .ZN(n9354) );
  NAND2_X1 U11372 ( .A1(n12042), .A2(n12043), .ZN(n8681) );
  NAND2_X1 U11373 ( .A1(n8683), .A2(n8682), .ZN(n8686) );
  NAND2_X1 U11374 ( .A1(n10875), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U11375 ( .A1(n10874), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8684) );
  OR2_X1 U11376 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  NAND2_X1 U11377 ( .A1(n8701), .A2(n8687), .ZN(n10793) );
  NAND2_X1 U11378 ( .A1(n10793), .A2(n9287), .ZN(n8692) );
  OAI21_X1 U11379 ( .B1(n8688), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8690) );
  INV_X1 U11380 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8689) );
  XNOR2_X1 U11381 ( .A(n8690), .B(n8689), .ZN(n11891) );
  INV_X1 U11382 ( .A(SI_9_), .ZN(n10794) );
  AOI22_X1 U11383 ( .A1(n11891), .A2(n8885), .B1(n8886), .B2(n10794), .ZN(
        n8691) );
  NAND2_X2 U11384 ( .A1(n8692), .A2(n8691), .ZN(n12485) );
  NAND2_X1 U11385 ( .A1(n9268), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8699) );
  INV_X1 U11386 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n12275) );
  OR2_X1 U11387 ( .A1(n8561), .A2(n12275), .ZN(n8698) );
  NAND2_X1 U11388 ( .A1(n8694), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8695) );
  AND2_X1 U11389 ( .A1(n8713), .A2(n8695), .ZN(n12484) );
  OR2_X1 U11390 ( .A1(n8744), .A2(n12484), .ZN(n8697) );
  INV_X1 U11391 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11892) );
  OR2_X1 U11392 ( .A1(n8969), .A2(n11892), .ZN(n8696) );
  NOR2_X1 U11393 ( .A1(n12485), .A2(n13099), .ZN(n9359) );
  NAND2_X1 U11394 ( .A1(n12485), .A2(n13099), .ZN(n9358) );
  NAND2_X1 U11395 ( .A1(n10919), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8720) );
  INV_X1 U11396 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10917) );
  NAND2_X1 U11397 ( .A1(n10917), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8702) );
  OR2_X1 U11398 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  NAND2_X1 U11399 ( .A1(n8721), .A2(n8705), .ZN(n10798) );
  NAND2_X1 U11400 ( .A1(n10798), .A2(n9287), .ZN(n8712) );
  INV_X1 U11401 ( .A(SI_10_), .ZN(n10799) );
  OAI21_X1 U11402 ( .B1(n8706), .B2(n8760), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8707) );
  MUX2_X1 U11403 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8707), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n8710) );
  NAND3_X1 U11404 ( .A1(n8709), .A2(n8708), .A3(n6508), .ZN(n8724) );
  NAND2_X1 U11405 ( .A1(n8710), .A2(n8724), .ZN(n10800) );
  AOI22_X1 U11406 ( .A1(n8886), .A2(n10799), .B1(n8885), .B2(n10800), .ZN(
        n8711) );
  NAND2_X1 U11407 ( .A1(n9279), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11408 ( .A1(n9268), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U11409 ( .A1(n8713), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8714) );
  AND2_X1 U11410 ( .A1(n8728), .A2(n8714), .ZN(n12341) );
  OR2_X1 U11411 ( .A1(n8744), .A2(n12341), .ZN(n8716) );
  INV_X1 U11412 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n15759) );
  NAND4_X1 U11413 ( .A1(n8718), .A2(n8717), .A3(n8716), .A4(n8715), .ZN(n13098) );
  NAND2_X1 U11414 ( .A1(n12955), .A2(n13098), .ZN(n9362) );
  INV_X1 U11415 ( .A(n9362), .ZN(n8719) );
  XNOR2_X1 U11416 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8722) );
  XNOR2_X1 U11417 ( .A(n8736), .B(n8722), .ZN(n10824) );
  NAND2_X1 U11418 ( .A1(n10824), .A2(n9287), .ZN(n8727) );
  NAND2_X1 U11419 ( .A1(n8724), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8723) );
  MUX2_X1 U11420 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8723), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n8725) );
  OR2_X1 U11421 ( .A1(n8724), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U11422 ( .A1(n8725), .A2(n8738), .ZN(n10826) );
  AOI22_X1 U11423 ( .A1(n8886), .A2(n10825), .B1(n8885), .B2(n10826), .ZN(
        n8726) );
  NAND2_X1 U11424 ( .A1(n9268), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11425 ( .A1(n8728), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8729) );
  AND2_X1 U11426 ( .A1(n8746), .A2(n8729), .ZN(n12534) );
  OR2_X1 U11427 ( .A1(n8744), .A2(n12534), .ZN(n8732) );
  NAND2_X1 U11428 ( .A1(n9279), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8731) );
  INV_X1 U11429 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12533) );
  OR2_X1 U11430 ( .A1(n8969), .A2(n12533), .ZN(n8730) );
  NAND4_X1 U11431 ( .A1(n8733), .A2(n8732), .A3(n8731), .A4(n8730), .ZN(n13097) );
  NAND2_X1 U11432 ( .A1(n12615), .A2(n13097), .ZN(n9365) );
  NAND2_X1 U11433 ( .A1(n9364), .A2(n9365), .ZN(n12523) );
  INV_X1 U11434 ( .A(n12523), .ZN(n12530) );
  INV_X1 U11435 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10944) );
  NAND2_X1 U11436 ( .A1(n10944), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8735) );
  INV_X1 U11437 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10945) );
  XNOR2_X1 U11438 ( .A(n11066), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n8752) );
  XNOR2_X1 U11439 ( .A(n8754), .B(n8752), .ZN(n10866) );
  NAND2_X1 U11440 ( .A1(n10866), .A2(n9287), .ZN(n8743) );
  NAND2_X1 U11441 ( .A1(n8738), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8737) );
  MUX2_X1 U11442 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8737), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8741) );
  INV_X1 U11443 ( .A(n8738), .ZN(n8740) );
  NAND2_X1 U11444 ( .A1(n8740), .A2(n8739), .ZN(n8757) );
  NAND2_X1 U11445 ( .A1(n8741), .A2(n8757), .ZN(n10869) );
  INV_X1 U11446 ( .A(n10869), .ZN(n13124) );
  AOI22_X1 U11447 ( .A1(n8886), .A2(SI_12_), .B1(n8885), .B2(n13124), .ZN(
        n8742) );
  INV_X1 U11448 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11449 ( .A1(n8746), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U11450 ( .A1(n8768), .A2(n8747), .ZN(n12631) );
  NAND2_X1 U11451 ( .A1(n9258), .A2(n12631), .ZN(n8751) );
  INV_X1 U11452 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12623) );
  OR2_X1 U11453 ( .A1(n8577), .A2(n12623), .ZN(n8750) );
  INV_X1 U11454 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n12626) );
  OR2_X1 U11455 ( .A1(n8561), .A2(n12626), .ZN(n8749) );
  INV_X1 U11456 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12629) );
  OR2_X1 U11457 ( .A1(n9068), .A2(n12629), .ZN(n8748) );
  NAND2_X1 U11458 ( .A1(n12632), .A2(n12589), .ZN(n9371) );
  INV_X1 U11459 ( .A(n8752), .ZN(n8753) );
  NAND2_X1 U11460 ( .A1(n11065), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8755) );
  XNOR2_X1 U11461 ( .A(n8798), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8775) );
  XNOR2_X1 U11462 ( .A(n8775), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10891) );
  NAND2_X1 U11463 ( .A1(n10891), .A2(n9287), .ZN(n8765) );
  NAND2_X1 U11464 ( .A1(n8757), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8758) );
  MUX2_X1 U11465 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8758), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8763) );
  NAND2_X1 U11466 ( .A1(n8763), .A2(n8781), .ZN(n13146) );
  AOI22_X1 U11467 ( .A1(n8886), .A2(n10892), .B1(n8885), .B2(n13146), .ZN(
        n8764) );
  INV_X1 U11468 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U11469 ( .A1(n8768), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U11470 ( .A1(n8785), .A2(n8769), .ZN(n12758) );
  NAND2_X1 U11471 ( .A1(n9258), .A2(n12758), .ZN(n8773) );
  INV_X1 U11472 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13134) );
  OR2_X1 U11473 ( .A1(n8577), .A2(n13134), .ZN(n8772) );
  INV_X1 U11474 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12747) );
  OR2_X1 U11475 ( .A1(n8561), .A2(n12747), .ZN(n8771) );
  INV_X1 U11476 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12755) );
  OR2_X1 U11477 ( .A1(n8969), .A2(n12755), .ZN(n8770) );
  NOR2_X1 U11478 ( .A1(n12757), .A2(n13095), .ZN(n9374) );
  NAND2_X1 U11479 ( .A1(n12757), .A2(n13095), .ZN(n9299) );
  NAND2_X1 U11480 ( .A1(n8775), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U11481 ( .A1(n8798), .A2(n11092), .ZN(n8776) );
  NAND2_X1 U11482 ( .A1(n8777), .A2(n8776), .ZN(n8779) );
  XNOR2_X1 U11483 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8778) );
  XNOR2_X1 U11484 ( .A(n8779), .B(n8778), .ZN(n10895) );
  NAND2_X1 U11485 ( .A1(n10895), .A2(n9287), .ZN(n8784) );
  NAND2_X1 U11486 ( .A1(n8781), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8780) );
  MUX2_X1 U11487 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8780), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n8782) );
  NAND2_X1 U11488 ( .A1(n8782), .A2(n9090), .ZN(n10897) );
  AOI22_X1 U11489 ( .A1(n8886), .A2(n10896), .B1(n8885), .B2(n10897), .ZN(
        n8783) );
  NAND2_X1 U11490 ( .A1(n8785), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U11491 ( .A1(n8807), .A2(n8786), .ZN(n13426) );
  NAND2_X1 U11492 ( .A1(n13426), .A2(n9258), .ZN(n8790) );
  NAND2_X1 U11493 ( .A1(n9268), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U11494 ( .A1(n9279), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8788) );
  NAND2_X1 U11495 ( .A1(n9278), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8787) );
  NAND4_X1 U11496 ( .A1(n8790), .A2(n8789), .A3(n8788), .A4(n8787), .ZN(n13094) );
  NAND2_X1 U11497 ( .A1(n13579), .A2(n13094), .ZN(n9382) );
  INV_X1 U11498 ( .A(n9382), .ZN(n8791) );
  NAND2_X1 U11499 ( .A1(n15740), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8792) );
  OAI21_X1 U11500 ( .B1(n11090), .B2(P2_DATAO_REG_13__SCAN_IN), .A(n8792), 
        .ZN(n8797) );
  NAND2_X1 U11501 ( .A1(n11090), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U11502 ( .A1(n8793), .A2(n15740), .ZN(n8795) );
  INV_X1 U11503 ( .A(n8793), .ZN(n8794) );
  AOI22_X1 U11504 ( .A1(n11349), .A2(n8795), .B1(n8794), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U11505 ( .A1(n15732), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U11506 ( .A1(n11517), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U11507 ( .A1(n8811), .A2(n8799), .ZN(n8800) );
  NAND2_X1 U11508 ( .A1(n8801), .A2(n8800), .ZN(n8802) );
  NAND2_X1 U11509 ( .A1(n8812), .A2(n8802), .ZN(n10893) );
  OR2_X1 U11510 ( .A1(n10893), .A2(n8905), .ZN(n8805) );
  NAND2_X1 U11511 ( .A1(n9090), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8803) );
  XNOR2_X1 U11512 ( .A(n8803), .B(P3_IR_REG_15__SCAN_IN), .ZN(n9227) );
  AOI22_X1 U11513 ( .A1(n8886), .A2(SI_15_), .B1(n8885), .B2(n9227), .ZN(n8804) );
  INV_X1 U11514 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13478) );
  INV_X1 U11515 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U11516 ( .A1(n8807), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U11517 ( .A1(n8819), .A2(n8808), .ZN(n13075) );
  NAND2_X1 U11518 ( .A1(n13075), .A2(n9258), .ZN(n8810) );
  AOI22_X1 U11519 ( .A1(n9278), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n9279), .B2(
        P3_REG0_REG_15__SCAN_IN), .ZN(n8809) );
  XNOR2_X1 U11520 ( .A(n13477), .B(n13093), .ZN(n9378) );
  INV_X1 U11521 ( .A(n13093), .ZN(n9379) );
  NAND2_X1 U11522 ( .A1(n13477), .A2(n9379), .ZN(n9385) );
  NAND2_X1 U11523 ( .A1(n11336), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U11524 ( .A1(n11337), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8813) );
  AND2_X1 U11525 ( .A1(n8824), .A2(n8813), .ZN(n8814) );
  OR2_X1 U11526 ( .A1(n8815), .A2(n8814), .ZN(n8816) );
  NAND2_X1 U11527 ( .A1(n8825), .A2(n8816), .ZN(n10922) );
  OR2_X1 U11528 ( .A1(n10922), .A2(n8905), .ZN(n8818) );
  NAND2_X1 U11529 ( .A1(n7502), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8828) );
  XNOR2_X1 U11530 ( .A(n8828), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U11531 ( .A1(n8886), .A2(SI_16_), .B1(n8885), .B2(n13182), .ZN(
        n8817) );
  INV_X1 U11532 ( .A(n8833), .ZN(n8834) );
  NAND2_X1 U11533 ( .A1(n8819), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U11534 ( .A1(n8834), .A2(n8820), .ZN(n13413) );
  NAND2_X1 U11535 ( .A1(n13413), .A2(n9258), .ZN(n8823) );
  AOI22_X1 U11536 ( .A1(n9268), .A2(P3_REG1_REG_16__SCAN_IN), .B1(n9279), .B2(
        P3_REG0_REG_16__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U11537 ( .A1(n9278), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8821) );
  OR2_X1 U11538 ( .A1(n13414), .A2(n13008), .ZN(n9381) );
  NAND2_X1 U11539 ( .A1(n13414), .A2(n13008), .ZN(n13391) );
  NAND2_X1 U11540 ( .A1(n9381), .A2(n13391), .ZN(n13409) );
  INV_X1 U11541 ( .A(n13409), .ZN(n13405) );
  NAND2_X1 U11542 ( .A1(n13406), .A2(n13405), .ZN(n13390) );
  NAND2_X1 U11543 ( .A1(n11510), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11544 ( .A1(n11509), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U11545 ( .A1(n8843), .A2(n8826), .ZN(n8840) );
  XNOR2_X1 U11546 ( .A(n8842), .B(n8840), .ZN(n11040) );
  NAND2_X1 U11547 ( .A1(n11040), .A2(n9287), .ZN(n8832) );
  INV_X1 U11548 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U11549 ( .A1(n8828), .A2(n8827), .ZN(n8829) );
  NAND2_X1 U11550 ( .A1(n8829), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8830) );
  XNOR2_X1 U11551 ( .A(n8830), .B(P3_IR_REG_17__SCAN_IN), .ZN(n9232) );
  AOI22_X1 U11552 ( .A1(n8886), .A2(SI_17_), .B1(n9232), .B2(n8885), .ZN(n8831) );
  INV_X1 U11553 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15748) );
  NAND2_X1 U11554 ( .A1(n8834), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11555 ( .A1(n8889), .A2(n8835), .ZN(n13402) );
  INV_X1 U11556 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13401) );
  NAND2_X1 U11557 ( .A1(n9279), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U11558 ( .A1(n9268), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8836) );
  OAI211_X1 U11559 ( .C1(n9068), .C2(n13401), .A(n8837), .B(n8836), .ZN(n8838)
         );
  AOI21_X1 U11560 ( .B1(n13402), .B2(n9258), .A(n8838), .ZN(n13049) );
  NAND2_X1 U11561 ( .A1(n13559), .A2(n13049), .ZN(n9392) );
  AND2_X1 U11562 ( .A1(n13391), .A2(n9392), .ZN(n8839) );
  OR2_X1 U11563 ( .A1(n13559), .A2(n13049), .ZN(n9389) );
  INV_X1 U11564 ( .A(n8840), .ZN(n8841) );
  NAND2_X1 U11565 ( .A1(n11744), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U11566 ( .A1(n11743), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8844) );
  AND2_X1 U11567 ( .A1(n8845), .A2(n8844), .ZN(n8879) );
  NAND2_X1 U11568 ( .A1(n8882), .A2(n8845), .ZN(n8862) );
  INV_X1 U11569 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12823) );
  NAND2_X1 U11570 ( .A1(n12823), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8847) );
  INV_X1 U11571 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12099) );
  NAND2_X1 U11572 ( .A1(n12099), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8846) );
  AND2_X1 U11573 ( .A1(n8847), .A2(n8846), .ZN(n8861) );
  INV_X1 U11574 ( .A(n8849), .ZN(n8848) );
  NAND2_X1 U11575 ( .A1(n8850), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11576 ( .A1(n8900), .A2(n8851), .ZN(n11525) );
  OR2_X1 U11577 ( .A1(n9288), .A2(n11524), .ZN(n8852) );
  INV_X1 U11578 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U11579 ( .A1(n8873), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U11580 ( .A1(n8908), .A2(n8855), .ZN(n13348) );
  NAND2_X1 U11581 ( .A1(n13348), .A2(n9258), .ZN(n8860) );
  INV_X1 U11582 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13356) );
  NAND2_X1 U11583 ( .A1(n9279), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8857) );
  NAND2_X1 U11584 ( .A1(n9268), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8856) );
  OAI211_X1 U11585 ( .C1(n9068), .C2(n13356), .A(n8857), .B(n8856), .ZN(n8858)
         );
  INV_X1 U11586 ( .A(n8858), .ZN(n8859) );
  OR2_X1 U11587 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  NAND2_X1 U11588 ( .A1(n8864), .A2(n8863), .ZN(n11178) );
  NAND2_X1 U11589 ( .A1(n11178), .A2(n9287), .ZN(n8871) );
  NAND2_X1 U11590 ( .A1(n8868), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8867) );
  MUX2_X1 U11591 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8867), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8869) );
  NAND2_X1 U11592 ( .A1(n8869), .A2(n9002), .ZN(n11176) );
  AOI22_X1 U11593 ( .A1(n11176), .A2(n8885), .B1(n8886), .B2(n11177), .ZN(
        n8870) );
  NAND2_X1 U11594 ( .A1(n8891), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U11595 ( .A1(n8873), .A2(n8872), .ZN(n13361) );
  NAND2_X1 U11596 ( .A1(n13361), .A2(n9258), .ZN(n8878) );
  INV_X1 U11597 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13372) );
  NAND2_X1 U11598 ( .A1(n9268), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U11599 ( .A1(n9279), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8874) );
  OAI211_X1 U11600 ( .C1(n13372), .C2(n9068), .A(n8875), .B(n8874), .ZN(n8876)
         );
  INV_X1 U11601 ( .A(n8876), .ZN(n8877) );
  NAND2_X1 U11602 ( .A1(n8878), .A2(n8877), .ZN(n13089) );
  NAND2_X1 U11603 ( .A1(n13546), .A2(n13089), .ZN(n9400) );
  NAND2_X1 U11604 ( .A1(n13327), .A2(n9400), .ZN(n8915) );
  OR2_X1 U11605 ( .A1(n8880), .A2(n8879), .ZN(n8881) );
  NAND2_X1 U11606 ( .A1(n8882), .A2(n8881), .ZN(n11068) );
  OR2_X1 U11607 ( .A1(n11068), .A2(n8905), .ZN(n8888) );
  NAND2_X1 U11608 ( .A1(n8883), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8884) );
  XNOR2_X1 U11609 ( .A(n8884), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13211) );
  AOI22_X1 U11610 ( .A1(n8886), .A2(SI_18_), .B1(n13211), .B2(n8885), .ZN(
        n8887) );
  NAND2_X1 U11611 ( .A1(n8889), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11612 ( .A1(n8891), .A2(n8890), .ZN(n13387) );
  NAND2_X1 U11613 ( .A1(n13387), .A2(n9258), .ZN(n8896) );
  INV_X1 U11614 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13386) );
  NAND2_X1 U11615 ( .A1(n9279), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8893) );
  NAND2_X1 U11616 ( .A1(n9268), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8892) );
  OAI211_X1 U11617 ( .C1(n9068), .C2(n13386), .A(n8893), .B(n8892), .ZN(n8894)
         );
  INV_X1 U11618 ( .A(n8894), .ZN(n8895) );
  INV_X1 U11619 ( .A(n13325), .ZN(n8897) );
  NAND2_X1 U11620 ( .A1(n13553), .A2(n13009), .ZN(n9391) );
  NAND2_X1 U11621 ( .A1(n6700), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U11622 ( .A1(n12210), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8901) );
  AND2_X1 U11623 ( .A1(n8918), .A2(n8901), .ZN(n8902) );
  INV_X1 U11624 ( .A(SI_21_), .ZN(n12826) );
  OR2_X1 U11625 ( .A1(n9288), .A2(n12826), .ZN(n8906) );
  INV_X1 U11626 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U11627 ( .A1(n8908), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8909) );
  NAND2_X1 U11628 ( .A1(n8922), .A2(n8909), .ZN(n13329) );
  INV_X1 U11629 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13343) );
  NAND2_X1 U11630 ( .A1(n9268), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U11631 ( .A1(n9279), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8910) );
  OAI211_X1 U11632 ( .C1(n13343), .C2(n8969), .A(n8911), .B(n8910), .ZN(n8912)
         );
  AOI21_X1 U11633 ( .B1(n13329), .B2(n9258), .A(n8912), .ZN(n13031) );
  NAND2_X1 U11634 ( .A1(n13538), .A2(n13031), .ZN(n9405) );
  NAND2_X1 U11635 ( .A1(n9399), .A2(n13088), .ZN(n8913) );
  INV_X1 U11636 ( .A(n9399), .ZN(n13326) );
  AOI22_X1 U11637 ( .A1(n13543), .A2(n8913), .B1(n13335), .B2(n13326), .ZN(
        n8914) );
  OAI211_X1 U11638 ( .C1(n8915), .C2(n9391), .A(n9405), .B(n8914), .ZN(n8916)
         );
  INV_X1 U11639 ( .A(n8916), .ZN(n8917) );
  XNOR2_X1 U11640 ( .A(n12220), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8930) );
  XNOR2_X1 U11641 ( .A(n8931), .B(n8930), .ZN(n11820) );
  NAND2_X1 U11642 ( .A1(n11820), .A2(n9287), .ZN(n8921) );
  OR2_X1 U11643 ( .A1(n9288), .A2(n8919), .ZN(n8920) );
  NAND2_X1 U11644 ( .A1(n8922), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U11645 ( .A1(n8933), .A2(n8923), .ZN(n13322) );
  NAND2_X1 U11646 ( .A1(n13322), .A2(n9258), .ZN(n8928) );
  INV_X1 U11647 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U11648 ( .A1(n9268), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8925) );
  NAND2_X1 U11649 ( .A1(n9279), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8924) );
  OAI211_X1 U11650 ( .C1(n13321), .C2(n9068), .A(n8925), .B(n8924), .ZN(n8926)
         );
  INV_X1 U11651 ( .A(n8926), .ZN(n8927) );
  NAND2_X1 U11652 ( .A1(n13532), .A2(n12941), .ZN(n9408) );
  NAND2_X1 U11653 ( .A1(n12220), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8929) );
  XNOR2_X1 U11654 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8942) );
  XNOR2_X1 U11655 ( .A(n8943), .B(n8942), .ZN(n12226) );
  INV_X1 U11656 ( .A(SI_23_), .ZN(n12229) );
  OR2_X1 U11657 ( .A1(n9288), .A2(n12229), .ZN(n8932) );
  NAND2_X1 U11658 ( .A1(n8933), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U11659 ( .A1(n13308), .A2(n9258), .ZN(n8939) );
  INV_X1 U11660 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13309) );
  NAND2_X1 U11661 ( .A1(n9279), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8936) );
  NAND2_X1 U11662 ( .A1(n9268), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8935) );
  OAI211_X1 U11663 ( .C1(n9068), .C2(n13309), .A(n8936), .B(n8935), .ZN(n8937)
         );
  INV_X1 U11664 ( .A(n8937), .ZN(n8938) );
  OR2_X1 U11665 ( .A1(n13452), .A2(n12942), .ZN(n8940) );
  AND2_X1 U11666 ( .A1(n13299), .A2(n8940), .ZN(n8941) );
  INV_X1 U11667 ( .A(n8940), .ZN(n9313) );
  INV_X1 U11668 ( .A(n8945), .ZN(n8944) );
  NAND2_X1 U11669 ( .A1(n8945), .A2(n12223), .ZN(n8946) );
  XNOR2_X1 U11670 ( .A(n8959), .B(n15734), .ZN(n12507) );
  NAND2_X1 U11671 ( .A1(n12507), .A2(n9287), .ZN(n8948) );
  INV_X1 U11672 ( .A(SI_24_), .ZN(n12508) );
  OR2_X1 U11673 ( .A1(n9288), .A2(n12508), .ZN(n8947) );
  INV_X1 U11674 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U11675 ( .A1(n8950), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U11676 ( .A1(n8965), .A2(n8951), .ZN(n13294) );
  NAND2_X1 U11677 ( .A1(n13294), .A2(n9258), .ZN(n8957) );
  INV_X1 U11678 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11679 ( .A1(n9279), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U11680 ( .A1(n9268), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8952) );
  OAI211_X1 U11681 ( .C1(n9068), .C2(n8954), .A(n8953), .B(n8952), .ZN(n8955)
         );
  INV_X1 U11682 ( .A(n8955), .ZN(n8956) );
  NAND2_X1 U11683 ( .A1(n13026), .A2(n8958), .ZN(n9315) );
  XNOR2_X1 U11684 ( .A(n12483), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8960) );
  XNOR2_X1 U11685 ( .A(n8974), .B(n8960), .ZN(n13606) );
  NAND2_X1 U11686 ( .A1(n13606), .A2(n9287), .ZN(n8962) );
  OR2_X1 U11687 ( .A1(n9288), .A2(n13608), .ZN(n8961) );
  INV_X1 U11688 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U11689 ( .A1(n8965), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11690 ( .A1(n8978), .A2(n8966), .ZN(n13283) );
  INV_X1 U11691 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U11692 ( .A1(n9268), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8968) );
  NAND2_X1 U11693 ( .A1(n9279), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8967) );
  OAI211_X1 U11694 ( .C1(n8970), .C2(n8969), .A(n8968), .B(n8967), .ZN(n8971)
         );
  AOI21_X1 U11695 ( .B1(n13283), .B2(n9258), .A(n8971), .ZN(n12927) );
  NAND2_X1 U11696 ( .A1(n12483), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8973) );
  INV_X1 U11697 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U11698 ( .A1(n12479), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8975) );
  XNOR2_X1 U11699 ( .A(n12670), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8976) );
  XNOR2_X1 U11700 ( .A(n8987), .B(n8976), .ZN(n13602) );
  OR2_X1 U11701 ( .A1(n9288), .A2(n13604), .ZN(n8977) );
  NAND2_X1 U11702 ( .A1(n8978), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U11703 ( .A1(n8991), .A2(n8979), .ZN(n13271) );
  NAND2_X1 U11704 ( .A1(n13271), .A2(n9258), .ZN(n8985) );
  INV_X1 U11705 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U11706 ( .A1(n9268), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8981) );
  NAND2_X1 U11707 ( .A1(n9279), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8980) );
  OAI211_X1 U11708 ( .C1(n8982), .C2(n9068), .A(n8981), .B(n8980), .ZN(n8983)
         );
  INV_X1 U11709 ( .A(n8983), .ZN(n8984) );
  NAND2_X1 U11710 ( .A1(n13270), .A2(n12928), .ZN(n9416) );
  AND2_X1 U11711 ( .A1(n12672), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8986) );
  XNOR2_X1 U11712 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8988) );
  XNOR2_X1 U11713 ( .A(n9247), .B(n8988), .ZN(n13597) );
  NAND2_X1 U11714 ( .A1(n13597), .A2(n9287), .ZN(n8990) );
  INV_X1 U11715 ( .A(SI_27_), .ZN(n13599) );
  OR2_X1 U11716 ( .A1(n9288), .A2(n13599), .ZN(n8989) );
  INV_X1 U11717 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15720) );
  NAND2_X1 U11718 ( .A1(n8991), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U11719 ( .A1(n9064), .A2(n8992), .ZN(n13258) );
  NAND2_X1 U11720 ( .A1(n13258), .A2(n9258), .ZN(n8998) );
  INV_X1 U11721 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8995) );
  NAND2_X1 U11722 ( .A1(n9268), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U11723 ( .A1(n9279), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8993) );
  OAI211_X1 U11724 ( .C1(n8995), .C2(n9068), .A(n8994), .B(n8993), .ZN(n8996)
         );
  INV_X1 U11725 ( .A(n8996), .ZN(n8997) );
  NAND2_X1 U11726 ( .A1(n12934), .A2(n12976), .ZN(n13249) );
  XNOR2_X2 U11727 ( .A(n9003), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9010) );
  NAND2_X1 U11728 ( .A1(n12825), .A2(n9075), .ZN(n9009) );
  INV_X1 U11729 ( .A(n9090), .ZN(n9005) );
  NAND2_X1 U11730 ( .A1(n9005), .A2(n9004), .ZN(n9007) );
  NAND2_X1 U11731 ( .A1(n9007), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9006) );
  MUX2_X1 U11732 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9006), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9008) );
  NAND2_X1 U11733 ( .A1(n9009), .A2(n11818), .ZN(n9013) );
  INV_X2 U11734 ( .A(n11176), .ZN(n9308) );
  OAI21_X1 U11735 ( .B1(n9010), .B2(n11818), .A(n9308), .ZN(n9011) );
  NAND2_X1 U11736 ( .A1(n9011), .A2(n12825), .ZN(n9012) );
  NAND2_X1 U11737 ( .A1(n9013), .A2(n9012), .ZN(n11316) );
  NAND2_X1 U11738 ( .A1(n9075), .A2(n11176), .ZN(n9127) );
  INV_X1 U11739 ( .A(n9127), .ZN(n9455) );
  AND2_X1 U11740 ( .A1(n15621), .A2(n9455), .ZN(n9014) );
  NAND2_X1 U11741 ( .A1(n11316), .A2(n9014), .ZN(n9016) );
  NAND2_X1 U11742 ( .A1(n11176), .A2(n9456), .ZN(n9079) );
  INV_X1 U11743 ( .A(n9079), .ZN(n9015) );
  NAND2_X1 U11744 ( .A1(n9015), .A2(n9010), .ZN(n9118) );
  NAND2_X1 U11745 ( .A1(n9016), .A2(n9118), .ZN(n15627) );
  NAND2_X1 U11746 ( .A1(n13262), .A2(n15627), .ZN(n9074) );
  NAND2_X1 U11747 ( .A1(n13108), .A2(n9017), .ZN(n13491) );
  NAND2_X1 U11748 ( .A1(n13496), .A2(n13491), .ZN(n9019) );
  NAND2_X1 U11749 ( .A1(n9018), .A2(n13500), .ZN(n11308) );
  NAND2_X1 U11750 ( .A1(n9019), .A2(n11308), .ZN(n11672) );
  NAND2_X1 U11751 ( .A1(n11672), .A2(n11671), .ZN(n9022) );
  NAND2_X1 U11752 ( .A1(n9020), .A2(n11679), .ZN(n9021) );
  NAND2_X1 U11753 ( .A1(n9024), .A2(n12038), .ZN(n9025) );
  NAND2_X1 U11754 ( .A1(n13104), .A2(n15613), .ZN(n9026) );
  NAND2_X1 U11755 ( .A1(n11863), .A2(n15616), .ZN(n12057) );
  AND2_X1 U11756 ( .A1(n12058), .A2(n12057), .ZN(n9027) );
  AOI22_X1 U11757 ( .A1(n9027), .A2(n12134), .B1(n13102), .B2(n12066), .ZN(
        n9028) );
  NAND2_X1 U11758 ( .A1(n9029), .A2(n9028), .ZN(n11716) );
  NAND2_X1 U11759 ( .A1(n11716), .A2(n12173), .ZN(n11715) );
  NAND2_X1 U11760 ( .A1(n13101), .A2(n12177), .ZN(n9030) );
  NAND2_X1 U11761 ( .A1(n11715), .A2(n9030), .ZN(n12044) );
  NAND2_X1 U11762 ( .A1(n13490), .A2(n12360), .ZN(n9031) );
  XNOR2_X1 U11763 ( .A(n12485), .B(n12559), .ZN(n9357) );
  NAND2_X1 U11764 ( .A1(n9361), .A2(n9362), .ZN(n12331) );
  INV_X1 U11765 ( .A(n13098), .ZN(n9033) );
  OR2_X1 U11766 ( .A1(n12955), .A2(n9033), .ZN(n12520) );
  INV_X1 U11767 ( .A(n13097), .ZN(n12579) );
  NAND2_X1 U11768 ( .A1(n12615), .A2(n12579), .ZN(n9034) );
  INV_X1 U11769 ( .A(n12589), .ZN(n13096) );
  NAND2_X1 U11770 ( .A1(n12632), .A2(n13096), .ZN(n9035) );
  NAND2_X1 U11771 ( .A1(n12620), .A2(n9035), .ZN(n12744) );
  NAND2_X1 U11772 ( .A1(n12757), .A2(n12687), .ZN(n9036) );
  NAND2_X1 U11773 ( .A1(n12744), .A2(n9036), .ZN(n13420) );
  OR2_X1 U11774 ( .A1(n12757), .A2(n12687), .ZN(n13419) );
  INV_X1 U11775 ( .A(n13094), .ZN(n12900) );
  OR2_X1 U11776 ( .A1(n13579), .A2(n12900), .ZN(n9038) );
  AND2_X1 U11777 ( .A1(n13419), .A2(n9038), .ZN(n12779) );
  AND2_X1 U11778 ( .A1(n13477), .A2(n13093), .ZN(n9040) );
  INV_X1 U11779 ( .A(n9040), .ZN(n9037) );
  AND2_X1 U11780 ( .A1(n12779), .A2(n9037), .ZN(n9041) );
  INV_X1 U11781 ( .A(n9038), .ZN(n9039) );
  NAND2_X1 U11782 ( .A1(n9377), .A2(n9382), .ZN(n13417) );
  OR2_X1 U11783 ( .A1(n9039), .A2(n13417), .ZN(n12780) );
  NAND2_X1 U11784 ( .A1(n9389), .A2(n9392), .ZN(n13395) );
  AND2_X1 U11785 ( .A1(n13395), .A2(n13409), .ZN(n9042) );
  INV_X1 U11786 ( .A(n13395), .ZN(n13379) );
  INV_X1 U11787 ( .A(n13008), .ZN(n13092) );
  NAND2_X1 U11788 ( .A1(n13414), .A2(n13092), .ZN(n13393) );
  NAND2_X1 U11789 ( .A1(n13325), .A2(n9391), .ZN(n13382) );
  INV_X1 U11790 ( .A(n13049), .ZN(n13091) );
  NAND2_X1 U11791 ( .A1(n13559), .A2(n13091), .ZN(n13380) );
  OAI211_X1 U11792 ( .C1(n13379), .C2(n13393), .A(n13382), .B(n13380), .ZN(
        n9043) );
  INV_X1 U11793 ( .A(n9043), .ZN(n9044) );
  NAND2_X1 U11794 ( .A1(n9399), .A2(n9400), .ZN(n13366) );
  INV_X1 U11795 ( .A(n13009), .ZN(n13090) );
  OR2_X1 U11796 ( .A1(n13553), .A2(n13090), .ZN(n13367) );
  NAND2_X1 U11797 ( .A1(n13366), .A2(n13367), .ZN(n13331) );
  AOI21_X1 U11798 ( .B1(n13334), .B2(n13335), .A(n13331), .ZN(n9045) );
  NAND2_X1 U11799 ( .A1(n9406), .A2(n9405), .ZN(n9291) );
  INV_X1 U11800 ( .A(n13089), .ZN(n13051) );
  NOR2_X1 U11801 ( .A1(n13546), .A2(n13051), .ZN(n9046) );
  INV_X1 U11802 ( .A(n9046), .ZN(n13333) );
  NAND2_X1 U11803 ( .A1(n13333), .A2(n13335), .ZN(n9047) );
  AOI22_X1 U11804 ( .A1(n13543), .A2(n9047), .B1(n9046), .B2(n13088), .ZN(
        n9048) );
  INV_X1 U11805 ( .A(n13031), .ZN(n13087) );
  OR2_X1 U11806 ( .A1(n13538), .A2(n13087), .ZN(n9050) );
  NOR2_X1 U11807 ( .A1(n13532), .A2(n13086), .ZN(n9052) );
  NAND2_X1 U11808 ( .A1(n13532), .A2(n13086), .ZN(n9051) );
  NAND2_X1 U11809 ( .A1(n13452), .A2(n13085), .ZN(n9053) );
  NAND2_X1 U11810 ( .A1(n9054), .A2(n9053), .ZN(n13288) );
  AND2_X1 U11811 ( .A1(n13026), .A2(n13084), .ZN(n9055) );
  OR2_X1 U11812 ( .A1(n13084), .A2(n13026), .ZN(n9056) );
  INV_X1 U11813 ( .A(n12927), .ZN(n13083) );
  NAND2_X1 U11814 ( .A1(n13270), .A2(n13082), .ZN(n9059) );
  NAND2_X1 U11815 ( .A1(n9061), .A2(n9059), .ZN(n9063) );
  INV_X1 U11816 ( .A(n9418), .ZN(n9306) );
  AND2_X1 U11817 ( .A1(n9306), .A2(n9059), .ZN(n9060) );
  INV_X1 U11818 ( .A(n10399), .ZN(n9062) );
  NAND2_X1 U11819 ( .A1(n9308), .A2(n9456), .ZN(n9125) );
  NAND2_X1 U11820 ( .A1(n9064), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U11821 ( .A1(n13231), .A2(n9065), .ZN(n13252) );
  INV_X1 U11822 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U11823 ( .A1(n9279), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U11824 ( .A1(n9268), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9066) );
  OAI211_X1 U11825 ( .C1(n9069), .C2(n9068), .A(n9067), .B(n9066), .ZN(n9070)
         );
  INV_X1 U11826 ( .A(n10403), .ZN(n13080) );
  INV_X1 U11827 ( .A(n12813), .ZN(n10401) );
  INV_X1 U11828 ( .A(n6983), .ZN(n9237) );
  NAND2_X1 U11829 ( .A1(n10401), .A2(n9237), .ZN(n9196) );
  NAND2_X1 U11830 ( .A1(n9168), .A2(n9196), .ZN(n9073) );
  AND2_X2 U11831 ( .A1(n9421), .A2(n9073), .ZN(n13060) );
  AOI22_X1 U11832 ( .A1(n13080), .A2(n13060), .B1(n13059), .B2(n13082), .ZN(
        n12932) );
  OAI21_X1 U11833 ( .B1(n15621), .B2(n9010), .A(n9079), .ZN(n9080) );
  NAND2_X1 U11834 ( .A1(n9080), .A2(n9127), .ZN(n9081) );
  NAND2_X1 U11835 ( .A1(n9081), .A2(n9393), .ZN(n9096) );
  INV_X1 U11836 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9082) );
  INV_X1 U11837 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9084) );
  XNOR2_X1 U11838 ( .A(n12510), .B(P3_B_REG_SCAN_IN), .ZN(n9088) );
  OAI21_X1 U11839 ( .B1(n9100), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9087) );
  INV_X1 U11840 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9086) );
  XNOR2_X1 U11841 ( .A(n9087), .B(n9086), .ZN(n13611) );
  NAND2_X1 U11842 ( .A1(n9088), .A2(n13611), .ZN(n9093) );
  OAI21_X1 U11843 ( .B1(n9090), .B2(n9089), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9091) );
  MUX2_X1 U11844 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9091), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9092) );
  OR2_X1 U11845 ( .A1(n10821), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9095) );
  INV_X1 U11846 ( .A(n9104), .ZN(n13605) );
  NAND2_X1 U11847 ( .A1(n13611), .A2(n13605), .ZN(n9094) );
  NAND2_X1 U11848 ( .A1(n9096), .A2(n11851), .ZN(n9121) );
  NAND2_X1 U11849 ( .A1(n13605), .A2(n12510), .ZN(n9097) );
  XNOR2_X1 U11850 ( .A(n9130), .B(n11851), .ZN(n9117) );
  NAND2_X1 U11851 ( .A1(n9098), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9099) );
  MUX2_X1 U11852 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9099), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n9101) );
  NAND2_X1 U11853 ( .A1(n9101), .A2(n9100), .ZN(n9170) );
  NAND2_X1 U11854 ( .A1(n9170), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13583) );
  INV_X1 U11855 ( .A(n12510), .ZN(n9103) );
  INV_X1 U11856 ( .A(n13611), .ZN(n9102) );
  NOR2_X1 U11857 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .ZN(
        n9108) );
  NOR4_X1 U11858 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n9107) );
  NOR4_X1 U11859 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9106) );
  NOR4_X1 U11860 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9105) );
  NAND4_X1 U11861 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(n9114)
         );
  NOR4_X1 U11862 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9112) );
  NOR4_X1 U11863 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9111) );
  NOR4_X1 U11864 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9110) );
  NOR4_X1 U11865 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9109) );
  NAND4_X1 U11866 ( .A1(n9112), .A2(n9111), .A3(n9110), .A4(n9109), .ZN(n9113)
         );
  NOR2_X1 U11867 ( .A1(n9114), .A2(n9113), .ZN(n9115) );
  OR2_X1 U11868 ( .A1(n10821), .A2(n9115), .ZN(n9129) );
  NAND2_X1 U11869 ( .A1(n11328), .A2(n9129), .ZN(n9116) );
  NOR2_X1 U11870 ( .A1(n9117), .A2(n9116), .ZN(n11854) );
  NAND2_X1 U11871 ( .A1(n9421), .A2(n9127), .ZN(n11852) );
  NAND2_X1 U11872 ( .A1(n9393), .A2(n9118), .ZN(n11856) );
  NAND2_X1 U11873 ( .A1(n11852), .A2(n11856), .ZN(n9119) );
  NAND2_X1 U11874 ( .A1(n9119), .A2(n13582), .ZN(n9120) );
  MUX2_X1 U11875 ( .A(n9122), .B(n9134), .S(n15639), .Z(n9124) );
  INV_X1 U11876 ( .A(n12934), .ZN(n13260) );
  NAND2_X1 U11877 ( .A1(n12934), .A2(n13471), .ZN(n9123) );
  NAND2_X1 U11878 ( .A1(n9124), .A2(n9123), .ZN(P3_U3486) );
  INV_X1 U11879 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n9135) );
  INV_X1 U11880 ( .A(n9125), .ZN(n9126) );
  NAND3_X1 U11881 ( .A1(n9126), .A2(n9010), .A3(n12825), .ZN(n11318) );
  OR2_X1 U11882 ( .A1(n9393), .A2(n9127), .ZN(n11846) );
  NAND2_X1 U11883 ( .A1(n11318), .A2(n11846), .ZN(n9128) );
  NAND2_X1 U11884 ( .A1(n9128), .A2(n11327), .ZN(n9132) );
  NAND2_X1 U11885 ( .A1(n11316), .A2(n11325), .ZN(n9131) );
  NAND2_X1 U11886 ( .A1(n9132), .A2(n9131), .ZN(n9133) );
  MUX2_X1 U11887 ( .A(n9135), .B(n9134), .S(n15631), .Z(n9138) );
  NAND2_X1 U11888 ( .A1(n9138), .A2(n9137), .ZN(P3_U3454) );
  INV_X1 U11889 ( .A(n13583), .ZN(n11306) );
  AND2_X2 U11890 ( .A1(n11306), .A2(n11298), .ZN(P3_U3897) );
  INV_X1 U11891 ( .A(n10897), .ZN(n10696) );
  INV_X1 U11892 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13481) );
  INV_X1 U11893 ( .A(n11236), .ZN(n9204) );
  NOR2_X1 U11894 ( .A1(n12834), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9139) );
  INV_X1 U11895 ( .A(n9140), .ZN(n9141) );
  NOR2_X1 U11896 ( .A1(n11210), .A2(n9141), .ZN(n11184) );
  NAND2_X1 U11897 ( .A1(n11138), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11137) );
  INV_X1 U11898 ( .A(n9143), .ZN(n11224) );
  INV_X1 U11899 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9144) );
  XNOR2_X1 U11900 ( .A(n11236), .B(n9144), .ZN(n11225) );
  INV_X1 U11901 ( .A(n9145), .ZN(n11476) );
  XNOR2_X1 U11902 ( .A(n11488), .B(P3_REG1_REG_6__SCAN_IN), .ZN(n11477) );
  XNOR2_X1 U11903 ( .A(n11460), .B(P3_REG1_REG_8__SCAN_IN), .ZN(n11453) );
  INV_X1 U11904 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U11905 ( .A1(n11457), .A2(n9149), .ZN(n9150) );
  INV_X1 U11906 ( .A(n9150), .ZN(n9152) );
  INV_X1 U11907 ( .A(n11891), .ZN(n9151) );
  XNOR2_X1 U11908 ( .A(n10800), .B(P3_REG1_REG_10__SCAN_IN), .ZN(n10711) );
  INV_X1 U11909 ( .A(n10826), .ZN(n12391) );
  XNOR2_X1 U11910 ( .A(n10869), .B(n12623), .ZN(n13110) );
  NAND2_X1 U11911 ( .A1(n10869), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9156) );
  XNOR2_X1 U11912 ( .A(n10897), .B(n13481), .ZN(n9224) );
  NAND2_X1 U11913 ( .A1(n9158), .A2(n9224), .ZN(n10687) );
  INV_X1 U11914 ( .A(n9227), .ZN(n13160) );
  INV_X1 U11915 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n9229) );
  OR2_X1 U11916 ( .A1(n13182), .A2(n9229), .ZN(n9161) );
  INV_X1 U11917 ( .A(n9232), .ZN(n13194) );
  OAI21_X1 U11918 ( .B1(n9162), .B2(n13194), .A(n13207), .ZN(n9163) );
  INV_X1 U11919 ( .A(n9163), .ZN(n13188) );
  INV_X1 U11920 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13470) );
  INV_X1 U11921 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13467) );
  OR2_X1 U11922 ( .A1(n13211), .A2(n13467), .ZN(n9165) );
  NAND2_X1 U11923 ( .A1(n13211), .A2(n13467), .ZN(n9164) );
  NAND2_X1 U11924 ( .A1(n9165), .A2(n9164), .ZN(n13206) );
  AOI21_X1 U11925 ( .B1(n13208), .B2(n13207), .A(n13206), .ZN(n13205) );
  INV_X1 U11926 ( .A(n9165), .ZN(n9166) );
  XNOR2_X1 U11927 ( .A(n9308), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n9235) );
  INV_X1 U11928 ( .A(n9170), .ZN(n9167) );
  OR2_X1 U11929 ( .A1(n9393), .A2(n9167), .ZN(n9169) );
  NAND2_X1 U11930 ( .A1(n9169), .A2(n9168), .ZN(n9243) );
  NOR2_X1 U11931 ( .A1(n9170), .A2(P3_U3151), .ZN(n9436) );
  OR2_X1 U11932 ( .A1(n11328), .A2(n9436), .ZN(n9242) );
  INV_X1 U11933 ( .A(n9242), .ZN(n9171) );
  NOR2_X1 U11934 ( .A1(n9243), .A2(n9171), .ZN(n9241) );
  INV_X1 U11935 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13425) );
  INV_X1 U11936 ( .A(n10800), .ZN(n9213) );
  INV_X1 U11937 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12050) );
  NOR2_X1 U11938 ( .A1(n11287), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9172) );
  OAI21_X1 U11939 ( .B1(n9173), .B2(n9172), .A(n9174), .ZN(n11215) );
  INV_X1 U11940 ( .A(n9174), .ZN(n9175) );
  NOR2_X1 U11941 ( .A1(n11188), .A2(n11189), .ZN(n11187) );
  INV_X1 U11942 ( .A(n9181), .ZN(n11230) );
  INV_X1 U11943 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n12022) );
  XNOR2_X1 U11944 ( .A(n11236), .B(n12022), .ZN(n11231) );
  INV_X1 U11945 ( .A(n9183), .ZN(n11481) );
  XNOR2_X1 U11946 ( .A(n11488), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n11482) );
  XNOR2_X1 U11947 ( .A(n11460), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U11948 ( .A1(n10703), .A2(n9186), .ZN(n11893) );
  NAND2_X1 U11949 ( .A1(n11895), .A2(n10703), .ZN(n9187) );
  XNOR2_X1 U11950 ( .A(n10800), .B(n15759), .ZN(n10702) );
  XNOR2_X1 U11951 ( .A(n10869), .B(n12629), .ZN(n13116) );
  NAND2_X1 U11952 ( .A1(n9189), .A2(n13146), .ZN(n10689) );
  XNOR2_X1 U11953 ( .A(n10897), .B(n13425), .ZN(n9225) );
  INV_X1 U11954 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12786) );
  XNOR2_X1 U11955 ( .A(n13182), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U11956 ( .A1(n9191), .A2(n13173), .ZN(n13177) );
  INV_X1 U11957 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n9230) );
  OR2_X1 U11958 ( .A1(n13182), .A2(n9230), .ZN(n9192) );
  OR2_X1 U11959 ( .A1(n13211), .A2(n13386), .ZN(n9195) );
  NAND2_X1 U11960 ( .A1(n13211), .A2(n13386), .ZN(n9194) );
  NAND2_X1 U11961 ( .A1(n9195), .A2(n9194), .ZN(n13219) );
  XNOR2_X1 U11962 ( .A(n11176), .B(n13372), .ZN(n9236) );
  INV_X1 U11963 ( .A(n9196), .ZN(n9197) );
  MUX2_X1 U11964 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6983), .Z(n9233) );
  MUX2_X1 U11965 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n6983), .Z(n9226) );
  MUX2_X1 U11966 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6983), .Z(n9223) );
  MUX2_X1 U11967 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6983), .Z(n9219) );
  INV_X1 U11968 ( .A(n9219), .ZN(n9220) );
  NOR2_X1 U11969 ( .A1(n9198), .A2(n10786), .ZN(n11286) );
  INV_X1 U11970 ( .A(n9173), .ZN(n9200) );
  MUX2_X1 U11971 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n13601), .Z(n9201) );
  XOR2_X1 U11972 ( .A(n9176), .B(n9201), .Z(n11182) );
  MUX2_X1 U11973 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13601), .Z(n9202) );
  XNOR2_X1 U11974 ( .A(n9202), .B(n11145), .ZN(n11135) );
  INV_X1 U11975 ( .A(n9202), .ZN(n9203) );
  MUX2_X1 U11976 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13601), .Z(n9205) );
  XOR2_X1 U11977 ( .A(n11236), .B(n9205), .Z(n11223) );
  MUX2_X1 U11978 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13601), .Z(n9206) );
  XNOR2_X1 U11979 ( .A(n9206), .B(n11160), .ZN(n11150) );
  INV_X1 U11980 ( .A(n9206), .ZN(n9207) );
  MUX2_X1 U11981 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n6983), .Z(n9208) );
  XNOR2_X1 U11982 ( .A(n9208), .B(n11488), .ZN(n11474) );
  MUX2_X1 U11983 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n6983), .Z(n9209) );
  XNOR2_X1 U11984 ( .A(n9209), .B(n11388), .ZN(n11382) );
  INV_X1 U11985 ( .A(n9209), .ZN(n9210) );
  MUX2_X1 U11986 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n6983), .Z(n9211) );
  XOR2_X1 U11987 ( .A(n11460), .B(n9211), .Z(n11447) );
  INV_X1 U11988 ( .A(n11460), .ZN(n10788) );
  MUX2_X1 U11989 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n6983), .Z(n9212) );
  NAND2_X1 U11990 ( .A1(n11891), .A2(n9212), .ZN(n11885) );
  OR2_X1 U11991 ( .A1(n9212), .A2(n11891), .ZN(n11887) );
  INV_X1 U11992 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12335) );
  MUX2_X1 U11993 ( .A(n15759), .B(n12335), .S(n6983), .Z(n9214) );
  NAND2_X1 U11994 ( .A1(n9214), .A2(n9213), .ZN(n9217) );
  INV_X1 U11995 ( .A(n9214), .ZN(n9215) );
  NAND2_X1 U11996 ( .A1(n9215), .A2(n10800), .ZN(n9216) );
  NAND2_X1 U11997 ( .A1(n9217), .A2(n9216), .ZN(n10708) );
  INV_X1 U11998 ( .A(n9217), .ZN(n9218) );
  XNOR2_X1 U11999 ( .A(n9219), .B(n10826), .ZN(n12386) );
  MUX2_X1 U12000 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6983), .Z(n9221) );
  XNOR2_X1 U12001 ( .A(n9221), .B(n13124), .ZN(n13125) );
  NAND2_X1 U12002 ( .A1(n9221), .A2(n10869), .ZN(n13138) );
  INV_X1 U12003 ( .A(n13146), .ZN(n9222) );
  XNOR2_X1 U12004 ( .A(n9223), .B(n9222), .ZN(n13137) );
  INV_X1 U12005 ( .A(n9224), .ZN(n10685) );
  INV_X1 U12006 ( .A(n9225), .ZN(n10690) );
  MUX2_X1 U12007 ( .A(n10685), .B(n10690), .S(n9237), .Z(n10694) );
  MUX2_X1 U12008 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6983), .Z(n13155) );
  MUX2_X1 U12009 ( .A(n9230), .B(n9229), .S(n6983), .Z(n9231) );
  NOR2_X1 U12010 ( .A1(n9231), .A2(n13182), .ZN(n13167) );
  XOR2_X1 U12011 ( .A(n9233), .B(n9232), .Z(n13191) );
  NOR2_X1 U12012 ( .A1(n13190), .A2(n13191), .ZN(n13189) );
  XNOR2_X1 U12013 ( .A(n9234), .B(n13211), .ZN(n13203) );
  MUX2_X1 U12014 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6983), .Z(n13204) );
  INV_X1 U12015 ( .A(n9235), .ZN(n9239) );
  INV_X1 U12016 ( .A(n9236), .ZN(n9238) );
  MUX2_X1 U12017 ( .A(n9239), .B(n9238), .S(n9237), .Z(n9240) );
  AND2_X1 U12018 ( .A1(P3_U3897), .A2(n12813), .ZN(n13140) );
  MUX2_X1 U12019 ( .A(P3_U3897), .B(n9241), .S(n12813), .Z(n13212) );
  NAND2_X1 U12020 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12965)
         );
  OAI21_X1 U12021 ( .B1(n13215), .B2(n15465), .A(n12965), .ZN(n9244) );
  AOI21_X1 U12022 ( .B1(n9308), .B2(n13212), .A(n9244), .ZN(n9245) );
  INV_X1 U12023 ( .A(n9247), .ZN(n9248) );
  INV_X1 U12024 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U12025 ( .A1(n9249), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9250) );
  INV_X1 U12026 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12883) );
  INV_X1 U12027 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14681) );
  NAND2_X1 U12028 ( .A1(n14681), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9252) );
  XNOR2_X1 U12029 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n9274) );
  INV_X1 U12030 ( .A(n9274), .ZN(n9253) );
  INV_X1 U12031 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12863) );
  INV_X1 U12032 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14675) );
  XNOR2_X1 U12033 ( .A(n14675), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n9264) );
  INV_X1 U12034 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12897) );
  XNOR2_X1 U12035 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n9254) );
  XNOR2_X1 U12036 ( .A(n9255), .B(n9254), .ZN(n13586) );
  NAND2_X1 U12037 ( .A1(n13586), .A2(n9287), .ZN(n9257) );
  INV_X1 U12038 ( .A(SI_31_), .ZN(n13592) );
  OR2_X1 U12039 ( .A1(n9288), .A2(n13592), .ZN(n9256) );
  INV_X1 U12040 ( .A(n13231), .ZN(n9259) );
  INV_X1 U12041 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13233) );
  NAND2_X1 U12042 ( .A1(n9279), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9261) );
  INV_X1 U12043 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13434) );
  OR2_X1 U12044 ( .A1(n8577), .A2(n13434), .ZN(n9260) );
  OAI211_X1 U12045 ( .C1(n13233), .C2(n9068), .A(n9261), .B(n9260), .ZN(n9262)
         );
  INV_X1 U12046 ( .A(n9262), .ZN(n9263) );
  XNOR2_X1 U12047 ( .A(n9265), .B(n9264), .ZN(n12808) );
  NAND2_X1 U12048 ( .A1(n12808), .A2(n9287), .ZN(n9267) );
  INV_X1 U12049 ( .A(SI_30_), .ZN(n12810) );
  OR2_X1 U12050 ( .A1(n9288), .A2(n12810), .ZN(n9266) );
  INV_X1 U12051 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n15744) );
  NAND2_X1 U12052 ( .A1(n9268), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U12053 ( .A1(n9279), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9269) );
  OAI211_X1 U12054 ( .C1(n15744), .C2(n9068), .A(n9270), .B(n9269), .ZN(n9271)
         );
  INV_X1 U12055 ( .A(n9271), .ZN(n9272) );
  NAND2_X1 U12056 ( .A1(n13234), .A2(n12348), .ZN(n9273) );
  XNOR2_X1 U12057 ( .A(n9275), .B(n9274), .ZN(n13593) );
  NAND2_X1 U12058 ( .A1(n13593), .A2(n9287), .ZN(n9277) );
  INV_X1 U12059 ( .A(SI_29_), .ZN(n13596) );
  OR2_X1 U12060 ( .A1(n9288), .A2(n13596), .ZN(n9276) );
  INV_X1 U12061 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n12887) );
  NAND2_X1 U12062 ( .A1(n9278), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U12063 ( .A1(n9279), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9280) );
  OAI211_X1 U12064 ( .C1(n12887), .C2(n8577), .A(n9281), .B(n9280), .ZN(n9282)
         );
  INV_X1 U12065 ( .A(n9282), .ZN(n9283) );
  XNOR2_X1 U12066 ( .A(n14681), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9285) );
  XNOR2_X1 U12067 ( .A(n9286), .B(n9285), .ZN(n12811) );
  NAND2_X1 U12068 ( .A1(n12811), .A2(n9287), .ZN(n9290) );
  INV_X1 U12069 ( .A(SI_28_), .ZN(n15760) );
  OR2_X1 U12070 ( .A1(n9288), .A2(n15760), .ZN(n9289) );
  NAND2_X1 U12071 ( .A1(n13253), .A2(n10403), .ZN(n9426) );
  NAND2_X1 U12072 ( .A1(n13299), .A2(n9408), .ZN(n13316) );
  INV_X1 U12073 ( .A(n13366), .ZN(n9302) );
  NOR2_X1 U12074 ( .A1(n13496), .A2(n11671), .ZN(n9294) );
  INV_X1 U12075 ( .A(n9316), .ZN(n9293) );
  NOR2_X1 U12076 ( .A1(n13495), .A2(n9293), .ZN(n11848) );
  NAND4_X1 U12077 ( .A1(n9294), .A2(n12134), .A3(n11848), .A4(n12030), .ZN(
        n9295) );
  NOR3_X1 U12078 ( .A1(n9295), .A2(n12058), .A3(n12018), .ZN(n9296) );
  NAND3_X1 U12079 ( .A1(n9296), .A2(n12043), .A3(n9347), .ZN(n9297) );
  NOR4_X1 U12080 ( .A1(n12523), .A2(n9297), .A3(n12331), .A4(n9032), .ZN(n9298) );
  NAND4_X1 U12081 ( .A1(n13405), .A2(n12617), .A3(n9298), .A4(n9378), .ZN(
        n9300) );
  OR2_X1 U12082 ( .A1(n9374), .A2(n7706), .ZN(n9369) );
  NOR3_X1 U12083 ( .A1(n9300), .A2(n13417), .A3(n9369), .ZN(n9301) );
  NOR2_X1 U12084 ( .A1(n13382), .A2(n13395), .ZN(n9397) );
  NAND4_X1 U12085 ( .A1(n13338), .A2(n9302), .A3(n9301), .A4(n9397), .ZN(n9303) );
  XNOR2_X1 U12086 ( .A(n13334), .B(n13088), .ZN(n13350) );
  NOR4_X1 U12087 ( .A1(n9412), .A2(n13316), .A3(n9303), .A4(n13350), .ZN(n9304) );
  NAND4_X1 U12088 ( .A1(n13266), .A2(n13282), .A3(n9304), .A4(n7010), .ZN(
        n9305) );
  NAND4_X1 U12089 ( .A1(n9435), .A2(n9307), .A3(n9448), .A4(n9433), .ZN(n9309)
         );
  NAND2_X1 U12090 ( .A1(n9443), .A2(n9421), .ZN(n9425) );
  INV_X1 U12091 ( .A(n13250), .ZN(n9424) );
  MUX2_X1 U12092 ( .A(n9311), .B(n9310), .S(n9421), .Z(n9312) );
  NAND2_X1 U12093 ( .A1(n13266), .A2(n9312), .ZN(n9420) );
  INV_X1 U12094 ( .A(n13026), .ZN(n13525) );
  AOI22_X1 U12095 ( .A1(n9313), .A2(n9315), .B1(n13525), .B2(n13084), .ZN(
        n9314) );
  MUX2_X1 U12096 ( .A(n9315), .B(n9314), .S(n9393), .Z(n9414) );
  OAI21_X1 U12097 ( .B1(n13495), .B2(n6432), .A(n9316), .ZN(n9317) );
  MUX2_X1 U12098 ( .A(n6571), .B(n9317), .S(n9393), .Z(n9318) );
  AOI21_X1 U12099 ( .B1(n9318), .B2(n11309), .A(n11671), .ZN(n9325) );
  AOI21_X1 U12100 ( .B1(n9329), .B2(n9319), .A(n9393), .ZN(n9324) );
  INV_X1 U12101 ( .A(n11309), .ZN(n9320) );
  NAND3_X1 U12102 ( .A1(n9320), .A2(n9329), .A3(n9319), .ZN(n9321) );
  MUX2_X1 U12103 ( .A(n9322), .B(n9321), .S(n9421), .Z(n9323) );
  OAI211_X1 U12104 ( .C1(n9325), .C2(n9324), .A(n9326), .B(n9323), .ZN(n9332)
         );
  NAND2_X1 U12105 ( .A1(n9326), .A2(n12027), .ZN(n9327) );
  NAND2_X1 U12106 ( .A1(n9327), .A2(n9393), .ZN(n9331) );
  OAI21_X1 U12107 ( .B1(n9421), .B2(n9329), .A(n9328), .ZN(n9330) );
  AOI21_X1 U12108 ( .B1(n9332), .B2(n9331), .A(n9330), .ZN(n9333) );
  INV_X1 U12109 ( .A(n12134), .ZN(n12131) );
  OR2_X1 U12110 ( .A1(n9333), .A2(n12131), .ZN(n9342) );
  NAND2_X1 U12111 ( .A1(n9345), .A2(n9334), .ZN(n9336) );
  NAND2_X1 U12112 ( .A1(n9336), .A2(n9393), .ZN(n9341) );
  NOR2_X1 U12113 ( .A1(n9336), .A2(n9335), .ZN(n9339) );
  AND2_X1 U12114 ( .A1(n13104), .A2(n9337), .ZN(n9338) );
  MUX2_X1 U12115 ( .A(n9339), .B(n9338), .S(n9421), .Z(n9340) );
  AOI21_X1 U12116 ( .B1(n9342), .B2(n9341), .A(n9340), .ZN(n9349) );
  AOI21_X1 U12117 ( .B1(n9344), .B2(n9343), .A(n9393), .ZN(n9348) );
  MUX2_X1 U12118 ( .A(n9345), .B(n9344), .S(n9393), .Z(n9346) );
  OAI211_X1 U12119 ( .C1(n9349), .C2(n9348), .A(n9347), .B(n9346), .ZN(n9353)
         );
  NAND2_X1 U12120 ( .A1(n13101), .A2(n12110), .ZN(n9351) );
  MUX2_X1 U12121 ( .A(n9351), .B(n9350), .S(n9421), .Z(n9352) );
  MUX2_X1 U12122 ( .A(n9355), .B(n9354), .S(n9393), .Z(n9356) );
  MUX2_X1 U12123 ( .A(n9359), .B(n7719), .S(n9393), .Z(n9360) );
  MUX2_X1 U12124 ( .A(n9362), .B(n9361), .S(n9421), .Z(n9363) );
  AND2_X1 U12125 ( .A1(n9371), .A2(n9364), .ZN(n9367) );
  AND2_X1 U12126 ( .A1(n9370), .A2(n9365), .ZN(n9366) );
  MUX2_X1 U12127 ( .A(n9367), .B(n9366), .S(n9421), .Z(n9368) );
  MUX2_X1 U12128 ( .A(n9371), .B(n9370), .S(n9393), .Z(n9372) );
  INV_X1 U12129 ( .A(n13417), .ZN(n13421) );
  MUX2_X1 U12130 ( .A(n9374), .B(n7706), .S(n9421), .Z(n9375) );
  INV_X1 U12131 ( .A(n9375), .ZN(n9376) );
  INV_X1 U12132 ( .A(n9378), .ZN(n12782) );
  OR2_X1 U12133 ( .A1(n13477), .A2(n9379), .ZN(n9380) );
  OAI211_X1 U12134 ( .C1(n12782), .C2(n9382), .A(n9381), .B(n9380), .ZN(n9383)
         );
  NAND2_X1 U12135 ( .A1(n9383), .A2(n9393), .ZN(n9384) );
  AOI21_X1 U12136 ( .B1(n13391), .B2(n9385), .A(n9393), .ZN(n9387) );
  OR2_X1 U12137 ( .A1(n13008), .A2(n9393), .ZN(n9386) );
  OAI22_X1 U12138 ( .A1(n9388), .A2(n9387), .B1(n13414), .B2(n9386), .ZN(n9398) );
  INV_X1 U12139 ( .A(n9391), .ZN(n9390) );
  OAI211_X1 U12140 ( .C1(n9390), .C2(n9389), .A(n9400), .B(n13325), .ZN(n9395)
         );
  OAI211_X1 U12141 ( .C1(n13382), .C2(n9392), .A(n9399), .B(n9391), .ZN(n9394)
         );
  MUX2_X1 U12142 ( .A(n9395), .B(n9394), .S(n9393), .Z(n9396) );
  AOI21_X1 U12143 ( .B1(n9398), .B2(n9397), .A(n9396), .ZN(n9402) );
  MUX2_X1 U12144 ( .A(n9400), .B(n9399), .S(n9421), .Z(n9401) );
  OR2_X1 U12145 ( .A1(n13334), .A2(n13088), .ZN(n9403) );
  MUX2_X1 U12146 ( .A(n9403), .B(n13327), .S(n9421), .Z(n9404) );
  MUX2_X1 U12147 ( .A(n9408), .B(n13299), .S(n9421), .Z(n9409) );
  NAND3_X1 U12148 ( .A1(n13452), .A2(n12942), .A3(n9421), .ZN(n9410) );
  MUX2_X1 U12149 ( .A(n9416), .B(n9415), .S(n9421), .Z(n9417) );
  OAI211_X1 U12150 ( .C1(n9420), .C2(n9419), .A(n9418), .B(n9417), .ZN(n9423)
         );
  OR3_X1 U12151 ( .A1(n12934), .A2(n12976), .A3(n9421), .ZN(n9422) );
  INV_X1 U12152 ( .A(n9425), .ZN(n9430) );
  AND2_X1 U12153 ( .A1(n9426), .A2(n13249), .ZN(n9441) );
  NOR2_X1 U12154 ( .A1(n9441), .A2(n9440), .ZN(n9429) );
  INV_X1 U12155 ( .A(n9444), .ZN(n9428) );
  AOI21_X1 U12156 ( .B1(n9430), .B2(n9429), .A(n9428), .ZN(n9431) );
  NAND2_X1 U12157 ( .A1(n9432), .A2(n9448), .ZN(n9434) );
  INV_X1 U12158 ( .A(n9436), .ZN(n12227) );
  NOR2_X1 U12159 ( .A1(n12227), .A2(n11176), .ZN(n9454) );
  AND2_X1 U12160 ( .A1(n9436), .A2(n11176), .ZN(n9462) );
  INV_X1 U12161 ( .A(n9462), .ZN(n9437) );
  NOR2_X1 U12162 ( .A1(n9437), .A2(n9010), .ZN(n9438) );
  NAND2_X1 U12163 ( .A1(n10409), .A2(n9443), .ZN(n9447) );
  INV_X1 U12164 ( .A(n13230), .ZN(n12468) );
  NAND2_X1 U12165 ( .A1(n9447), .A2(n9446), .ZN(n9453) );
  INV_X1 U12166 ( .A(n13228), .ZN(n13505) );
  NAND2_X1 U12167 ( .A1(n9455), .A2(n11328), .ZN(n11324) );
  NOR2_X1 U12168 ( .A1(n11324), .A2(n12813), .ZN(n9458) );
  OAI21_X1 U12169 ( .B1(n12227), .B2(n9456), .A(P3_B_REG_SCAN_IN), .ZN(n9457)
         );
  AOI21_X1 U12170 ( .B1(n9458), .B2(n13059), .A(n9457), .ZN(n9459) );
  INV_X1 U12171 ( .A(n9459), .ZN(n9460) );
  NAND3_X1 U12172 ( .A1(n6432), .A2(n9010), .A3(n9462), .ZN(n9463) );
  NOR2_X1 U12173 ( .A1(n9464), .A2(n9463), .ZN(n9465) );
  NOR2_X1 U12174 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n9469) );
  NAND4_X1 U12175 ( .A1(n9675), .A2(n9676), .A3(n9674), .A4(n9469), .ZN(n9472)
         );
  NAND4_X1 U12176 ( .A1(n9470), .A2(n9623), .A3(n9551), .A4(n9565), .ZN(n9471)
         );
  NAND2_X1 U12177 ( .A1(n9865), .A2(n9474), .ZN(n9868) );
  INV_X1 U12178 ( .A(n9868), .ZN(n9477) );
  INV_X1 U12179 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9481) );
  INV_X1 U12180 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9482) );
  AND2_X2 U12181 ( .A1(n9487), .A2(n9485), .ZN(n9527) );
  NAND2_X1 U12182 ( .A1(n10254), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9492) );
  INV_X1 U12183 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n15727) );
  NAND2_X4 U12184 ( .A1(n9486), .A2(n15401), .ZN(n10255) );
  INV_X1 U12185 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11993) );
  INV_X1 U12186 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9488) );
  OR2_X1 U12187 ( .A1(n9528), .A2(n9488), .ZN(n9489) );
  XNOR2_X2 U12188 ( .A(n9494), .B(n9493), .ZN(n12885) );
  AND2_X4 U12189 ( .A1(n9516), .A2(n7007), .ZN(n10318) );
  NAND2_X2 U12190 ( .A1(n9516), .A2(n10801), .ZN(n9695) );
  INV_X1 U12191 ( .A(n10929), .ZN(n10924) );
  NAND2_X1 U12192 ( .A1(n9534), .A2(n10924), .ZN(n9503) );
  INV_X1 U12193 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9508) );
  OR2_X1 U12194 ( .A1(n9519), .A2(n9508), .ZN(n9511) );
  INV_X1 U12195 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9509) );
  AND2_X1 U12196 ( .A1(n9511), .A2(n9510), .ZN(n9514) );
  INV_X1 U12197 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10845) );
  OR2_X1 U12198 ( .A1(n9915), .A2(n10845), .ZN(n9513) );
  NAND2_X1 U12199 ( .A1(n9782), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9512) );
  NAND3_X2 U12200 ( .A1(n9514), .A2(n9513), .A3(n9512), .ZN(n10460) );
  INV_X1 U12201 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n11244) );
  NOR2_X1 U12202 ( .A1(n10801), .A2(n10784), .ZN(n9515) );
  XNOR2_X1 U12203 ( .A(n9515), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15404) );
  NAND2_X1 U12204 ( .A1(n10460), .A2(n11203), .ZN(n11164) );
  INV_X1 U12205 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9518) );
  INV_X1 U12206 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n12146) );
  OR2_X1 U12207 ( .A1(n9519), .A2(n12146), .ZN(n9523) );
  INV_X1 U12208 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10925) );
  INV_X1 U12209 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9520) );
  OR2_X1 U12210 ( .A1(n9528), .A2(n9520), .ZN(n9521) );
  NAND2_X1 U12211 ( .A1(n10254), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9533) );
  OR2_X1 U12212 ( .A1(n9519), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9532) );
  INV_X1 U12213 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n12124) );
  OR2_X1 U12214 ( .A1(n10255), .A2(n12124), .ZN(n9531) );
  INV_X1 U12215 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9529) );
  OR2_X1 U12216 ( .A1(n9528), .A2(n9529), .ZN(n9530) );
  NAND4_X1 U12217 ( .A1(n9533), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(n14852) );
  NAND2_X1 U12218 ( .A1(n10318), .A2(n10823), .ZN(n9540) );
  NAND2_X1 U12219 ( .A1(n9534), .A2(n10931), .ZN(n9538) );
  NAND2_X1 U12220 ( .A1(n14852), .A2(n10469), .ZN(n10146) );
  OR2_X1 U12221 ( .A1(n14852), .A2(n7106), .ZN(n9541) );
  INV_X1 U12222 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9542) );
  INV_X1 U12223 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11970) );
  OR2_X1 U12224 ( .A1(n10255), .A2(n11970), .ZN(n9546) );
  OAI21_X1 U12225 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n9556), .ZN(n11971) );
  OR2_X1 U12226 ( .A1(n9519), .A2(n11971), .ZN(n9545) );
  INV_X1 U12227 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9543) );
  OR2_X1 U12228 ( .A1(n9915), .A2(n9543), .ZN(n9544) );
  NAND4_X2 U12229 ( .A1(n9547), .A2(n9546), .A3(n9545), .A4(n9544), .ZN(n14851) );
  OR2_X1 U12230 ( .A1(n9536), .A2(n9863), .ZN(n9548) );
  AOI22_X1 U12231 ( .A1(n10319), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9534), 
        .B2(n14868), .ZN(n9550) );
  NAND2_X1 U12232 ( .A1(n10795), .A2(n10318), .ZN(n9549) );
  XNOR2_X1 U12233 ( .A(n14851), .B(n11276), .ZN(n11280) );
  INV_X1 U12234 ( .A(n11280), .ZN(n11274) );
  OR2_X1 U12235 ( .A1(n14851), .A2(n11276), .ZN(n11797) );
  NAND2_X1 U12236 ( .A1(n10840), .A2(n10318), .ZN(n9554) );
  NAND2_X1 U12237 ( .A1(n9536), .A2(n9551), .ZN(n9562) );
  NAND2_X1 U12238 ( .A1(n9562), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9552) );
  XNOR2_X1 U12239 ( .A(n9552), .B(P1_IR_REG_5__SCAN_IN), .ZN(n14879) );
  AOI22_X1 U12240 ( .A1(n6431), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9534), .B2(
        n14879), .ZN(n9553) );
  INV_X1 U12241 ( .A(n11952), .ZN(n15496) );
  INV_X1 U12242 ( .A(n9528), .ZN(n9612) );
  NAND2_X1 U12243 ( .A1(n9612), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9561) );
  INV_X1 U12244 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11948) );
  OR2_X1 U12245 ( .A1(n10255), .A2(n11948), .ZN(n9560) );
  INV_X1 U12246 ( .A(n9570), .ZN(n9572) );
  NAND2_X1 U12247 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  NAND2_X1 U12248 ( .A1(n9572), .A2(n9557), .ZN(n11951) );
  OR2_X1 U12249 ( .A1(n9519), .A2(n11951), .ZN(n9559) );
  INV_X1 U12250 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10926) );
  OR2_X1 U12251 ( .A1(n9915), .A2(n10926), .ZN(n9558) );
  OR2_X1 U12252 ( .A1(n15496), .A2(n14850), .ZN(n11799) );
  NAND3_X1 U12253 ( .A1(n11798), .A2(n11797), .A3(n11799), .ZN(n9582) );
  NAND2_X1 U12254 ( .A1(n10838), .A2(n10318), .ZN(n9569) );
  NAND2_X1 U12255 ( .A1(n9564), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9563) );
  MUX2_X1 U12256 ( .A(n9563), .B(P1_IR_REG_31__SCAN_IN), .S(n9565), .Z(n9567)
         );
  NAND2_X1 U12257 ( .A1(n9567), .A2(n9594), .ZN(n10939) );
  AOI22_X1 U12258 ( .A1(n6431), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9534), .B2(
        n10983), .ZN(n9568) );
  AND2_X2 U12259 ( .A1(n9569), .A2(n9568), .ZN(n11922) );
  INV_X1 U12260 ( .A(n11922), .ZN(n11424) );
  NAND2_X1 U12261 ( .A1(n9612), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9578) );
  INV_X1 U12262 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11907) );
  OR2_X1 U12263 ( .A1(n10255), .A2(n11907), .ZN(n9577) );
  INV_X1 U12264 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9571) );
  NAND2_X1 U12265 ( .A1(n9572), .A2(n9571), .ZN(n9573) );
  NAND2_X1 U12266 ( .A1(n9585), .A2(n9573), .ZN(n11910) );
  OR2_X1 U12267 ( .A1(n9519), .A2(n11910), .ZN(n9576) );
  INV_X1 U12268 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9574) );
  OR2_X1 U12269 ( .A1(n9915), .A2(n9574), .ZN(n9575) );
  NAND4_X4 U12270 ( .A1(n9578), .A2(n9577), .A3(n9576), .A4(n9575), .ZN(n14849) );
  XNOR2_X1 U12271 ( .A(n11424), .B(n11938), .ZN(n10337) );
  NAND2_X1 U12272 ( .A1(n9582), .A2(n9581), .ZN(n11917) );
  OR2_X1 U12273 ( .A1(n11424), .A2(n14849), .ZN(n11916) );
  NAND2_X1 U12274 ( .A1(n9594), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9625) );
  XNOR2_X1 U12275 ( .A(n9625), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U12276 ( .A1(n6431), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9534), .B2(
        n11262), .ZN(n9583) );
  NAND2_X1 U12277 ( .A1(n9612), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9590) );
  INV_X1 U12278 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11928) );
  OR2_X1 U12279 ( .A1(n10255), .A2(n11928), .ZN(n9589) );
  NAND2_X1 U12280 ( .A1(n9585), .A2(n9584), .ZN(n9586) );
  NAND2_X1 U12281 ( .A1(n9600), .A2(n9586), .ZN(n11931) );
  OR2_X1 U12282 ( .A1(n9519), .A2(n11931), .ZN(n9588) );
  INV_X1 U12283 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10980) );
  OR2_X1 U12284 ( .A1(n9915), .A2(n10980), .ZN(n9587) );
  NAND4_X1 U12285 ( .A1(n9590), .A2(n9589), .A3(n9588), .A4(n9587), .ZN(n14848) );
  OR2_X1 U12286 ( .A1(n15503), .A2(n14848), .ZN(n9591) );
  AND2_X1 U12287 ( .A1(n11916), .A2(n9591), .ZN(n9593) );
  INV_X1 U12288 ( .A(n9591), .ZN(n9592) );
  XNOR2_X1 U12289 ( .A(n15503), .B(n14848), .ZN(n10339) );
  INV_X1 U12290 ( .A(n10339), .ZN(n11920) );
  NAND2_X1 U12291 ( .A1(n10870), .A2(n10318), .ZN(n9598) );
  NAND2_X1 U12292 ( .A1(n9678), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9595) );
  INV_X1 U12293 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U12294 ( .A1(n9595), .A2(n9622), .ZN(n9608) );
  OR2_X1 U12295 ( .A1(n9595), .A2(n9622), .ZN(n9596) );
  AOI22_X1 U12296 ( .A1(n6431), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9534), .B2(
        n14901), .ZN(n9597) );
  NAND2_X1 U12297 ( .A1(n9782), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9606) );
  OR2_X1 U12298 ( .A1(n9915), .A2(n7435), .ZN(n9605) );
  NAND2_X1 U12299 ( .A1(n9600), .A2(n9599), .ZN(n9601) );
  NAND2_X1 U12300 ( .A1(n9614), .A2(n9601), .ZN(n11962) );
  OR2_X1 U12301 ( .A1(n9519), .A2(n11962), .ZN(n9604) );
  INV_X1 U12302 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9602) );
  OR2_X1 U12303 ( .A1(n9528), .A2(n9602), .ZN(n9603) );
  XNOR2_X1 U12304 ( .A(n11961), .B(n12075), .ZN(n11733) );
  INV_X1 U12305 ( .A(n12075), .ZN(n14847) );
  OR2_X1 U12306 ( .A1(n11961), .A2(n14847), .ZN(n9607) );
  NAND2_X1 U12307 ( .A1(n9608), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9609) );
  XNOR2_X1 U12308 ( .A(n9609), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U12309 ( .A1(n11266), .A2(n9534), .B1(n6431), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U12310 ( .A1(n9912), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9619) );
  INV_X1 U12311 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n12082) );
  OR2_X1 U12312 ( .A1(n10255), .A2(n12082), .ZN(n9618) );
  NAND2_X1 U12313 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  NAND2_X1 U12314 ( .A1(n9630), .A2(n9615), .ZN(n12102) );
  OR2_X1 U12315 ( .A1(n9519), .A2(n12102), .ZN(n9617) );
  INV_X1 U12316 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15666) );
  OR2_X1 U12317 ( .A1(n9915), .A2(n15666), .ZN(n9616) );
  XNOR2_X1 U12318 ( .A(n12217), .B(n12162), .ZN(n12074) );
  INV_X1 U12319 ( .A(n12162), .ZN(n14846) );
  OR2_X1 U12320 ( .A1(n12217), .A2(n14846), .ZN(n9620) );
  NAND2_X1 U12321 ( .A1(n12069), .A2(n9620), .ZN(n12156) );
  NAND2_X1 U12322 ( .A1(n10916), .A2(n10318), .ZN(n9628) );
  INV_X1 U12323 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9621) );
  AND3_X1 U12324 ( .A1(n9623), .A2(n9622), .A3(n9621), .ZN(n9624) );
  NAND2_X1 U12325 ( .A1(n9625), .A2(n9624), .ZN(n9636) );
  NAND2_X1 U12326 ( .A1(n9636), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9626) );
  XNOR2_X1 U12327 ( .A(n9626), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U12328 ( .A1(n6431), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11620), 
        .B2(n9534), .ZN(n9627) );
  NAND2_X1 U12329 ( .A1(n9912), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9635) );
  INV_X1 U12330 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12204) );
  OR2_X1 U12331 ( .A1(n10255), .A2(n12204), .ZN(n9634) );
  INV_X1 U12332 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U12333 ( .A1(n9630), .A2(n9629), .ZN(n9631) );
  NAND2_X1 U12334 ( .A1(n9640), .A2(n9631), .ZN(n12197) );
  OR2_X1 U12335 ( .A1(n9519), .A2(n12197), .ZN(n9633) );
  INV_X1 U12336 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11614) );
  OR2_X1 U12337 ( .A1(n9915), .A2(n11614), .ZN(n9632) );
  NAND4_X1 U12338 ( .A1(n9635), .A2(n9634), .A3(n9633), .A4(n9632), .ZN(n14845) );
  XNOR2_X1 U12339 ( .A(n12166), .B(n14845), .ZN(n12160) );
  INV_X1 U12340 ( .A(n12160), .ZN(n12157) );
  NAND2_X1 U12341 ( .A1(n10943), .A2(n10318), .ZN(n9639) );
  NAND2_X1 U12342 ( .A1(n9649), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9637) );
  XNOR2_X1 U12343 ( .A(n9637), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U12344 ( .A1(n11826), .A2(n9534), .B1(n6431), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U12345 ( .A1(n9912), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9645) );
  INV_X1 U12346 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n12235) );
  OR2_X1 U12347 ( .A1(n10255), .A2(n12235), .ZN(n9644) );
  NAND2_X1 U12348 ( .A1(n9640), .A2(n15650), .ZN(n9641) );
  NAND2_X1 U12349 ( .A1(n9654), .A2(n9641), .ZN(n12516) );
  OR2_X1 U12350 ( .A1(n9519), .A2(n12516), .ZN(n9643) );
  INV_X1 U12351 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11823) );
  OR2_X1 U12352 ( .A1(n9915), .A2(n11823), .ZN(n9642) );
  NAND4_X1 U12353 ( .A1(n9645), .A2(n9644), .A3(n9643), .A4(n9642), .ZN(n14844) );
  XNOR2_X1 U12354 ( .A(n15349), .B(n14844), .ZN(n10342) );
  INV_X1 U12355 ( .A(n10342), .ZN(n12243) );
  AND2_X1 U12356 ( .A1(n12157), .A2(n12243), .ZN(n9646) );
  OR2_X1 U12357 ( .A1(n15349), .A2(n14844), .ZN(n9647) );
  OR2_X1 U12358 ( .A1(n12166), .A2(n14845), .ZN(n12238) );
  OR2_X1 U12359 ( .A1(n10342), .A2(n12238), .ZN(n12240) );
  NAND2_X1 U12360 ( .A1(n11064), .A2(n10318), .ZN(n9652) );
  NAND2_X1 U12361 ( .A1(n9650), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9661) );
  XNOR2_X1 U12362 ( .A(n9661), .B(P1_IR_REG_12__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U12363 ( .A1(n12283), .A2(n9534), .B1(n6431), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U12364 ( .A1(n9912), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9659) );
  INV_X1 U12365 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12323) );
  OR2_X1 U12366 ( .A1(n10255), .A2(n12323), .ZN(n9658) );
  INV_X1 U12367 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U12368 ( .A1(n9654), .A2(n9653), .ZN(n9655) );
  NAND2_X1 U12369 ( .A1(n9666), .A2(n9655), .ZN(n12700) );
  OR2_X1 U12370 ( .A1(n9519), .A2(n12700), .ZN(n9657) );
  INV_X1 U12371 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n12601) );
  OR2_X1 U12372 ( .A1(n9915), .A2(n12601), .ZN(n9656) );
  NAND4_X1 U12373 ( .A1(n9659), .A2(n9658), .A3(n9657), .A4(n9656), .ZN(n14843) );
  XNOR2_X1 U12374 ( .A(n12322), .B(n14843), .ZN(n12317) );
  INV_X1 U12375 ( .A(n12317), .ZN(n12314) );
  NAND2_X1 U12376 ( .A1(n11089), .A2(n10318), .ZN(n9664) );
  INV_X1 U12377 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9660) );
  NAND2_X1 U12378 ( .A1(n9661), .A2(n9660), .ZN(n9662) );
  NAND2_X1 U12379 ( .A1(n9662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9692) );
  XNOR2_X1 U12380 ( .A(n9692), .B(P1_IR_REG_13__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U12381 ( .A1(n12432), .A2(n9534), .B1(n6431), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9663) );
  INV_X1 U12382 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U12383 ( .A1(n9666), .A2(n9665), .ZN(n9667) );
  NAND2_X1 U12384 ( .A1(n9699), .A2(n9667), .ZN(n12544) );
  OR2_X1 U12385 ( .A1(n12544), .A2(n9519), .ZN(n9672) );
  INV_X1 U12386 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15772) );
  OR2_X1 U12387 ( .A1(n9528), .A2(n15772), .ZN(n9671) );
  INV_X1 U12388 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9668) );
  OR2_X1 U12389 ( .A1(n10255), .A2(n9668), .ZN(n9670) );
  INV_X1 U12390 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n12667) );
  OR2_X1 U12391 ( .A1(n9915), .A2(n12667), .ZN(n9669) );
  NAND4_X1 U12392 ( .A1(n9672), .A2(n9671), .A3(n9670), .A4(n9669), .ZN(n14842) );
  XNOR2_X1 U12393 ( .A(n12552), .B(n14842), .ZN(n12546) );
  INV_X1 U12394 ( .A(n12546), .ZN(n12550) );
  NAND2_X1 U12395 ( .A1(n12551), .A2(n12550), .ZN(n12549) );
  OR2_X1 U12396 ( .A1(n12552), .A2(n14842), .ZN(n9673) );
  INV_X1 U12397 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9691) );
  NAND4_X1 U12398 ( .A1(n9676), .A2(n9674), .A3(n9675), .A4(n9691), .ZN(n9677)
         );
  OR2_X1 U12399 ( .A1(n9678), .A2(n9677), .ZN(n9680) );
  NAND2_X1 U12400 ( .A1(n9680), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9679) );
  MUX2_X1 U12401 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9679), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9681) );
  OR2_X1 U12402 ( .A1(n9680), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n9708) );
  NAND2_X1 U12403 ( .A1(n9681), .A2(n9708), .ZN(n12797) );
  OAI22_X1 U12404 ( .A1(n12797), .A2(n9779), .B1(n9695), .B2(n15732), .ZN(
        n9682) );
  INV_X1 U12405 ( .A(n9682), .ZN(n9683) );
  INV_X1 U12406 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n12442) );
  INV_X1 U12407 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n15692) );
  NAND2_X1 U12408 ( .A1(n9701), .A2(n15692), .ZN(n9685) );
  NAND2_X1 U12409 ( .A1(n9712), .A2(n9685), .ZN(n15209) );
  OR2_X1 U12410 ( .A1(n15209), .A2(n9519), .ZN(n9690) );
  INV_X1 U12411 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15210) );
  OR2_X1 U12412 ( .A1(n10255), .A2(n15210), .ZN(n9687) );
  INV_X1 U12413 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15336) );
  OR2_X1 U12414 ( .A1(n9915), .A2(n15336), .ZN(n9686) );
  AND2_X1 U12415 ( .A1(n9687), .A2(n9686), .ZN(n9689) );
  NAND2_X1 U12416 ( .A1(n9912), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U12417 ( .A1(n15213), .A2(n14746), .ZN(n10199) );
  NAND2_X1 U12418 ( .A1(n11348), .A2(n10318), .ZN(n9698) );
  NAND2_X1 U12419 ( .A1(n9692), .A2(n9691), .ZN(n9693) );
  NAND2_X1 U12420 ( .A1(n9693), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9694) );
  XNOR2_X1 U12421 ( .A(n9694), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12676) );
  NOR2_X1 U12422 ( .A1(n9695), .A2(n15740), .ZN(n9696) );
  AOI21_X1 U12423 ( .B1(n12676), .B2(n9534), .A(n9696), .ZN(n9697) );
  NAND2_X2 U12424 ( .A1(n9698), .A2(n9697), .ZN(n15338) );
  NAND2_X1 U12425 ( .A1(n9699), .A2(n12442), .ZN(n9700) );
  AND2_X1 U12426 ( .A1(n9701), .A2(n9700), .ZN(n14692) );
  NAND2_X1 U12427 ( .A1(n14692), .A2(n9911), .ZN(n9705) );
  NAND2_X1 U12428 ( .A1(n9782), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9704) );
  INV_X1 U12429 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15730) );
  OR2_X1 U12430 ( .A1(n9528), .A2(n15730), .ZN(n9703) );
  INV_X1 U12431 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15344) );
  OR2_X1 U12432 ( .A1(n9915), .A2(n15344), .ZN(n9702) );
  NAND4_X1 U12433 ( .A1(n9705), .A2(n9704), .A3(n9703), .A4(n9702), .ZN(n14841) );
  INV_X1 U12434 ( .A(n14841), .ZN(n14820) );
  NAND2_X1 U12435 ( .A1(n15338), .A2(n14820), .ZN(n10198) );
  NAND2_X1 U12436 ( .A1(n15338), .A2(n14841), .ZN(n15203) );
  INV_X1 U12437 ( .A(n14746), .ZN(n15191) );
  OR2_X1 U12438 ( .A1(n15213), .A2(n15191), .ZN(n9706) );
  AND2_X1 U12439 ( .A1(n15218), .A2(n15203), .ZN(n15179) );
  NAND2_X1 U12440 ( .A1(n11335), .A2(n10318), .ZN(n9711) );
  NAND2_X1 U12441 ( .A1(n9708), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9709) );
  XNOR2_X1 U12442 ( .A(n9709), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14922) );
  AOI22_X1 U12443 ( .A1(n14922), .A2(n9534), .B1(n6431), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n9710) );
  INV_X1 U12444 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12803) );
  NAND2_X1 U12445 ( .A1(n9712), .A2(n12803), .ZN(n9713) );
  AND2_X1 U12446 ( .A1(n9723), .A2(n9713), .ZN(n15194) );
  NAND2_X1 U12447 ( .A1(n15194), .A2(n9911), .ZN(n9716) );
  AOI22_X1 U12448 ( .A1(n9912), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n9782), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U12449 ( .A1(n10254), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9714) );
  XNOR2_X1 U12450 ( .A(n15188), .B(n15167), .ZN(n15183) );
  INV_X1 U12451 ( .A(n15167), .ZN(n14840) );
  OR2_X1 U12452 ( .A1(n15188), .A2(n14840), .ZN(n9718) );
  NAND2_X1 U12453 ( .A1(n11508), .A2(n10318), .ZN(n9721) );
  NAND2_X1 U12454 ( .A1(n9932), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9719) );
  XNOR2_X1 U12455 ( .A(n9719), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14939) );
  AOI22_X1 U12456 ( .A1(n6431), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9534), 
        .B2(n14939), .ZN(n9720) );
  INV_X1 U12457 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n15731) );
  NAND2_X1 U12458 ( .A1(n9723), .A2(n15731), .ZN(n9724) );
  NAND2_X1 U12459 ( .A1(n9747), .A2(n9724), .ZN(n15160) );
  OR2_X1 U12460 ( .A1(n15160), .A2(n9519), .ZN(n9730) );
  INV_X1 U12461 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U12462 ( .A1(n9912), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9726) );
  INV_X1 U12463 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14928) );
  OR2_X1 U12464 ( .A1(n10255), .A2(n14928), .ZN(n9725) );
  OAI211_X1 U12465 ( .C1(n9727), .C2(n9915), .A(n9726), .B(n9725), .ZN(n9728)
         );
  INV_X1 U12466 ( .A(n9728), .ZN(n9729) );
  NAND2_X1 U12467 ( .A1(n9730), .A2(n9729), .ZN(n15193) );
  NAND2_X1 U12468 ( .A1(n15319), .A2(n15193), .ZN(n10221) );
  NAND2_X1 U12469 ( .A1(n9731), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9732) );
  XNOR2_X1 U12470 ( .A(n9732), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14956) );
  AOI22_X1 U12471 ( .A1(n6431), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9534), 
        .B2(n14956), .ZN(n9733) );
  XNOR2_X1 U12472 ( .A(n9747), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n15150) );
  NAND2_X1 U12473 ( .A1(n15150), .A2(n9911), .ZN(n9740) );
  INV_X1 U12474 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15316) );
  NAND2_X1 U12475 ( .A1(n9912), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9737) );
  INV_X1 U12476 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9735) );
  OR2_X1 U12477 ( .A1(n10255), .A2(n9735), .ZN(n9736) );
  OAI211_X1 U12478 ( .C1(n15316), .C2(n9915), .A(n9737), .B(n9736), .ZN(n9738)
         );
  INV_X1 U12479 ( .A(n9738), .ZN(n9739) );
  NAND2_X1 U12480 ( .A1(n9740), .A2(n9739), .ZN(n15125) );
  OR2_X1 U12481 ( .A1(n15149), .A2(n15125), .ZN(n9898) );
  AND2_X1 U12482 ( .A1(n15136), .A2(n9898), .ZN(n9741) );
  NAND2_X1 U12483 ( .A1(n15149), .A2(n15125), .ZN(n10201) );
  NAND2_X1 U12484 ( .A1(n12098), .A2(n10318), .ZN(n9745) );
  AOI22_X1 U12485 ( .A1(n6431), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9877), 
        .B2(n9534), .ZN(n9744) );
  INV_X1 U12486 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n14803) );
  INV_X1 U12487 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9746) );
  OAI21_X1 U12488 ( .B1(n9747), .B2(n14803), .A(n9746), .ZN(n9748) );
  AND2_X1 U12489 ( .A1(n9748), .A2(n9758), .ZN(n15129) );
  NAND2_X1 U12490 ( .A1(n15129), .A2(n9911), .ZN(n9753) );
  INV_X1 U12491 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14954) );
  NAND2_X1 U12492 ( .A1(n9912), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U12493 ( .A1(n9782), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9749) );
  OAI211_X1 U12494 ( .C1(n14954), .C2(n9915), .A(n9750), .B(n9749), .ZN(n9751)
         );
  INV_X1 U12495 ( .A(n9751), .ZN(n9752) );
  NAND2_X1 U12496 ( .A1(n9753), .A2(n9752), .ZN(n14839) );
  OR2_X1 U12497 ( .A1(n15307), .A2(n14839), .ZN(n9754) );
  NAND2_X1 U12498 ( .A1(n6431), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9755) );
  INV_X1 U12499 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14771) );
  NAND2_X1 U12500 ( .A1(n9758), .A2(n14771), .ZN(n9759) );
  AND2_X1 U12501 ( .A1(n9768), .A2(n9759), .ZN(n15108) );
  NAND2_X1 U12502 ( .A1(n15108), .A2(n9911), .ZN(n9764) );
  INV_X1 U12503 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15304) );
  NAND2_X1 U12504 ( .A1(n9912), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U12505 ( .A1(n9782), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9760) );
  OAI211_X1 U12506 ( .C1(n15304), .C2(n9915), .A(n9761), .B(n9760), .ZN(n9762)
         );
  INV_X1 U12507 ( .A(n9762), .ZN(n9763) );
  INV_X1 U12508 ( .A(n15104), .ZN(n15107) );
  INV_X1 U12509 ( .A(n15089), .ZN(n15126) );
  NAND2_X1 U12510 ( .A1(n15115), .A2(n15126), .ZN(n9765) );
  NAND2_X1 U12511 ( .A1(n6431), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9766) );
  INV_X1 U12512 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14726) );
  NAND2_X1 U12513 ( .A1(n9768), .A2(n14726), .ZN(n9769) );
  NAND2_X1 U12514 ( .A1(n9780), .A2(n9769), .ZN(n15097) );
  OR2_X1 U12515 ( .A1(n15097), .A2(n9519), .ZN(n9775) );
  INV_X1 U12516 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U12517 ( .A1(n9782), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U12518 ( .A1(n9912), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9770) );
  OAI211_X1 U12519 ( .C1(n9772), .C2(n9915), .A(n9771), .B(n9770), .ZN(n9773)
         );
  INV_X1 U12520 ( .A(n9773), .ZN(n9774) );
  XNOR2_X1 U12521 ( .A(n15099), .B(n15069), .ZN(n15086) );
  OR2_X1 U12522 ( .A1(n15099), .A2(n15069), .ZN(n9776) );
  INV_X1 U12523 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14792) );
  NAND2_X1 U12524 ( .A1(n9780), .A2(n14792), .ZN(n9781) );
  AND2_X1 U12525 ( .A1(n9791), .A2(n9781), .ZN(n15079) );
  NAND2_X1 U12526 ( .A1(n15079), .A2(n9911), .ZN(n9787) );
  INV_X1 U12527 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15291) );
  NAND2_X1 U12528 ( .A1(n9912), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U12529 ( .A1(n9782), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9783) );
  OAI211_X1 U12530 ( .C1(n15291), .C2(n9915), .A(n9784), .B(n9783), .ZN(n9785)
         );
  INV_X1 U12531 ( .A(n9785), .ZN(n9786) );
  XNOR2_X1 U12532 ( .A(n15370), .B(n15090), .ZN(n9900) );
  NAND2_X1 U12533 ( .A1(n15370), .A2(n15090), .ZN(n9788) );
  NAND2_X1 U12534 ( .A1(n6431), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9789) );
  INV_X1 U12535 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9790) );
  NAND2_X1 U12536 ( .A1(n9791), .A2(n9790), .ZN(n9792) );
  NAND2_X1 U12537 ( .A1(n9803), .A2(n9792), .ZN(n15064) );
  INV_X1 U12538 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9795) );
  NAND2_X1 U12539 ( .A1(n9782), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U12540 ( .A1(n9912), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9793) );
  OAI211_X1 U12541 ( .C1(n9915), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9796)
         );
  INV_X1 U12542 ( .A(n9796), .ZN(n9797) );
  INV_X1 U12543 ( .A(n15059), .ZN(n10347) );
  NAND2_X1 U12544 ( .A1(n15282), .A2(n14837), .ZN(n9799) );
  NAND2_X1 U12545 ( .A1(n6431), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9800) );
  INV_X1 U12546 ( .A(n9803), .ZN(n9802) );
  INV_X1 U12547 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n15757) );
  NAND2_X1 U12548 ( .A1(n9803), .A2(n15757), .ZN(n9804) );
  NAND2_X1 U12549 ( .A1(n15050), .A2(n9911), .ZN(n9809) );
  INV_X1 U12550 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n15279) );
  NAND2_X1 U12551 ( .A1(n9912), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U12552 ( .A1(n9782), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9805) );
  OAI211_X1 U12553 ( .C1(n15279), .C2(n9915), .A(n9806), .B(n9805), .ZN(n9807)
         );
  INV_X1 U12554 ( .A(n9807), .ZN(n9808) );
  AND2_X2 U12555 ( .A1(n9809), .A2(n9808), .ZN(n10609) );
  XNOR2_X1 U12556 ( .A(n15049), .B(n14836), .ZN(n15042) );
  NAND2_X1 U12557 ( .A1(n12669), .A2(n10318), .ZN(n9812) );
  NAND2_X1 U12558 ( .A1(n6431), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9811) );
  INV_X1 U12559 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9814) );
  OR2_X2 U12560 ( .A1(n9828), .A2(n9814), .ZN(n9840) );
  NAND2_X1 U12561 ( .A1(n9828), .A2(n9814), .ZN(n9815) );
  NAND2_X1 U12562 ( .A1(n14811), .A2(n9911), .ZN(n9821) );
  INV_X1 U12563 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9818) );
  NAND2_X1 U12564 ( .A1(n9912), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U12565 ( .A1(n9782), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9816) );
  OAI211_X1 U12566 ( .C1(n9818), .C2(n9915), .A(n9817), .B(n9816), .ZN(n9819)
         );
  INV_X1 U12567 ( .A(n9819), .ZN(n9820) );
  NAND2_X1 U12568 ( .A1(n15264), .A2(n15012), .ZN(n15004) );
  OR2_X1 U12569 ( .A1(n15264), .A2(n15012), .ZN(n9822) );
  NAND2_X1 U12570 ( .A1(n12478), .A2(n10318), .ZN(n9824) );
  NAND2_X1 U12571 ( .A1(n6431), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9823) );
  INV_X1 U12572 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U12573 ( .A1(n9826), .A2(n9825), .ZN(n9827) );
  NAND2_X1 U12574 ( .A1(n9828), .A2(n9827), .ZN(n14733) );
  INV_X1 U12575 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U12576 ( .A1(n9912), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U12577 ( .A1(n9782), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9829) );
  OAI211_X1 U12578 ( .C1(n9831), .C2(n9915), .A(n9830), .B(n9829), .ZN(n9832)
         );
  INV_X1 U12579 ( .A(n9832), .ZN(n9833) );
  NOR2_X1 U12580 ( .A1(n15035), .A2(n15045), .ZN(n9901) );
  INV_X1 U12581 ( .A(n9901), .ZN(n9835) );
  NAND2_X1 U12582 ( .A1(n15035), .A2(n15045), .ZN(n12873) );
  NAND2_X1 U12583 ( .A1(n12872), .A2(n15029), .ZN(n9837) );
  AND2_X1 U12584 ( .A1(n15035), .A2(n14835), .ZN(n12865) );
  AOI22_X1 U12585 ( .A1(n12872), .A2(n12865), .B1(n14834), .B2(n15264), .ZN(
        n9836) );
  NAND2_X1 U12586 ( .A1(n6431), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9838) );
  INV_X1 U12587 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n12816) );
  NAND2_X1 U12588 ( .A1(n9840), .A2(n12816), .ZN(n9841) );
  NAND2_X1 U12589 ( .A1(n14991), .A2(n9841), .ZN(n12817) );
  NAND2_X1 U12590 ( .A1(n15020), .A2(n9911), .ZN(n9846) );
  INV_X1 U12591 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n15729) );
  NAND2_X1 U12592 ( .A1(n9912), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U12593 ( .A1(n10254), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9842) );
  OAI211_X1 U12594 ( .C1(n10255), .C2(n15729), .A(n9843), .B(n9842), .ZN(n9844) );
  INV_X1 U12595 ( .A(n9844), .ZN(n9845) );
  OR2_X1 U12596 ( .A1(n15258), .A2(n14833), .ZN(n9847) );
  INV_X1 U12597 ( .A(n9848), .ZN(n9849) );
  NAND2_X1 U12598 ( .A1(n9849), .A2(n13599), .ZN(n9850) );
  MUX2_X1 U12599 ( .A(n12883), .B(n14681), .S(n10801), .Z(n10015) );
  XNOR2_X1 U12600 ( .A(n10015), .B(SI_28_), .ZN(n10013) );
  NAND2_X1 U12601 ( .A1(n6431), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U12602 ( .A1(n12889), .A2(n9911), .ZN(n9858) );
  INV_X1 U12603 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U12604 ( .A1(n9782), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U12605 ( .A1(n9912), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9853) );
  OAI211_X1 U12606 ( .C1(n9915), .C2(n9855), .A(n9854), .B(n9853), .ZN(n9856)
         );
  INV_X1 U12607 ( .A(n9856), .ZN(n9857) );
  AND2_X2 U12608 ( .A1(n9858), .A2(n9857), .ZN(n15013) );
  AND2_X2 U12609 ( .A1(n14982), .A2(n9859), .ZN(n10349) );
  INV_X1 U12610 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9863) );
  INV_X1 U12611 ( .A(n9870), .ZN(n9867) );
  NAND3_X1 U12612 ( .A1(n9867), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n9876) );
  NOR2_X1 U12613 ( .A1(n9868), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n9869) );
  INV_X1 U12614 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U12615 ( .A1(n9868), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n9871) );
  NAND2_X1 U12616 ( .A1(n9871), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9872) );
  OAI21_X1 U12617 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(n9873), .A(n9872), .ZN(
        n9874) );
  NAND2_X1 U12618 ( .A1(n10419), .A2(n10125), .ZN(n9879) );
  INV_X1 U12619 ( .A(n10125), .ZN(n9878) );
  INV_X2 U12620 ( .A(n10449), .ZN(n10427) );
  NAND2_X1 U12621 ( .A1(n11957), .A2(n14967), .ZN(n15147) );
  NAND2_X1 U12622 ( .A1(n6435), .A2(n9927), .ZN(n10321) );
  OR2_X1 U12623 ( .A1(n10321), .A2(n14967), .ZN(n15507) );
  INV_X1 U12624 ( .A(n10460), .ZN(n11166) );
  NAND2_X1 U12625 ( .A1(n11166), .A2(n11203), .ZN(n10128) );
  NAND2_X1 U12626 ( .A1(n10133), .A2(n10128), .ZN(n9881) );
  AND2_X1 U12627 ( .A1(n9881), .A2(n10132), .ZN(n11113) );
  OR2_X1 U12628 ( .A1(n14853), .A2(n6845), .ZN(n12118) );
  NAND2_X1 U12629 ( .A1(n12120), .A2(n12118), .ZN(n9882) );
  NAND2_X1 U12630 ( .A1(n9882), .A2(n10335), .ZN(n12122) );
  NAND2_X1 U12631 ( .A1(n12122), .A2(n10147), .ZN(n11281) );
  INV_X1 U12632 ( .A(n11276), .ZN(n11972) );
  OR2_X1 U12633 ( .A1(n11972), .A2(n14851), .ZN(n9883) );
  AOI22_X1 U12634 ( .A1(n11922), .A2(n14849), .B1(n11952), .B2(n14850), .ZN(
        n9884) );
  NAND2_X1 U12635 ( .A1(n15496), .A2(n11805), .ZN(n11802) );
  NAND2_X1 U12636 ( .A1(n11802), .A2(n14849), .ZN(n9886) );
  NOR2_X1 U12637 ( .A1(n14849), .A2(n14850), .ZN(n9885) );
  AOI22_X1 U12638 ( .A1(n9886), .A2(n11424), .B1(n9885), .B2(n15496), .ZN(
        n9887) );
  INV_X1 U12639 ( .A(n14848), .ZN(n11806) );
  NAND2_X1 U12640 ( .A1(n15503), .A2(n11806), .ZN(n9888) );
  OR2_X1 U12641 ( .A1(n11961), .A2(n12075), .ZN(n9889) );
  NAND2_X1 U12642 ( .A1(n12217), .A2(n12162), .ZN(n9890) );
  INV_X1 U12643 ( .A(n14845), .ZN(n10423) );
  OR2_X1 U12644 ( .A1(n12166), .A2(n10423), .ZN(n9891) );
  NAND2_X1 U12645 ( .A1(n12159), .A2(n9891), .ZN(n12230) );
  INV_X1 U12646 ( .A(n14844), .ZN(n12702) );
  OR2_X1 U12647 ( .A1(n15349), .A2(n12702), .ZN(n9892) );
  INV_X1 U12648 ( .A(n14843), .ZN(n10515) );
  OR2_X1 U12649 ( .A1(n12322), .A2(n10515), .ZN(n9893) );
  INV_X1 U12650 ( .A(n14842), .ZN(n12701) );
  NAND2_X1 U12651 ( .A1(n12647), .A2(n12648), .ZN(n15217) );
  AND2_X1 U12652 ( .A1(n10209), .A2(n15216), .ZN(n9895) );
  INV_X1 U12653 ( .A(n10199), .ZN(n9894) );
  OR2_X2 U12654 ( .A1(n15182), .A2(n15183), .ZN(n15184) );
  INV_X1 U12655 ( .A(n15164), .ZN(n9896) );
  NAND2_X1 U12656 ( .A1(n15188), .A2(n15167), .ZN(n15163) );
  AND2_X1 U12657 ( .A1(n9896), .A2(n15163), .ZN(n9897) );
  INV_X1 U12658 ( .A(n15193), .ZN(n15142) );
  NOR2_X1 U12659 ( .A1(n15319), .A2(n15142), .ZN(n15119) );
  INV_X1 U12660 ( .A(n15125), .ZN(n15169) );
  NOR2_X1 U12661 ( .A1(n15149), .A2(n15169), .ZN(n15121) );
  INV_X1 U12662 ( .A(n14839), .ZN(n15143) );
  NAND2_X1 U12663 ( .A1(n15307), .A2(n15143), .ZN(n10219) );
  NAND2_X1 U12664 ( .A1(n15282), .A2(n15072), .ZN(n12869) );
  OAI211_X1 U12665 ( .C1(n15365), .C2(n14836), .A(n12873), .B(n12869), .ZN(
        n9903) );
  NOR2_X1 U12666 ( .A1(n15049), .A2(n10609), .ZN(n12871) );
  OAI21_X1 U12667 ( .B1(n9901), .B2(n12871), .A(n12873), .ZN(n9902) );
  NOR2_X1 U12668 ( .A1(n15023), .A2(n14833), .ZN(n9904) );
  INV_X1 U12669 ( .A(n9904), .ZN(n9905) );
  NAND2_X1 U12670 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  OR2_X1 U12671 ( .A1(n15003), .A2(n9907), .ZN(n9908) );
  NAND2_X1 U12672 ( .A1(n14983), .A2(n9908), .ZN(n9922) );
  INV_X1 U12673 ( .A(n9909), .ZN(n10124) );
  NAND2_X1 U12674 ( .A1(n10324), .A2(n10124), .ZN(n10123) );
  NAND2_X1 U12675 ( .A1(n15403), .A2(n9877), .ZN(n9910) );
  NAND2_X1 U12676 ( .A1(n10123), .A2(n9910), .ZN(n15327) );
  NAND2_X1 U12677 ( .A1(n10324), .A2(n15403), .ZN(n10654) );
  INV_X1 U12678 ( .A(n10654), .ZN(n10721) );
  INV_X1 U12679 ( .A(n12885), .ZN(n10844) );
  NAND2_X1 U12680 ( .A1(n9911), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9919) );
  INV_X1 U12681 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U12682 ( .A1(n9782), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9914) );
  NAND2_X1 U12683 ( .A1(n9912), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9913) );
  OAI211_X1 U12684 ( .C1(n9916), .C2(n9915), .A(n9914), .B(n9913), .ZN(n9917)
         );
  INV_X1 U12685 ( .A(n9917), .ZN(n9918) );
  INV_X1 U12686 ( .A(n12166), .ZN(n12357) );
  INV_X1 U12687 ( .A(n15349), .ZN(n12234) );
  INV_X1 U12688 ( .A(n15282), .ZN(n10599) );
  NAND2_X1 U12689 ( .A1(n15077), .A2(n10599), .ZN(n15063) );
  OR2_X4 U12690 ( .A1(n10121), .A2(n10124), .ZN(n15187) );
  INV_X1 U12691 ( .A(n15187), .ZN(n15283) );
  OAI211_X1 U12692 ( .C1(n15018), .C2(n14997), .A(n15283), .B(n14985), .ZN(
        n12888) );
  AND2_X1 U12693 ( .A1(n6435), .A2(n14967), .ZN(n9963) );
  OR2_X1 U12694 ( .A1(n10654), .A2(n9963), .ZN(n10665) );
  NAND2_X1 U12695 ( .A1(n9928), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9930) );
  XNOR2_X1 U12696 ( .A(n9930), .B(n9929), .ZN(n10833) );
  NAND2_X1 U12697 ( .A1(n9942), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9936) );
  INV_X1 U12698 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9935) );
  AND2_X1 U12699 ( .A1(n10833), .A2(n10421), .ZN(n9943) );
  NOR4_X1 U12700 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n15725) );
  NOR2_X1 U12701 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n9946) );
  NOR4_X1 U12702 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n9945) );
  NOR4_X1 U12703 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9944) );
  NAND4_X1 U12704 ( .A1(n15725), .A2(n9946), .A3(n9945), .A4(n9944), .ZN(n9956) );
  NOR4_X1 U12705 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9950) );
  NOR4_X1 U12706 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n9949) );
  NOR4_X1 U12707 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n9948) );
  NOR4_X1 U12708 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9947) );
  NAND4_X1 U12709 ( .A1(n9950), .A2(n9949), .A3(n9948), .A4(n9947), .ZN(n9955)
         );
  NAND2_X1 U12710 ( .A1(n12480), .A2(P1_B_REG_SCAN_IN), .ZN(n9952) );
  MUX2_X1 U12711 ( .A(P1_B_REG_SCAN_IN), .B(n9952), .S(n12222), .Z(n9954) );
  INV_X1 U12712 ( .A(n12674), .ZN(n9953) );
  OAI21_X1 U12713 ( .B1(n9956), .B2(n9955), .A(n10830), .ZN(n10651) );
  NAND3_X1 U12714 ( .A1(n10670), .A2(P1_STATE_REG_SCAN_IN), .A3(n10651), .ZN(
        n11901) );
  INV_X1 U12715 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n15792) );
  NAND2_X1 U12716 ( .A1(n10830), .A2(n15792), .ZN(n9958) );
  NAND2_X1 U12717 ( .A1(n12674), .A2(n12480), .ZN(n9957) );
  NAND2_X1 U12718 ( .A1(n9958), .A2(n9957), .ZN(n15791) );
  NAND2_X1 U12719 ( .A1(n15791), .A2(n10668), .ZN(n9959) );
  INV_X1 U12720 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10835) );
  AND2_X1 U12721 ( .A1(n12222), .A2(n12674), .ZN(n10832) );
  INV_X1 U12722 ( .A(n9965), .ZN(n11071) );
  NAND2_X1 U12723 ( .A1(n11120), .A2(n11121), .ZN(n9967) );
  XNOR2_X1 U12724 ( .A(n14109), .B(n13774), .ZN(n10048) );
  NAND2_X1 U12725 ( .A1(n11079), .A2(n10048), .ZN(n9969) );
  INV_X1 U12726 ( .A(n13774), .ZN(n11081) );
  NAND2_X1 U12727 ( .A1(n9969), .A2(n9968), .ZN(n11369) );
  XNOR2_X1 U12728 ( .A(n14108), .B(n13783), .ZN(n11431) );
  NAND2_X1 U12729 ( .A1(n11369), .A2(n11431), .ZN(n11428) );
  OR2_X1 U12730 ( .A1(n14108), .A2(n15563), .ZN(n11427) );
  OR2_X1 U12731 ( .A1(n13791), .A2(n14107), .ZN(n11630) );
  NAND2_X1 U12732 ( .A1(n11428), .A2(n7789), .ZN(n9974) );
  INV_X1 U12733 ( .A(n14107), .ZN(n9971) );
  NAND2_X1 U12734 ( .A1(n11429), .A2(n11630), .ZN(n9972) );
  NAND2_X1 U12735 ( .A1(n13806), .A2(n13808), .ZN(n11573) );
  NAND2_X1 U12736 ( .A1(n10053), .A2(n11573), .ZN(n11572) );
  NAND2_X1 U12737 ( .A1(n9974), .A2(n9973), .ZN(n9976) );
  INV_X1 U12738 ( .A(n13808), .ZN(n14106) );
  OR2_X1 U12739 ( .A1(n13806), .A2(n14106), .ZN(n9975) );
  NAND2_X1 U12740 ( .A1(n9976), .A2(n9975), .ZN(n11568) );
  NAND2_X1 U12741 ( .A1(n11568), .A2(n14048), .ZN(n9978) );
  INV_X1 U12742 ( .A(n13815), .ZN(n14105) );
  OR2_X1 U12743 ( .A1(n13813), .A2(n14105), .ZN(n9977) );
  NAND2_X1 U12744 ( .A1(n9978), .A2(n9977), .ZN(n11534) );
  XNOR2_X1 U12745 ( .A(n14614), .B(n13820), .ZN(n14049) );
  INV_X1 U12746 ( .A(n13820), .ZN(n14104) );
  OR2_X1 U12747 ( .A1(n14614), .A2(n14104), .ZN(n9979) );
  NAND2_X1 U12748 ( .A1(n13840), .A2(n14103), .ZN(n9981) );
  XNOR2_X1 U12749 ( .A(n14610), .B(n13837), .ZN(n11779) );
  INV_X1 U12750 ( .A(n13837), .ZN(n14101) );
  NAND2_X1 U12751 ( .A1(n14610), .A2(n14101), .ZN(n9982) );
  NAND2_X1 U12752 ( .A1(n9983), .A2(n9982), .ZN(n12002) );
  XNOR2_X1 U12753 ( .A(n14604), .B(n13848), .ZN(n14054) );
  INV_X1 U12754 ( .A(n13848), .ZN(n14100) );
  NAND2_X1 U12755 ( .A1(n14604), .A2(n14100), .ZN(n9984) );
  OR2_X1 U12756 ( .A1(n13860), .A2(n14099), .ZN(n9985) );
  XNOR2_X1 U12757 ( .A(n14599), .B(n14098), .ZN(n14055) );
  OR2_X1 U12758 ( .A1(n14599), .A2(n14098), .ZN(n9987) );
  NAND2_X1 U12759 ( .A1(n12290), .A2(n9987), .ZN(n12405) );
  NAND2_X1 U12760 ( .A1(n14594), .A2(n14097), .ZN(n9988) );
  NAND2_X1 U12761 ( .A1(n12405), .A2(n9988), .ZN(n9990) );
  OR2_X1 U12762 ( .A1(n14594), .A2(n14097), .ZN(n9989) );
  NOR2_X1 U12763 ( .A1(n13880), .A2(n14096), .ZN(n12493) );
  NAND2_X1 U12764 ( .A1(n13880), .A2(n14096), .ZN(n12492) );
  XNOR2_X1 U12765 ( .A(n13887), .B(n14095), .ZN(n14060) );
  NAND2_X1 U12766 ( .A1(n14655), .A2(n14094), .ZN(n14465) );
  INV_X1 U12767 ( .A(n14465), .ZN(n9995) );
  XNOR2_X1 U12768 ( .A(n14651), .B(n13896), .ZN(n14466) );
  NOR2_X1 U12769 ( .A1(n13887), .A2(n14095), .ZN(n14462) );
  INV_X1 U12770 ( .A(n14094), .ZN(n12713) );
  INV_X1 U12771 ( .A(n14655), .ZN(n9992) );
  AOI22_X1 U12772 ( .A1(n14462), .A2(n14465), .B1(n12713), .B2(n9992), .ZN(
        n9993) );
  NAND2_X1 U12773 ( .A1(n14651), .A2(n14093), .ZN(n9996) );
  XNOR2_X1 U12774 ( .A(n14450), .B(n14092), .ZN(n14445) );
  AND2_X1 U12775 ( .A1(n14433), .A2(n14091), .ZN(n9998) );
  OR2_X1 U12776 ( .A1(n14450), .A2(n14092), .ZN(n14421) );
  OR2_X1 U12777 ( .A1(n9998), .A2(n14421), .ZN(n9999) );
  OR2_X1 U12778 ( .A1(n14557), .A2(n14090), .ZN(n10000) );
  OR2_X1 U12779 ( .A1(n14433), .A2(n14091), .ZN(n14413) );
  NAND2_X1 U12780 ( .A1(n14557), .A2(n14090), .ZN(n10001) );
  XNOR2_X1 U12781 ( .A(n14638), .B(n14089), .ZN(n14394) );
  NAND2_X1 U12782 ( .A1(n14634), .A2(n13960), .ZN(n10003) );
  INV_X1 U12783 ( .A(n13960), .ZN(n14088) );
  NAND2_X1 U12784 ( .A1(n14634), .A2(n14088), .ZN(n10005) );
  NAND2_X1 U12785 ( .A1(n14629), .A2(n14085), .ZN(n10006) );
  NAND2_X1 U12786 ( .A1(n10007), .A2(n10006), .ZN(n14326) );
  NAND2_X1 U12787 ( .A1(n14519), .A2(n14083), .ZN(n10008) );
  NAND2_X1 U12788 ( .A1(n14293), .A2(n14082), .ZN(n10012) );
  INV_X1 U12789 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15398) );
  MUX2_X1 U12790 ( .A(n15398), .B(n12863), .S(n10801), .Z(n10262) );
  XNOR2_X1 U12791 ( .A(n10262), .B(SI_29_), .ZN(n10260) );
  NAND2_X1 U12792 ( .A1(n10274), .A2(n7072), .ZN(n10017) );
  OR2_X1 U12793 ( .A1(n10042), .A2(n7091), .ZN(n10024) );
  INV_X1 U12794 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10021) );
  NAND2_X1 U12795 ( .A1(n10379), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n10020) );
  NAND2_X1 U12796 ( .A1(n7904), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n10019) );
  OAI211_X1 U12797 ( .C1(n10021), .C2(n10380), .A(n10020), .B(n10019), .ZN(
        n10022) );
  INV_X1 U12798 ( .A(n10022), .ZN(n10023) );
  NAND2_X1 U12799 ( .A1(n10024), .A2(n10023), .ZN(n14081) );
  NAND2_X1 U12800 ( .A1(n15557), .A2(n15558), .ZN(n10029) );
  NAND2_X1 U12801 ( .A1(n10028), .A2(n10027), .ZN(n10116) );
  NOR2_X1 U12802 ( .A1(n10029), .A2(n10116), .ZN(n10385) );
  INV_X1 U12803 ( .A(n10114), .ZN(n10030) );
  NAND2_X1 U12804 ( .A1(n10385), .A2(n10030), .ZN(n10031) );
  OR2_X1 U12805 ( .A1(n14033), .A2(n14031), .ZN(n11633) );
  NAND2_X1 U12806 ( .A1(n14426), .A2(n11633), .ZN(n10033) );
  OR2_X1 U12807 ( .A1(n14518), .A2(n14497), .ZN(n10102) );
  AND2_X1 U12808 ( .A1(n10034), .A2(n13755), .ZN(n11128) );
  INV_X1 U12809 ( .A(n13806), .ZN(n11701) );
  INV_X1 U12810 ( .A(n13813), .ZN(n11663) );
  INV_X1 U12811 ( .A(n14604), .ZN(n10038) );
  INV_X1 U12812 ( .A(n14594), .ZN(n12412) );
  NAND2_X2 U12813 ( .A1(n14311), .A2(n10415), .ZN(n10107) );
  INV_X1 U12814 ( .A(n14516), .ZN(n10045) );
  INV_X1 U12815 ( .A(n10042), .ZN(n10043) );
  INV_X1 U12816 ( .A(n14485), .ZN(n14510) );
  AOI22_X1 U12817 ( .A1(n10043), .A2(n14510), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14490), .ZN(n10044) );
  OAI21_X1 U12818 ( .B1(n10045), .B2(n14455), .A(n10044), .ZN(n10046) );
  INV_X1 U12819 ( .A(n10048), .ZN(n14043) );
  NAND2_X1 U12820 ( .A1(n11434), .A2(n15563), .ZN(n11430) );
  OR2_X1 U12821 ( .A1(n14109), .A2(n13774), .ZN(n11370) );
  NAND2_X1 U12822 ( .A1(n14108), .A2(n13783), .ZN(n10050) );
  INV_X1 U12823 ( .A(n11570), .ZN(n10052) );
  INV_X1 U12824 ( .A(n14048), .ZN(n11569) );
  NAND2_X1 U12825 ( .A1(n13813), .A2(n13815), .ZN(n10054) );
  OR2_X1 U12826 ( .A1(n14614), .A2(n13820), .ZN(n10055) );
  NAND2_X1 U12827 ( .A1(n14614), .A2(n13820), .ZN(n11749) );
  INV_X1 U12828 ( .A(n14103), .ZN(n10056) );
  OR2_X1 U12829 ( .A1(n13840), .A2(n10056), .ZN(n10057) );
  NAND2_X1 U12830 ( .A1(n11753), .A2(n10057), .ZN(n11782) );
  INV_X1 U12831 ( .A(n11779), .ZN(n14052) );
  OR2_X1 U12832 ( .A1(n14610), .A2(n13837), .ZN(n10058) );
  INV_X1 U12833 ( .A(n14054), .ZN(n10059) );
  OR2_X1 U12834 ( .A1(n14604), .A2(n13848), .ZN(n10060) );
  INV_X1 U12835 ( .A(n14099), .ZN(n10062) );
  XNOR2_X1 U12836 ( .A(n13860), .B(n10062), .ZN(n12185) );
  NAND2_X1 U12837 ( .A1(n13860), .A2(n10062), .ZN(n10063) );
  INV_X1 U12838 ( .A(n14098), .ZN(n12186) );
  OR2_X1 U12839 ( .A1(n14599), .A2(n12186), .ZN(n12407) );
  XNOR2_X1 U12840 ( .A(n14594), .B(n14097), .ZN(n14057) );
  INV_X1 U12841 ( .A(n14097), .ZN(n13869) );
  OR2_X1 U12842 ( .A1(n14594), .A2(n13869), .ZN(n12491) );
  INV_X1 U12843 ( .A(n14096), .ZN(n13882) );
  OR2_X1 U12844 ( .A1(n13880), .A2(n13882), .ZN(n10064) );
  AND2_X1 U12845 ( .A1(n12491), .A2(n10064), .ZN(n10065) );
  INV_X1 U12846 ( .A(n14095), .ZN(n13657) );
  OR2_X1 U12847 ( .A1(n13887), .A2(n13657), .ZN(n10066) );
  XNOR2_X1 U12848 ( .A(n14655), .B(n14094), .ZN(n14493) );
  NAND2_X1 U12849 ( .A1(n14651), .A2(n13896), .ZN(n10067) );
  OR2_X1 U12850 ( .A1(n14651), .A2(n13896), .ZN(n10068) );
  INV_X1 U12851 ( .A(n14092), .ZN(n10070) );
  OR2_X1 U12852 ( .A1(n14450), .A2(n10070), .ZN(n10071) );
  INV_X1 U12853 ( .A(n14091), .ZN(n13708) );
  NOR2_X1 U12854 ( .A1(n14433), .A2(n13708), .ZN(n14038) );
  INV_X1 U12855 ( .A(n14090), .ZN(n14039) );
  NOR2_X1 U12856 ( .A1(n14557), .A2(n14039), .ZN(n10072) );
  INV_X1 U12857 ( .A(n10072), .ZN(n10073) );
  AOI22_X1 U12858 ( .A1(n10073), .A2(n14404), .B1(n14039), .B2(n14557), .ZN(
        n10074) );
  INV_X1 U12859 ( .A(n14089), .ZN(n13709) );
  OR2_X1 U12860 ( .A1(n14638), .A2(n13709), .ZN(n10075) );
  NAND2_X1 U12861 ( .A1(n14638), .A2(n13709), .ZN(n10076) );
  NAND2_X1 U12862 ( .A1(n14541), .A2(n14064), .ZN(n10078) );
  NAND2_X1 U12863 ( .A1(n14360), .A2(n10078), .ZN(n10080) );
  OR2_X1 U12864 ( .A1(n14541), .A2(n14064), .ZN(n10079) );
  INV_X1 U12865 ( .A(n14347), .ZN(n10081) );
  INV_X1 U12866 ( .A(n14086), .ZN(n10082) );
  NAND2_X1 U12867 ( .A1(n14536), .A2(n10082), .ZN(n10083) );
  INV_X1 U12868 ( .A(n14085), .ZN(n13733) );
  NAND2_X1 U12869 ( .A1(n14629), .A2(n13733), .ZN(n14318) );
  NAND2_X1 U12870 ( .A1(n14527), .A2(n13986), .ZN(n14062) );
  AND2_X1 U12871 ( .A1(n14318), .A2(n14062), .ZN(n10085) );
  OR2_X1 U12872 ( .A1(n14527), .A2(n13986), .ZN(n14063) );
  INV_X1 U12873 ( .A(n14063), .ZN(n10084) );
  NAND2_X1 U12874 ( .A1(n14519), .A2(n13735), .ZN(n10086) );
  NAND2_X1 U12875 ( .A1(n13756), .A2(n14041), .ZN(n10088) );
  NAND2_X1 U12876 ( .A1(n14076), .A2(n14280), .ZN(n10087) );
  INV_X1 U12877 ( .A(n14481), .ZN(n14443) );
  AOI211_X1 U12878 ( .C1(n10415), .C2(n14082), .A(n14443), .B(n10025), .ZN(
        n10089) );
  NAND3_X1 U12879 ( .A1(n10415), .A2(n14082), .A3(n14481), .ZN(n10094) );
  INV_X1 U12880 ( .A(n14683), .ZN(n14074) );
  NAND2_X1 U12881 ( .A1(n14074), .A2(P2_B_REG_SCAN_IN), .ZN(n10090) );
  AND2_X1 U12882 ( .A1(n13725), .A2(n10090), .ZN(n10384) );
  INV_X1 U12883 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U12884 ( .A1(n10379), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n10092) );
  INV_X1 U12885 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n15651) );
  OR2_X1 U12886 ( .A1(n10380), .A2(n15651), .ZN(n10091) );
  OAI211_X1 U12887 ( .C1(n7040), .C2(n12843), .A(n10092), .B(n10091), .ZN(
        n14080) );
  AOI22_X1 U12888 ( .A1(n14082), .A2(n14073), .B1(n10384), .B2(n14080), .ZN(
        n10093) );
  OAI21_X1 U12889 ( .B1(n10098), .B2(n10094), .A(n10093), .ZN(n10095) );
  INV_X1 U12890 ( .A(n10095), .ZN(n10096) );
  OR2_X1 U12891 ( .A1(n10098), .A2(n14443), .ZN(n10099) );
  INV_X2 U12892 ( .A(n14490), .ZN(n14502) );
  INV_X1 U12893 ( .A(n14068), .ZN(n10103) );
  NAND2_X1 U12894 ( .A1(n10105), .A2(n10104), .ZN(n14292) );
  INV_X1 U12895 ( .A(n14564), .ZN(n11698) );
  INV_X1 U12896 ( .A(n14311), .ZN(n10106) );
  AOI21_X1 U12897 ( .B1(n10106), .B2(n14293), .A(n14486), .ZN(n10108) );
  NAND2_X1 U12898 ( .A1(n10108), .A2(n10107), .ZN(n14295) );
  NAND2_X1 U12899 ( .A1(n14081), .A2(n13725), .ZN(n10112) );
  NAND2_X1 U12900 ( .A1(n14083), .A2(n14073), .ZN(n10111) );
  AND2_X1 U12901 ( .A1(n10112), .A2(n10111), .ZN(n12855) );
  NOR2_X1 U12902 ( .A1(n10116), .A2(n15557), .ZN(n10117) );
  NAND2_X1 U12903 ( .A1(n10413), .A2(n14618), .ZN(n10120) );
  NOR2_X1 U12904 ( .A1(n15403), .A2(n14967), .ZN(n10126) );
  OAI21_X1 U12905 ( .B1(n10126), .B2(n10125), .A(n10124), .ZN(n10127) );
  MUX2_X1 U12906 ( .A(n14848), .B(n15503), .S(n10139), .Z(n10163) );
  XNOR2_X1 U12907 ( .A(n10139), .B(n10128), .ZN(n10131) );
  OR2_X1 U12908 ( .A1(n10460), .A2(n11203), .ZN(n10129) );
  NAND2_X1 U12909 ( .A1(n11164), .A2(n10129), .ZN(n15476) );
  NAND2_X1 U12910 ( .A1(n15476), .A2(n10419), .ZN(n10130) );
  MUX2_X1 U12911 ( .A(n10133), .B(n10132), .S(n10139), .Z(n10134) );
  NAND2_X1 U12912 ( .A1(n10139), .A2(n6845), .ZN(n10136) );
  OAI211_X1 U12913 ( .C1(n10139), .C2(n14853), .A(n10136), .B(n10135), .ZN(
        n10137) );
  NAND3_X1 U12914 ( .A1(n10139), .A2(n10146), .A3(n12148), .ZN(n10140) );
  OAI21_X1 U12915 ( .B1(n6844), .B2(n10139), .A(n10140), .ZN(n10141) );
  NAND2_X1 U12916 ( .A1(n10141), .A2(n10147), .ZN(n10144) );
  NAND2_X1 U12917 ( .A1(n10335), .A2(n10142), .ZN(n10143) );
  NAND2_X1 U12918 ( .A1(n10144), .A2(n10143), .ZN(n10145) );
  MUX2_X1 U12919 ( .A(n10147), .B(n10146), .S(n10206), .Z(n10148) );
  NAND2_X1 U12920 ( .A1(n10149), .A2(n10148), .ZN(n10152) );
  INV_X1 U12921 ( .A(n14851), .ZN(n11939) );
  MUX2_X1 U12922 ( .A(n11972), .B(n11939), .S(n10139), .Z(n10151) );
  MUX2_X1 U12923 ( .A(n14851), .B(n11276), .S(n10139), .Z(n10150) );
  NAND2_X1 U12924 ( .A1(n10152), .A2(n10151), .ZN(n10153) );
  MUX2_X1 U12925 ( .A(n14850), .B(n15496), .S(n10139), .Z(n10156) );
  MUX2_X1 U12926 ( .A(n14849), .B(n11424), .S(n10206), .Z(n10158) );
  MUX2_X1 U12927 ( .A(n11938), .B(n11922), .S(n10139), .Z(n10157) );
  MUX2_X1 U12928 ( .A(n14848), .B(n15503), .S(n10281), .Z(n10160) );
  MUX2_X1 U12929 ( .A(n14847), .B(n11961), .S(n10281), .Z(n10167) );
  NAND2_X1 U12930 ( .A1(n10166), .A2(n10167), .ZN(n10165) );
  MUX2_X1 U12931 ( .A(n14847), .B(n11961), .S(n7046), .Z(n10164) );
  MUX2_X1 U12932 ( .A(n12217), .B(n14846), .S(n10281), .Z(n10170) );
  MUX2_X1 U12933 ( .A(n12217), .B(n14846), .S(n10139), .Z(n10169) );
  INV_X1 U12934 ( .A(n10170), .ZN(n10171) );
  MUX2_X1 U12935 ( .A(n14845), .B(n12166), .S(n10281), .Z(n10174) );
  MUX2_X1 U12936 ( .A(n14845), .B(n12166), .S(n7046), .Z(n10172) );
  INV_X1 U12937 ( .A(n10174), .ZN(n10175) );
  MUX2_X1 U12938 ( .A(n14844), .B(n15349), .S(n10139), .Z(n10179) );
  MUX2_X1 U12939 ( .A(n14844), .B(n15349), .S(n10281), .Z(n10176) );
  NAND2_X1 U12940 ( .A1(n10177), .A2(n10176), .ZN(n10182) );
  INV_X1 U12941 ( .A(n10178), .ZN(n10180) );
  NAND2_X1 U12942 ( .A1(n10180), .A2(n6878), .ZN(n10181) );
  MUX2_X1 U12943 ( .A(n14843), .B(n12322), .S(n10281), .Z(n10184) );
  MUX2_X1 U12944 ( .A(n14843), .B(n12322), .S(n10139), .Z(n10183) );
  INV_X1 U12945 ( .A(n10184), .ZN(n10185) );
  MUX2_X1 U12946 ( .A(n14842), .B(n12552), .S(n10139), .Z(n10186) );
  NAND4_X1 U12947 ( .A1(n12648), .A2(n14842), .A3(n10199), .A4(n10139), .ZN(
        n10195) );
  INV_X1 U12948 ( .A(n10186), .ZN(n10187) );
  AOI21_X1 U12949 ( .B1(n15216), .B2(n14746), .A(n10281), .ZN(n10188) );
  INV_X1 U12950 ( .A(n10188), .ZN(n10191) );
  OAI21_X1 U12951 ( .B1(n15216), .B2(n14746), .A(n15213), .ZN(n10189) );
  INV_X1 U12952 ( .A(n10189), .ZN(n10190) );
  OAI22_X1 U12953 ( .A1(n10192), .A2(n6480), .B1(n10191), .B2(n10190), .ZN(
        n10193) );
  INV_X1 U12954 ( .A(n10193), .ZN(n10194) );
  OAI21_X1 U12955 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10213) );
  OAI21_X1 U12956 ( .B1(n10281), .B2(n15149), .A(n10201), .ZN(n10202) );
  NAND2_X1 U12957 ( .A1(n10219), .A2(n10202), .ZN(n10204) );
  OR2_X1 U12958 ( .A1(n15121), .A2(n7046), .ZN(n10203) );
  NAND2_X1 U12959 ( .A1(n10204), .A2(n10203), .ZN(n10225) );
  OR2_X1 U12960 ( .A1(n15307), .A2(n15143), .ZN(n10224) );
  NAND2_X1 U12961 ( .A1(n15319), .A2(n10281), .ZN(n10205) );
  OAI211_X1 U12962 ( .C1(n15142), .C2(n10206), .A(n15136), .B(n10205), .ZN(
        n10207) );
  AND2_X1 U12963 ( .A1(n10224), .A2(n10207), .ZN(n10208) );
  AND2_X1 U12964 ( .A1(n10225), .A2(n10208), .ZN(n10214) );
  INV_X1 U12965 ( .A(n10209), .ZN(n10210) );
  INV_X1 U12966 ( .A(n15188), .ZN(n15325) );
  MUX2_X1 U12967 ( .A(n15167), .B(n15325), .S(n10281), .Z(n10216) );
  MUX2_X1 U12968 ( .A(n14840), .B(n15188), .S(n7046), .Z(n10215) );
  AOI22_X1 U12969 ( .A1(n10210), .A2(n10281), .B1(n10216), .B2(n10215), .ZN(
        n10211) );
  INV_X1 U12970 ( .A(n10214), .ZN(n10229) );
  INV_X1 U12971 ( .A(n10215), .ZN(n10218) );
  INV_X1 U12972 ( .A(n10216), .ZN(n10217) );
  NAND2_X1 U12973 ( .A1(n10218), .A2(n10217), .ZN(n10228) );
  MUX2_X1 U12974 ( .A(n10219), .B(n10224), .S(n7046), .Z(n10227) );
  NAND2_X1 U12975 ( .A1(n15142), .A2(n7046), .ZN(n10220) );
  OAI211_X1 U12976 ( .C1(n15319), .C2(n10139), .A(n10221), .B(n10220), .ZN(
        n10222) );
  NAND2_X1 U12977 ( .A1(n15138), .A2(n10222), .ZN(n10223) );
  NAND3_X1 U12978 ( .A1(n10225), .A2(n10224), .A3(n10223), .ZN(n10226) );
  OAI211_X1 U12979 ( .C1(n10229), .C2(n10228), .A(n10227), .B(n10226), .ZN(
        n10230) );
  INV_X1 U12980 ( .A(n10230), .ZN(n10231) );
  MUX2_X1 U12981 ( .A(n15089), .B(n15375), .S(n7046), .Z(n10234) );
  MUX2_X1 U12982 ( .A(n15126), .B(n15115), .S(n10281), .Z(n10233) );
  MUX2_X1 U12983 ( .A(n15069), .B(n15099), .S(n10206), .Z(n10236) );
  MUX2_X1 U12984 ( .A(n15069), .B(n15099), .S(n10139), .Z(n10235) );
  INV_X1 U12985 ( .A(n10236), .ZN(n10237) );
  INV_X1 U12986 ( .A(n15090), .ZN(n14838) );
  MUX2_X1 U12987 ( .A(n14838), .B(n15078), .S(n7046), .Z(n10238) );
  NAND2_X1 U12988 ( .A1(n10239), .A2(n10238), .ZN(n10242) );
  MUX2_X1 U12989 ( .A(n15090), .B(n15370), .S(n10281), .Z(n10240) );
  INV_X1 U12990 ( .A(n10240), .ZN(n10241) );
  NAND2_X1 U12991 ( .A1(n10242), .A2(n10241), .ZN(n10243) );
  MUX2_X1 U12992 ( .A(n14837), .B(n15282), .S(n10281), .Z(n10244) );
  MUX2_X1 U12993 ( .A(n14837), .B(n15282), .S(n10139), .Z(n10245) );
  MUX2_X1 U12994 ( .A(n14836), .B(n15049), .S(n7046), .Z(n10247) );
  INV_X1 U12995 ( .A(n15035), .ZN(n15270) );
  MUX2_X1 U12996 ( .A(n15045), .B(n15270), .S(n10281), .Z(n10249) );
  MUX2_X1 U12997 ( .A(n14835), .B(n15035), .S(n7046), .Z(n10248) );
  MUX2_X1 U12998 ( .A(n10609), .B(n15365), .S(n10281), .Z(n10246) );
  NAND2_X1 U12999 ( .A1(n10249), .A2(n10248), .ZN(n10283) );
  NAND2_X1 U13000 ( .A1(n10254), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n10253) );
  INV_X1 U13001 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10250) );
  OR2_X1 U13002 ( .A1(n10255), .A2(n10250), .ZN(n10252) );
  INV_X1 U13003 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10394) );
  OR2_X1 U13004 ( .A1(n9528), .A2(n10394), .ZN(n10251) );
  AND3_X1 U13005 ( .A1(n10253), .A2(n10252), .A3(n10251), .ZN(n10393) );
  NAND2_X1 U13006 ( .A1(n10254), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n10258) );
  INV_X1 U13007 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14978) );
  OR2_X1 U13008 ( .A1(n10255), .A2(n14978), .ZN(n10257) );
  INV_X1 U13009 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15355) );
  OR2_X1 U13010 ( .A1(n9528), .A2(n15355), .ZN(n10256) );
  AND3_X1 U13011 ( .A1(n10258), .A2(n10257), .A3(n10256), .ZN(n14988) );
  AOI21_X1 U13012 ( .B1(n10393), .B2(n10259), .A(n14988), .ZN(n10271) );
  NAND2_X1 U13013 ( .A1(n10262), .A2(n13596), .ZN(n10263) );
  MUX2_X1 U13014 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10801), .Z(n10265) );
  NAND2_X1 U13015 ( .A1(n10265), .A2(SI_30_), .ZN(n10313) );
  OAI21_X1 U13016 ( .B1(n10265), .B2(SI_30_), .A(n10313), .ZN(n10266) );
  NAND2_X1 U13017 ( .A1(n10267), .A2(n10266), .ZN(n10268) );
  NAND2_X1 U13018 ( .A1(n6431), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n10269) );
  MUX2_X1 U13019 ( .A(n10271), .B(n10333), .S(n10281), .Z(n10288) );
  INV_X1 U13020 ( .A(n10393), .ZN(n14832) );
  NAND2_X1 U13021 ( .A1(n10281), .A2(n14832), .ZN(n10327) );
  AOI21_X1 U13022 ( .B1(n10327), .B2(n10272), .A(n14988), .ZN(n10273) );
  AOI21_X1 U13023 ( .B1(n10333), .B2(n7046), .A(n10273), .ZN(n10294) );
  NAND2_X1 U13024 ( .A1(n10288), .A2(n10294), .ZN(n10278) );
  INV_X1 U13025 ( .A(n15242), .ZN(n15237) );
  NAND2_X1 U13026 ( .A1(n10274), .A2(n10318), .ZN(n10276) );
  NAND2_X1 U13027 ( .A1(n6431), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n10275) );
  INV_X1 U13028 ( .A(n15246), .ZN(n14986) );
  MUX2_X1 U13029 ( .A(n15242), .B(n15246), .S(n10281), .Z(n10289) );
  NAND2_X1 U13030 ( .A1(n10290), .A2(n10289), .ZN(n10277) );
  NAND2_X1 U13031 ( .A1(n10278), .A2(n10277), .ZN(n10304) );
  MUX2_X1 U13032 ( .A(n15243), .B(n15244), .S(n10281), .Z(n10305) );
  AND2_X1 U13033 ( .A1(n10306), .A2(n10305), .ZN(n10279) );
  MUX2_X1 U13034 ( .A(n14816), .B(n15023), .S(n10139), .Z(n10300) );
  MUX2_X1 U13035 ( .A(n14833), .B(n15258), .S(n10281), .Z(n10299) );
  NAND2_X1 U13036 ( .A1(n10300), .A2(n10299), .ZN(n10280) );
  MUX2_X1 U13037 ( .A(n15012), .B(n12868), .S(n10139), .Z(n10286) );
  MUX2_X1 U13038 ( .A(n14834), .B(n15264), .S(n10281), .Z(n10285) );
  AND2_X1 U13039 ( .A1(n10286), .A2(n10285), .ZN(n10282) );
  INV_X1 U13040 ( .A(n10288), .ZN(n10298) );
  INV_X1 U13041 ( .A(n10289), .ZN(n10292) );
  INV_X1 U13042 ( .A(n10290), .ZN(n10291) );
  NAND2_X1 U13043 ( .A1(n10292), .A2(n10291), .ZN(n10293) );
  NAND2_X1 U13044 ( .A1(n10293), .A2(n10294), .ZN(n10297) );
  INV_X1 U13045 ( .A(n10293), .ZN(n10296) );
  INV_X1 U13046 ( .A(n10294), .ZN(n10295) );
  AOI22_X1 U13047 ( .A1(n10298), .A2(n10297), .B1(n10296), .B2(n10295), .ZN(
        n10312) );
  INV_X1 U13048 ( .A(n10299), .ZN(n10302) );
  INV_X1 U13049 ( .A(n10300), .ZN(n10301) );
  NAND3_X1 U13050 ( .A1(n10303), .A2(n10302), .A3(n10301), .ZN(n10311) );
  INV_X1 U13051 ( .A(n10304), .ZN(n10309) );
  INV_X1 U13052 ( .A(n10305), .ZN(n10308) );
  INV_X1 U13053 ( .A(n10306), .ZN(n10307) );
  NAND3_X1 U13054 ( .A1(n10309), .A2(n10308), .A3(n10307), .ZN(n10310) );
  MUX2_X1 U13055 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10801), .Z(n10315) );
  XNOR2_X1 U13056 ( .A(n10315), .B(SI_31_), .ZN(n10316) );
  NAND2_X1 U13057 ( .A1(n6431), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10320) );
  XNOR2_X1 U13058 ( .A(n10395), .B(n14832), .ZN(n10352) );
  NAND2_X1 U13059 ( .A1(n10419), .A2(n9877), .ZN(n11905) );
  NAND2_X1 U13060 ( .A1(n10654), .A2(n10321), .ZN(n10322) );
  NAND2_X1 U13061 ( .A1(n11905), .A2(n10322), .ZN(n10332) );
  INV_X1 U13062 ( .A(n10332), .ZN(n10323) );
  INV_X1 U13063 ( .A(n10352), .ZN(n10326) );
  OR2_X1 U13064 ( .A1(n10324), .A2(n6435), .ZN(n10354) );
  NAND2_X1 U13065 ( .A1(n10332), .A2(n10354), .ZN(n10358) );
  INV_X1 U13066 ( .A(n10358), .ZN(n10325) );
  NAND2_X1 U13067 ( .A1(n10326), .A2(n10325), .ZN(n10331) );
  INV_X1 U13068 ( .A(n10327), .ZN(n10328) );
  NOR2_X1 U13069 ( .A1(n10329), .A2(n10328), .ZN(n10359) );
  INV_X1 U13070 ( .A(n10359), .ZN(n10330) );
  MUX2_X1 U13071 ( .A(n10332), .B(n10331), .S(n10330), .Z(n10357) );
  XNOR2_X1 U13072 ( .A(n10333), .B(n14988), .ZN(n10351) );
  XNOR2_X1 U13073 ( .A(n15246), .B(n15242), .ZN(n15235) );
  INV_X1 U13074 ( .A(n15235), .ZN(n15252) );
  INV_X1 U13075 ( .A(n12648), .ZN(n12651) );
  NAND4_X1 U13076 ( .A1(n7392), .A2(n10335), .A3(n10334), .A4(n15476), .ZN(
        n10336) );
  NOR2_X1 U13077 ( .A1(n10336), .A2(n11274), .ZN(n10338) );
  INV_X1 U13078 ( .A(n10337), .ZN(n11803) );
  XNOR2_X1 U13079 ( .A(n11952), .B(n11805), .ZN(n11801) );
  NAND4_X1 U13080 ( .A1(n10339), .A2(n10338), .A3(n11803), .A4(n11801), .ZN(
        n10340) );
  NOR2_X1 U13081 ( .A1(n12074), .A2(n10340), .ZN(n10341) );
  AND4_X1 U13082 ( .A1(n10342), .A2(n10341), .A3(n12160), .A4(n6861), .ZN(
        n10343) );
  NAND3_X1 U13083 ( .A1(n12546), .A2(n10343), .A3(n12317), .ZN(n10344) );
  OR4_X1 U13084 ( .A1(n15164), .A2(n12651), .A3(n15183), .A4(n10344), .ZN(
        n10345) );
  NOR4_X1 U13085 ( .A1(n15029), .A2(n7424), .A3(n15075), .A4(n10346), .ZN(
        n10348) );
  NAND4_X1 U13086 ( .A1(n10348), .A2(n12866), .A3(n10349), .A4(n10347), .ZN(
        n10350) );
  NOR4_X1 U13087 ( .A1(n10351), .A2(n15252), .A3(n15010), .A4(n10350), .ZN(
        n10353) );
  INV_X1 U13088 ( .A(n10354), .ZN(n10355) );
  INV_X1 U13089 ( .A(n10833), .ZN(n10361) );
  NAND2_X1 U13090 ( .A1(n10361), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12375) );
  INV_X1 U13091 ( .A(n12375), .ZN(n10362) );
  NOR2_X1 U13092 ( .A1(n10363), .A2(P1_U3086), .ZN(n12710) );
  NAND3_X1 U13093 ( .A1(n10670), .A2(n15190), .A3(n12710), .ZN(n10364) );
  OAI211_X1 U13094 ( .C1(n15403), .C2(n12375), .A(n10364), .B(P1_B_REG_SCAN_IN), .ZN(n10365) );
  INV_X1 U13095 ( .A(n11902), .ZN(n10366) );
  INV_X1 U13096 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10369) );
  NOR2_X1 U13097 ( .A1(n15512), .A2(n10369), .ZN(n10370) );
  INV_X1 U13098 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10387) );
  NAND2_X1 U13099 ( .A1(n14666), .A2(n7072), .ZN(n10378) );
  INV_X1 U13100 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14669) );
  INV_X1 U13101 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10383) );
  NAND2_X1 U13102 ( .A1(n10379), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n10382) );
  INV_X1 U13103 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n12829) );
  OR2_X1 U13104 ( .A1(n10380), .A2(n12829), .ZN(n10381) );
  OAI211_X1 U13105 ( .C1(n7040), .C2(n10383), .A(n10382), .B(n10381), .ZN(
        n14079) );
  AND2_X1 U13106 ( .A1(n14079), .A2(n10384), .ZN(n12839) );
  NOR2_X1 U13107 ( .A1(n14284), .A2(n12839), .ZN(n12828) );
  AND2_X2 U13108 ( .A1(n10386), .A2(n10385), .ZN(n15572) );
  MUX2_X1 U13109 ( .A(n10387), .B(n12828), .S(n15572), .Z(n10390) );
  NAND2_X1 U13110 ( .A1(n15572), .A2(n15564), .ZN(n14660) );
  NAND2_X1 U13111 ( .A1(n14023), .A2(n10388), .ZN(n10389) );
  NAND2_X1 U13112 ( .A1(n10390), .A2(n10389), .ZN(P2_U3498) );
  XNOR2_X1 U13113 ( .A(n14977), .B(n10395), .ZN(n10391) );
  INV_X1 U13114 ( .A(n10363), .ZN(n10842) );
  NAND2_X1 U13115 ( .A1(n10842), .A2(P1_B_REG_SCAN_IN), .ZN(n10392) );
  NAND2_X1 U13116 ( .A1(n15192), .A2(n10392), .ZN(n14987) );
  NOR2_X1 U13117 ( .A1(n10393), .A2(n14987), .ZN(n14974) );
  NOR2_X1 U13118 ( .A1(n14973), .A2(n14974), .ZN(n15226) );
  MUX2_X1 U13119 ( .A(n10394), .B(n15226), .S(n15512), .Z(n10397) );
  NAND2_X1 U13120 ( .A1(n10395), .A2(n10371), .ZN(n10396) );
  NAND2_X1 U13121 ( .A1(n10397), .A2(n10396), .ZN(P1_U3527) );
  INV_X1 U13122 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10411) );
  OR2_X1 U13123 ( .A1(n12934), .A2(n13081), .ZN(n10398) );
  INV_X1 U13124 ( .A(n13253), .ZN(n13510) );
  NAND2_X1 U13125 ( .A1(n13253), .A2(n13080), .ZN(n10400) );
  NAND2_X1 U13126 ( .A1(n10401), .A2(P3_B_REG_SCAN_IN), .ZN(n10402) );
  NAND2_X1 U13127 ( .A1(n13060), .A2(n10402), .ZN(n13229) );
  NOR2_X1 U13128 ( .A1(n13242), .A2(n10410), .ZN(n12886) );
  NAND2_X1 U13129 ( .A1(n15570), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n10414) );
  INV_X2 U13130 ( .A(n10627), .ZN(n10648) );
  AND2_X4 U13131 ( .A1(n12878), .A2(n6439), .ZN(n10585) );
  NOR2_X1 U13132 ( .A1(n10423), .A2(n10473), .ZN(n10424) );
  AOI21_X1 U13133 ( .B1(n12166), .B2(n10641), .A(n10424), .ZN(n10503) );
  NAND2_X1 U13134 ( .A1(n12166), .A2(n10643), .ZN(n10426) );
  INV_X2 U13135 ( .A(n10627), .ZN(n10641) );
  NAND2_X1 U13136 ( .A1(n14845), .A2(n10641), .ZN(n10425) );
  NAND2_X1 U13137 ( .A1(n10426), .A2(n10425), .ZN(n10428) );
  INV_X2 U13138 ( .A(n10427), .ZN(n10631) );
  XNOR2_X1 U13139 ( .A(n10428), .B(n10631), .ZN(n10502) );
  AOI22_X1 U13140 ( .A1(n11961), .A2(n10641), .B1(n6430), .B2(n14847), .ZN(
        n10495) );
  AOI22_X1 U13141 ( .A1(n11961), .A2(n10643), .B1(n10641), .B2(n14847), .ZN(
        n10429) );
  XNOR2_X1 U13142 ( .A(n10429), .B(n10631), .ZN(n10494) );
  OR2_X1 U13143 ( .A1(n11952), .A2(n10627), .ZN(n10431) );
  NAND2_X1 U13144 ( .A1(n10585), .A2(n14850), .ZN(n10430) );
  NAND2_X1 U13145 ( .A1(n6439), .A2(n11276), .ZN(n10433) );
  NAND2_X1 U13146 ( .A1(n14851), .A2(n6438), .ZN(n10432) );
  NAND2_X1 U13147 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  NAND2_X1 U13148 ( .A1(n10585), .A2(n14851), .ZN(n10436) );
  NAND2_X1 U13149 ( .A1(n11276), .A2(n6438), .ZN(n10435) );
  NAND2_X1 U13150 ( .A1(n10436), .A2(n10435), .ZN(n11604) );
  NAND2_X1 U13151 ( .A1(n10445), .A2(n11604), .ZN(n10438) );
  INV_X1 U13152 ( .A(n10438), .ZN(n10437) );
  NAND2_X1 U13153 ( .A1(n11602), .A2(n10437), .ZN(n10443) );
  NAND2_X1 U13154 ( .A1(n10438), .A2(n10444), .ZN(n10441) );
  OAI22_X1 U13155 ( .A1(n11952), .A2(n10588), .B1(n11805), .B2(n10627), .ZN(
        n10440) );
  XNOR2_X1 U13156 ( .A(n10440), .B(n10449), .ZN(n11601) );
  NAND2_X1 U13157 ( .A1(n10441), .A2(n11601), .ZN(n10442) );
  NOR2_X1 U13158 ( .A1(n11601), .A2(n11602), .ZN(n11600) );
  INV_X1 U13159 ( .A(n10445), .ZN(n10446) );
  INV_X1 U13160 ( .A(n11604), .ZN(n11519) );
  OAI22_X1 U13161 ( .A1(n11922), .A2(n10588), .B1(n11938), .B2(n10628), .ZN(
        n10450) );
  XNOR2_X1 U13162 ( .A(n10450), .B(n10427), .ZN(n10484) );
  OR2_X1 U13163 ( .A1(n11922), .A2(n10627), .ZN(n10452) );
  NAND2_X1 U13164 ( .A1(n6430), .A2(n14849), .ZN(n10451) );
  NAND2_X1 U13165 ( .A1(n10452), .A2(n10451), .ZN(n10485) );
  XNOR2_X1 U13166 ( .A(n10484), .B(n10485), .ZN(n11420) );
  NOR2_X1 U13167 ( .A1(n11987), .A2(n10627), .ZN(n10453) );
  NAND2_X1 U13168 ( .A1(n14855), .A2(n6438), .ZN(n10455) );
  OR2_X1 U13169 ( .A1(n10439), .A2(n11987), .ZN(n10454) );
  OR2_X1 U13170 ( .A1(n10457), .A2(n10458), .ZN(n10459) );
  NAND2_X1 U13171 ( .A1(n10460), .A2(n6438), .ZN(n10462) );
  NAND2_X1 U13172 ( .A1(n10643), .A2(n11203), .ZN(n10461) );
  OAI211_X1 U13173 ( .C1(n10845), .C2(n10421), .A(n10462), .B(n10461), .ZN(
        n11053) );
  OR2_X1 U13174 ( .A1(n11053), .A2(n10427), .ZN(n10463) );
  NAND2_X1 U13175 ( .A1(n14853), .A2(n6438), .ZN(n10466) );
  NAND2_X1 U13176 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  XNOR2_X1 U13177 ( .A(n10467), .B(n10449), .ZN(n10474) );
  NOR2_X1 U13178 ( .A1(n6845), .A2(n10627), .ZN(n10468) );
  AOI21_X1 U13179 ( .B1(n6430), .B2(n14853), .A(n10468), .ZN(n10475) );
  XNOR2_X1 U13180 ( .A(n10474), .B(n10475), .ZN(n11362) );
  NAND2_X1 U13181 ( .A1(n14852), .A2(n6438), .ZN(n10471) );
  OR2_X1 U13182 ( .A1(n10439), .A2(n10469), .ZN(n10470) );
  NAND2_X1 U13183 ( .A1(n10471), .A2(n10470), .ZN(n10472) );
  XNOR2_X1 U13184 ( .A(n10472), .B(n10427), .ZN(n10478) );
  INV_X1 U13185 ( .A(n14852), .ZN(n11364) );
  OAI22_X1 U13186 ( .A1(n6436), .A2(n11364), .B1(n10469), .B2(n10627), .ZN(
        n10479) );
  XNOR2_X1 U13187 ( .A(n10478), .B(n10479), .ZN(n11353) );
  INV_X1 U13188 ( .A(n10474), .ZN(n10476) );
  NAND2_X1 U13189 ( .A1(n10476), .A2(n10475), .ZN(n11354) );
  INV_X1 U13190 ( .A(n10478), .ZN(n10480) );
  NAND2_X1 U13191 ( .A1(n10480), .A2(n10479), .ZN(n11415) );
  NAND2_X1 U13192 ( .A1(n11355), .A2(n10481), .ZN(n10482) );
  NAND2_X1 U13193 ( .A1(n10483), .A2(n10482), .ZN(n11419) );
  INV_X1 U13194 ( .A(n10484), .ZN(n10486) );
  NAND2_X1 U13195 ( .A1(n10486), .A2(n10485), .ZN(n10487) );
  NOR2_X1 U13196 ( .A1(n11806), .A2(n10473), .ZN(n10488) );
  AOI21_X1 U13197 ( .B1(n15503), .B2(n10641), .A(n10488), .ZN(n10491) );
  AOI22_X1 U13198 ( .A1(n15503), .A2(n10643), .B1(n10648), .B2(n14848), .ZN(
        n10489) );
  XNOR2_X1 U13199 ( .A(n10489), .B(n10631), .ZN(n10490) );
  XOR2_X1 U13200 ( .A(n10491), .B(n10490), .Z(n11527) );
  NOR2_X1 U13201 ( .A1(n10491), .A2(n10490), .ZN(n10492) );
  XNOR2_X1 U13202 ( .A(n10494), .B(n10495), .ZN(n11709) );
  AOI22_X1 U13203 ( .A1(n12217), .A2(n10641), .B1(n10585), .B2(n14846), .ZN(
        n10500) );
  NAND2_X1 U13204 ( .A1(n12217), .A2(n10643), .ZN(n10497) );
  OR2_X1 U13205 ( .A1(n12162), .A2(n10627), .ZN(n10496) );
  NAND2_X1 U13206 ( .A1(n10497), .A2(n10496), .ZN(n10498) );
  XNOR2_X1 U13207 ( .A(n10498), .B(n10631), .ZN(n10499) );
  XOR2_X1 U13208 ( .A(n10500), .B(n10499), .Z(n12101) );
  INV_X1 U13209 ( .A(n10499), .ZN(n10501) );
  XNOR2_X1 U13210 ( .A(n10502), .B(n10503), .ZN(n12350) );
  NAND2_X1 U13211 ( .A1(n15349), .A2(n10643), .ZN(n10505) );
  NAND2_X1 U13212 ( .A1(n14844), .A2(n10648), .ZN(n10504) );
  NAND2_X1 U13213 ( .A1(n10505), .A2(n10504), .ZN(n10506) );
  XNOR2_X1 U13214 ( .A(n10506), .B(n10449), .ZN(n10507) );
  OAI22_X1 U13215 ( .A1(n12234), .A2(n10627), .B1(n12702), .B2(n10473), .ZN(
        n10508) );
  XNOR2_X1 U13216 ( .A(n10507), .B(n10508), .ZN(n12513) );
  INV_X1 U13217 ( .A(n10507), .ZN(n10510) );
  INV_X1 U13218 ( .A(n10508), .ZN(n10509) );
  NAND2_X1 U13219 ( .A1(n10510), .A2(n10509), .ZN(n10511) );
  NAND2_X1 U13220 ( .A1(n12322), .A2(n10643), .ZN(n10513) );
  NAND2_X1 U13221 ( .A1(n14843), .A2(n10641), .ZN(n10512) );
  NAND2_X1 U13222 ( .A1(n10513), .A2(n10512), .ZN(n10514) );
  XNOR2_X1 U13223 ( .A(n10514), .B(n10631), .ZN(n10519) );
  NOR2_X1 U13224 ( .A1(n10515), .A2(n10473), .ZN(n10516) );
  AOI21_X1 U13225 ( .B1(n12322), .B2(n10641), .A(n10516), .ZN(n10517) );
  XNOR2_X1 U13226 ( .A(n10519), .B(n10517), .ZN(n12698) );
  INV_X1 U13227 ( .A(n10517), .ZN(n10518) );
  NAND2_X1 U13228 ( .A1(n10519), .A2(n10518), .ZN(n10520) );
  NOR2_X1 U13229 ( .A1(n12701), .A2(n10473), .ZN(n10521) );
  AOI21_X1 U13230 ( .B1(n12552), .B2(n10648), .A(n10521), .ZN(n10524) );
  AOI22_X1 U13231 ( .A1(n12552), .A2(n10643), .B1(n10648), .B2(n14842), .ZN(
        n10522) );
  XNOR2_X1 U13232 ( .A(n10522), .B(n10449), .ZN(n10523) );
  XOR2_X1 U13233 ( .A(n10524), .B(n10523), .Z(n14776) );
  INV_X1 U13234 ( .A(n10523), .ZN(n10526) );
  INV_X1 U13235 ( .A(n10524), .ZN(n10525) );
  NAND2_X1 U13236 ( .A1(n10526), .A2(n10525), .ZN(n10527) );
  AOI22_X1 U13237 ( .A1(n15338), .A2(n10641), .B1(n6430), .B2(n14841), .ZN(
        n10531) );
  NAND2_X1 U13238 ( .A1(n15338), .A2(n10643), .ZN(n10529) );
  NAND2_X1 U13239 ( .A1(n14841), .A2(n10641), .ZN(n10528) );
  NAND2_X1 U13240 ( .A1(n10529), .A2(n10528), .ZN(n10530) );
  XNOR2_X1 U13241 ( .A(n10530), .B(n10449), .ZN(n10533) );
  XOR2_X1 U13242 ( .A(n10531), .B(n10533), .Z(n14691) );
  INV_X1 U13243 ( .A(n10531), .ZN(n10532) );
  OR2_X1 U13244 ( .A1(n10533), .A2(n10532), .ZN(n10534) );
  NAND2_X1 U13245 ( .A1(n15213), .A2(n10643), .ZN(n10536) );
  NAND2_X1 U13246 ( .A1(n15191), .A2(n10641), .ZN(n10535) );
  NAND2_X1 U13247 ( .A1(n10536), .A2(n10535), .ZN(n10537) );
  XNOR2_X1 U13248 ( .A(n10537), .B(n10631), .ZN(n14741) );
  NAND2_X1 U13249 ( .A1(n15213), .A2(n10648), .ZN(n10539) );
  NAND2_X1 U13250 ( .A1(n15191), .A2(n10585), .ZN(n10538) );
  NAND2_X1 U13251 ( .A1(n10539), .A2(n10538), .ZN(n10547) );
  NAND2_X1 U13252 ( .A1(n15188), .A2(n10643), .ZN(n10541) );
  OR2_X1 U13253 ( .A1(n15167), .A2(n10627), .ZN(n10540) );
  NAND2_X1 U13254 ( .A1(n10541), .A2(n10540), .ZN(n10542) );
  XNOR2_X1 U13255 ( .A(n10542), .B(n10631), .ZN(n14739) );
  NAND2_X1 U13256 ( .A1(n15188), .A2(n10648), .ZN(n10544) );
  OR2_X1 U13257 ( .A1(n15167), .A2(n10473), .ZN(n10543) );
  NAND2_X1 U13258 ( .A1(n10544), .A2(n10543), .ZN(n10549) );
  AND2_X1 U13259 ( .A1(n14739), .A2(n10549), .ZN(n10546) );
  AOI21_X1 U13260 ( .B1(n14741), .B2(n10547), .A(n10546), .ZN(n10545) );
  NAND2_X1 U13261 ( .A1(n14740), .A2(n10545), .ZN(n10554) );
  INV_X1 U13262 ( .A(n10546), .ZN(n10548) );
  INV_X1 U13263 ( .A(n10547), .ZN(n14828) );
  NAND2_X1 U13264 ( .A1(n10548), .A2(n14828), .ZN(n10551) );
  INV_X1 U13265 ( .A(n14739), .ZN(n10550) );
  INV_X1 U13266 ( .A(n10549), .ZN(n14738) );
  NAND2_X1 U13267 ( .A1(n10550), .A2(n14738), .ZN(n14754) );
  OAI21_X1 U13268 ( .B1(n14741), .B2(n10551), .A(n14754), .ZN(n10552) );
  INV_X1 U13269 ( .A(n10552), .ZN(n10553) );
  NAND2_X1 U13270 ( .A1(n10554), .A2(n10553), .ZN(n10560) );
  NAND2_X1 U13271 ( .A1(n15319), .A2(n10643), .ZN(n10556) );
  NAND2_X1 U13272 ( .A1(n15193), .A2(n10641), .ZN(n10555) );
  NAND2_X1 U13273 ( .A1(n10556), .A2(n10555), .ZN(n10557) );
  XNOR2_X1 U13274 ( .A(n10557), .B(n10427), .ZN(n10562) );
  AND2_X1 U13275 ( .A1(n15193), .A2(n6430), .ZN(n10558) );
  AOI21_X1 U13276 ( .B1(n15319), .B2(n10648), .A(n10558), .ZN(n10561) );
  XNOR2_X1 U13277 ( .A(n10562), .B(n10561), .ZN(n14753) );
  NAND2_X1 U13278 ( .A1(n10562), .A2(n10561), .ZN(n10563) );
  NAND2_X1 U13279 ( .A1(n15149), .A2(n10643), .ZN(n10565) );
  NAND2_X1 U13280 ( .A1(n15125), .A2(n10648), .ZN(n10564) );
  NAND2_X1 U13281 ( .A1(n10565), .A2(n10564), .ZN(n10566) );
  XNOR2_X1 U13282 ( .A(n10566), .B(n10631), .ZN(n10567) );
  AOI22_X1 U13283 ( .A1(n15149), .A2(n10641), .B1(n6430), .B2(n15125), .ZN(
        n10568) );
  XNOR2_X1 U13284 ( .A(n10567), .B(n10568), .ZN(n14799) );
  INV_X1 U13285 ( .A(n10567), .ZN(n10569) );
  NAND2_X1 U13286 ( .A1(n10569), .A2(n10568), .ZN(n10570) );
  AND2_X1 U13287 ( .A1(n14839), .A2(n10585), .ZN(n10571) );
  AOI21_X1 U13288 ( .B1(n15307), .B2(n10641), .A(n10571), .ZN(n10575) );
  NAND2_X1 U13289 ( .A1(n15307), .A2(n10643), .ZN(n10573) );
  NAND2_X1 U13290 ( .A1(n14839), .A2(n10641), .ZN(n10572) );
  NAND2_X1 U13291 ( .A1(n10573), .A2(n10572), .ZN(n10574) );
  XNOR2_X1 U13292 ( .A(n10574), .B(n10631), .ZN(n10577) );
  XOR2_X1 U13293 ( .A(n10575), .B(n10577), .Z(n14706) );
  INV_X1 U13294 ( .A(n10575), .ZN(n10576) );
  OAI22_X1 U13295 ( .A1(n15375), .A2(n10439), .B1(n15089), .B2(n10627), .ZN(
        n10578) );
  XNOR2_X1 U13296 ( .A(n10578), .B(n10631), .ZN(n10580) );
  NOR2_X1 U13297 ( .A1(n15089), .A2(n10473), .ZN(n10579) );
  AOI21_X1 U13298 ( .B1(n15115), .B2(n10648), .A(n10579), .ZN(n10581) );
  XNOR2_X1 U13299 ( .A(n10580), .B(n10581), .ZN(n14770) );
  INV_X1 U13300 ( .A(n10580), .ZN(n10582) );
  OR2_X1 U13301 ( .A1(n10582), .A2(n10581), .ZN(n10583) );
  AOI22_X1 U13302 ( .A1(n15099), .A2(n10643), .B1(n10648), .B2(n15069), .ZN(
        n10584) );
  XNOR2_X1 U13303 ( .A(n10584), .B(n10631), .ZN(n10591) );
  AOI22_X1 U13304 ( .A1(n15099), .A2(n10648), .B1(n10585), .B2(n15069), .ZN(
        n10590) );
  XNOR2_X1 U13305 ( .A(n10591), .B(n10590), .ZN(n14725) );
  OR2_X1 U13306 ( .A1(n15370), .A2(n10628), .ZN(n10587) );
  NAND2_X1 U13307 ( .A1(n14838), .A2(n6430), .ZN(n10586) );
  NAND2_X1 U13308 ( .A1(n10587), .A2(n10586), .ZN(n10596) );
  OAI22_X1 U13309 ( .A1(n15370), .A2(n10588), .B1(n15090), .B2(n10627), .ZN(
        n10589) );
  XNOR2_X1 U13310 ( .A(n10589), .B(n10631), .ZN(n10595) );
  XOR2_X1 U13311 ( .A(n10596), .B(n10595), .Z(n14790) );
  INV_X1 U13312 ( .A(n14790), .ZN(n10592) );
  NAND2_X1 U13313 ( .A1(n10591), .A2(n10590), .ZN(n14786) );
  OR2_X1 U13314 ( .A1(n10592), .A2(n14786), .ZN(n10593) );
  INV_X1 U13315 ( .A(n10595), .ZN(n10598) );
  INV_X1 U13316 ( .A(n10596), .ZN(n10597) );
  OAI22_X1 U13317 ( .A1(n10599), .A2(n10628), .B1(n15072), .B2(n10473), .ZN(
        n10604) );
  NAND2_X1 U13318 ( .A1(n15282), .A2(n10643), .ZN(n10601) );
  NAND2_X1 U13319 ( .A1(n14837), .A2(n10641), .ZN(n10600) );
  NAND2_X1 U13320 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  XNOR2_X1 U13321 ( .A(n10602), .B(n10631), .ZN(n10603) );
  XOR2_X1 U13322 ( .A(n10604), .B(n10603), .Z(n14700) );
  NAND2_X1 U13323 ( .A1(n14699), .A2(n14700), .ZN(n10608) );
  INV_X1 U13324 ( .A(n10603), .ZN(n10606) );
  INV_X1 U13325 ( .A(n10604), .ZN(n10605) );
  NAND2_X1 U13326 ( .A1(n10606), .A2(n10605), .ZN(n10607) );
  OAI22_X1 U13327 ( .A1(n15365), .A2(n10627), .B1(n10609), .B2(n10473), .ZN(
        n10614) );
  NAND2_X1 U13328 ( .A1(n15049), .A2(n6439), .ZN(n10611) );
  NAND2_X1 U13329 ( .A1(n14836), .A2(n10641), .ZN(n10610) );
  NAND2_X1 U13330 ( .A1(n10611), .A2(n10610), .ZN(n10612) );
  XNOR2_X1 U13331 ( .A(n10612), .B(n10631), .ZN(n10613) );
  XOR2_X1 U13332 ( .A(n10614), .B(n10613), .Z(n14762) );
  INV_X1 U13333 ( .A(n10613), .ZN(n10616) );
  INV_X1 U13334 ( .A(n10614), .ZN(n10615) );
  NAND2_X1 U13335 ( .A1(n10616), .A2(n10615), .ZN(n10617) );
  OAI22_X1 U13336 ( .A1(n15270), .A2(n10627), .B1(n15045), .B2(n10473), .ZN(
        n10623) );
  NAND2_X1 U13337 ( .A1(n15035), .A2(n6439), .ZN(n10620) );
  NAND2_X1 U13338 ( .A1(n14835), .A2(n10648), .ZN(n10619) );
  NAND2_X1 U13339 ( .A1(n10620), .A2(n10619), .ZN(n10621) );
  XNOR2_X1 U13340 ( .A(n10621), .B(n10631), .ZN(n10622) );
  XOR2_X1 U13341 ( .A(n10623), .B(n10622), .Z(n14732) );
  INV_X1 U13342 ( .A(n10622), .ZN(n10625) );
  INV_X1 U13343 ( .A(n10623), .ZN(n10624) );
  NAND2_X1 U13344 ( .A1(n10625), .A2(n10624), .ZN(n10626) );
  OAI22_X1 U13345 ( .A1(n12868), .A2(n10627), .B1(n15012), .B2(n10473), .ZN(
        n10634) );
  NAND2_X1 U13346 ( .A1(n15264), .A2(n10643), .ZN(n10630) );
  OR2_X1 U13347 ( .A1(n15012), .A2(n10627), .ZN(n10629) );
  NAND2_X1 U13348 ( .A1(n10630), .A2(n10629), .ZN(n10632) );
  XNOR2_X1 U13349 ( .A(n10632), .B(n10631), .ZN(n10633) );
  XOR2_X1 U13350 ( .A(n10634), .B(n10633), .Z(n14809) );
  INV_X1 U13351 ( .A(n10633), .ZN(n10636) );
  INV_X1 U13352 ( .A(n10634), .ZN(n10635) );
  NAND2_X1 U13353 ( .A1(n15258), .A2(n10643), .ZN(n10638) );
  NAND2_X1 U13354 ( .A1(n14833), .A2(n6438), .ZN(n10637) );
  NAND2_X1 U13355 ( .A1(n10638), .A2(n10637), .ZN(n10639) );
  XNOR2_X1 U13356 ( .A(n10639), .B(n10427), .ZN(n10660) );
  NOR2_X1 U13357 ( .A1(n14816), .A2(n10473), .ZN(n10640) );
  AOI21_X1 U13358 ( .B1(n15258), .B2(n10648), .A(n10640), .ZN(n10659) );
  XNOR2_X1 U13359 ( .A(n10660), .B(n10659), .ZN(n12814) );
  INV_X1 U13360 ( .A(n12814), .ZN(n10642) );
  INV_X1 U13361 ( .A(n10661), .ZN(n10658) );
  NAND2_X1 U13362 ( .A1(n15244), .A2(n10643), .ZN(n10645) );
  NAND2_X1 U13363 ( .A1(n15243), .A2(n10648), .ZN(n10644) );
  NAND2_X1 U13364 ( .A1(n10645), .A2(n10644), .ZN(n10646) );
  XNOR2_X1 U13365 ( .A(n10646), .B(n10427), .ZN(n10650) );
  NOR2_X1 U13366 ( .A1(n15013), .A2(n10473), .ZN(n10647) );
  AOI21_X1 U13367 ( .B1(n15244), .B2(n6438), .A(n10647), .ZN(n10649) );
  XNOR2_X1 U13368 ( .A(n10650), .B(n10649), .ZN(n10675) );
  INV_X1 U13369 ( .A(n10675), .ZN(n10657) );
  INV_X1 U13370 ( .A(n15791), .ZN(n10652) );
  NAND3_X1 U13371 ( .A1(n10652), .A2(n11902), .A3(n10651), .ZN(n10669) );
  AND2_X1 U13372 ( .A1(n10421), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10653) );
  INV_X1 U13373 ( .A(n15790), .ZN(n10720) );
  OR2_X1 U13374 ( .A1(n10669), .A2(n10720), .ZN(n10667) );
  INV_X1 U13375 ( .A(n10667), .ZN(n10656) );
  AND2_X1 U13376 ( .A1(n15489), .A2(n10654), .ZN(n10655) );
  NAND2_X1 U13377 ( .A1(n10658), .A2(n7801), .ZN(n10680) );
  NAND2_X1 U13378 ( .A1(n10660), .A2(n10659), .ZN(n10674) );
  NAND4_X1 U13379 ( .A1(n10661), .A2(n14801), .A3(n10675), .A4(n10674), .ZN(
        n10679) );
  NOR2_X1 U13380 ( .A1(n9962), .A2(n6435), .ZN(n11909) );
  INV_X1 U13381 ( .A(n11909), .ZN(n10663) );
  INV_X1 U13382 ( .A(n10668), .ZN(n10662) );
  INV_X1 U13383 ( .A(n10665), .ZN(n10666) );
  INV_X1 U13384 ( .A(n14812), .ZN(n14804) );
  NAND2_X1 U13385 ( .A1(n14822), .A2(n15192), .ZN(n14815) );
  INV_X1 U13386 ( .A(n14815), .ZN(n14751) );
  AOI22_X1 U13387 ( .A1(n15242), .A2(n14751), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10673) );
  NAND2_X1 U13388 ( .A1(n10669), .A2(n10668), .ZN(n10671) );
  NAND2_X1 U13389 ( .A1(n10671), .A2(n10670), .ZN(n11051) );
  NAND2_X1 U13390 ( .A1(n11051), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14824) );
  NAND2_X1 U13391 ( .A1(n12889), .A2(n14810), .ZN(n10672) );
  OAI211_X1 U13392 ( .C1(n14816), .C2(n14804), .A(n10673), .B(n10672), .ZN(
        n10677) );
  NOR3_X1 U13393 ( .A1(n10675), .A2(n14826), .A3(n10674), .ZN(n10676) );
  AOI211_X1 U13394 ( .C1(n10664), .C2(n15244), .A(n10677), .B(n10676), .ZN(
        n10678) );
  NAND3_X1 U13395 ( .A1(n10680), .A2(n10679), .A3(n10678), .ZN(P1_U3220) );
  INV_X1 U13396 ( .A(n12399), .ZN(n10681) );
  NOR2_X1 U13397 ( .A1(n10682), .A2(n10681), .ZN(n10901) );
  NOR2_X1 U13398 ( .A1(n10421), .A2(P1_U3086), .ZN(n10683) );
  NAND3_X1 U13399 ( .A1(n13131), .A2(n10685), .A3(n10684), .ZN(n10686) );
  AOI21_X1 U13400 ( .B1(n10687), .B2(n10686), .A(n13165), .ZN(n10701) );
  NAND3_X1 U13401 ( .A1(n10688), .A2(n10690), .A3(n10689), .ZN(n10691) );
  AOI21_X1 U13402 ( .B1(n10692), .B2(n10691), .A(n13200), .ZN(n10700) );
  AOI211_X1 U13403 ( .C1(n10695), .C2(n10694), .A(n13226), .B(n10693), .ZN(
        n10699) );
  INV_X1 U13404 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15413) );
  NAND2_X1 U13405 ( .A1(n13212), .A2(n10696), .ZN(n10697) );
  NAND2_X1 U13406 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12692)
         );
  OAI211_X1 U13407 ( .C1(n13215), .C2(n15413), .A(n10697), .B(n12692), .ZN(
        n10698) );
  INV_X1 U13408 ( .A(n10702), .ZN(n10704) );
  NAND3_X1 U13409 ( .A1(n11895), .A2(n10704), .A3(n10703), .ZN(n10705) );
  AOI21_X1 U13410 ( .B1(n10706), .B2(n10705), .A(n13200), .ZN(n10718) );
  INV_X1 U13411 ( .A(n10707), .ZN(n10710) );
  NAND3_X1 U13412 ( .A1(n11883), .A2(n11887), .A3(n10708), .ZN(n10709) );
  AOI21_X1 U13413 ( .B1(n10710), .B2(n10709), .A(n13226), .ZN(n10717) );
  NAND3_X1 U13414 ( .A1(n11889), .A2(n10711), .A3(n7346), .ZN(n10712) );
  AOI21_X1 U13415 ( .B1(n6836), .B2(n10712), .A(n13165), .ZN(n10716) );
  INV_X1 U13416 ( .A(n13212), .ZN(n13195) );
  NAND2_X1 U13417 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n10714)
         );
  NAND2_X1 U13418 ( .A1(n15575), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n10713) );
  OAI211_X1 U13419 ( .C1(n13195), .C2(n10800), .A(n10714), .B(n10713), .ZN(
        n10715) );
  OR4_X1 U13420 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        P3_U3192) );
  NAND2_X1 U13421 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10723) );
  INV_X1 U13422 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10719) );
  XNOR2_X1 U13423 ( .A(n10929), .B(n10719), .ZN(n10722) );
  NAND2_X1 U13424 ( .A1(n10720), .A2(n12375), .ZN(n10730) );
  AOI21_X1 U13425 ( .B1(n10721), .B2(n10833), .A(n9534), .ZN(n10728) );
  NAND2_X1 U13426 ( .A1(n10730), .A2(n10728), .ZN(n10727) );
  INV_X1 U13427 ( .A(n10727), .ZN(n10848) );
  AND2_X1 U13428 ( .A1(n10848), .A2(n10363), .ZN(n14965) );
  AOI211_X1 U13429 ( .C1(n10723), .C2(n10722), .A(n10923), .B(n14940), .ZN(
        n10734) );
  NAND2_X1 U13430 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n11240) );
  MUX2_X1 U13431 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n11993), .S(n10929), .Z(
        n10726) );
  INV_X1 U13432 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10724) );
  NOR3_X1 U13433 ( .A1(n10726), .A2(n10724), .A3(n11244), .ZN(n11245) );
  NAND2_X1 U13434 ( .A1(n10844), .A2(n10842), .ZN(n10725) );
  OR2_X1 U13435 ( .A1(n10727), .A2(n10725), .ZN(n14960) );
  AOI211_X1 U13436 ( .C1(n11240), .C2(n10726), .A(n11245), .B(n14960), .ZN(
        n10733) );
  NOR2_X1 U13437 ( .A1(n14959), .A2(n10929), .ZN(n10732) );
  INV_X1 U13438 ( .A(n10728), .ZN(n10729) );
  NAND2_X1 U13439 ( .A1(n10730), .A2(n10729), .ZN(n14972) );
  OAI22_X1 U13440 ( .A1(n14972), .A2(n10747), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15727), .ZN(n10731) );
  OR4_X1 U13441 ( .A1(n10734), .A2(n10733), .A3(n10732), .A4(n10731), .ZN(
        P1_U3244) );
  INV_X1 U13442 ( .A(n10745), .ZN(n10737) );
  XNOR2_X1 U13443 ( .A(n10746), .B(n10737), .ZN(n10741) );
  XNOR2_X1 U13444 ( .A(n10741), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n10739) );
  INV_X1 U13445 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10735) );
  NAND2_X1 U13446 ( .A1(n10735), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n10736) );
  NAND2_X1 U13447 ( .A1(n10737), .A2(n10736), .ZN(n15406) );
  AND2_X1 U13448 ( .A1(n15406), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n10738) );
  NAND2_X1 U13449 ( .A1(n10739), .A2(n10738), .ZN(n10744) );
  OAI21_X1 U13450 ( .B1(n10739), .B2(n10738), .A(n10744), .ZN(n10740) );
  INV_X1 U13451 ( .A(n10740), .ZN(SUB_1596_U5) );
  INV_X1 U13452 ( .A(n10741), .ZN(n10742) );
  NAND2_X1 U13453 ( .A1(n10742), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10743) );
  NAND2_X1 U13454 ( .A1(n10744), .A2(n10743), .ZN(n10755) );
  NAND2_X1 U13455 ( .A1(n10746), .A2(n10745), .ZN(n10749) );
  NAND2_X1 U13456 ( .A1(n10747), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10748) );
  NAND2_X1 U13457 ( .A1(n10749), .A2(n10748), .ZN(n10762) );
  NAND2_X1 U13458 ( .A1(n10750), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10763) );
  INV_X1 U13459 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10751) );
  NAND2_X1 U13460 ( .A1(n10751), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10752) );
  XNOR2_X1 U13461 ( .A(n10762), .B(n10761), .ZN(n10756) );
  XNOR2_X1 U13462 ( .A(n10756), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(n10753) );
  XNOR2_X1 U13463 ( .A(n10755), .B(n10753), .ZN(SUB_1596_U61) );
  AND2_X1 U13464 ( .A1(n10756), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10754) );
  OR2_X1 U13465 ( .A1(n10755), .A2(n10754), .ZN(n10760) );
  INV_X1 U13466 ( .A(n10756), .ZN(n10758) );
  INV_X1 U13467 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10757) );
  NAND2_X1 U13468 ( .A1(n10758), .A2(n10757), .ZN(n10759) );
  NAND2_X1 U13469 ( .A1(n10760), .A2(n10759), .ZN(n10771) );
  INV_X1 U13470 ( .A(n10771), .ZN(n10769) );
  NAND2_X1 U13471 ( .A1(n10762), .A2(n10761), .ZN(n10764) );
  NAND2_X1 U13472 ( .A1(n10764), .A2(n10763), .ZN(n10765) );
  NAND2_X1 U13473 ( .A1(n10765), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10773) );
  INV_X1 U13474 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10767) );
  XNOR2_X1 U13475 ( .A(n10774), .B(n10767), .ZN(n10770) );
  INV_X1 U13476 ( .A(n10770), .ZN(n10768) );
  NAND2_X1 U13477 ( .A1(n10769), .A2(n10768), .ZN(n10779) );
  NAND2_X1 U13478 ( .A1(n10771), .A2(n10770), .ZN(n10778) );
  NAND2_X1 U13479 ( .A1(n10779), .A2(n10778), .ZN(n10772) );
  XNOR2_X1 U13480 ( .A(n10772), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  NAND2_X1 U13481 ( .A1(n10775), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10814) );
  INV_X1 U13482 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10777) );
  NAND2_X1 U13483 ( .A1(n10778), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n10780) );
  NAND2_X1 U13484 ( .A1(n10780), .A2(n10779), .ZN(n10781) );
  NAND2_X1 U13485 ( .A1(n10782), .A2(n10781), .ZN(n10813) );
  OAI21_X1 U13486 ( .B1(n10782), .B2(n10781), .A(n10813), .ZN(n10783) );
  INV_X1 U13487 ( .A(n10783), .ZN(SUB_1596_U59) );
  NOR2_X1 U13488 ( .A1(n10801), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13585) );
  INV_X1 U13489 ( .A(n13585), .ZN(n13610) );
  NAND2_X1 U13490 ( .A1(n10801), .A2(P3_U3151), .ZN(n13598) );
  OAI222_X1 U13491 ( .A1(P3_U3151), .A2(n10786), .B1(n13610), .B2(n10785), 
        .C1(n10784), .C2(n13598), .ZN(P3_U3295) );
  OAI222_X1 U13492 ( .A1(P3_U3151), .A2(n10788), .B1(n13598), .B2(n6998), .C1(
        n13610), .C2(n10787), .ZN(P3_U3287) );
  INV_X1 U13493 ( .A(SI_7_), .ZN(n10790) );
  OAI222_X1 U13494 ( .A1(P3_U3151), .A2(n6916), .B1(n13598), .B2(n10790), .C1(
        n13610), .C2(n10789), .ZN(P3_U3288) );
  OAI222_X1 U13495 ( .A1(P3_U3151), .A2(n9173), .B1(n13598), .B2(n10792), .C1(
        n13610), .C2(n10791), .ZN(P3_U3294) );
  OAI222_X1 U13496 ( .A1(P3_U3151), .A2(n11891), .B1(n13598), .B2(n10794), 
        .C1(n13610), .C2(n10793), .ZN(P3_U3286) );
  INV_X1 U13497 ( .A(n14868), .ZN(n10797) );
  INV_X1 U13498 ( .A(n10795), .ZN(n10855) );
  OAI222_X1 U13499 ( .A1(P1_U3086), .A2(n10797), .B1(n15400), .B2(n10855), 
        .C1(n10796), .C2(n15397), .ZN(P1_U3351) );
  OAI222_X1 U13500 ( .A1(P3_U3151), .A2(n10800), .B1(n13598), .B2(n10799), 
        .C1(n13610), .C2(n10798), .ZN(P3_U3285) );
  NAND2_X1 U13501 ( .A1(n10801), .A2(P2_U3088), .ZN(n14673) );
  INV_X1 U13502 ( .A(n10802), .ZN(n10822) );
  OAI222_X1 U13503 ( .A1(n14682), .A2(n10803), .B1(n14673), .B2(n10822), .C1(
        n14113), .C2(P2_U3088), .ZN(P2_U3326) );
  INV_X1 U13504 ( .A(n13598), .ZN(n10920) );
  AOI222_X1 U13505 ( .A1(n10804), .A2(n13585), .B1(SI_4_), .B2(n10920), .C1(
        n11236), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10805) );
  INV_X1 U13506 ( .A(n10805), .ZN(P3_U3291) );
  AOI222_X1 U13507 ( .A1(n10806), .A2(n13585), .B1(n11145), .B2(
        P3_STATE_REG_SCAN_IN), .C1(n10920), .C2(SI_3_), .ZN(n10807) );
  INV_X1 U13508 ( .A(n10807), .ZN(P3_U3292) );
  AOI222_X1 U13509 ( .A1(n10808), .A2(n13585), .B1(n10920), .B2(SI_2_), .C1(
        n9176), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10809) );
  INV_X1 U13510 ( .A(n10809), .ZN(P3_U3293) );
  INV_X1 U13511 ( .A(n10810), .ZN(n10811) );
  NAND2_X1 U13512 ( .A1(n10811), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U13513 ( .A1(n10813), .A2(n10812), .ZN(n10881) );
  NAND2_X1 U13514 ( .A1(n10816), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10885) );
  INV_X1 U13515 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14877) );
  XNOR2_X1 U13516 ( .A(n10881), .B(n10879), .ZN(n10878) );
  INV_X1 U13517 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10877) );
  XNOR2_X1 U13518 ( .A(n10878), .B(n10877), .ZN(SUB_1596_U58) );
  AOI222_X1 U13519 ( .A1(n10817), .A2(n13585), .B1(n11160), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_5_), .C2(n10920), .ZN(n10818) );
  INV_X1 U13520 ( .A(n10818), .ZN(P3_U3290) );
  INV_X1 U13521 ( .A(n10819), .ZN(n10853) );
  INV_X1 U13522 ( .A(n11247), .ZN(n11257) );
  OAI222_X1 U13523 ( .A1(n15397), .A2(n10820), .B1(n15400), .B2(n10853), .C1(
        n11257), .C2(P1_U3086), .ZN(P1_U3353) );
  NAND2_X1 U13524 ( .A1(n11306), .A2(n10821), .ZN(n10827) );
  AND2_X1 U13525 ( .A1(n10827), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13526 ( .A1(n10827), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U13527 ( .A1(n10827), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13528 ( .A1(n10827), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13529 ( .A1(n10827), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13530 ( .A1(n10827), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13531 ( .A1(n10827), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U13532 ( .A1(n10827), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13533 ( .A1(n10827), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13534 ( .A1(n10827), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U13535 ( .A1(n10827), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13536 ( .A1(n10827), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U13537 ( .A1(n10827), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U13538 ( .A1(n10827), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U13539 ( .A1(n10827), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U13540 ( .A1(n10827), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U13541 ( .A1(n10827), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U13542 ( .A1(n10827), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U13543 ( .A1(n10827), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U13544 ( .A1(n10827), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U13545 ( .A1(n10827), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13546 ( .A1(n10827), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13547 ( .A1(n10827), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13548 ( .A1(n10827), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U13549 ( .A1(n10827), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U13550 ( .A1(n10827), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U13551 ( .A1(n10827), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  OAI222_X1 U13552 ( .A1(P1_U3086), .A2(n10929), .B1(n15400), .B2(n10822), 
        .C1(n7075), .C2(n15397), .ZN(P1_U3354) );
  INV_X1 U13553 ( .A(n10931), .ZN(n10958) );
  INV_X1 U13554 ( .A(n10823), .ZN(n10863) );
  OAI222_X1 U13555 ( .A1(P1_U3086), .A2(n10958), .B1(n15400), .B2(n10863), 
        .C1(n7822), .C2(n15397), .ZN(P1_U3352) );
  AND2_X1 U13556 ( .A1(n14972), .A2(n14854), .ZN(P1_U3085) );
  OAI222_X1 U13557 ( .A1(P3_U3151), .A2(n10826), .B1(n13598), .B2(n10825), 
        .C1(n13610), .C2(n10824), .ZN(P3_U3284) );
  INV_X1 U13558 ( .A(n10827), .ZN(n10828) );
  INV_X1 U13559 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n15754) );
  NOR2_X1 U13560 ( .A1(n10828), .A2(n15754), .ZN(P3_U3243) );
  INV_X1 U13561 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n15668) );
  NOR2_X1 U13562 ( .A1(n10828), .A2(n15668), .ZN(P3_U3236) );
  INV_X1 U13563 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15693) );
  NOR2_X1 U13564 ( .A1(n10828), .A2(n15693), .ZN(P3_U3253) );
  NAND2_X1 U13565 ( .A1(n14854), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10829) );
  OAI21_X1 U13566 ( .B1(n14988), .B2(n14854), .A(n10829), .ZN(P1_U3590) );
  INV_X1 U13567 ( .A(n10830), .ZN(n10831) );
  AND2_X1 U13568 ( .A1(n10832), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13569 ( .A1(n15487), .A2(n10835), .B1(n10834), .B2(n10833), .ZN(
        P1_U3445) );
  INV_X1 U13570 ( .A(n10920), .ZN(n13607) );
  OAI222_X1 U13571 ( .A1(n11488), .A2(P3_U3151), .B1(n13610), .B2(n10837), 
        .C1(n10836), .C2(n13607), .ZN(P3_U3289) );
  INV_X1 U13572 ( .A(n10838), .ZN(n10859) );
  OAI222_X1 U13573 ( .A1(n10939), .A2(P1_U3086), .B1(n15400), .B2(n10859), 
        .C1(n10839), .C2(n15397), .ZN(P1_U3349) );
  INV_X1 U13574 ( .A(n10840), .ZN(n10861) );
  INV_X1 U13575 ( .A(n14879), .ZN(n10932) );
  OAI222_X1 U13576 ( .A1(n15397), .A2(n10841), .B1(n15400), .B2(n10861), .C1(
        n10932), .C2(P1_U3086), .ZN(P1_U3350) );
  NAND2_X1 U13577 ( .A1(n10842), .A2(n10724), .ZN(n10843) );
  NAND2_X1 U13578 ( .A1(n10844), .A2(n10843), .ZN(n11243) );
  AOI21_X1 U13579 ( .B1(n10363), .B2(n10845), .A(n11243), .ZN(n10846) );
  XNOR2_X1 U13580 ( .A(n10846), .B(n11244), .ZN(n10847) );
  AOI22_X1 U13581 ( .A1(n10848), .A2(n10847), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10849) );
  OAI21_X1 U13582 ( .B1(n10850), .B2(n14972), .A(n10849), .ZN(P1_U3243) );
  INV_X1 U13583 ( .A(n10851), .ZN(n10857) );
  INV_X1 U13584 ( .A(n11262), .ZN(n11264) );
  OAI222_X1 U13585 ( .A1(n15397), .A2(n10852), .B1(n15400), .B2(n10857), .C1(
        n11264), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U13586 ( .A(n14673), .ZN(n14677) );
  INV_X1 U13587 ( .A(n14677), .ZN(n14685) );
  OAI222_X1 U13588 ( .A1(n14682), .A2(n10854), .B1(n14685), .B2(n10853), .C1(
        P2_U3088), .C2(n15523), .ZN(P2_U3325) );
  INV_X1 U13589 ( .A(n14144), .ZN(n14138) );
  OAI222_X1 U13590 ( .A1(n14682), .A2(n10856), .B1(n14685), .B2(n10855), .C1(
        n14138), .C2(P2_U3088), .ZN(P2_U3323) );
  INV_X1 U13591 ( .A(n11018), .ZN(n15542) );
  OAI222_X1 U13592 ( .A1(n14682), .A2(n10858), .B1(n14685), .B2(n10857), .C1(
        P2_U3088), .C2(n15542), .ZN(P2_U3320) );
  OAI222_X1 U13593 ( .A1(n14682), .A2(n10860), .B1(n14685), .B2(n10859), .C1(
        P2_U3088), .C2(n14172), .ZN(P2_U3321) );
  INV_X1 U13594 ( .A(n14159), .ZN(n14153) );
  OAI222_X1 U13595 ( .A1(n14682), .A2(n10862), .B1(n14685), .B2(n10861), .C1(
        P2_U3088), .C2(n14153), .ZN(P2_U3322) );
  INV_X1 U13596 ( .A(n14130), .ZN(n14124) );
  OAI222_X1 U13597 ( .A1(n14682), .A2(n10864), .B1(n14685), .B2(n10863), .C1(
        n14124), .C2(P2_U3088), .ZN(P2_U3324) );
  INV_X1 U13598 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n15769) );
  NAND2_X1 U13599 ( .A1(n9024), .A2(P3_U3897), .ZN(n10865) );
  OAI21_X1 U13600 ( .B1(P3_U3897), .B2(n15769), .A(n10865), .ZN(P3_U3494) );
  INV_X1 U13601 ( .A(n10866), .ZN(n10867) );
  OAI222_X1 U13602 ( .A1(P3_U3151), .A2(n10869), .B1(n13598), .B2(n10868), 
        .C1(n13610), .C2(n10867), .ZN(P3_U3283) );
  INV_X1 U13603 ( .A(n10870), .ZN(n10873) );
  OAI222_X1 U13604 ( .A1(n14682), .A2(n10871), .B1(n14685), .B2(n10873), .C1(
        P2_U3088), .C2(n14187), .ZN(P2_U3319) );
  OAI222_X1 U13605 ( .A1(n7436), .A2(P1_U3086), .B1(n15400), .B2(n10873), .C1(
        n10872), .C2(n15397), .ZN(P1_U3347) );
  INV_X1 U13606 ( .A(n11396), .ZN(n11406) );
  OAI222_X1 U13607 ( .A1(P2_U3088), .A2(n11406), .B1(n14685), .B2(n10876), 
        .C1(n10874), .C2(n14682), .ZN(P2_U3318) );
  INV_X1 U13608 ( .A(n11266), .ZN(n11619) );
  OAI222_X1 U13609 ( .A1(P1_U3086), .A2(n11619), .B1(n15400), .B2(n10876), 
        .C1(n10875), .C2(n15397), .ZN(P1_U3346) );
  NAND2_X1 U13610 ( .A1(n10878), .A2(n10877), .ZN(n10883) );
  INV_X1 U13611 ( .A(n10879), .ZN(n10880) );
  OR2_X1 U13612 ( .A1(n10881), .A2(n10880), .ZN(n10882) );
  NAND2_X1 U13613 ( .A1(n10886), .A2(n10885), .ZN(n10961) );
  XNOR2_X1 U13614 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n10887) );
  XNOR2_X1 U13615 ( .A(n10961), .B(n10887), .ZN(n10888) );
  OAI21_X1 U13616 ( .B1(n10889), .B2(n10888), .A(n10969), .ZN(n10890) );
  INV_X1 U13617 ( .A(n10890), .ZN(SUB_1596_U57) );
  OAI222_X1 U13618 ( .A1(P3_U3151), .A2(n13146), .B1(n13598), .B2(n10892), 
        .C1(n13610), .C2(n10891), .ZN(P3_U3282) );
  OAI222_X1 U13619 ( .A1(P3_U3151), .A2(n13160), .B1(n13598), .B2(n10894), 
        .C1(n13610), .C2(n10893), .ZN(P3_U3280) );
  OAI222_X1 U13620 ( .A1(P3_U3151), .A2(n10897), .B1(n13598), .B2(n10896), 
        .C1(n13610), .C2(n10895), .ZN(P3_U3281) );
  AOI21_X1 U13621 ( .B1(n10899), .B2(n12399), .A(n10898), .ZN(n10900) );
  OR2_X1 U13622 ( .A1(n10901), .A2(n10900), .ZN(n10911) );
  OR2_X1 U13623 ( .A1(n10904), .A2(P2_U3088), .ZN(n14679) );
  INV_X1 U13624 ( .A(n14679), .ZN(n10902) );
  AND2_X1 U13625 ( .A1(n10911), .A2(n10902), .ZN(n10903) );
  NAND2_X1 U13626 ( .A1(n10903), .A2(n14683), .ZN(n15529) );
  NAND2_X1 U13627 ( .A1(n15546), .A2(n10908), .ZN(n10906) );
  AND2_X1 U13628 ( .A1(n10904), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10905) );
  NAND2_X1 U13629 ( .A1(n10911), .A2(n10905), .ZN(n15543) );
  OAI211_X1 U13630 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15529), .A(n10906), .B(
        n15543), .ZN(n10910) );
  INV_X1 U13631 ( .A(n15546), .ZN(n14269) );
  OAI22_X1 U13632 ( .A1(n14269), .A2(n10908), .B1(n10907), .B2(n15529), .ZN(
        n10909) );
  MUX2_X1 U13633 ( .A(n10910), .B(n10909), .S(n7134), .Z(n10915) );
  NOR2_X2 U13634 ( .A1(n10911), .A2(P2_U3088), .ZN(n15525) );
  INV_X1 U13635 ( .A(n15525), .ZN(n15552) );
  INV_X1 U13636 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10913) );
  OAI22_X1 U13637 ( .A1(n15552), .A2(n10913), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10912), .ZN(n10914) );
  OR2_X1 U13638 ( .A1(n10915), .A2(n10914), .ZN(P2_U3214) );
  INV_X1 U13639 ( .A(n10916), .ZN(n10918) );
  INV_X1 U13640 ( .A(n11407), .ZN(n14198) );
  OAI222_X1 U13641 ( .A1(n14682), .A2(n10917), .B1(n14673), .B2(n10918), .C1(
        P2_U3088), .C2(n14198), .ZN(P2_U3317) );
  INV_X1 U13642 ( .A(n11620), .ZN(n14910) );
  OAI222_X1 U13643 ( .A1(n15397), .A2(n10919), .B1(n15400), .B2(n10918), .C1(
        n14910), .C2(P1_U3086), .ZN(P1_U3345) );
  AOI22_X1 U13644 ( .A1(n13182), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_16_), .B2(
        n10920), .ZN(n10921) );
  OAI21_X1 U13645 ( .B1(n10922), .B2(n13610), .A(n10921), .ZN(P3_U3279) );
  XNOR2_X1 U13646 ( .A(n10983), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10928) );
  XNOR2_X1 U13647 ( .A(n10931), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n10948) );
  XNOR2_X1 U13648 ( .A(n14868), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n14865) );
  MUX2_X1 U13649 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10926), .S(n14879), .Z(
        n14873) );
  AOI211_X1 U13650 ( .C1(n10928), .C2(n10927), .A(n14940), .B(n10979), .ZN(
        n10942) );
  NOR2_X1 U13651 ( .A1(n10929), .A2(n11993), .ZN(n11246) );
  MUX2_X1 U13652 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9518), .S(n11247), .Z(
        n10930) );
  OAI21_X1 U13653 ( .B1(n11245), .B2(n11246), .A(n10930), .ZN(n11252) );
  NAND2_X1 U13654 ( .A1(n11247), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10951) );
  MUX2_X1 U13655 ( .A(n12124), .B(P1_REG2_REG_3__SCAN_IN), .S(n10931), .Z(
        n10950) );
  NOR2_X1 U13656 ( .A1(n10958), .A2(n12124), .ZN(n14858) );
  MUX2_X1 U13657 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11970), .S(n14868), .Z(
        n14857) );
  OAI21_X1 U13658 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14883) );
  NAND2_X1 U13659 ( .A1(n14868), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14882) );
  MUX2_X1 U13660 ( .A(n11948), .B(P1_REG2_REG_5__SCAN_IN), .S(n14879), .Z(
        n14881) );
  AOI21_X1 U13661 ( .B1(n14883), .B2(n14882), .A(n14881), .ZN(n14880) );
  NOR2_X1 U13662 ( .A1(n10932), .A2(n11948), .ZN(n10934) );
  MUX2_X1 U13663 ( .A(n11907), .B(P1_REG2_REG_6__SCAN_IN), .S(n10939), .Z(
        n10933) );
  INV_X1 U13664 ( .A(n10986), .ZN(n10936) );
  NOR3_X1 U13665 ( .A1(n14880), .A2(n10934), .A3(n10933), .ZN(n10935) );
  NOR3_X1 U13666 ( .A1(n10936), .A2(n10935), .A3(n14960), .ZN(n10941) );
  NOR2_X1 U13667 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9571), .ZN(n10937) );
  AOI21_X1 U13668 ( .B1(n14945), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10937), .ZN(
        n10938) );
  OAI21_X1 U13669 ( .B1(n10939), .B2(n14959), .A(n10938), .ZN(n10940) );
  OR3_X1 U13670 ( .A1(n10942), .A2(n10941), .A3(n10940), .ZN(P1_U3249) );
  INV_X1 U13671 ( .A(n10943), .ZN(n10946) );
  INV_X1 U13672 ( .A(n11589), .ZN(n11584) );
  OAI222_X1 U13673 ( .A1(n14682), .A2(n10944), .B1(n14673), .B2(n10946), .C1(
        P2_U3088), .C2(n11584), .ZN(P2_U3316) );
  INV_X1 U13674 ( .A(n11826), .ZN(n11824) );
  OAI222_X1 U13675 ( .A1(n11824), .A2(P1_U3086), .B1(n15400), .B2(n10946), 
        .C1(n10945), .C2(n15397), .ZN(P1_U3344) );
  AOI211_X1 U13676 ( .C1(n10949), .C2(n10948), .A(n10947), .B(n14940), .ZN(
        n10954) );
  AND3_X1 U13677 ( .A1(n11252), .A2(n10951), .A3(n10950), .ZN(n10952) );
  NOR3_X1 U13678 ( .A1(n14960), .A2(n14859), .A3(n10952), .ZN(n10953) );
  NOR2_X1 U13679 ( .A1(n10954), .A2(n10953), .ZN(n10957) );
  AND2_X1 U13680 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10955) );
  AOI21_X1 U13681 ( .B1(n14945), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n10955), .ZN(
        n10956) );
  OAI211_X1 U13682 ( .C1(n10958), .C2(n14959), .A(n10957), .B(n10956), .ZN(
        P1_U3246) );
  INV_X1 U13683 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10959) );
  NAND2_X1 U13684 ( .A1(n10959), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10960) );
  NAND2_X1 U13685 ( .A1(n10961), .A2(n10960), .ZN(n10964) );
  INV_X1 U13686 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U13687 ( .A1(n10962), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10963) );
  INV_X1 U13688 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n11390) );
  XNOR2_X1 U13689 ( .A(n11097), .B(n11390), .ZN(n11096) );
  INV_X1 U13690 ( .A(n11096), .ZN(n10965) );
  XNOR2_X1 U13691 ( .A(n10965), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n10971) );
  INV_X1 U13692 ( .A(n10966), .ZN(n10967) );
  NAND2_X1 U13693 ( .A1(n10967), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10968) );
  INV_X1 U13694 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15551) );
  OAI21_X1 U13695 ( .B1(n10971), .B2(n10970), .A(n11095), .ZN(n10972) );
  INV_X1 U13696 ( .A(n10972), .ZN(SUB_1596_U56) );
  INV_X1 U13697 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U13698 ( .A1(n11121), .A2(n10973), .ZN(n14040) );
  AOI21_X1 U13699 ( .B1(n14443), .B2(n14426), .A(n14040), .ZN(n10975) );
  NAND2_X1 U13700 ( .A1(n14110), .A2(n13725), .ZN(n11036) );
  INV_X1 U13701 ( .A(n11036), .ZN(n10974) );
  NOR2_X1 U13702 ( .A1(n10975), .A2(n10974), .ZN(n11654) );
  NAND2_X1 U13703 ( .A1(n13763), .A2(n10976), .ZN(n11655) );
  OAI211_X1 U13704 ( .C1(n14040), .C2(n11698), .A(n11654), .B(n11655), .ZN(
        n14619) );
  NAND2_X1 U13705 ( .A1(n15572), .A2(n14619), .ZN(n10977) );
  OAI21_X1 U13706 ( .B1(n15572), .B2(n10978), .A(n10977), .ZN(P2_U3430) );
  MUX2_X1 U13707 ( .A(n10980), .B(P1_REG1_REG_7__SCAN_IN), .S(n11262), .Z(
        n10981) );
  AOI211_X1 U13708 ( .C1(n10982), .C2(n10981), .A(n14940), .B(n11261), .ZN(
        n10992) );
  NAND2_X1 U13709 ( .A1(n10983), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10985) );
  MUX2_X1 U13710 ( .A(n11928), .B(P1_REG2_REG_7__SCAN_IN), .S(n11262), .Z(
        n10984) );
  INV_X1 U13711 ( .A(n14900), .ZN(n10988) );
  NAND3_X1 U13712 ( .A1(n10986), .A2(n10985), .A3(n10984), .ZN(n10987) );
  NAND3_X1 U13713 ( .A1(n10988), .A2(n14964), .A3(n10987), .ZN(n10990) );
  AND2_X1 U13714 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11530) );
  AOI21_X1 U13715 ( .B1(n14945), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n11530), .ZN(
        n10989) );
  OAI211_X1 U13716 ( .C1(n14959), .C2(n11264), .A(n10990), .B(n10989), .ZN(
        n10991) );
  OR2_X1 U13717 ( .A1(n10992), .A2(n10991), .ZN(P1_U3250) );
  XNOR2_X1 U13718 ( .A(n11396), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n11002) );
  XNOR2_X1 U13719 ( .A(n14113), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n14119) );
  AND2_X1 U13720 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14118) );
  NAND2_X1 U13721 ( .A1(n14119), .A2(n14118), .ZN(n14117) );
  INV_X1 U13722 ( .A(n14113), .ZN(n11006) );
  NAND2_X1 U13723 ( .A1(n11006), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10993) );
  NAND2_X1 U13724 ( .A1(n14117), .A2(n10993), .ZN(n15520) );
  XNOR2_X1 U13725 ( .A(n15523), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n15521) );
  NAND2_X1 U13726 ( .A1(n15520), .A2(n15521), .ZN(n15519) );
  XOR2_X1 U13727 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n14159), .Z(n14158) );
  XNOR2_X1 U13728 ( .A(n14172), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n14171) );
  XOR2_X1 U13729 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n11018), .Z(n15539) );
  XNOR2_X1 U13730 ( .A(n14187), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n14186) );
  OAI21_X1 U13731 ( .B1(n11000), .B2(n14187), .A(n14184), .ZN(n11001) );
  AOI21_X1 U13732 ( .B1(n11002), .B2(n11001), .A(n11404), .ZN(n11032) );
  AND2_X1 U13733 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11838) );
  NOR2_X1 U13734 ( .A1(n15543), .A2(n11406), .ZN(n11003) );
  AOI211_X1 U13735 ( .C1(n15525), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n11838), .B(
        n11003), .ZN(n11031) );
  INV_X1 U13736 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n14504) );
  MUX2_X1 U13737 ( .A(n14504), .B(P2_REG2_REG_1__SCAN_IN), .S(n14113), .Z(
        n11005) );
  AND2_X1 U13738 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n11004) );
  NAND2_X1 U13739 ( .A1(n11006), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U13740 ( .A1(n11008), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n14131) );
  MUX2_X1 U13741 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11374), .S(n14130), .Z(
        n11009) );
  NAND2_X1 U13742 ( .A1(n11010), .A2(n11009), .ZN(n14147) );
  NAND2_X1 U13743 ( .A1(n14130), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n14146) );
  NAND2_X1 U13744 ( .A1(n14147), .A2(n14146), .ZN(n11012) );
  MUX2_X1 U13745 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11436), .S(n14144), .Z(
        n11011) );
  NAND2_X1 U13746 ( .A1(n14144), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n14160) );
  MUX2_X1 U13747 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11640), .S(n14159), .Z(
        n11013) );
  NAND2_X1 U13748 ( .A1(n14159), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n14173) );
  MUX2_X1 U13749 ( .A(n11660), .B(P2_REG2_REG_6__SCAN_IN), .S(n14172), .Z(
        n11014) );
  NAND2_X1 U13750 ( .A1(n11015), .A2(n11014), .ZN(n14177) );
  NAND2_X1 U13751 ( .A1(n11016), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n11017) );
  NAND2_X1 U13752 ( .A1(n14177), .A2(n11017), .ZN(n15547) );
  INV_X1 U13753 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11539) );
  MUX2_X1 U13754 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11539), .S(n11018), .Z(
        n15548) );
  NAND2_X1 U13755 ( .A1(n11018), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n14189) );
  NAND2_X1 U13756 ( .A1(n15545), .A2(n14189), .ZN(n11021) );
  MUX2_X1 U13757 ( .A(n11019), .B(P2_REG2_REG_8__SCAN_IN), .S(n14187), .Z(
        n11020) );
  NAND2_X1 U13758 ( .A1(n11021), .A2(n11020), .ZN(n14191) );
  NAND2_X1 U13759 ( .A1(n11022), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11023) );
  INV_X1 U13760 ( .A(n11026), .ZN(n11028) );
  INV_X1 U13761 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11024) );
  MUX2_X1 U13762 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11024), .S(n11396), .Z(
        n11027) );
  MUX2_X1 U13763 ( .A(n11024), .B(P2_REG2_REG_9__SCAN_IN), .S(n11396), .Z(
        n11025) );
  OAI21_X1 U13764 ( .B1(n11028), .B2(n11027), .A(n11398), .ZN(n11029) );
  NAND2_X1 U13765 ( .A1(n11029), .A2(n15546), .ZN(n11030) );
  OAI211_X1 U13766 ( .C1(n11032), .C2(n15529), .A(n11031), .B(n11030), .ZN(
        P2_U3223) );
  AOI21_X1 U13767 ( .B1(n13714), .B2(n11033), .A(n13751), .ZN(n11039) );
  OR2_X1 U13768 ( .A1(n11034), .A2(P2_U3088), .ZN(n11072) );
  OAI21_X1 U13769 ( .B1(n13726), .B2(n11036), .A(n11035), .ZN(n11037) );
  AOI21_X1 U13770 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n11072), .A(n11037), .ZN(
        n11038) );
  OAI21_X1 U13771 ( .B1(n11039), .B2(n13755), .A(n11038), .ZN(P2_U3204) );
  INV_X1 U13772 ( .A(n11040), .ZN(n11041) );
  OAI222_X1 U13773 ( .A1(n13607), .A2(n11042), .B1(n13610), .B2(n11041), .C1(
        P3_U3151), .C2(n13194), .ZN(P3_U3278) );
  OAI21_X1 U13774 ( .B1(n11045), .B2(n11044), .A(n11043), .ZN(n11046) );
  AOI22_X1 U13775 ( .A1(n7087), .A2(n13751), .B1(n13714), .B2(n11046), .ZN(
        n11050) );
  NAND2_X1 U13776 ( .A1(n14109), .A2(n13725), .ZN(n11048) );
  NAND2_X1 U13777 ( .A1(n11048), .A2(n11047), .ZN(n11126) );
  AOI22_X1 U13778 ( .A1(n13746), .A2(n11126), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n11072), .ZN(n11049) );
  NAND2_X1 U13779 ( .A1(n11050), .A2(n11049), .ZN(P2_U3194) );
  NOR2_X1 U13780 ( .A1(n11051), .A2(P1_U3086), .ZN(n11363) );
  INV_X1 U13781 ( .A(n11363), .ZN(n14719) );
  AOI22_X1 U13782 ( .A1(n14719), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n11203), 
        .B2(n10664), .ZN(n11056) );
  OAI21_X1 U13783 ( .B1(n11054), .B2(n11053), .A(n11052), .ZN(n11239) );
  NOR2_X1 U13784 ( .A1(n9507), .A2(n15168), .ZN(n15475) );
  AOI22_X1 U13785 ( .A1(n14801), .A2(n11239), .B1(n14822), .B2(n15475), .ZN(
        n11055) );
  NAND2_X1 U13786 ( .A1(n11056), .A2(n11055), .ZN(P1_U3232) );
  AND2_X1 U13787 ( .A1(n11073), .A2(n11057), .ZN(n13693) );
  XNOR2_X1 U13788 ( .A(n13693), .B(n13692), .ZN(n11063) );
  NAND2_X1 U13789 ( .A1(n14107), .A2(n13725), .ZN(n11059) );
  NAND2_X1 U13790 ( .A1(n14109), .A2(n14073), .ZN(n11058) );
  AND2_X1 U13791 ( .A1(n11059), .A2(n11058), .ZN(n11371) );
  INV_X1 U13792 ( .A(n11371), .ZN(n11060) );
  AOI22_X1 U13793 ( .A1(n13746), .A2(n11060), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11062) );
  INV_X1 U13794 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U13795 ( .A1(n13751), .A2(n15563), .B1(n13700), .B2(n14123), .ZN(
        n11061) );
  OAI211_X1 U13796 ( .C1(n11063), .C2(n13753), .A(n11062), .B(n11061), .ZN(
        P2_U3190) );
  INV_X1 U13797 ( .A(n11064), .ZN(n11067) );
  INV_X1 U13798 ( .A(n12283), .ZN(n11830) );
  OAI222_X1 U13799 ( .A1(n15397), .A2(n11065), .B1(n15400), .B2(n11067), .C1(
        P1_U3086), .C2(n11830), .ZN(P1_U3343) );
  OAI222_X1 U13800 ( .A1(P2_U3088), .A2(n12261), .B1(n14673), .B2(n11067), 
        .C1(n11066), .C2(n14682), .ZN(P2_U3315) );
  INV_X1 U13801 ( .A(n13211), .ZN(n11070) );
  OAI222_X1 U13802 ( .A1(P3_U3151), .A2(n11070), .B1(n13607), .B2(n11069), 
        .C1(n13610), .C2(n11068), .ZN(P3_U3277) );
  OAI22_X1 U13803 ( .A1(n11071), .A2(n13732), .B1(n11434), .B2(n13734), .ZN(
        n11084) );
  AOI22_X1 U13804 ( .A1(n13746), .A2(n11084), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n11072), .ZN(n11078) );
  OAI21_X1 U13805 ( .B1(n11075), .B2(n11074), .A(n11073), .ZN(n11076) );
  NAND2_X1 U13806 ( .A1(n13714), .A2(n11076), .ZN(n11077) );
  OAI211_X1 U13807 ( .C1(n13774), .C2(n13738), .A(n11078), .B(n11077), .ZN(
        P2_U3209) );
  INV_X1 U13808 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11088) );
  XNOR2_X1 U13809 ( .A(n14043), .B(n11079), .ZN(n11652) );
  INV_X1 U13810 ( .A(n11128), .ZN(n11080) );
  AOI211_X1 U13811 ( .C1(n11081), .C2(n11080), .A(n7907), .B(n10035), .ZN(
        n11647) );
  AOI21_X1 U13812 ( .B1(n15564), .B2(n11081), .A(n11647), .ZN(n11086) );
  OAI21_X1 U13813 ( .B1(n11083), .B2(n14043), .A(n11082), .ZN(n11085) );
  AOI21_X1 U13814 ( .B1(n11085), .B2(n14481), .A(n11084), .ZN(n11649) );
  OAI211_X1 U13815 ( .C1(n15567), .C2(n11652), .A(n11086), .B(n11649), .ZN(
        n11179) );
  NAND2_X1 U13816 ( .A1(n11179), .A2(n15572), .ZN(n11087) );
  OAI21_X1 U13817 ( .B1(n15572), .B2(n11088), .A(n11087), .ZN(P2_U3436) );
  INV_X1 U13818 ( .A(n12263), .ZN(n14211) );
  INV_X1 U13819 ( .A(n11089), .ZN(n11091) );
  OAI222_X1 U13820 ( .A1(P2_U3088), .A2(n14211), .B1(n14673), .B2(n11091), 
        .C1(n11090), .C2(n14682), .ZN(P2_U3314) );
  INV_X1 U13821 ( .A(n12432), .ZN(n12435) );
  OAI222_X1 U13822 ( .A1(n15397), .A2(n11092), .B1(n15400), .B2(n11091), .C1(
        P1_U3086), .C2(n12435), .ZN(P1_U3342) );
  NAND2_X1 U13823 ( .A1(n11093), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n11094) );
  NAND2_X1 U13824 ( .A1(n11096), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n11099) );
  INV_X1 U13825 ( .A(n11105), .ZN(n11103) );
  INV_X1 U13826 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11452) );
  NAND2_X1 U13827 ( .A1(n11452), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n11766) );
  INV_X1 U13828 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n11100) );
  NAND2_X1 U13829 ( .A1(n11100), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n11101) );
  AND2_X1 U13830 ( .A1(n11766), .A2(n11101), .ZN(n11104) );
  INV_X1 U13831 ( .A(n11104), .ZN(n11102) );
  NAND2_X1 U13832 ( .A1(n11103), .A2(n11102), .ZN(n11106) );
  NAND2_X1 U13833 ( .A1(n11106), .A2(n11767), .ZN(n11762) );
  INV_X1 U13834 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n11760) );
  XNOR2_X1 U13835 ( .A(n11761), .B(n11760), .ZN(SUB_1596_U55) );
  INV_X1 U13836 ( .A(n15507), .ZN(n15314) );
  OAI21_X1 U13837 ( .B1(n11109), .B2(n11108), .A(n11107), .ZN(n12150) );
  OR2_X1 U13838 ( .A1(n11111), .A2(n6845), .ZN(n11112) );
  AND3_X1 U13839 ( .A1(n11110), .A2(n15283), .A3(n11112), .ZN(n12149) );
  INV_X1 U13840 ( .A(n12150), .ZN(n11117) );
  OAI21_X1 U13841 ( .B1(n11113), .B2(n7392), .A(n12120), .ZN(n11115) );
  OAI22_X1 U13842 ( .A1(n11364), .A2(n15168), .B1(n9507), .B2(n15166), .ZN(
        n11114) );
  AOI21_X1 U13843 ( .B1(n11115), .B2(n15327), .A(n11114), .ZN(n11116) );
  OAI21_X1 U13844 ( .B1(n11117), .B2(n15147), .A(n11116), .ZN(n12145) );
  AOI211_X1 U13845 ( .C1(n15314), .C2(n12150), .A(n12149), .B(n12145), .ZN(
        n11380) );
  OAI22_X1 U13846 ( .A1(n15389), .A2(n6845), .B1(n15512), .B2(n9520), .ZN(
        n11118) );
  INV_X1 U13847 ( .A(n11118), .ZN(n11119) );
  OAI21_X1 U13848 ( .B1(n11380), .B2(n15510), .A(n11119), .ZN(P1_U3465) );
  INV_X1 U13849 ( .A(n11121), .ZN(n11122) );
  XNOR2_X1 U13850 ( .A(n11120), .B(n11122), .ZN(n14505) );
  OAI21_X1 U13851 ( .B1(n14042), .B2(n11124), .A(n11123), .ZN(n11127) );
  NOR2_X1 U13852 ( .A1(n14505), .A2(n14426), .ZN(n11125) );
  AOI211_X1 U13853 ( .C1(n14481), .C2(n11127), .A(n11126), .B(n11125), .ZN(
        n14503) );
  OAI21_X1 U13854 ( .B1(n10034), .B2(n13755), .A(n14469), .ZN(n11129) );
  NOR2_X1 U13855 ( .A1(n11129), .A2(n11128), .ZN(n14506) );
  INV_X1 U13856 ( .A(n14506), .ZN(n11130) );
  OAI211_X1 U13857 ( .C1(n14505), .C2(n11698), .A(n14503), .B(n11130), .ZN(
        n11795) );
  INV_X1 U13858 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11131) );
  OAI22_X1 U13859 ( .A1(n14660), .A2(n10034), .B1(n15572), .B2(n11131), .ZN(
        n11132) );
  AOI21_X1 U13860 ( .B1(n11795), .B2(n15572), .A(n11132), .ZN(n11133) );
  INV_X1 U13861 ( .A(n11133), .ZN(P2_U3433) );
  XOR2_X1 U13862 ( .A(n11134), .B(n11135), .Z(n11148) );
  OAI21_X1 U13863 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n11136), .A(n11232), .ZN(
        n11144) );
  INV_X1 U13864 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n11142) );
  OAI21_X1 U13865 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n11138), .A(n11137), .ZN(
        n11139) );
  NAND2_X1 U13866 ( .A1(n13217), .A2(n11139), .ZN(n11141) );
  NAND2_X1 U13867 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n11140) );
  OAI211_X1 U13868 ( .C1(n13215), .C2(n11142), .A(n11141), .B(n11140), .ZN(
        n11143) );
  AOI21_X1 U13869 ( .B1(n13222), .B2(n11144), .A(n11143), .ZN(n11147) );
  NAND2_X1 U13870 ( .A1(n13212), .A2(n11145), .ZN(n11146) );
  OAI211_X1 U13871 ( .C1(n11148), .C2(n13226), .A(n11147), .B(n11146), .ZN(
        P3_U3185) );
  XOR2_X1 U13872 ( .A(n11149), .B(n11150), .Z(n11163) );
  OAI21_X1 U13873 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11151), .A(n11483), .ZN(
        n11159) );
  INV_X1 U13874 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n11157) );
  OAI21_X1 U13875 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n11153), .A(n11152), .ZN(
        n11154) );
  NAND2_X1 U13876 ( .A1(n11154), .A2(n13217), .ZN(n11156) );
  NAND2_X1 U13877 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n11155) );
  OAI211_X1 U13878 ( .C1(n13215), .C2(n11157), .A(n11156), .B(n11155), .ZN(
        n11158) );
  AOI21_X1 U13879 ( .B1(n13222), .B2(n11159), .A(n11158), .ZN(n11162) );
  NAND2_X1 U13880 ( .A1(n13212), .A2(n11160), .ZN(n11161) );
  OAI211_X1 U13881 ( .C1(n11163), .C2(n13226), .A(n11162), .B(n11161), .ZN(
        P3_U3187) );
  INV_X1 U13882 ( .A(n11164), .ZN(n11165) );
  XNOR2_X1 U13883 ( .A(n11167), .B(n11165), .ZN(n11988) );
  OAI21_X1 U13884 ( .B1(n11167), .B2(n11166), .A(n15327), .ZN(n11170) );
  AOI21_X1 U13885 ( .B1(n11168), .B2(n15327), .A(n10460), .ZN(n11169) );
  AOI21_X1 U13886 ( .B1(n15166), .B2(n11170), .A(n11169), .ZN(n11171) );
  NOR2_X1 U13887 ( .A1(n6844), .A2(n15168), .ZN(n14718) );
  NOR2_X1 U13888 ( .A1(n11171), .A2(n14718), .ZN(n11992) );
  XNOR2_X1 U13889 ( .A(n11987), .B(n11203), .ZN(n11172) );
  AND2_X1 U13890 ( .A1(n11172), .A2(n15283), .ZN(n11991) );
  INV_X1 U13891 ( .A(n11991), .ZN(n11173) );
  OAI211_X1 U13892 ( .C1(n15353), .C2(n11988), .A(n11992), .B(n11173), .ZN(
        n11506) );
  OAI22_X1 U13893 ( .A1(n15389), .A2(n11987), .B1(n15512), .B2(n9488), .ZN(
        n11174) );
  AOI21_X1 U13894 ( .B1(n11506), .B2(n15512), .A(n11174), .ZN(n11175) );
  INV_X1 U13895 ( .A(n11175), .ZN(P1_U3462) );
  OAI222_X1 U13896 ( .A1(n13610), .A2(n11178), .B1(n13598), .B2(n11177), .C1(
        P3_U3151), .C2(n11176), .ZN(P3_U3276) );
  NAND2_X1 U13897 ( .A1(n11179), .A2(n14618), .ZN(n11180) );
  OAI21_X1 U13898 ( .B1(n14618), .B2(n10994), .A(n11180), .ZN(P2_U3501) );
  XOR2_X1 U13899 ( .A(n11181), .B(n11182), .Z(n11195) );
  AOI21_X1 U13900 ( .B1(n11185), .B2(n11184), .A(n11183), .ZN(n11186) );
  NOR2_X1 U13901 ( .A1(n13165), .A2(n11186), .ZN(n11193) );
  AOI21_X1 U13902 ( .B1(n11189), .B2(n11188), .A(n11187), .ZN(n11191) );
  AOI22_X1 U13903 ( .A1(n15575), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11190) );
  OAI21_X1 U13904 ( .B1(n13200), .B2(n11191), .A(n11190), .ZN(n11192) );
  AOI211_X1 U13905 ( .C1(n13212), .C2(n9176), .A(n11193), .B(n11192), .ZN(
        n11194) );
  OAI21_X1 U13906 ( .B1(n11195), .B2(n13226), .A(n11194), .ZN(P3_U3184) );
  XNOR2_X1 U13907 ( .A(n11197), .B(n11196), .ZN(n11202) );
  OR2_X1 U13908 ( .A1(n13808), .A2(n13732), .ZN(n11199) );
  OR2_X1 U13909 ( .A1(n13820), .A2(n13734), .ZN(n11198) );
  NAND2_X1 U13910 ( .A1(n11199), .A2(n11198), .ZN(n11576) );
  AND2_X1 U13911 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14168) );
  OAI22_X1 U13912 ( .A1(n13738), .A2(n11663), .B1(n13748), .B2(n11662), .ZN(
        n11200) );
  AOI211_X1 U13913 ( .C1(n13746), .C2(n11576), .A(n14168), .B(n11200), .ZN(
        n11201) );
  OAI21_X1 U13914 ( .B1(n11202), .B2(n13753), .A(n11201), .ZN(P2_U3211) );
  NOR2_X1 U13915 ( .A1(n15494), .A2(n15327), .ZN(n11205) );
  INV_X1 U13916 ( .A(n15475), .ZN(n11204) );
  NAND2_X1 U13917 ( .A1(n11203), .A2(n7518), .ZN(n15473) );
  OAI211_X1 U13918 ( .C1(n11205), .C2(n15476), .A(n11204), .B(n15473), .ZN(
        n11207) );
  NAND2_X1 U13919 ( .A1(n11207), .A2(n15512), .ZN(n11206) );
  OAI21_X1 U13920 ( .B1(n15512), .B2(n9509), .A(n11206), .ZN(P1_U3459) );
  NAND2_X1 U13921 ( .A1(n11207), .A2(n15518), .ZN(n11208) );
  OAI21_X1 U13922 ( .B1(n15518), .B2(n10845), .A(n11208), .ZN(P1_U3528) );
  XNOR2_X1 U13923 ( .A(n11209), .B(n11286), .ZN(n11220) );
  AOI21_X1 U13924 ( .B1(n11212), .B2(n11211), .A(n11210), .ZN(n11213) );
  NOR2_X1 U13925 ( .A1(n13165), .A2(n11213), .ZN(n11219) );
  AOI21_X1 U13926 ( .B1(n15596), .B2(n11215), .A(n11214), .ZN(n11217) );
  AOI22_X1 U13927 ( .A1(n15575), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11216) );
  OAI21_X1 U13928 ( .B1(n13200), .B2(n11217), .A(n11216), .ZN(n11218) );
  AOI211_X1 U13929 ( .C1(n11220), .C2(n13140), .A(n11219), .B(n11218), .ZN(
        n11221) );
  OAI21_X1 U13930 ( .B1(n9173), .B2(n13195), .A(n11221), .ZN(P3_U3183) );
  XOR2_X1 U13931 ( .A(n11222), .B(n11223), .Z(n11238) );
  AND3_X1 U13932 ( .A1(n11137), .A2(n11225), .A3(n11224), .ZN(n11226) );
  OAI21_X1 U13933 ( .B1(n11227), .B2(n11226), .A(n13217), .ZN(n11229) );
  NAND2_X1 U13934 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n11228) );
  OAI211_X1 U13935 ( .C1(n13215), .C2(n7022), .A(n11229), .B(n11228), .ZN(
        n11235) );
  NAND3_X1 U13936 ( .A1(n11232), .A2(n11231), .A3(n11230), .ZN(n11233) );
  AOI21_X1 U13937 ( .B1(n6633), .B2(n11233), .A(n13200), .ZN(n11234) );
  AOI211_X1 U13938 ( .C1(n13212), .C2(n11236), .A(n11235), .B(n11234), .ZN(
        n11237) );
  OAI21_X1 U13939 ( .B1(n11238), .B2(n13226), .A(n11237), .ZN(P3_U3186) );
  MUX2_X1 U13940 ( .A(n11240), .B(n11239), .S(n10363), .Z(n11241) );
  NOR2_X1 U13941 ( .A1(n11241), .A2(n12885), .ZN(n11242) );
  INV_X1 U13942 ( .A(n11245), .ZN(n11250) );
  INV_X1 U13943 ( .A(n11246), .ZN(n11249) );
  MUX2_X1 U13944 ( .A(n9518), .B(P1_REG2_REG_2__SCAN_IN), .S(n11247), .Z(
        n11248) );
  NAND3_X1 U13945 ( .A1(n11250), .A2(n11249), .A3(n11248), .ZN(n11251) );
  AND3_X1 U13946 ( .A1(n14964), .A2(n11252), .A3(n11251), .ZN(n11260) );
  AOI211_X1 U13947 ( .C1(n11255), .C2(n11254), .A(n11253), .B(n14940), .ZN(
        n11259) );
  AOI22_X1 U13948 ( .A1(n14945), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n11256) );
  OAI21_X1 U13949 ( .B1(n11257), .B2(n14959), .A(n11256), .ZN(n11258) );
  OR4_X1 U13950 ( .A1(n14856), .A2(n11260), .A3(n11259), .A4(n11258), .ZN(
        P1_U3245) );
  MUX2_X1 U13951 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7435), .S(n14901), .Z(
        n14890) );
  XOR2_X1 U13952 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n11266), .Z(n11612) );
  XOR2_X1 U13953 ( .A(n11613), .B(n11612), .Z(n11273) );
  INV_X1 U13954 ( .A(n14959), .ZN(n14902) );
  INV_X1 U13955 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n11773) );
  NAND2_X1 U13956 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n12103) );
  OAI21_X1 U13957 ( .B1(n14972), .B2(n11773), .A(n12103), .ZN(n11263) );
  AOI21_X1 U13958 ( .B1(n14902), .B2(n11266), .A(n11263), .ZN(n11272) );
  NOR2_X1 U13959 ( .A1(n11264), .A2(n11928), .ZN(n14895) );
  INV_X1 U13960 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11960) );
  MUX2_X1 U13961 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11960), .S(n14901), .Z(
        n11265) );
  NAND2_X1 U13962 ( .A1(n14901), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11268) );
  MUX2_X1 U13963 ( .A(n12082), .B(P1_REG2_REG_9__SCAN_IN), .S(n11266), .Z(
        n11267) );
  INV_X1 U13964 ( .A(n14915), .ZN(n11270) );
  NAND3_X1 U13965 ( .A1(n14898), .A2(n11268), .A3(n11267), .ZN(n11269) );
  NAND3_X1 U13966 ( .A1(n11270), .A2(n14964), .A3(n11269), .ZN(n11271) );
  OAI211_X1 U13967 ( .C1(n11273), .C2(n14940), .A(n11272), .B(n11271), .ZN(
        P1_U3252) );
  OAI21_X1 U13968 ( .B1(n11275), .B2(n11274), .A(n11798), .ZN(n11968) );
  NAND2_X1 U13969 ( .A1(n12125), .A2(n11276), .ZN(n11277) );
  NAND2_X1 U13970 ( .A1(n11277), .A2(n15283), .ZN(n11278) );
  NOR2_X1 U13971 ( .A1(n11949), .A2(n11278), .ZN(n11974) );
  OAI21_X1 U13972 ( .B1(n11281), .B2(n11280), .A(n11279), .ZN(n11282) );
  OAI22_X1 U13973 ( .A1(n11805), .A2(n15168), .B1(n11364), .B2(n15166), .ZN(
        n11521) );
  AOI21_X1 U13974 ( .B1(n11282), .B2(n15327), .A(n11521), .ZN(n11969) );
  INV_X1 U13975 ( .A(n11969), .ZN(n11283) );
  AOI211_X1 U13976 ( .C1(n15494), .C2(n11968), .A(n11974), .B(n11283), .ZN(
        n11504) );
  OAI22_X1 U13977 ( .A1(n15389), .A2(n11972), .B1(n15512), .B2(n9542), .ZN(
        n11284) );
  INV_X1 U13978 ( .A(n11284), .ZN(n11285) );
  OAI21_X1 U13979 ( .B1(n11504), .B2(n15510), .A(n11285), .ZN(P1_U3471) );
  NOR3_X1 U13980 ( .A1(n13222), .A2(n13217), .A3(n13140), .ZN(n11296) );
  INV_X1 U13981 ( .A(n11286), .ZN(n11295) );
  MUX2_X1 U13982 ( .A(n11287), .B(n12834), .S(n6983), .Z(n11290) );
  NAND2_X1 U13983 ( .A1(n13222), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U13984 ( .A1(n13217), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11288) );
  OAI211_X1 U13985 ( .C1(n11290), .C2(n13226), .A(n11289), .B(n11288), .ZN(
        n11291) );
  MUX2_X1 U13986 ( .A(n11291), .B(n13212), .S(P3_IR_REG_0__SCAN_IN), .Z(n11292) );
  INV_X1 U13987 ( .A(n11292), .ZN(n11294) );
  AOI22_X1 U13988 ( .A1(n15575), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11293) );
  OAI211_X1 U13989 ( .C1(n11296), .C2(n11295), .A(n11294), .B(n11293), .ZN(
        P3_U3182) );
  INV_X1 U13990 ( .A(n11327), .ZN(n11297) );
  NAND2_X1 U13991 ( .A1(n11297), .A2(n11316), .ZN(n11301) );
  INV_X1 U13992 ( .A(n11298), .ZN(n11300) );
  OR2_X1 U13993 ( .A1(n11325), .A2(n11318), .ZN(n11299) );
  NAND4_X1 U13994 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11852), .ZN(
        n11302) );
  NAND2_X1 U13995 ( .A1(n11302), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11305) );
  INV_X1 U13996 ( .A(n11846), .ZN(n11303) );
  INV_X1 U13997 ( .A(n11325), .ZN(n11319) );
  NAND3_X1 U13998 ( .A1(n11303), .A2(n11328), .A3(n11319), .ZN(n11304) );
  AND2_X1 U13999 ( .A1(n11544), .A2(n11306), .ZN(n11515) );
  NAND3_X1 U14000 ( .A1(n13106), .A2(n11331), .A3(n12906), .ZN(n11310) );
  INV_X1 U14001 ( .A(n13495), .ZN(n11313) );
  OAI211_X1 U14002 ( .C1(n11315), .C2(n13491), .A(n11339), .B(n11314), .ZN(
        n11321) );
  NAND3_X1 U14003 ( .A1(n11327), .A2(n11316), .A3(n15621), .ZN(n11317) );
  OAI21_X1 U14004 ( .B1(n11319), .B2(n11318), .A(n11317), .ZN(n11320) );
  NAND2_X1 U14005 ( .A1(n11320), .A2(n11328), .ZN(n13066) );
  NAND2_X1 U14006 ( .A1(n11321), .A2(n13044), .ZN(n11333) );
  NAND2_X1 U14007 ( .A1(n13105), .A2(n13060), .ZN(n11323) );
  NAND2_X1 U14008 ( .A1(n13059), .A2(n13108), .ZN(n11322) );
  NAND2_X1 U14009 ( .A1(n11323), .A2(n11322), .ZN(n13492) );
  INV_X1 U14010 ( .A(n11324), .ZN(n11326) );
  INV_X1 U14011 ( .A(n13071), .ZN(n13034) );
  NAND3_X1 U14012 ( .A1(n11327), .A2(n15614), .A3(n11328), .ZN(n11330) );
  AND2_X1 U14013 ( .A1(n15579), .A2(n11328), .ZN(n11329) );
  AOI22_X1 U14014 ( .A1(n13492), .A2(n13034), .B1(n13063), .B2(n11331), .ZN(
        n11332) );
  OAI211_X1 U14015 ( .C1(n11515), .C2(n11334), .A(n11333), .B(n11332), .ZN(
        P3_U3162) );
  INV_X1 U14016 ( .A(n14922), .ZN(n14927) );
  INV_X1 U14017 ( .A(n11335), .ZN(n11338) );
  OAI222_X1 U14018 ( .A1(P1_U3086), .A2(n14927), .B1(n15400), .B2(n11338), 
        .C1(n11336), .C2(n15397), .ZN(P1_U3339) );
  OAI222_X1 U14019 ( .A1(P2_U3088), .A2(n14237), .B1(n14673), .B2(n11338), 
        .C1(n11337), .C2(n14682), .ZN(P2_U3311) );
  XNOR2_X1 U14020 ( .A(n12906), .B(n11345), .ZN(n11545) );
  XNOR2_X1 U14021 ( .A(n11545), .B(n9020), .ZN(n11341) );
  OAI21_X1 U14022 ( .B1(n11341), .B2(n11340), .A(n11548), .ZN(n11342) );
  NAND2_X1 U14023 ( .A1(n11342), .A2(n13044), .ZN(n11347) );
  NAND2_X1 U14024 ( .A1(n9024), .A2(n13060), .ZN(n11344) );
  NAND2_X1 U14025 ( .A1(n13106), .A2(n13059), .ZN(n11343) );
  NAND2_X1 U14026 ( .A1(n11344), .A2(n11343), .ZN(n11673) );
  AOI22_X1 U14027 ( .A1(n11673), .A2(n13034), .B1(n13063), .B2(n11345), .ZN(
        n11346) );
  OAI211_X1 U14028 ( .C1(n11515), .C2(n15577), .A(n11347), .B(n11346), .ZN(
        P3_U3177) );
  INV_X1 U14029 ( .A(n12676), .ZN(n12678) );
  INV_X1 U14030 ( .A(n11348), .ZN(n11350) );
  OAI222_X1 U14031 ( .A1(P1_U3086), .A2(n12678), .B1(n15400), .B2(n11350), 
        .C1(n15740), .C2(n15397), .ZN(P1_U3341) );
  INV_X1 U14032 ( .A(n12764), .ZN(n12771) );
  OAI222_X1 U14033 ( .A1(P2_U3088), .A2(n12771), .B1(n14673), .B2(n11350), 
        .C1(n11349), .C2(n14682), .ZN(P2_U3313) );
  AOI21_X1 U14034 ( .B1(n11352), .B2(n11354), .A(n11353), .ZN(n11360) );
  NAND2_X1 U14035 ( .A1(n11355), .A2(n14801), .ZN(n11359) );
  MUX2_X1 U14036 ( .A(n14810), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n11357) );
  OAI22_X1 U14037 ( .A1(n14804), .A2(n6844), .B1(n10469), .B2(n14808), .ZN(
        n11356) );
  AOI211_X1 U14038 ( .C1(n14751), .C2(n14851), .A(n11357), .B(n11356), .ZN(
        n11358) );
  OAI21_X1 U14039 ( .B1(n11360), .B2(n11359), .A(n11358), .ZN(P1_U3218) );
  OAI21_X1 U14040 ( .B1(n11362), .B2(n11361), .A(n11352), .ZN(n11367) );
  OAI22_X1 U14041 ( .A1(n14808), .A2(n6845), .B1(n11363), .B2(n12146), .ZN(
        n11366) );
  OAI22_X1 U14042 ( .A1(n14804), .A2(n9507), .B1(n11364), .B2(n14815), .ZN(
        n11365) );
  AOI211_X1 U14043 ( .C1(n14801), .C2(n11367), .A(n11366), .B(n11365), .ZN(
        n11368) );
  INV_X1 U14044 ( .A(n11368), .ZN(P1_U3237) );
  INV_X1 U14045 ( .A(n11431), .ZN(n14044) );
  XNOR2_X1 U14046 ( .A(n11369), .B(n14044), .ZN(n15566) );
  AND2_X1 U14047 ( .A1(n11082), .A2(n11370), .ZN(n11432) );
  XNOR2_X1 U14048 ( .A(n11432), .B(n14044), .ZN(n11372) );
  OAI21_X1 U14049 ( .B1(n11372), .B2(n14443), .A(n11371), .ZN(n15568) );
  AOI21_X1 U14050 ( .B1(n14510), .B2(n14123), .A(n15568), .ZN(n11373) );
  MUX2_X1 U14051 ( .A(n11374), .B(n11373), .S(n14502), .Z(n11378) );
  INV_X1 U14052 ( .A(n11437), .ZN(n11375) );
  AOI211_X1 U14053 ( .C1(n15563), .C2(n11376), .A(n7907), .B(n11375), .ZN(
        n15562) );
  AOI22_X1 U14054 ( .A1(n14511), .A2(n15563), .B1(n14507), .B2(n15562), .ZN(
        n11377) );
  OAI211_X1 U14055 ( .C1(n14497), .C2(n15566), .A(n11378), .B(n11377), .ZN(
        P2_U3262) );
  AOI22_X1 U14056 ( .A1(n12215), .A2(n12148), .B1(n15516), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n11379) );
  OAI21_X1 U14057 ( .B1(n11380), .B2(n15516), .A(n11379), .ZN(P1_U3530) );
  XOR2_X1 U14058 ( .A(n11381), .B(n11382), .Z(n11395) );
  INV_X1 U14059 ( .A(n11383), .ZN(n11384) );
  OAI21_X1 U14060 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n11385), .A(n11384), .ZN(
        n11393) );
  AOI21_X1 U14061 ( .B1(n15659), .B2(n11386), .A(n11454), .ZN(n11387) );
  NOR2_X1 U14062 ( .A1(n11387), .A2(n13165), .ZN(n11392) );
  NAND2_X1 U14063 ( .A1(n13212), .A2(n11388), .ZN(n11389) );
  NAND2_X1 U14064 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n12174) );
  OAI211_X1 U14065 ( .C1(n13215), .C2(n11390), .A(n11389), .B(n12174), .ZN(
        n11391) );
  AOI211_X1 U14066 ( .C1(n11393), .C2(n13222), .A(n11392), .B(n11391), .ZN(
        n11394) );
  OAI21_X1 U14067 ( .B1(n11395), .B2(n13226), .A(n11394), .ZN(P3_U3189) );
  OR2_X1 U14068 ( .A1(n11396), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11397) );
  MUX2_X1 U14069 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n11399), .S(n11407), .Z(
        n14202) );
  NAND2_X1 U14070 ( .A1(n11407), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11400) );
  NAND2_X1 U14071 ( .A1(n14201), .A2(n11400), .ZN(n11403) );
  INV_X1 U14072 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n12191) );
  MUX2_X1 U14073 ( .A(n12191), .B(P2_REG2_REG_11__SCAN_IN), .S(n11589), .Z(
        n11402) );
  OR2_X2 U14074 ( .A1(n11403), .A2(n11402), .ZN(n11594) );
  INV_X1 U14075 ( .A(n11594), .ZN(n11401) );
  AOI21_X1 U14076 ( .B1(n11403), .B2(n11402), .A(n11401), .ZN(n11414) );
  INV_X1 U14077 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11408) );
  XOR2_X1 U14078 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n11407), .Z(n14196) );
  XOR2_X1 U14079 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11589), .Z(n11409) );
  OAI211_X1 U14080 ( .C1(n11410), .C2(n11409), .A(n11582), .B(n15537), .ZN(
        n11413) );
  NAND2_X1 U14081 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12251)
         );
  OAI21_X1 U14082 ( .B1(n15543), .B2(n11584), .A(n12251), .ZN(n11411) );
  AOI21_X1 U14083 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(n15525), .A(n11411), 
        .ZN(n11412) );
  OAI211_X1 U14084 ( .C1(n11414), .C2(n14269), .A(n11413), .B(n11412), .ZN(
        P2_U3225) );
  NAND2_X1 U14085 ( .A1(n11355), .A2(n11415), .ZN(n11603) );
  INV_X1 U14086 ( .A(n11603), .ZN(n11418) );
  OAI21_X1 U14087 ( .B1(n11418), .B2(n11417), .A(n11416), .ZN(n11421) );
  OAI211_X1 U14088 ( .C1(n11421), .C2(n11420), .A(n14801), .B(n11419), .ZN(
        n11426) );
  OAI22_X1 U14089 ( .A1(n14824), .A2(n11910), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9571), .ZN(n11423) );
  OAI22_X1 U14090 ( .A1(n14804), .A2(n11805), .B1(n11806), .B2(n14815), .ZN(
        n11422) );
  AOI211_X1 U14091 ( .C1(n11424), .C2(n10664), .A(n11423), .B(n11422), .ZN(
        n11425) );
  NAND2_X1 U14092 ( .A1(n11426), .A2(n11425), .ZN(P1_U3239) );
  NAND2_X1 U14093 ( .A1(n11428), .A2(n11427), .ZN(n11629) );
  XNOR2_X1 U14094 ( .A(n11629), .B(n11429), .ZN(n11497) );
  OAI21_X1 U14095 ( .B1(n11432), .B2(n11431), .A(n11430), .ZN(n11433) );
  NAND2_X1 U14096 ( .A1(n11433), .A2(n11429), .ZN(n11571) );
  OAI21_X1 U14097 ( .B1(n11429), .B2(n11433), .A(n11571), .ZN(n11435) );
  OAI22_X1 U14098 ( .A1(n11434), .A2(n13732), .B1(n13808), .B2(n13734), .ZN(
        n13701) );
  AOI21_X1 U14099 ( .B1(n11435), .B2(n14481), .A(n13701), .ZN(n11496) );
  MUX2_X1 U14100 ( .A(n11436), .B(n11496), .S(n14502), .Z(n11445) );
  NAND2_X1 U14101 ( .A1(n11437), .A2(n13791), .ZN(n11438) );
  NAND2_X1 U14102 ( .A1(n11438), .A2(n14469), .ZN(n11439) );
  NOR2_X1 U14103 ( .A1(n11641), .A2(n11439), .ZN(n11494) );
  NAND2_X1 U14104 ( .A1(n14507), .A2(n11494), .ZN(n11442) );
  INV_X1 U14105 ( .A(n11440), .ZN(n13699) );
  NAND2_X1 U14106 ( .A1(n14510), .A2(n13699), .ZN(n11441) );
  OAI211_X1 U14107 ( .C1(n9970), .C2(n14455), .A(n11442), .B(n11441), .ZN(
        n11443) );
  INV_X1 U14108 ( .A(n11443), .ZN(n11444) );
  OAI211_X1 U14109 ( .C1(n14497), .C2(n11497), .A(n11445), .B(n11444), .ZN(
        P2_U3261) );
  XOR2_X1 U14110 ( .A(n11446), .B(n11447), .Z(n11463) );
  NOR3_X1 U14111 ( .A1(n11383), .A2(n11449), .A3(n11448), .ZN(n11450) );
  OAI21_X1 U14112 ( .B1(n6628), .B2(n11450), .A(n13222), .ZN(n11462) );
  NAND2_X1 U14113 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n11451) );
  OAI21_X1 U14114 ( .B1(n13215), .B2(n11452), .A(n11451), .ZN(n11459) );
  OR3_X1 U14115 ( .A1(n11455), .A2(n11454), .A3(n11453), .ZN(n11456) );
  AOI21_X1 U14116 ( .B1(n11457), .B2(n11456), .A(n13165), .ZN(n11458) );
  AOI211_X1 U14117 ( .C1(n13212), .C2(n11460), .A(n11459), .B(n11458), .ZN(
        n11461) );
  OAI211_X1 U14118 ( .C1(n11463), .C2(n13226), .A(n11462), .B(n11461), .ZN(
        P3_U3190) );
  XNOR2_X1 U14119 ( .A(n11464), .B(n11465), .ZN(n11472) );
  OR2_X1 U14120 ( .A1(n13815), .A2(n13732), .ZN(n11467) );
  NAND2_X1 U14121 ( .A1(n14103), .A2(n13725), .ZN(n11466) );
  AND2_X1 U14122 ( .A1(n11467), .A2(n11466), .ZN(n11536) );
  INV_X1 U14123 ( .A(n11540), .ZN(n11468) );
  NAND2_X1 U14124 ( .A1(n13700), .A2(n11468), .ZN(n11469) );
  NAND2_X1 U14125 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15540) );
  OAI211_X1 U14126 ( .C1(n13726), .C2(n11536), .A(n11469), .B(n15540), .ZN(
        n11470) );
  AOI21_X1 U14127 ( .B1(n14614), .B2(n13751), .A(n11470), .ZN(n11471) );
  OAI21_X1 U14128 ( .B1(n11472), .B2(n13753), .A(n11471), .ZN(P2_U3185) );
  XOR2_X1 U14129 ( .A(n11473), .B(n11474), .Z(n11493) );
  INV_X1 U14130 ( .A(n11475), .ZN(n11479) );
  NAND3_X1 U14131 ( .A1(n11152), .A2(n11477), .A3(n11476), .ZN(n11478) );
  AOI21_X1 U14132 ( .B1(n11479), .B2(n11478), .A(n13165), .ZN(n11491) );
  INV_X1 U14133 ( .A(n11480), .ZN(n11485) );
  NAND3_X1 U14134 ( .A1(n11483), .A2(n11482), .A3(n11481), .ZN(n11484) );
  AOI21_X1 U14135 ( .B1(n11485), .B2(n11484), .A(n13200), .ZN(n11490) );
  NAND2_X1 U14136 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n11487) );
  NAND2_X1 U14137 ( .A1(n15575), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n11486) );
  OAI211_X1 U14138 ( .C1(n13195), .C2(n11488), .A(n11487), .B(n11486), .ZN(
        n11489) );
  NOR3_X1 U14139 ( .A1(n11491), .A2(n11490), .A3(n11489), .ZN(n11492) );
  OAI21_X1 U14140 ( .B1(n11493), .B2(n13226), .A(n11492), .ZN(P3_U3188) );
  INV_X1 U14141 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11499) );
  AOI21_X1 U14142 ( .B1(n15564), .B2(n13791), .A(n11494), .ZN(n11495) );
  OAI211_X1 U14143 ( .C1(n15567), .C2(n11497), .A(n11496), .B(n11495), .ZN(
        n11500) );
  NAND2_X1 U14144 ( .A1(n11500), .A2(n15572), .ZN(n11498) );
  OAI21_X1 U14145 ( .B1(n15572), .B2(n11499), .A(n11498), .ZN(P2_U3442) );
  NAND2_X1 U14146 ( .A1(n11500), .A2(n14618), .ZN(n11501) );
  OAI21_X1 U14147 ( .B1(n14618), .B2(n10996), .A(n11501), .ZN(P2_U3503) );
  OAI22_X1 U14148 ( .A1(n15346), .A2(n11972), .B1(n15518), .B2(n9543), .ZN(
        n11502) );
  INV_X1 U14149 ( .A(n11502), .ZN(n11503) );
  OAI21_X1 U14150 ( .B1(n11504), .B2(n15516), .A(n11503), .ZN(P1_U3532) );
  OAI22_X1 U14151 ( .A1(n15346), .A2(n11987), .B1(n15518), .B2(n10719), .ZN(
        n11505) );
  AOI21_X1 U14152 ( .B1(n11506), .B2(n15518), .A(n11505), .ZN(n11507) );
  INV_X1 U14153 ( .A(n11507), .ZN(P1_U3529) );
  INV_X1 U14154 ( .A(n11508), .ZN(n11511) );
  INV_X1 U14155 ( .A(n14261), .ZN(n14236) );
  OAI222_X1 U14156 ( .A1(n14682), .A2(n11509), .B1(n14673), .B2(n11511), .C1(
        n14236), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U14157 ( .A(n14939), .ZN(n14947) );
  OAI222_X1 U14158 ( .A1(P1_U3086), .A2(n14947), .B1(n15400), .B2(n11511), 
        .C1(n11510), .C2(n15397), .ZN(P1_U3338) );
  INV_X1 U14159 ( .A(n11848), .ZN(n11513) );
  NAND2_X1 U14160 ( .A1(n13106), .A2(n13060), .ZN(n11849) );
  OAI22_X1 U14161 ( .A1(n13078), .A2(n9292), .B1(n11849), .B2(n13071), .ZN(
        n11512) );
  AOI21_X1 U14162 ( .B1(n13044), .B2(n11513), .A(n11512), .ZN(n11514) );
  OAI21_X1 U14163 ( .B1(n11515), .B2(n11859), .A(n11514), .ZN(P3_U3172) );
  INV_X1 U14164 ( .A(n11516), .ZN(n11518) );
  OAI222_X1 U14165 ( .A1(P1_U3086), .A2(n12797), .B1(n15400), .B2(n11518), 
        .C1(n15732), .C2(n15397), .ZN(P1_U3340) );
  OAI222_X1 U14166 ( .A1(P2_U3088), .A2(n7272), .B1(n14673), .B2(n11518), .C1(
        n11517), .C2(n14682), .ZN(P2_U3312) );
  XNOR2_X1 U14167 ( .A(n11603), .B(n11519), .ZN(n11605) );
  XNOR2_X1 U14168 ( .A(n10445), .B(n11605), .ZN(n11523) );
  AND2_X1 U14169 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n14863) );
  OAI22_X1 U14170 ( .A1(n14808), .A2(n11972), .B1(n11971), .B2(n14824), .ZN(
        n11520) );
  AOI211_X1 U14171 ( .C1(n14822), .C2(n11521), .A(n14863), .B(n11520), .ZN(
        n11522) );
  OAI21_X1 U14172 ( .B1(n11523), .B2(n14826), .A(n11522), .ZN(P1_U3230) );
  OAI222_X1 U14173 ( .A1(n13610), .A2(n11525), .B1(n13607), .B2(n11524), .C1(
        P3_U3151), .C2(n9075), .ZN(P3_U3275) );
  INV_X1 U14174 ( .A(n15503), .ZN(n11932) );
  OAI211_X1 U14175 ( .C1(n11528), .C2(n11527), .A(n11526), .B(n14801), .ZN(
        n11533) );
  INV_X1 U14176 ( .A(n11931), .ZN(n11531) );
  OAI22_X1 U14177 ( .A1(n14804), .A2(n11938), .B1(n12075), .B2(n14815), .ZN(
        n11529) );
  AOI211_X1 U14178 ( .C1(n14810), .C2(n11531), .A(n11530), .B(n11529), .ZN(
        n11532) );
  OAI211_X1 U14179 ( .C1(n11932), .C2(n14808), .A(n11533), .B(n11532), .ZN(
        P1_U3213) );
  XOR2_X1 U14180 ( .A(n14049), .B(n11534), .Z(n14617) );
  XOR2_X1 U14181 ( .A(n11535), .B(n14049), .Z(n11538) );
  INV_X1 U14182 ( .A(n11536), .ZN(n11537) );
  AOI21_X1 U14183 ( .B1(n11538), .B2(n14481), .A(n11537), .ZN(n14615) );
  MUX2_X1 U14184 ( .A(n14615), .B(n11539), .S(n14490), .Z(n11543) );
  AOI211_X1 U14185 ( .C1(n14614), .C2(n11579), .A(n14486), .B(n6624), .ZN(
        n14613) );
  OAI22_X1 U14186 ( .A1(n14455), .A2(n10036), .B1(n14485), .B2(n11540), .ZN(
        n11541) );
  AOI21_X1 U14187 ( .B1(n14613), .B2(n14507), .A(n11541), .ZN(n11542) );
  OAI211_X1 U14188 ( .C1(n14497), .C2(n14617), .A(n11543), .B(n11542), .ZN(
        P2_U3258) );
  INV_X1 U14189 ( .A(n11545), .ZN(n11546) );
  NAND2_X1 U14190 ( .A1(n11546), .A2(n9020), .ZN(n11547) );
  XNOR2_X1 U14191 ( .A(n12906), .B(n12038), .ZN(n11550) );
  XNOR2_X1 U14192 ( .A(n11550), .B(n9024), .ZN(n11564) );
  NAND2_X1 U14193 ( .A1(n11550), .A2(n9024), .ZN(n11551) );
  XNOR2_X1 U14194 ( .A(n12906), .B(n15613), .ZN(n11683) );
  XNOR2_X1 U14195 ( .A(n11683), .B(n11684), .ZN(n11552) );
  OAI21_X1 U14196 ( .B1(n11553), .B2(n11552), .A(n11687), .ZN(n11554) );
  NAND2_X1 U14197 ( .A1(n11554), .A2(n13044), .ZN(n11560) );
  NAND2_X1 U14198 ( .A1(n13103), .A2(n13060), .ZN(n11556) );
  NAND2_X1 U14199 ( .A1(n9024), .A2(n13059), .ZN(n11555) );
  AND2_X1 U14200 ( .A1(n11556), .A2(n11555), .ZN(n12020) );
  OAI22_X1 U14201 ( .A1(n12020), .A2(n13071), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11557), .ZN(n11558) );
  AOI21_X1 U14202 ( .B1(n15613), .B2(n13063), .A(n11558), .ZN(n11559) );
  OAI211_X1 U14203 ( .C1(n12023), .C2(n13011), .A(n11560), .B(n11559), .ZN(
        P3_U3170) );
  INV_X1 U14204 ( .A(n11561), .ZN(n11562) );
  AOI211_X1 U14205 ( .C1(n11564), .C2(n11563), .A(n13066), .B(n11562), .ZN(
        n11567) );
  MUX2_X1 U14206 ( .A(n13074), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n11566) );
  AOI22_X1 U14207 ( .A1(n13105), .A2(n13059), .B1(n13060), .B2(n13104), .ZN(
        n12032) );
  OAI22_X1 U14208 ( .A1(n12032), .A2(n13071), .B1(n13078), .B2(n15603), .ZN(
        n11565) );
  OR3_X1 U14209 ( .A1(n11567), .A2(n11566), .A3(n11565), .ZN(P3_U3158) );
  XNOR2_X1 U14210 ( .A(n11569), .B(n11568), .ZN(n11668) );
  NAND2_X1 U14211 ( .A1(n11571), .A2(n11570), .ZN(n11635) );
  INV_X1 U14212 ( .A(n11572), .ZN(n14046) );
  NAND2_X1 U14213 ( .A1(n11635), .A2(n14046), .ZN(n11634) );
  NAND3_X1 U14214 ( .A1(n11634), .A2(n14048), .A3(n11573), .ZN(n11575) );
  AOI21_X1 U14215 ( .B1(n11575), .B2(n11574), .A(n14443), .ZN(n11577) );
  NOR2_X1 U14216 ( .A1(n11577), .A2(n11576), .ZN(n11659) );
  OAI211_X1 U14217 ( .C1(n11578), .C2(n11663), .A(n14469), .B(n11579), .ZN(
        n11661) );
  OAI211_X1 U14218 ( .C1(n15567), .C2(n11668), .A(n11659), .B(n11661), .ZN(
        n11580) );
  INV_X1 U14219 ( .A(n11580), .ZN(n11670) );
  AOI22_X1 U14220 ( .A1(n10388), .A2(n13813), .B1(P2_REG0_REG_6__SCAN_IN), 
        .B2(n15570), .ZN(n11581) );
  OAI21_X1 U14221 ( .B1(n11670), .B2(n15570), .A(n11581), .ZN(P2_U3448) );
  XNOR2_X1 U14222 ( .A(n12261), .B(n12262), .ZN(n11586) );
  AOI21_X1 U14223 ( .B1(n11586), .B2(n11585), .A(n12260), .ZN(n11599) );
  NOR2_X1 U14224 ( .A1(n11587), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12428) );
  INV_X1 U14225 ( .A(n12428), .ZN(n11588) );
  OAI21_X1 U14226 ( .B1(n15543), .B2(n12261), .A(n11588), .ZN(n11597) );
  OR2_X1 U14227 ( .A1(n11589), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11592) );
  NAND2_X1 U14228 ( .A1(n11594), .A2(n11592), .ZN(n11590) );
  MUX2_X1 U14229 ( .A(n12298), .B(P2_REG2_REG_12__SCAN_IN), .S(n12261), .Z(
        n11591) );
  NAND2_X1 U14230 ( .A1(n11590), .A2(n11591), .ZN(n12257) );
  INV_X1 U14231 ( .A(n11591), .ZN(n11593) );
  NAND3_X1 U14232 ( .A1(n11594), .A2(n11593), .A3(n11592), .ZN(n11595) );
  AOI21_X1 U14233 ( .B1(n12257), .B2(n11595), .A(n14269), .ZN(n11596) );
  AOI211_X1 U14234 ( .C1(n15525), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n11597), 
        .B(n11596), .ZN(n11598) );
  OAI21_X1 U14235 ( .B1(n11599), .B2(n15529), .A(n11598), .ZN(P2_U3226) );
  AOI21_X1 U14236 ( .B1(n11602), .B2(n11601), .A(n11600), .ZN(n11607) );
  AOI22_X1 U14237 ( .A1(n11605), .A2(n10445), .B1(n11604), .B2(n11603), .ZN(
        n11606) );
  XOR2_X1 U14238 ( .A(n11607), .B(n11606), .Z(n11611) );
  NAND2_X1 U14239 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n14876) );
  OAI21_X1 U14240 ( .B1(n14824), .B2(n11951), .A(n14876), .ZN(n11609) );
  OAI22_X1 U14241 ( .A1(n14804), .A2(n11939), .B1(n11952), .B2(n14808), .ZN(
        n11608) );
  AOI211_X1 U14242 ( .C1(n14751), .C2(n14849), .A(n11609), .B(n11608), .ZN(
        n11610) );
  OAI21_X1 U14243 ( .B1(n11611), .B2(n14826), .A(n11610), .ZN(P1_U3227) );
  XNOR2_X1 U14244 ( .A(n11826), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n11616) );
  XOR2_X1 U14245 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n11620), .Z(n14908) );
  NAND2_X1 U14246 ( .A1(n14909), .A2(n14908), .ZN(n14907) );
  AOI21_X1 U14247 ( .B1(n11616), .B2(n11615), .A(n11822), .ZN(n11627) );
  NAND2_X1 U14248 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12514)
         );
  INV_X1 U14249 ( .A(n12514), .ZN(n11618) );
  NOR2_X1 U14250 ( .A1(n14959), .A2(n11824), .ZN(n11617) );
  AOI211_X1 U14251 ( .C1(n14945), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11618), 
        .B(n11617), .ZN(n11626) );
  NOR2_X1 U14252 ( .A1(n11619), .A2(n12082), .ZN(n14914) );
  MUX2_X1 U14253 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n12204), .S(n11620), .Z(
        n14913) );
  OAI21_X1 U14254 ( .B1(n14915), .B2(n14914), .A(n14913), .ZN(n14917) );
  NAND2_X1 U14255 ( .A1(n11620), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11622) );
  MUX2_X1 U14256 ( .A(n12235), .B(P1_REG2_REG_11__SCAN_IN), .S(n11826), .Z(
        n11621) );
  INV_X1 U14257 ( .A(n11825), .ZN(n11624) );
  NAND3_X1 U14258 ( .A1(n14917), .A2(n11622), .A3(n11621), .ZN(n11623) );
  NAND3_X1 U14259 ( .A1(n11624), .A2(n14964), .A3(n11623), .ZN(n11625) );
  OAI211_X1 U14260 ( .C1(n11627), .C2(n14940), .A(n11626), .B(n11625), .ZN(
        P1_U3254) );
  INV_X1 U14261 ( .A(n11429), .ZN(n11628) );
  NAND2_X1 U14262 ( .A1(n11629), .A2(n11628), .ZN(n11631) );
  NAND2_X1 U14263 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  XNOR2_X1 U14264 ( .A(n11632), .B(n14046), .ZN(n11699) );
  OR2_X1 U14265 ( .A1(n14473), .A2(n11633), .ZN(n14439) );
  OAI21_X1 U14266 ( .B1(n14046), .B2(n11635), .A(n11634), .ZN(n11639) );
  OR2_X1 U14267 ( .A1(n13815), .A2(n13734), .ZN(n11637) );
  NAND2_X1 U14268 ( .A1(n14107), .A2(n14073), .ZN(n11636) );
  NAND2_X1 U14269 ( .A1(n11637), .A2(n11636), .ZN(n13669) );
  NOR2_X1 U14270 ( .A1(n11699), .A2(n14426), .ZN(n11638) );
  AOI211_X1 U14271 ( .C1(n14481), .C2(n11639), .A(n13669), .B(n11638), .ZN(
        n11697) );
  MUX2_X1 U14272 ( .A(n11640), .B(n11697), .S(n14502), .Z(n11645) );
  INV_X1 U14273 ( .A(n11641), .ZN(n11642) );
  AOI211_X1 U14274 ( .C1(n13806), .C2(n11642), .A(n14486), .B(n11578), .ZN(
        n11695) );
  OAI22_X1 U14275 ( .A1(n14455), .A2(n11701), .B1(n13667), .B2(n14485), .ZN(
        n11643) );
  AOI21_X1 U14276 ( .B1(n14507), .B2(n11695), .A(n11643), .ZN(n11644) );
  OAI211_X1 U14277 ( .C1(n11699), .C2(n14439), .A(n11645), .B(n11644), .ZN(
        P2_U3260) );
  OAI22_X1 U14278 ( .A1(n14455), .A2(n13774), .B1(n14485), .B2(n15522), .ZN(
        n11646) );
  AOI21_X1 U14279 ( .B1(n14507), .B2(n11647), .A(n11646), .ZN(n11651) );
  MUX2_X1 U14280 ( .A(n11649), .B(n11648), .S(n14473), .Z(n11650) );
  OAI211_X1 U14281 ( .C1(n14497), .C2(n11652), .A(n11651), .B(n11650), .ZN(
        P2_U3263) );
  INV_X1 U14282 ( .A(n14439), .ZN(n14509) );
  INV_X1 U14283 ( .A(n14040), .ZN(n11653) );
  NAND2_X1 U14284 ( .A1(n14509), .A2(n11653), .ZN(n11658) );
  OAI21_X1 U14285 ( .B1(n14070), .B2(n11655), .A(n11654), .ZN(n11656) );
  AOI22_X1 U14286 ( .A1(n14502), .A2(n11656), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n14510), .ZN(n11657) );
  OAI211_X1 U14287 ( .C1(n10908), .C2(n14502), .A(n11658), .B(n11657), .ZN(
        P2_U3265) );
  MUX2_X1 U14288 ( .A(n11660), .B(n11659), .S(n14502), .Z(n11667) );
  INV_X1 U14289 ( .A(n11661), .ZN(n11665) );
  OAI22_X1 U14290 ( .A1(n14455), .A2(n11663), .B1(n14485), .B2(n11662), .ZN(
        n11664) );
  AOI21_X1 U14291 ( .B1(n14507), .B2(n11665), .A(n11664), .ZN(n11666) );
  OAI211_X1 U14292 ( .C1(n14497), .C2(n11668), .A(n11667), .B(n11666), .ZN(
        P2_U3259) );
  AOI22_X1 U14293 ( .A1(n14584), .A2(n13813), .B1(n15573), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11669) );
  OAI21_X1 U14294 ( .B1(n11670), .B2(n15573), .A(n11669), .ZN(P2_U3505) );
  XNOR2_X1 U14295 ( .A(n11672), .B(n11671), .ZN(n11674) );
  AOI21_X1 U14296 ( .B1(n11674), .B2(n13493), .A(n11673), .ZN(n11678) );
  XNOR2_X1 U14297 ( .A(n11676), .B(n11675), .ZN(n15584) );
  NAND2_X1 U14298 ( .A1(n15584), .A2(n15627), .ZN(n11677) );
  AND2_X1 U14299 ( .A1(n11678), .A2(n11677), .ZN(n15581) );
  NOR2_X1 U14300 ( .A1(n15621), .A2(n11679), .ZN(n15576) );
  AOI21_X1 U14301 ( .B1(n15584), .B2(n15607), .A(n15576), .ZN(n11680) );
  AND2_X1 U14302 ( .A1(n15581), .A2(n11680), .ZN(n15600) );
  MUX2_X1 U14303 ( .A(n9142), .B(n15600), .S(n15639), .Z(n11681) );
  INV_X1 U14304 ( .A(n11681), .ZN(P3_U3461) );
  XNOR2_X1 U14305 ( .A(n12972), .B(n11682), .ZN(n11862) );
  XNOR2_X1 U14306 ( .A(n11862), .B(n11863), .ZN(n11866) );
  INV_X1 U14307 ( .A(n11683), .ZN(n11685) );
  NAND2_X1 U14308 ( .A1(n11685), .A2(n11684), .ZN(n11686) );
  XOR2_X1 U14309 ( .A(n11867), .B(n11866), .Z(n11694) );
  INV_X1 U14310 ( .A(n12133), .ZN(n11692) );
  NAND2_X1 U14311 ( .A1(n13102), .A2(n13060), .ZN(n11689) );
  NAND2_X1 U14312 ( .A1(n13059), .A2(n13104), .ZN(n11688) );
  NAND2_X1 U14313 ( .A1(n11689), .A2(n11688), .ZN(n12138) );
  AOI22_X1 U14314 ( .A1(n12138), .A2(n13034), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11690) );
  OAI21_X1 U14315 ( .B1(n13078), .B2(n15616), .A(n11690), .ZN(n11691) );
  AOI21_X1 U14316 ( .B1(n13074), .B2(n11692), .A(n11691), .ZN(n11693) );
  OAI21_X1 U14317 ( .B1(n11694), .B2(n13066), .A(n11693), .ZN(P3_U3167) );
  INV_X1 U14318 ( .A(n11695), .ZN(n11696) );
  OAI211_X1 U14319 ( .C1(n11699), .C2(n11698), .A(n11697), .B(n11696), .ZN(
        n11704) );
  INV_X1 U14320 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11700) );
  OAI22_X1 U14321 ( .A1(n14660), .A2(n11701), .B1(n15572), .B2(n11700), .ZN(
        n11702) );
  AOI21_X1 U14322 ( .B1(n11704), .B2(n15572), .A(n11702), .ZN(n11703) );
  INV_X1 U14323 ( .A(n11703), .ZN(P2_U3445) );
  NAND2_X1 U14324 ( .A1(n11704), .A2(n14618), .ZN(n11706) );
  NAND2_X1 U14325 ( .A1(n14584), .A2(n13806), .ZN(n11705) );
  OAI211_X1 U14326 ( .C1(n14618), .C2(n10997), .A(n11706), .B(n11705), .ZN(
        P2_U3504) );
  AOI21_X1 U14327 ( .B1(n11709), .B2(n11708), .A(n11707), .ZN(n11713) );
  AOI22_X1 U14328 ( .A1(n14751), .A2(n14846), .B1(n14812), .B2(n14848), .ZN(
        n11710) );
  NAND2_X1 U14329 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n14893) );
  OAI211_X1 U14330 ( .C1(n11962), .C2(n14824), .A(n11710), .B(n14893), .ZN(
        n11711) );
  AOI21_X1 U14331 ( .B1(n11961), .B2(n10664), .A(n11711), .ZN(n11712) );
  OAI21_X1 U14332 ( .B1(n11713), .B2(n14826), .A(n11712), .ZN(P1_U3221) );
  XNOR2_X1 U14333 ( .A(n11714), .B(n12173), .ZN(n11718) );
  INV_X1 U14334 ( .A(n11718), .ZN(n12114) );
  INV_X1 U14335 ( .A(n15627), .ZN(n15609) );
  AOI22_X1 U14336 ( .A1(n13102), .A2(n13059), .B1(n13060), .B2(n13100), .ZN(
        n12175) );
  OAI211_X1 U14337 ( .C1(n11716), .C2(n12173), .A(n11715), .B(n13493), .ZN(
        n11717) );
  OAI211_X1 U14338 ( .C1(n11718), .C2(n15609), .A(n12175), .B(n11717), .ZN(
        n12111) );
  AOI21_X1 U14339 ( .B1(n15607), .B2(n12114), .A(n12111), .ZN(n11873) );
  NAND2_X1 U14340 ( .A1(n15629), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n11720) );
  OR2_X1 U14341 ( .A1(n13580), .A2(n12110), .ZN(n11719) );
  OAI211_X1 U14342 ( .C1(n11873), .C2(n15629), .A(n11720), .B(n11719), .ZN(
        P3_U3411) );
  INV_X1 U14343 ( .A(n11721), .ZN(n11722) );
  AOI21_X1 U14344 ( .B1(n11724), .B2(n11723), .A(n11722), .ZN(n11731) );
  OR2_X1 U14345 ( .A1(n13837), .A2(n13734), .ZN(n11726) );
  OR2_X1 U14346 ( .A1(n13820), .A2(n13732), .ZN(n11725) );
  AND2_X1 U14347 ( .A1(n11726), .A2(n11725), .ZN(n11754) );
  INV_X1 U14348 ( .A(n11727), .ZN(n11875) );
  NAND2_X1 U14349 ( .A1(n13700), .A2(n11875), .ZN(n11728) );
  NAND2_X1 U14350 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14181) );
  OAI211_X1 U14351 ( .C1(n13726), .C2(n11754), .A(n11728), .B(n14181), .ZN(
        n11729) );
  AOI21_X1 U14352 ( .B1(n13840), .B2(n13751), .A(n11729), .ZN(n11730) );
  OAI21_X1 U14353 ( .B1(n11731), .B2(n13753), .A(n11730), .ZN(P2_U3193) );
  OAI21_X1 U14354 ( .B1(n11734), .B2(n11733), .A(n11732), .ZN(n11956) );
  INV_X1 U14355 ( .A(n11735), .ZN(n11929) );
  INV_X1 U14356 ( .A(n12081), .ZN(n11736) );
  AOI211_X1 U14357 ( .C1(n11961), .C2(n11929), .A(n15187), .B(n11736), .ZN(
        n11964) );
  OAI211_X1 U14358 ( .C1(n6622), .C2(n6861), .A(n15327), .B(n11737), .ZN(
        n11739) );
  AOI22_X1 U14359 ( .A1(n14846), .A2(n15192), .B1(n15190), .B2(n14848), .ZN(
        n11738) );
  NAND2_X1 U14360 ( .A1(n11739), .A2(n11738), .ZN(n11958) );
  AOI211_X1 U14361 ( .C1(n15494), .C2(n11956), .A(n11964), .B(n11958), .ZN(
        n11742) );
  AOI22_X1 U14362 ( .A1(n12215), .A2(n11961), .B1(n15516), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n11740) );
  OAI21_X1 U14363 ( .B1(n11742), .B2(n15516), .A(n11740), .ZN(P1_U3536) );
  AOI22_X1 U14364 ( .A1(n10371), .A2(n11961), .B1(n15510), .B2(
        P1_REG0_REG_8__SCAN_IN), .ZN(n11741) );
  OAI21_X1 U14365 ( .B1(n11742), .B2(n15510), .A(n11741), .ZN(P1_U3483) );
  INV_X1 U14366 ( .A(n14255), .ZN(n14264) );
  OAI222_X1 U14367 ( .A1(P2_U3088), .A2(n14264), .B1(n14673), .B2(n11745), 
        .C1(n11743), .C2(n14682), .ZN(P2_U3309) );
  INV_X1 U14368 ( .A(n14956), .ZN(n14952) );
  OAI222_X1 U14369 ( .A1(P1_U3086), .A2(n14952), .B1(n15400), .B2(n11745), 
        .C1(n11744), .C2(n15397), .ZN(P1_U3337) );
  INV_X1 U14370 ( .A(n11746), .ZN(n11747) );
  AOI21_X1 U14371 ( .B1(n14050), .B2(n11748), .A(n11747), .ZN(n11881) );
  INV_X1 U14372 ( .A(n15567), .ZN(n14589) );
  NAND2_X1 U14373 ( .A1(n11750), .A2(n11749), .ZN(n11751) );
  NAND2_X1 U14374 ( .A1(n11751), .A2(n9980), .ZN(n11752) );
  NAND3_X1 U14375 ( .A1(n11753), .A2(n14481), .A3(n11752), .ZN(n11755) );
  NAND2_X1 U14376 ( .A1(n11755), .A2(n11754), .ZN(n11878) );
  INV_X1 U14377 ( .A(n15564), .ZN(n12726) );
  OAI211_X1 U14378 ( .C1(n7119), .C2(n6624), .A(n14469), .B(n11788), .ZN(
        n11877) );
  OAI21_X1 U14379 ( .B1(n7119), .B2(n12726), .A(n11877), .ZN(n11756) );
  AOI211_X1 U14380 ( .C1(n11881), .C2(n14589), .A(n11878), .B(n11756), .ZN(
        n11759) );
  NAND2_X1 U14381 ( .A1(n15573), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n11757) );
  OAI21_X1 U14382 ( .B1(n11759), .B2(n15573), .A(n11757), .ZN(P2_U3507) );
  NAND2_X1 U14383 ( .A1(n15570), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n11758) );
  OAI21_X1 U14384 ( .B1(n11759), .B2(n15570), .A(n11758), .ZN(P2_U3454) );
  INV_X1 U14385 ( .A(n11762), .ZN(n11763) );
  OR2_X1 U14386 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  XNOR2_X1 U14387 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), 
        .ZN(n11771) );
  XNOR2_X1 U14388 ( .A(n11770), .B(n11771), .ZN(n11769) );
  NAND2_X1 U14389 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n11774), .ZN(n12089) );
  NAND2_X1 U14390 ( .A1(n12091), .A2(n12089), .ZN(n11775) );
  XNOR2_X1 U14391 ( .A(n11775), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n11776) );
  OAI21_X1 U14392 ( .B1(n11777), .B2(n12088), .A(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n11778) );
  OAI21_X1 U14393 ( .B1(n6968), .B2(n12088), .A(n11778), .ZN(SUB_1596_U70) );
  XNOR2_X1 U14394 ( .A(n11780), .B(n11779), .ZN(n14612) );
  OAI211_X1 U14395 ( .C1(n11782), .C2(n14052), .A(n11781), .B(n14481), .ZN(
        n11786) );
  OR2_X1 U14396 ( .A1(n13848), .A2(n13734), .ZN(n11784) );
  NAND2_X1 U14397 ( .A1(n14103), .A2(n14073), .ZN(n11783) );
  NAND2_X1 U14398 ( .A1(n11784), .A2(n11783), .ZN(n11839) );
  INV_X1 U14399 ( .A(n11839), .ZN(n11785) );
  NAND2_X1 U14400 ( .A1(n11786), .A2(n11785), .ZN(n14608) );
  MUX2_X1 U14401 ( .A(n14608), .B(P2_REG2_REG_9__SCAN_IN), .S(n14473), .Z(
        n11787) );
  INV_X1 U14402 ( .A(n11787), .ZN(n11792) );
  AOI211_X1 U14403 ( .C1(n14610), .C2(n11788), .A(n14486), .B(n12006), .ZN(
        n14609) );
  INV_X1 U14404 ( .A(n14610), .ZN(n11789) );
  OAI22_X1 U14405 ( .A1(n11789), .A2(n14455), .B1(n14485), .B2(n11842), .ZN(
        n11790) );
  AOI21_X1 U14406 ( .B1(n14609), .B2(n14507), .A(n11790), .ZN(n11791) );
  OAI211_X1 U14407 ( .C1(n14612), .C2(n14497), .A(n11792), .B(n11791), .ZN(
        P2_U3256) );
  INV_X1 U14408 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n11793) );
  OAI22_X1 U14409 ( .A1(n7043), .A2(n10034), .B1(n14618), .B2(n11793), .ZN(
        n11794) );
  AOI21_X1 U14410 ( .B1(n14618), .B2(n11795), .A(n11794), .ZN(n11796) );
  INV_X1 U14411 ( .A(n11796), .ZN(P2_U3500) );
  NAND2_X1 U14412 ( .A1(n11798), .A2(n11797), .ZN(n11937) );
  INV_X1 U14413 ( .A(n11801), .ZN(n11941) );
  NAND2_X1 U14414 ( .A1(n11937), .A2(n11941), .ZN(n11936) );
  NAND3_X1 U14415 ( .A1(n11936), .A2(n11803), .A3(n11799), .ZN(n11800) );
  AND2_X1 U14416 ( .A1(n11917), .A2(n11800), .ZN(n11915) );
  NAND2_X1 U14417 ( .A1(n11940), .A2(n11801), .ZN(n11943) );
  NAND2_X1 U14418 ( .A1(n11943), .A2(n11802), .ZN(n11804) );
  NAND2_X1 U14419 ( .A1(n11804), .A2(n11803), .ZN(n11921) );
  OAI21_X1 U14420 ( .B1(n11804), .B2(n11803), .A(n11921), .ZN(n11809) );
  OAI22_X1 U14421 ( .A1(n11806), .A2(n15168), .B1(n11805), .B2(n15166), .ZN(
        n11808) );
  NOR2_X1 U14422 ( .A1(n11915), .A2(n15147), .ZN(n11807) );
  AOI211_X1 U14423 ( .C1(n15327), .C2(n11809), .A(n11808), .B(n11807), .ZN(
        n11906) );
  OAI211_X1 U14424 ( .C1(n11810), .C2(n11922), .A(n15283), .B(n11930), .ZN(
        n11908) );
  OAI211_X1 U14425 ( .C1(n11915), .C2(n15507), .A(n11906), .B(n11908), .ZN(
        n11815) );
  INV_X1 U14426 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11811) );
  OAI22_X1 U14427 ( .A1(n15389), .A2(n11922), .B1(n15512), .B2(n11811), .ZN(
        n11812) );
  AOI21_X1 U14428 ( .B1(n11815), .B2(n15512), .A(n11812), .ZN(n11813) );
  INV_X1 U14429 ( .A(n11813), .ZN(P1_U3477) );
  OAI22_X1 U14430 ( .A1(n15346), .A2(n11922), .B1(n15518), .B2(n9574), .ZN(
        n11814) );
  AOI21_X1 U14431 ( .B1(n11815), .B2(n15518), .A(n11814), .ZN(n11816) );
  INV_X1 U14432 ( .A(n11816), .ZN(P1_U3534) );
  NOR2_X1 U14433 ( .A1(n13607), .A2(SI_22_), .ZN(n11817) );
  AOI21_X1 U14434 ( .B1(n11818), .B2(P3_STATE_REG_SCAN_IN), .A(n11817), .ZN(
        n11819) );
  OAI21_X1 U14435 ( .B1(n11820), .B2(n13610), .A(n11819), .ZN(n11821) );
  INV_X1 U14436 ( .A(n11821), .ZN(P3_U3273) );
  XNOR2_X1 U14437 ( .A(n12283), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n12278) );
  XOR2_X1 U14438 ( .A(n12278), .B(n12279), .Z(n11834) );
  MUX2_X1 U14439 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n12323), .S(n12283), .Z(
        n11828) );
  AOI21_X1 U14440 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n11826), .A(n11825), 
        .ZN(n11827) );
  NAND2_X1 U14441 ( .A1(n11827), .A2(n11828), .ZN(n12282) );
  OAI21_X1 U14442 ( .B1(n11828), .B2(n11827), .A(n12282), .ZN(n11832) );
  AND2_X1 U14443 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n12704) );
  AOI21_X1 U14444 ( .B1(n14945), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n12704), 
        .ZN(n11829) );
  OAI21_X1 U14445 ( .B1(n11830), .B2(n14959), .A(n11829), .ZN(n11831) );
  AOI21_X1 U14446 ( .B1(n11832), .B2(n14964), .A(n11831), .ZN(n11833) );
  OAI21_X1 U14447 ( .B1(n11834), .B2(n14940), .A(n11833), .ZN(P1_U3255) );
  OAI21_X1 U14448 ( .B1(n11837), .B2(n11836), .A(n11835), .ZN(n11844) );
  AOI21_X1 U14449 ( .B1(n13746), .B2(n11839), .A(n11838), .ZN(n11841) );
  NAND2_X1 U14450 ( .A1(n14610), .A2(n13751), .ZN(n11840) );
  OAI211_X1 U14451 ( .C1(n13748), .C2(n11842), .A(n11841), .B(n11840), .ZN(
        n11843) );
  AOI21_X1 U14452 ( .B1(n11844), .B2(n13714), .A(n11843), .ZN(n11845) );
  INV_X1 U14453 ( .A(n11845), .ZN(P2_U3203) );
  NAND2_X1 U14454 ( .A1(n11846), .A2(n15621), .ZN(n11847) );
  OR2_X1 U14455 ( .A1(n11848), .A2(n11847), .ZN(n11850) );
  NAND2_X1 U14456 ( .A1(n11850), .A2(n11849), .ZN(n12831) );
  NAND2_X1 U14457 ( .A1(n11852), .A2(n11851), .ZN(n11853) );
  NAND2_X1 U14458 ( .A1(n11853), .A2(n11856), .ZN(n11855) );
  OAI211_X1 U14459 ( .C1(n13582), .C2(n11856), .A(n11855), .B(n11854), .ZN(
        n11858) );
  AND2_X2 U14460 ( .A1(n11858), .A2(n15578), .ZN(n15587) );
  MUX2_X1 U14461 ( .A(n12831), .B(P3_REG2_REG_0__SCAN_IN), .S(n15587), .Z(
        n11861) );
  INV_X1 U14462 ( .A(n15579), .ZN(n15590) );
  NAND2_X1 U14463 ( .A1(n15614), .A2(n15590), .ZN(n11857) );
  OAI22_X1 U14464 ( .A1(n13363), .A2(n9292), .B1(n15578), .B2(n11859), .ZN(
        n11860) );
  OR2_X1 U14465 ( .A1(n11861), .A2(n11860), .ZN(P3_U3233) );
  INV_X1 U14466 ( .A(n11862), .ZN(n11864) );
  AND2_X1 U14467 ( .A1(n11864), .A2(n11863), .ZN(n11865) );
  XNOR2_X1 U14468 ( .A(n12972), .B(n15622), .ZN(n12169) );
  XNOR2_X1 U14469 ( .A(n12169), .B(n13102), .ZN(n11868) );
  OAI211_X1 U14470 ( .C1(n11869), .C2(n11868), .A(n12172), .B(n13044), .ZN(
        n11872) );
  AOI22_X1 U14471 ( .A1(n13103), .A2(n13059), .B1(n13060), .B2(n13101), .ZN(
        n12060) );
  OAI22_X1 U14472 ( .A1(n12060), .A2(n13071), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n7124), .ZN(n11870) );
  AOI21_X1 U14473 ( .B1(n12066), .B2(n13063), .A(n11870), .ZN(n11871) );
  OAI211_X1 U14474 ( .C1(n12064), .C2(n13011), .A(n11872), .B(n11871), .ZN(
        P3_U3179) );
  MUX2_X1 U14475 ( .A(n15659), .B(n11873), .S(n15639), .Z(n11874) );
  OAI21_X1 U14476 ( .B1(n13485), .B2(n12110), .A(n11874), .ZN(P3_U3466) );
  AOI22_X1 U14477 ( .A1(n14511), .A2(n13840), .B1(n14510), .B2(n11875), .ZN(
        n11876) );
  OAI21_X1 U14478 ( .B1(n11877), .B2(n14492), .A(n11876), .ZN(n11880) );
  MUX2_X1 U14479 ( .A(n11878), .B(P2_REG2_REG_8__SCAN_IN), .S(n14473), .Z(
        n11879) );
  AOI211_X1 U14480 ( .C1(n11881), .C2(n14477), .A(n11880), .B(n11879), .ZN(
        n11882) );
  INV_X1 U14481 ( .A(n11882), .ZN(P2_U3257) );
  INV_X1 U14482 ( .A(n11883), .ZN(n11888) );
  AOI21_X1 U14483 ( .B1(n11887), .B2(n11885), .A(n11884), .ZN(n11886) );
  AOI21_X1 U14484 ( .B1(n11888), .B2(n11887), .A(n11886), .ZN(n11900) );
  NAND2_X1 U14485 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n12369) );
  NAND2_X1 U14486 ( .A1(n15575), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11890) );
  OAI211_X1 U14487 ( .C1(n13195), .C2(n11891), .A(n12369), .B(n11890), .ZN(
        n11897) );
  NAND2_X1 U14488 ( .A1(n11893), .A2(n11892), .ZN(n11894) );
  AOI21_X1 U14489 ( .B1(n11895), .B2(n11894), .A(n13200), .ZN(n11896) );
  AOI211_X1 U14490 ( .C1(n13217), .C2(n11898), .A(n11897), .B(n11896), .ZN(
        n11899) );
  OAI21_X1 U14491 ( .B1(n11900), .B2(n13226), .A(n11899), .ZN(P3_U3191) );
  INV_X1 U14492 ( .A(n11901), .ZN(n11904) );
  NOR2_X1 U14493 ( .A1(n11902), .A2(n15791), .ZN(n11903) );
  NAND2_X1 U14494 ( .A1(n11904), .A2(n11903), .ZN(n14989) );
  INV_X2 U14495 ( .A(n15482), .ZN(n15484) );
  NOR2_X1 U14496 ( .A1(n15484), .A2(n11905), .ZN(n15025) );
  INV_X1 U14497 ( .A(n15025), .ZN(n15155) );
  MUX2_X1 U14498 ( .A(n11907), .B(n11906), .S(n15482), .Z(n11914) );
  INV_X1 U14499 ( .A(n11908), .ZN(n11912) );
  OAI22_X1 U14500 ( .A1(n15196), .A2(n11922), .B1(n15208), .B2(n11910), .ZN(
        n11911) );
  AOI21_X1 U14501 ( .B1(n11912), .B2(n15175), .A(n11911), .ZN(n11913) );
  OAI211_X1 U14502 ( .C1(n11915), .C2(n15155), .A(n11914), .B(n11913), .ZN(
        P1_U3287) );
  NAND2_X1 U14503 ( .A1(n11917), .A2(n11916), .ZN(n11919) );
  NAND2_X1 U14504 ( .A1(n11919), .A2(n11920), .ZN(n11918) );
  OAI21_X1 U14505 ( .B1(n11919), .B2(n11920), .A(n11918), .ZN(n11927) );
  INV_X1 U14506 ( .A(n11927), .ZN(n15508) );
  INV_X1 U14507 ( .A(n15147), .ZN(n15015) );
  OAI22_X1 U14508 ( .A1(n11938), .A2(n15166), .B1(n12075), .B2(n15168), .ZN(
        n11926) );
  OAI211_X1 U14509 ( .C1(n11922), .C2(n14849), .A(n11921), .B(n11920), .ZN(
        n11924) );
  AOI21_X1 U14510 ( .B1(n11924), .B2(n11923), .A(n15300), .ZN(n11925) );
  AOI211_X1 U14511 ( .C1(n15015), .C2(n11927), .A(n11926), .B(n11925), .ZN(
        n15506) );
  MUX2_X1 U14512 ( .A(n11928), .B(n15506), .S(n15482), .Z(n11935) );
  AOI211_X1 U14513 ( .C1(n15503), .C2(n11930), .A(n15187), .B(n11735), .ZN(
        n15502) );
  OAI22_X1 U14514 ( .A1(n15196), .A2(n11932), .B1(n11931), .B2(n15208), .ZN(
        n11933) );
  AOI21_X1 U14515 ( .B1(n15502), .B2(n15175), .A(n11933), .ZN(n11934) );
  OAI211_X1 U14516 ( .C1(n15508), .C2(n15155), .A(n11935), .B(n11934), .ZN(
        P1_U3286) );
  OAI21_X1 U14517 ( .B1(n11937), .B2(n11941), .A(n11936), .ZN(n11947) );
  INV_X1 U14518 ( .A(n11947), .ZN(n15499) );
  OAI22_X1 U14519 ( .A1(n11939), .A2(n15166), .B1(n11938), .B2(n15168), .ZN(
        n11946) );
  INV_X1 U14520 ( .A(n11940), .ZN(n11942) );
  NAND2_X1 U14521 ( .A1(n11942), .A2(n11941), .ZN(n11944) );
  AOI21_X1 U14522 ( .B1(n11944), .B2(n11943), .A(n15300), .ZN(n11945) );
  AOI211_X1 U14523 ( .C1(n15015), .C2(n11947), .A(n11946), .B(n11945), .ZN(
        n15498) );
  MUX2_X1 U14524 ( .A(n11948), .B(n15498), .S(n15482), .Z(n11955) );
  INV_X1 U14525 ( .A(n11949), .ZN(n11950) );
  AOI211_X1 U14526 ( .C1(n15496), .C2(n11950), .A(n15187), .B(n11810), .ZN(
        n15495) );
  OAI22_X1 U14527 ( .A1(n15196), .A2(n11952), .B1(n11951), .B2(n15208), .ZN(
        n11953) );
  AOI21_X1 U14528 ( .B1(n15495), .B2(n15175), .A(n11953), .ZN(n11954) );
  OAI211_X1 U14529 ( .C1(n15499), .C2(n15155), .A(n11955), .B(n11954), .ZN(
        P1_U3288) );
  INV_X1 U14530 ( .A(n11956), .ZN(n11967) );
  INV_X1 U14531 ( .A(n11958), .ZN(n11959) );
  MUX2_X1 U14532 ( .A(n11960), .B(n11959), .S(n15482), .Z(n11966) );
  OAI22_X1 U14533 ( .A1(n9924), .A2(n15196), .B1(n15208), .B2(n11962), .ZN(
        n11963) );
  AOI21_X1 U14534 ( .B1(n11964), .B2(n15175), .A(n11963), .ZN(n11965) );
  OAI211_X1 U14535 ( .C1(n11967), .C2(n15478), .A(n11966), .B(n11965), .ZN(
        P1_U3285) );
  INV_X1 U14536 ( .A(n11968), .ZN(n11977) );
  MUX2_X1 U14537 ( .A(n11970), .B(n11969), .S(n15482), .Z(n11976) );
  OAI22_X1 U14538 ( .A1(n15196), .A2(n11972), .B1(n11971), .B2(n15208), .ZN(
        n11973) );
  AOI21_X1 U14539 ( .B1(n15175), .B2(n11974), .A(n11973), .ZN(n11975) );
  OAI211_X1 U14540 ( .C1(n11977), .C2(n15478), .A(n11976), .B(n11975), .ZN(
        P1_U3289) );
  XNOR2_X1 U14541 ( .A(n11978), .B(n11979), .ZN(n11986) );
  OR2_X1 U14542 ( .A1(n13837), .A2(n13732), .ZN(n11981) );
  NAND2_X1 U14543 ( .A1(n14099), .A2(n13725), .ZN(n11980) );
  NAND2_X1 U14544 ( .A1(n11981), .A2(n11980), .ZN(n11998) );
  NOR2_X1 U14545 ( .A1(n11982), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14200) );
  AOI21_X1 U14546 ( .B1(n13746), .B2(n11998), .A(n14200), .ZN(n11983) );
  OAI21_X1 U14547 ( .B1(n12004), .B2(n13748), .A(n11983), .ZN(n11984) );
  AOI21_X1 U14548 ( .B1(n14604), .B2(n13751), .A(n11984), .ZN(n11985) );
  OAI21_X1 U14549 ( .B1(n11986), .B2(n13753), .A(n11985), .ZN(P2_U3189) );
  OAI22_X1 U14550 ( .A1(n15196), .A2(n11987), .B1(n15208), .B2(n15727), .ZN(
        n11990) );
  NOR2_X1 U14551 ( .A1(n15478), .A2(n11988), .ZN(n11989) );
  AOI211_X1 U14552 ( .C1(n15175), .C2(n11991), .A(n11990), .B(n11989), .ZN(
        n11995) );
  MUX2_X1 U14553 ( .A(n11993), .B(n11992), .S(n15482), .Z(n11994) );
  NAND2_X1 U14554 ( .A1(n11995), .A2(n11994), .ZN(P1_U3292) );
  INV_X1 U14555 ( .A(n11996), .ZN(n11997) );
  AOI21_X1 U14556 ( .B1(n11997), .B2(n14054), .A(n14443), .ZN(n12000) );
  AOI21_X1 U14557 ( .B1(n12000), .B2(n11999), .A(n11998), .ZN(n14606) );
  OAI21_X1 U14558 ( .B1(n12002), .B2(n14054), .A(n12001), .ZN(n14607) );
  NAND2_X1 U14559 ( .A1(n14473), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n12003) );
  OAI21_X1 U14560 ( .B1(n14485), .B2(n12004), .A(n12003), .ZN(n12005) );
  AOI21_X1 U14561 ( .B1(n14604), .B2(n14511), .A(n12005), .ZN(n12010) );
  INV_X1 U14562 ( .A(n12006), .ZN(n12007) );
  NAND2_X1 U14563 ( .A1(n12007), .A2(n14604), .ZN(n12008) );
  AND3_X1 U14564 ( .A1(n12008), .A2(n12189), .A3(n14469), .ZN(n14603) );
  NAND2_X1 U14565 ( .A1(n14603), .A2(n14507), .ZN(n12009) );
  OAI211_X1 U14566 ( .C1(n14607), .C2(n14497), .A(n12010), .B(n12009), .ZN(
        n12011) );
  INV_X1 U14567 ( .A(n12011), .ZN(n12012) );
  OAI21_X1 U14568 ( .B1(n14606), .B2(n14490), .A(n12012), .ZN(P2_U3255) );
  OAI222_X1 U14569 ( .A1(P2_U3088), .A2(n12014), .B1(n14685), .B2(n12155), 
        .C1(n12013), .C2(n14682), .ZN(P2_U3307) );
  AND2_X1 U14570 ( .A1(n6432), .A2(n15579), .ZN(n15585) );
  NOR2_X1 U14571 ( .A1(n15627), .A2(n15585), .ZN(n12015) );
  XNOR2_X1 U14572 ( .A(n12016), .B(n12018), .ZN(n15608) );
  OAI211_X1 U14573 ( .C1(n12019), .C2(n12018), .A(n12017), .B(n13493), .ZN(
        n12021) );
  AND2_X1 U14574 ( .A1(n12021), .A2(n12020), .ZN(n15610) );
  MUX2_X1 U14575 ( .A(n15610), .B(n12022), .S(n15587), .Z(n12026) );
  INV_X1 U14576 ( .A(n12023), .ZN(n12024) );
  AOI22_X1 U14577 ( .A1(n13427), .A2(n15613), .B1(n15592), .B2(n12024), .ZN(
        n12025) );
  OAI211_X1 U14578 ( .C1(n13431), .C2(n15608), .A(n12026), .B(n12025), .ZN(
        P3_U3229) );
  NAND2_X1 U14579 ( .A1(n12028), .A2(n12027), .ZN(n12029) );
  XNOR2_X1 U14580 ( .A(n12029), .B(n12030), .ZN(n15605) );
  INV_X1 U14581 ( .A(n15605), .ZN(n12041) );
  AOI21_X1 U14582 ( .B1(n12031), .B2(n12030), .A(n13397), .ZN(n12035) );
  INV_X1 U14583 ( .A(n12032), .ZN(n12033) );
  AOI21_X1 U14584 ( .B1(n12035), .B2(n12034), .A(n12033), .ZN(n15602) );
  MUX2_X1 U14585 ( .A(n15602), .B(n12036), .S(n15587), .Z(n12040) );
  AOI22_X1 U14586 ( .A1(n13427), .A2(n12038), .B1(n15592), .B2(n12037), .ZN(
        n12039) );
  OAI211_X1 U14587 ( .C1(n13431), .C2(n12041), .A(n12040), .B(n12039), .ZN(
        P3_U3230) );
  XNOR2_X1 U14588 ( .A(n12042), .B(n12043), .ZN(n13487) );
  INV_X1 U14589 ( .A(n13487), .ZN(n12054) );
  NAND2_X1 U14590 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  NAND2_X1 U14591 ( .A1(n7792), .A2(n12045), .ZN(n12049) );
  NAND2_X1 U14592 ( .A1(n13099), .A2(n13060), .ZN(n12047) );
  NAND2_X1 U14593 ( .A1(n13059), .A2(n13101), .ZN(n12046) );
  AND2_X1 U14594 ( .A1(n12047), .A2(n12046), .ZN(n12307) );
  INV_X1 U14595 ( .A(n12307), .ZN(n12048) );
  AOI21_X1 U14596 ( .B1(n12049), .B2(n13493), .A(n12048), .ZN(n13489) );
  MUX2_X1 U14597 ( .A(n12050), .B(n13489), .S(n15597), .Z(n12053) );
  INV_X1 U14598 ( .A(n12312), .ZN(n12051) );
  AOI22_X1 U14599 ( .A1(n13427), .A2(n12309), .B1(n15592), .B2(n12051), .ZN(
        n12052) );
  OAI211_X1 U14600 ( .C1(n13431), .C2(n12054), .A(n12053), .B(n12052), .ZN(
        P3_U3225) );
  XNOR2_X1 U14601 ( .A(n12055), .B(n12058), .ZN(n15623) );
  OR2_X1 U14602 ( .A1(n12056), .A2(n12134), .ZN(n12136) );
  NAND2_X1 U14603 ( .A1(n12136), .A2(n12057), .ZN(n12059) );
  XNOR2_X1 U14604 ( .A(n12059), .B(n12058), .ZN(n12062) );
  INV_X1 U14605 ( .A(n12060), .ZN(n12061) );
  AOI21_X1 U14606 ( .B1(n12062), .B2(n13493), .A(n12061), .ZN(n15624) );
  MUX2_X1 U14607 ( .A(n15624), .B(n12063), .S(n15587), .Z(n12068) );
  INV_X1 U14608 ( .A(n12064), .ZN(n12065) );
  AOI22_X1 U14609 ( .A1(n13427), .A2(n12066), .B1(n15592), .B2(n12065), .ZN(
        n12067) );
  OAI211_X1 U14610 ( .C1(n13431), .C2(n15623), .A(n12068), .B(n12067), .ZN(
        P3_U3227) );
  OAI21_X1 U14611 ( .B1(n12070), .B2(n12074), .A(n12069), .ZN(n12214) );
  INV_X1 U14612 ( .A(n12214), .ZN(n12087) );
  INV_X1 U14613 ( .A(n12071), .ZN(n12072) );
  AOI21_X1 U14614 ( .B1(n12074), .B2(n12073), .A(n12072), .ZN(n12079) );
  OR2_X1 U14615 ( .A1(n12075), .A2(n15166), .ZN(n12077) );
  NAND2_X1 U14616 ( .A1(n14845), .A2(n15192), .ZN(n12076) );
  AND2_X1 U14617 ( .A1(n12077), .A2(n12076), .ZN(n12104) );
  NAND2_X1 U14618 ( .A1(n12214), .A2(n15015), .ZN(n12078) );
  OAI211_X1 U14619 ( .C1(n12079), .C2(n15300), .A(n12104), .B(n12078), .ZN(
        n12212) );
  NAND2_X1 U14620 ( .A1(n12212), .A2(n15482), .ZN(n12086) );
  AOI211_X1 U14621 ( .C1(n12217), .C2(n12081), .A(n15187), .B(n12080), .ZN(
        n12213) );
  NOR2_X1 U14622 ( .A1(n7455), .A2(n15196), .ZN(n12084) );
  OAI22_X1 U14623 ( .A1(n15482), .A2(n12082), .B1(n12102), .B2(n15208), .ZN(
        n12083) );
  AOI211_X1 U14624 ( .C1(n12213), .C2(n15175), .A(n12084), .B(n12083), .ZN(
        n12085) );
  OAI211_X1 U14625 ( .C1(n12087), .C2(n15155), .A(n12086), .B(n12085), .ZN(
        P1_U3284) );
  NAND2_X1 U14626 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n12089), .ZN(n12090) );
  NAND2_X1 U14627 ( .A1(n12091), .A2(n12090), .ZN(n12095) );
  INV_X1 U14628 ( .A(n12095), .ZN(n12092) );
  XNOR2_X1 U14629 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n12093) );
  INV_X1 U14630 ( .A(n12093), .ZN(n12094) );
  NAND2_X1 U14631 ( .A1(n12095), .A2(n12094), .ZN(n12096) );
  NAND2_X1 U14632 ( .A1(n12455), .A2(n12096), .ZN(n12449) );
  INV_X1 U14633 ( .A(n12449), .ZN(n12450) );
  XNOR2_X1 U14634 ( .A(n12450), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(n12097) );
  XNOR2_X1 U14635 ( .A(n12452), .B(n12097), .ZN(SUB_1596_U69) );
  INV_X1 U14636 ( .A(n12098), .ZN(n12824) );
  OAI222_X1 U14637 ( .A1(n14682), .A2(n12099), .B1(n14685), .B2(n12824), .C1(
        P2_U3088), .C2(n14031), .ZN(P2_U3308) );
  AOI21_X1 U14638 ( .B1(n6609), .B2(n12101), .A(n12100), .ZN(n12108) );
  NOR2_X1 U14639 ( .A1(n14824), .A2(n12102), .ZN(n12106) );
  INV_X1 U14640 ( .A(n14822), .ZN(n14780) );
  OAI21_X1 U14641 ( .B1(n14780), .B2(n12104), .A(n12103), .ZN(n12105) );
  AOI211_X1 U14642 ( .C1(n12217), .C2(n10664), .A(n12106), .B(n12105), .ZN(
        n12107) );
  OAI21_X1 U14643 ( .B1(n12108), .B2(n14826), .A(n12107), .ZN(P1_U3231) );
  INV_X1 U14644 ( .A(n15585), .ZN(n12109) );
  OR2_X1 U14645 ( .A1(n15587), .A2(n12109), .ZN(n13314) );
  OAI22_X1 U14646 ( .A1(n13363), .A2(n12110), .B1(n12180), .B2(n15578), .ZN(
        n12113) );
  MUX2_X1 U14647 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n12111), .S(n15597), .Z(
        n12112) );
  AOI211_X1 U14648 ( .C1(n12114), .C2(n15594), .A(n12113), .B(n12112), .ZN(
        n12115) );
  INV_X1 U14649 ( .A(n12115), .ZN(P3_U3226) );
  OAI21_X1 U14650 ( .B1(n12117), .B2(n12119), .A(n12116), .ZN(n15493) );
  INV_X1 U14651 ( .A(n15493), .ZN(n12130) );
  NAND3_X1 U14652 ( .A1(n12120), .A2(n12119), .A3(n12118), .ZN(n12121) );
  NAND2_X1 U14653 ( .A1(n12122), .A2(n12121), .ZN(n12123) );
  AOI222_X1 U14654 ( .A1(n15327), .A2(n12123), .B1(n14853), .B2(n15190), .C1(
        n14851), .C2(n15192), .ZN(n15490) );
  MUX2_X1 U14655 ( .A(n12124), .B(n15490), .S(n15482), .Z(n12129) );
  INV_X1 U14656 ( .A(n11110), .ZN(n12126) );
  OAI211_X1 U14657 ( .C1(n12126), .C2(n10469), .A(n15283), .B(n12125), .ZN(
        n15488) );
  OAI22_X1 U14658 ( .A1(n15215), .A2(n15488), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15208), .ZN(n12127) );
  AOI21_X1 U14659 ( .B1(n15212), .B2(n7106), .A(n12127), .ZN(n12128) );
  OAI211_X1 U14660 ( .C1(n12130), .C2(n15478), .A(n12129), .B(n12128), .ZN(
        P1_U3290) );
  XNOR2_X1 U14661 ( .A(n12132), .B(n12131), .ZN(n15617) );
  INV_X1 U14662 ( .A(n15617), .ZN(n12143) );
  OAI22_X1 U14663 ( .A1(n13363), .A2(n15616), .B1(n12133), .B2(n15578), .ZN(
        n12142) );
  NAND2_X1 U14664 ( .A1(n12056), .A2(n12134), .ZN(n12135) );
  NAND2_X1 U14665 ( .A1(n12136), .A2(n12135), .ZN(n12137) );
  NAND2_X1 U14666 ( .A1(n12137), .A2(n13493), .ZN(n12140) );
  INV_X1 U14667 ( .A(n12138), .ZN(n12139) );
  OAI211_X1 U14668 ( .C1(n15609), .C2(n15617), .A(n12140), .B(n12139), .ZN(
        n15619) );
  MUX2_X1 U14669 ( .A(n15619), .B(P3_REG2_REG_5__SCAN_IN), .S(n15587), .Z(
        n12141) );
  AOI211_X1 U14670 ( .C1(n12143), .C2(n15594), .A(n12142), .B(n12141), .ZN(
        n12144) );
  INV_X1 U14671 ( .A(n12144), .ZN(P3_U3228) );
  INV_X1 U14672 ( .A(n12145), .ZN(n12153) );
  OAI22_X1 U14673 ( .A1(n15482), .A2(n9518), .B1(n12146), .B2(n15208), .ZN(
        n12147) );
  AOI21_X1 U14674 ( .B1(n15212), .B2(n12148), .A(n12147), .ZN(n12152) );
  AOI22_X1 U14675 ( .A1(n15025), .A2(n12150), .B1(n15175), .B2(n12149), .ZN(
        n12151) );
  OAI211_X1 U14676 ( .C1(n12153), .C2(n15484), .A(n12152), .B(n12151), .ZN(
        P1_U3291) );
  OAI222_X1 U14677 ( .A1(P1_U3086), .A2(n6435), .B1(n15400), .B2(n12155), .C1(
        n12154), .C2(n15397), .ZN(P1_U3335) );
  NAND2_X1 U14678 ( .A1(n12158), .A2(n12157), .ZN(n12239) );
  OAI21_X1 U14679 ( .B1(n12158), .B2(n12157), .A(n12239), .ZN(n12207) );
  OAI211_X1 U14680 ( .C1(n12161), .C2(n12160), .A(n15327), .B(n12159), .ZN(
        n12198) );
  NOR2_X1 U14681 ( .A1(n12702), .A2(n15168), .ZN(n12201) );
  NOR2_X1 U14682 ( .A1(n12162), .A2(n15166), .ZN(n12200) );
  NOR2_X1 U14683 ( .A1(n12201), .A2(n12200), .ZN(n12352) );
  INV_X1 U14684 ( .A(n12163), .ZN(n12233) );
  OAI211_X1 U14685 ( .C1(n12357), .C2(n12080), .A(n12233), .B(n15283), .ZN(
        n12203) );
  NAND3_X1 U14686 ( .A1(n12198), .A2(n12352), .A3(n12203), .ZN(n12164) );
  AOI21_X1 U14687 ( .B1(n15494), .B2(n12207), .A(n12164), .ZN(n12168) );
  AOI22_X1 U14688 ( .A1(n12166), .A2(n10371), .B1(P1_REG0_REG_10__SCAN_IN), 
        .B2(n15510), .ZN(n12165) );
  OAI21_X1 U14689 ( .B1(n12168), .B2(n15510), .A(n12165), .ZN(P1_U3489) );
  AOI22_X1 U14690 ( .A1(n12166), .A2(n12215), .B1(P1_REG1_REG_10__SCAN_IN), 
        .B2(n15516), .ZN(n12167) );
  OAI21_X1 U14691 ( .B1(n12168), .B2(n15516), .A(n12167), .ZN(P1_U3538) );
  INV_X1 U14692 ( .A(n12169), .ZN(n12170) );
  NAND2_X1 U14693 ( .A1(n12170), .A2(n13102), .ZN(n12171) );
  INV_X1 U14694 ( .A(n12303), .ZN(n12363) );
  NAND2_X1 U14695 ( .A1(n12558), .A2(n12363), .ZN(n12304) );
  OAI211_X1 U14696 ( .C1(n12558), .C2(n12363), .A(n12304), .B(n13044), .ZN(
        n12179) );
  OAI21_X1 U14697 ( .B1(n12175), .B2(n13071), .A(n12174), .ZN(n12176) );
  AOI21_X1 U14698 ( .B1(n12177), .B2(n13063), .A(n12176), .ZN(n12178) );
  OAI211_X1 U14699 ( .C1(n12180), .C2(n13011), .A(n12179), .B(n12178), .ZN(
        P3_U3153) );
  XNOR2_X1 U14700 ( .A(n12181), .B(n10061), .ZN(n12380) );
  INV_X1 U14701 ( .A(n12380), .ZN(n12196) );
  INV_X1 U14702 ( .A(n12182), .ZN(n12183) );
  AOI21_X1 U14703 ( .B1(n12185), .B2(n12184), .A(n12183), .ZN(n12188) );
  OAI22_X1 U14704 ( .A1(n12186), .A2(n13734), .B1(n13848), .B2(n13732), .ZN(
        n12249) );
  INV_X1 U14705 ( .A(n12249), .ZN(n12187) );
  OAI21_X1 U14706 ( .B1(n12188), .B2(n14443), .A(n12187), .ZN(n12378) );
  NAND2_X1 U14707 ( .A1(n12378), .A2(n14502), .ZN(n12195) );
  AOI211_X1 U14708 ( .C1(n13860), .C2(n12189), .A(n14486), .B(n7118), .ZN(
        n12379) );
  INV_X1 U14709 ( .A(n13860), .ZN(n12190) );
  NOR2_X1 U14710 ( .A1(n12190), .A2(n14455), .ZN(n12193) );
  OAI22_X1 U14711 ( .A1(n14502), .A2(n12191), .B1(n12252), .B2(n14485), .ZN(
        n12192) );
  AOI211_X1 U14712 ( .C1(n12379), .C2(n14507), .A(n12193), .B(n12192), .ZN(
        n12194) );
  OAI211_X1 U14713 ( .C1(n14497), .C2(n12196), .A(n12195), .B(n12194), .ZN(
        P2_U3254) );
  INV_X1 U14714 ( .A(n15208), .ZN(n15480) );
  INV_X1 U14715 ( .A(n12197), .ZN(n12354) );
  INV_X1 U14716 ( .A(n12198), .ZN(n12199) );
  AOI211_X1 U14717 ( .C1(n15480), .C2(n12354), .A(n12200), .B(n12199), .ZN(
        n12209) );
  INV_X1 U14718 ( .A(n12201), .ZN(n12202) );
  AOI21_X1 U14719 ( .B1(n12203), .B2(n12202), .A(n15215), .ZN(n12206) );
  OAI22_X1 U14720 ( .A1(n12357), .A2(n15196), .B1(n12204), .B2(n15482), .ZN(
        n12205) );
  AOI211_X1 U14721 ( .C1(n12207), .C2(n15224), .A(n12206), .B(n12205), .ZN(
        n12208) );
  OAI21_X1 U14722 ( .B1(n12209), .B2(n15484), .A(n12208), .ZN(P1_U3283) );
  OAI222_X1 U14723 ( .A1(P2_U3088), .A2(n8505), .B1(n14685), .B2(n12211), .C1(
        n12210), .C2(n14682), .ZN(P2_U3306) );
  AOI211_X1 U14724 ( .C1(n15314), .C2(n12214), .A(n12213), .B(n12212), .ZN(
        n12219) );
  AOI22_X1 U14725 ( .A1(n12217), .A2(n12215), .B1(P1_REG1_REG_9__SCAN_IN), 
        .B2(n15516), .ZN(n12216) );
  OAI21_X1 U14726 ( .B1(n12219), .B2(n15516), .A(n12216), .ZN(P1_U3537) );
  AOI22_X1 U14727 ( .A1(n12217), .A2(n10371), .B1(P1_REG0_REG_9__SCAN_IN), 
        .B2(n15510), .ZN(n12218) );
  OAI21_X1 U14728 ( .B1(n12219), .B2(n15510), .A(n12218), .ZN(P1_U3486) );
  OAI222_X1 U14729 ( .A1(P2_U3088), .A2(n13757), .B1(n14685), .B2(n12221), 
        .C1(n12220), .C2(n14682), .ZN(P2_U3305) );
  OAI222_X1 U14730 ( .A1(P1_U3086), .A2(n12222), .B1(n15400), .B2(n12224), 
        .C1(n15734), .C2(n15397), .ZN(P1_U3331) );
  OAI222_X1 U14731 ( .A1(n12225), .A2(P2_U3088), .B1(n14685), .B2(n12224), 
        .C1(n12223), .C2(n14682), .ZN(P2_U3303) );
  NAND2_X1 U14732 ( .A1(n12226), .A2(n13585), .ZN(n12228) );
  OAI211_X1 U14733 ( .C1(n12229), .C2(n13607), .A(n12228), .B(n12227), .ZN(
        P3_U3272) );
  XNOR2_X1 U14734 ( .A(n12230), .B(n12243), .ZN(n12231) );
  AOI222_X1 U14735 ( .A1(n15327), .A2(n12231), .B1(n14843), .B2(n15192), .C1(
        n14845), .C2(n15190), .ZN(n15351) );
  AOI211_X1 U14736 ( .C1(n15349), .C2(n12233), .A(n15187), .B(n12232), .ZN(
        n15348) );
  NOR2_X1 U14737 ( .A1(n12234), .A2(n15196), .ZN(n12237) );
  OAI22_X1 U14738 ( .A1(n15482), .A2(n12235), .B1(n12516), .B2(n15208), .ZN(
        n12236) );
  AOI211_X1 U14739 ( .C1(n15348), .C2(n15175), .A(n12237), .B(n12236), .ZN(
        n12246) );
  NAND2_X1 U14740 ( .A1(n12239), .A2(n12238), .ZN(n12244) );
  AND2_X1 U14741 ( .A1(n12241), .A2(n12240), .ZN(n12242) );
  OAI21_X1 U14742 ( .B1(n12244), .B2(n12243), .A(n12242), .ZN(n15347) );
  NAND2_X1 U14743 ( .A1(n15347), .A2(n15224), .ZN(n12245) );
  OAI211_X1 U14744 ( .C1(n15351), .C2(n15484), .A(n12246), .B(n12245), .ZN(
        P1_U3282) );
  XNOR2_X1 U14745 ( .A(n12248), .B(n12247), .ZN(n12255) );
  NAND2_X1 U14746 ( .A1(n13746), .A2(n12249), .ZN(n12250) );
  OAI211_X1 U14747 ( .C1(n13748), .C2(n12252), .A(n12251), .B(n12250), .ZN(
        n12253) );
  AOI21_X1 U14748 ( .B1(n13860), .B2(n13751), .A(n12253), .ZN(n12254) );
  OAI21_X1 U14749 ( .B1(n12255), .B2(n13753), .A(n12254), .ZN(P2_U3208) );
  NAND2_X1 U14750 ( .A1(n12261), .A2(n12298), .ZN(n12256) );
  AND2_X1 U14751 ( .A1(n12257), .A2(n12256), .ZN(n14215) );
  MUX2_X1 U14752 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n12258), .S(n12263), .Z(
        n14214) );
  NAND2_X1 U14753 ( .A1(n12263), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12259) );
  XNOR2_X1 U14754 ( .A(n12763), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n12270) );
  INV_X1 U14755 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12264) );
  XOR2_X1 U14756 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n12263), .Z(n14208) );
  XOR2_X1 U14757 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n12764), .Z(n12265) );
  OAI211_X1 U14758 ( .C1(n12266), .C2(n12265), .A(n12770), .B(n15537), .ZN(
        n12269) );
  NAND2_X1 U14759 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n12739)
         );
  OAI21_X1 U14760 ( .B1(n15543), .B2(n12771), .A(n12739), .ZN(n12267) );
  AOI21_X1 U14761 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(n15525), .A(n12267), 
        .ZN(n12268) );
  OAI211_X1 U14762 ( .C1(n12270), .C2(n14269), .A(n12269), .B(n12268), .ZN(
        P2_U3228) );
  XNOR2_X1 U14763 ( .A(n12271), .B(n9032), .ZN(n12274) );
  INV_X1 U14764 ( .A(n12274), .ZN(n12489) );
  AOI22_X1 U14765 ( .A1(n13059), .A2(n13100), .B1(n13060), .B2(n13098), .ZN(
        n12370) );
  OAI211_X1 U14766 ( .C1(n6620), .C2(n9032), .A(n13493), .B(n12272), .ZN(
        n12273) );
  OAI211_X1 U14767 ( .C1(n12274), .C2(n15609), .A(n12370), .B(n12273), .ZN(
        n12486) );
  AOI21_X1 U14768 ( .B1(n15607), .B2(n12489), .A(n12486), .ZN(n12402) );
  OAI22_X1 U14769 ( .A1(n13580), .A2(n12485), .B1(n15631), .B2(n12275), .ZN(
        n12276) );
  INV_X1 U14770 ( .A(n12276), .ZN(n12277) );
  OAI21_X1 U14771 ( .B1(n12402), .B2(n15629), .A(n12277), .ZN(P3_U3417) );
  XNOR2_X1 U14772 ( .A(n12432), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n12281) );
  NOR2_X1 U14773 ( .A1(n12280), .A2(n12281), .ZN(n12431) );
  AOI211_X1 U14774 ( .C1(n12281), .C2(n12280), .A(n14940), .B(n12431), .ZN(
        n12289) );
  OAI21_X1 U14775 ( .B1(n12283), .B2(P1_REG2_REG_12__SCAN_IN), .A(n12282), 
        .ZN(n12285) );
  MUX2_X1 U14776 ( .A(n9668), .B(P1_REG2_REG_13__SCAN_IN), .S(n12432), .Z(
        n12284) );
  AOI211_X1 U14777 ( .C1(n12285), .C2(n12284), .A(n14960), .B(n12441), .ZN(
        n12288) );
  NAND2_X1 U14778 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14778)
         );
  NAND2_X1 U14779 ( .A1(n14945), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n12286) );
  OAI211_X1 U14780 ( .C1(n14959), .C2(n12435), .A(n14778), .B(n12286), .ZN(
        n12287) );
  OR3_X1 U14781 ( .A1(n12289), .A2(n12288), .A3(n12287), .ZN(P1_U3256) );
  INV_X1 U14782 ( .A(n12290), .ZN(n12291) );
  AOI21_X1 U14783 ( .B1(n14055), .B2(n12292), .A(n12291), .ZN(n14602) );
  OAI211_X1 U14784 ( .C1(n12294), .C2(n14055), .A(n12293), .B(n14481), .ZN(
        n14600) );
  INV_X1 U14785 ( .A(n14600), .ZN(n12297) );
  NAND2_X1 U14786 ( .A1(n14097), .A2(n13725), .ZN(n12296) );
  NAND2_X1 U14787 ( .A1(n14099), .A2(n14073), .ZN(n12295) );
  NAND2_X1 U14788 ( .A1(n12296), .A2(n12295), .ZN(n14598) );
  OAI21_X1 U14789 ( .B1(n12297), .B2(n14598), .A(n14502), .ZN(n12302) );
  AOI211_X1 U14790 ( .C1(n14599), .C2(n7807), .A(n14486), .B(n12411), .ZN(
        n14597) );
  NOR2_X1 U14791 ( .A1(n7117), .A2(n14455), .ZN(n12300) );
  OAI22_X1 U14792 ( .A1(n14502), .A2(n12298), .B1(n12426), .B2(n14485), .ZN(
        n12299) );
  AOI211_X1 U14793 ( .C1(n14597), .C2(n14507), .A(n12300), .B(n12299), .ZN(
        n12301) );
  OAI211_X1 U14794 ( .C1(n14602), .C2(n14497), .A(n12302), .B(n12301), .ZN(
        P2_U3253) );
  NAND2_X1 U14795 ( .A1(n12303), .A2(n13101), .ZN(n12367) );
  NAND2_X1 U14796 ( .A1(n12304), .A2(n12367), .ZN(n12306) );
  XNOR2_X1 U14797 ( .A(n12359), .B(n12360), .ZN(n12305) );
  NAND2_X1 U14798 ( .A1(n12306), .A2(n12305), .ZN(n12358) );
  OAI211_X1 U14799 ( .C1(n12306), .C2(n12305), .A(n12358), .B(n13044), .ZN(
        n12311) );
  OAI22_X1 U14800 ( .A1(n12307), .A2(n13071), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n6985), .ZN(n12308) );
  AOI21_X1 U14801 ( .B1(n12309), .B2(n13063), .A(n12308), .ZN(n12310) );
  OAI211_X1 U14802 ( .C1(n12312), .C2(n13011), .A(n12311), .B(n12310), .ZN(
        P3_U3161) );
  OAI21_X1 U14803 ( .B1(n12315), .B2(n12314), .A(n12313), .ZN(n12597) );
  INV_X1 U14804 ( .A(n12597), .ZN(n12328) );
  XNOR2_X1 U14805 ( .A(n12316), .B(n12317), .ZN(n12320) );
  OAI22_X1 U14806 ( .A1(n12702), .A2(n15166), .B1(n12701), .B2(n15168), .ZN(
        n12318) );
  AOI21_X1 U14807 ( .B1(n12597), .B2(n15015), .A(n12318), .ZN(n12319) );
  OAI21_X1 U14808 ( .B1(n15300), .B2(n12320), .A(n12319), .ZN(n12595) );
  NAND2_X1 U14809 ( .A1(n12595), .A2(n15482), .ZN(n12327) );
  INV_X1 U14810 ( .A(n12232), .ZN(n12321) );
  AOI211_X1 U14811 ( .C1(n12322), .C2(n12321), .A(n15187), .B(n6602), .ZN(
        n12596) );
  NOR2_X1 U14812 ( .A1(n12708), .A2(n15196), .ZN(n12325) );
  OAI22_X1 U14813 ( .A1(n15482), .A2(n12323), .B1(n12700), .B2(n15208), .ZN(
        n12324) );
  AOI211_X1 U14814 ( .C1(n12596), .C2(n15175), .A(n12325), .B(n12324), .ZN(
        n12326) );
  OAI211_X1 U14815 ( .C1(n12328), .C2(n15155), .A(n12327), .B(n12326), .ZN(
        P1_U3281) );
  XOR2_X1 U14816 ( .A(n12329), .B(n12331), .Z(n12346) );
  NAND2_X1 U14817 ( .A1(n15639), .A2(n13486), .ZN(n13480) );
  OAI211_X1 U14818 ( .C1(n12331), .C2(n12330), .A(n12521), .B(n13493), .ZN(
        n12334) );
  NAND2_X1 U14819 ( .A1(n13060), .A2(n13097), .ZN(n12332) );
  OAI21_X1 U14820 ( .B1(n12559), .B2(n13048), .A(n12332), .ZN(n12954) );
  INV_X1 U14821 ( .A(n12954), .ZN(n12333) );
  NAND2_X1 U14822 ( .A1(n12334), .A2(n12333), .ZN(n12344) );
  OAI22_X1 U14823 ( .A1(n13485), .A2(n12955), .B1(n15639), .B2(n12335), .ZN(
        n12336) );
  AOI21_X1 U14824 ( .B1(n12344), .B2(n15639), .A(n12336), .ZN(n12337) );
  OAI21_X1 U14825 ( .B1(n12346), .B2(n13480), .A(n12337), .ZN(P3_U3469) );
  NAND2_X1 U14826 ( .A1(n15631), .A2(n13486), .ZN(n13571) );
  INV_X1 U14827 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n12338) );
  OAI22_X1 U14828 ( .A1(n13580), .A2(n12955), .B1(n15631), .B2(n12338), .ZN(
        n12339) );
  AOI21_X1 U14829 ( .B1(n12344), .B2(n15631), .A(n12339), .ZN(n12340) );
  OAI21_X1 U14830 ( .B1(n12346), .B2(n13571), .A(n12340), .ZN(P3_U3420) );
  INV_X1 U14831 ( .A(n12341), .ZN(n12956) );
  AOI22_X1 U14832 ( .A1(n15587), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15592), 
        .B2(n12956), .ZN(n12342) );
  OAI21_X1 U14833 ( .B1(n12955), .B2(n13363), .A(n12342), .ZN(n12343) );
  AOI21_X1 U14834 ( .B1(n12344), .B2(n15597), .A(n12343), .ZN(n12345) );
  OAI21_X1 U14835 ( .B1(n12346), .B2(n13431), .A(n12345), .ZN(P3_U3223) );
  INV_X1 U14836 ( .A(P3_U3897), .ZN(n13107) );
  NAND2_X1 U14837 ( .A1(n13107), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n12347) );
  OAI21_X1 U14838 ( .B1(n12348), .B2(n13107), .A(n12347), .ZN(P3_U3521) );
  OAI211_X1 U14839 ( .C1(n12351), .C2(n12350), .A(n12349), .B(n14801), .ZN(
        n12356) );
  OAI22_X1 U14840 ( .A1(n14780), .A2(n12352), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9629), .ZN(n12353) );
  AOI21_X1 U14841 ( .B1(n12354), .B2(n14810), .A(n12353), .ZN(n12355) );
  OAI211_X1 U14842 ( .C1(n12357), .C2(n14808), .A(n12356), .B(n12355), .ZN(
        P1_U3217) );
  NAND2_X1 U14843 ( .A1(n12359), .A2(n13100), .ZN(n12364) );
  XNOR2_X1 U14844 ( .A(n12485), .B(n12972), .ZN(n12560) );
  XNOR2_X1 U14845 ( .A(n12560), .B(n13099), .ZN(n12365) );
  AOI21_X1 U14846 ( .B1(n12358), .B2(n12364), .A(n12365), .ZN(n12368) );
  INV_X1 U14847 ( .A(n12359), .ZN(n12361) );
  AND2_X1 U14848 ( .A1(n12361), .A2(n12360), .ZN(n12366) );
  INV_X1 U14849 ( .A(n12366), .ZN(n12362) );
  AND2_X1 U14850 ( .A1(n12363), .A2(n12362), .ZN(n12561) );
  AOI21_X1 U14851 ( .B1(n12558), .B2(n12561), .A(n12562), .ZN(n12950) );
  OAI21_X1 U14852 ( .B1(n12368), .B2(n12950), .A(n13044), .ZN(n12374) );
  INV_X1 U14853 ( .A(n12485), .ZN(n12372) );
  OAI21_X1 U14854 ( .B1(n12370), .B2(n13071), .A(n12369), .ZN(n12371) );
  AOI21_X1 U14855 ( .B1(n12372), .B2(n13063), .A(n12371), .ZN(n12373) );
  OAI211_X1 U14856 ( .C1(n12484), .C2(n13011), .A(n12374), .B(n12373), .ZN(
        P3_U3171) );
  INV_X1 U14857 ( .A(n12398), .ZN(n12377) );
  INV_X1 U14858 ( .A(n15397), .ZN(n15394) );
  NAND2_X1 U14859 ( .A1(n15394), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12376) );
  OAI211_X1 U14860 ( .C1(n12377), .C2(n15400), .A(n12376), .B(n12375), .ZN(
        P1_U3332) );
  AOI211_X1 U14861 ( .C1(n14589), .C2(n12380), .A(n12379), .B(n12378), .ZN(
        n12383) );
  AOI22_X1 U14862 ( .A1(n13860), .A2(n14584), .B1(P2_REG1_REG_11__SCAN_IN), 
        .B2(n15573), .ZN(n12381) );
  OAI21_X1 U14863 ( .B1(n12383), .B2(n15573), .A(n12381), .ZN(P2_U3510) );
  AOI22_X1 U14864 ( .A1(n13860), .A2(n10388), .B1(P2_REG0_REG_11__SCAN_IN), 
        .B2(n15570), .ZN(n12382) );
  OAI21_X1 U14865 ( .B1(n12383), .B2(n15570), .A(n12382), .ZN(P2_U3463) );
  AOI21_X1 U14866 ( .B1(n12533), .B2(n12384), .A(n6601), .ZN(n12397) );
  INV_X1 U14867 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n12453) );
  NAND2_X1 U14868 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12609)
         );
  OAI21_X1 U14869 ( .B1(n13215), .B2(n12453), .A(n12609), .ZN(n12390) );
  AOI21_X1 U14870 ( .B1(n12387), .B2(n12386), .A(n12385), .ZN(n12388) );
  NOR2_X1 U14871 ( .A1(n12388), .A2(n13226), .ZN(n12389) );
  AOI211_X1 U14872 ( .C1(n13212), .C2(n12391), .A(n12390), .B(n12389), .ZN(
        n12396) );
  NOR2_X1 U14873 ( .A1(n12392), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n12394) );
  OAI21_X1 U14874 ( .B1(n12394), .B2(n13112), .A(n13217), .ZN(n12395) );
  OAI211_X1 U14875 ( .C1(n12397), .C2(n13200), .A(n12396), .B(n12395), .ZN(
        P3_U3193) );
  NAND2_X1 U14876 ( .A1(n12398), .A2(n14677), .ZN(n12400) );
  OR2_X1 U14877 ( .A1(n12399), .A2(P2_U3088), .ZN(n14078) );
  OAI211_X1 U14878 ( .C1(n12401), .C2(n14682), .A(n12400), .B(n14078), .ZN(
        P2_U3304) );
  INV_X1 U14879 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12403) );
  MUX2_X1 U14880 ( .A(n12403), .B(n12402), .S(n15639), .Z(n12404) );
  OAI21_X1 U14881 ( .B1(n13485), .B2(n12485), .A(n12404), .ZN(P3_U3468) );
  XNOR2_X1 U14882 ( .A(n12405), .B(n14057), .ZN(n14596) );
  NAND3_X1 U14883 ( .A1(n12293), .A2(n6759), .A3(n12407), .ZN(n12408) );
  NAND3_X1 U14884 ( .A1(n12406), .A2(n14481), .A3(n12408), .ZN(n12410) );
  AND2_X1 U14885 ( .A1(n14098), .A2(n14073), .ZN(n12409) );
  AOI21_X1 U14886 ( .B1(n14096), .B2(n13725), .A(n12409), .ZN(n12473) );
  NAND2_X1 U14887 ( .A1(n12410), .A2(n12473), .ZN(n14592) );
  OR2_X1 U14888 ( .A1(n12412), .A2(n12411), .ZN(n12413) );
  AND3_X1 U14889 ( .A1(n12413), .A2(n12499), .A3(n14469), .ZN(n14593) );
  NAND2_X1 U14890 ( .A1(n14593), .A2(n14507), .ZN(n12417) );
  NAND2_X1 U14891 ( .A1(n14473), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12414) );
  OAI21_X1 U14892 ( .B1(n14485), .B2(n12472), .A(n12414), .ZN(n12415) );
  AOI21_X1 U14893 ( .B1(n14594), .B2(n14511), .A(n12415), .ZN(n12416) );
  NAND2_X1 U14894 ( .A1(n12417), .A2(n12416), .ZN(n12418) );
  AOI21_X1 U14895 ( .B1(n14592), .B2(n14502), .A(n12418), .ZN(n12419) );
  OAI21_X1 U14896 ( .B1(n14497), .B2(n14596), .A(n12419), .ZN(P2_U3252) );
  INV_X1 U14897 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n15733) );
  INV_X1 U14898 ( .A(n12975), .ZN(n12420) );
  NAND2_X1 U14899 ( .A1(n12420), .A2(P3_U3897), .ZN(n12421) );
  OAI21_X1 U14900 ( .B1(P3_U3897), .B2(n15733), .A(n12421), .ZN(P3_U3520) );
  OAI21_X1 U14901 ( .B1(n12424), .B2(n12422), .A(n12423), .ZN(n12425) );
  NAND2_X1 U14902 ( .A1(n12425), .A2(n13714), .ZN(n12430) );
  NOR2_X1 U14903 ( .A1(n13748), .A2(n12426), .ZN(n12427) );
  AOI211_X1 U14904 ( .C1(n13746), .C2(n14598), .A(n12428), .B(n12427), .ZN(
        n12429) );
  OAI211_X1 U14905 ( .C1(n7117), .C2(n13738), .A(n12430), .B(n12429), .ZN(
        P2_U3196) );
  XNOR2_X1 U14906 ( .A(n12676), .B(n15344), .ZN(n12434) );
  OAI21_X1 U14907 ( .B1(n12434), .B2(n12433), .A(n12675), .ZN(n12446) );
  INV_X1 U14908 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12679) );
  MUX2_X1 U14909 ( .A(n12679), .B(P1_REG2_REG_14__SCAN_IN), .S(n12676), .Z(
        n12437) );
  NOR2_X1 U14910 ( .A1(n12435), .A2(n9668), .ZN(n12439) );
  INV_X1 U14911 ( .A(n12439), .ZN(n12436) );
  NAND2_X1 U14912 ( .A1(n12437), .A2(n12436), .ZN(n12440) );
  MUX2_X1 U14913 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n12679), .S(n12676), .Z(
        n12438) );
  OAI211_X1 U14914 ( .C1(n12441), .C2(n12440), .A(n12677), .B(n14964), .ZN(
        n12444) );
  NOR2_X1 U14915 ( .A1(n12442), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14693) );
  AOI21_X1 U14916 ( .B1(n14945), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n14693), 
        .ZN(n12443) );
  OAI211_X1 U14917 ( .C1(n14959), .C2(n12678), .A(n12444), .B(n12443), .ZN(
        n12445) );
  AOI21_X1 U14918 ( .B1(n12446), .B2(n14965), .A(n12445), .ZN(n12447) );
  INV_X1 U14919 ( .A(n12447), .ZN(P1_U3257) );
  INV_X1 U14920 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n12448) );
  NOR2_X1 U14921 ( .A1(n12449), .A2(n12448), .ZN(n12451) );
  NAND2_X1 U14922 ( .A1(n12453), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n12454) );
  INV_X1 U14923 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n13122) );
  XNOR2_X1 U14924 ( .A(n13122), .B(P1_ADDR_REG_12__SCAN_IN), .ZN(n12459) );
  INV_X1 U14925 ( .A(n12459), .ZN(n12456) );
  XNOR2_X1 U14926 ( .A(n12460), .B(n12456), .ZN(n12457) );
  NAND2_X1 U14927 ( .A1(n12458), .A2(n12457), .ZN(n12466) );
  INV_X1 U14928 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n12461) );
  NAND2_X1 U14929 ( .A1(n12461), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n12642) );
  INV_X1 U14930 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U14931 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n12462), .ZN(n12640) );
  AND2_X1 U14932 ( .A1(n12642), .A2(n12640), .ZN(n12463) );
  XNOR2_X1 U14933 ( .A(n12641), .B(n12463), .ZN(n12636) );
  INV_X1 U14934 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15665) );
  XNOR2_X1 U14935 ( .A(n12636), .B(n15665), .ZN(n12464) );
  XNOR2_X1 U14936 ( .A(n12639), .B(n12464), .ZN(SUB_1596_U67) );
  NAND2_X1 U14937 ( .A1(n6967), .A2(n12466), .ZN(n12467) );
  XNOR2_X1 U14938 ( .A(n12467), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  INV_X1 U14939 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n15704) );
  NAND2_X1 U14940 ( .A1(n12468), .A2(P3_U3897), .ZN(n12469) );
  OAI21_X1 U14941 ( .B1(P3_U3897), .B2(n15704), .A(n12469), .ZN(P3_U3522) );
  XNOR2_X1 U14942 ( .A(n12470), .B(n12471), .ZN(n12477) );
  NOR2_X1 U14943 ( .A1(n13748), .A2(n12472), .ZN(n12475) );
  NAND2_X1 U14944 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n14210)
         );
  OAI21_X1 U14945 ( .B1(n13726), .B2(n12473), .A(n14210), .ZN(n12474) );
  AOI211_X1 U14946 ( .C1(n14594), .C2(n13751), .A(n12475), .B(n12474), .ZN(
        n12476) );
  OAI21_X1 U14947 ( .B1(n12477), .B2(n13753), .A(n12476), .ZN(P2_U3206) );
  INV_X1 U14948 ( .A(n12478), .ZN(n12482) );
  OAI222_X1 U14949 ( .A1(n12480), .A2(P1_U3086), .B1(n15400), .B2(n12482), 
        .C1(n12479), .C2(n15397), .ZN(P1_U3330) );
  OAI222_X1 U14950 ( .A1(n14682), .A2(n12483), .B1(n14685), .B2(n12482), .C1(
        n12481), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI22_X1 U14951 ( .A1(n13363), .A2(n12485), .B1(n12484), .B2(n15578), .ZN(
        n12488) );
  MUX2_X1 U14952 ( .A(n12486), .B(P3_REG2_REG_9__SCAN_IN), .S(n15587), .Z(
        n12487) );
  AOI211_X1 U14953 ( .C1(n12489), .C2(n15594), .A(n12488), .B(n12487), .ZN(
        n12490) );
  INV_X1 U14954 ( .A(n12490), .ZN(P3_U3224) );
  NAND2_X1 U14955 ( .A1(n12406), .A2(n12491), .ZN(n12494) );
  NOR2_X1 U14956 ( .A1(n12493), .A2(n7772), .ZN(n14059) );
  XNOR2_X1 U14957 ( .A(n12494), .B(n14059), .ZN(n12497) );
  NAND2_X1 U14958 ( .A1(n14095), .A2(n13725), .ZN(n12496) );
  NAND2_X1 U14959 ( .A1(n14097), .A2(n14073), .ZN(n12495) );
  NAND2_X1 U14960 ( .A1(n12496), .A2(n12495), .ZN(n12737) );
  AOI21_X1 U14961 ( .B1(n12497), .B2(n14481), .A(n12737), .ZN(n12731) );
  XNOR2_X1 U14962 ( .A(n12498), .B(n14059), .ZN(n12729) );
  AOI21_X1 U14963 ( .B1(n13880), .B2(n12499), .A(n14486), .ZN(n12501) );
  NAND2_X1 U14964 ( .A1(n12501), .A2(n12718), .ZN(n12725) );
  INV_X1 U14965 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12502) );
  OAI22_X1 U14966 ( .A1(n14502), .A2(n12502), .B1(n12740), .B2(n14485), .ZN(
        n12503) );
  AOI21_X1 U14967 ( .B1(n13880), .B2(n14511), .A(n12503), .ZN(n12504) );
  OAI21_X1 U14968 ( .B1(n12725), .B2(n14492), .A(n12504), .ZN(n12505) );
  AOI21_X1 U14969 ( .B1(n12729), .B2(n14477), .A(n12505), .ZN(n12506) );
  OAI21_X1 U14970 ( .B1(n12731), .B2(n14490), .A(n12506), .ZN(P2_U3251) );
  INV_X1 U14971 ( .A(n12507), .ZN(n12509) );
  OAI222_X1 U14972 ( .A1(n12510), .A2(P3_U3151), .B1(n13610), .B2(n12509), 
        .C1(n12508), .C2(n13607), .ZN(P3_U3271) );
  AOI21_X1 U14973 ( .B1(n12513), .B2(n12512), .A(n12511), .ZN(n12519) );
  AOI22_X1 U14974 ( .A1(n14751), .A2(n14843), .B1(n14812), .B2(n14845), .ZN(
        n12515) );
  OAI211_X1 U14975 ( .C1(n14824), .C2(n12516), .A(n12515), .B(n12514), .ZN(
        n12517) );
  AOI21_X1 U14976 ( .B1(n15349), .B2(n10664), .A(n12517), .ZN(n12518) );
  OAI21_X1 U14977 ( .B1(n12519), .B2(n14826), .A(n12518), .ZN(P1_U3236) );
  INV_X1 U14978 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12528) );
  AND2_X1 U14979 ( .A1(n12521), .A2(n12520), .ZN(n12524) );
  OAI21_X1 U14980 ( .B1(n12524), .B2(n12523), .A(n12522), .ZN(n12527) );
  NAND2_X1 U14981 ( .A1(n13096), .A2(n13060), .ZN(n12526) );
  NAND2_X1 U14982 ( .A1(n13059), .A2(n13098), .ZN(n12525) );
  NAND2_X1 U14983 ( .A1(n12526), .A2(n12525), .ZN(n12608) );
  AOI21_X1 U14984 ( .B1(n12527), .B2(n13493), .A(n12608), .ZN(n12539) );
  MUX2_X1 U14985 ( .A(n12528), .B(n12539), .S(n15631), .Z(n12532) );
  XNOR2_X1 U14986 ( .A(n12529), .B(n12530), .ZN(n12541) );
  INV_X1 U14987 ( .A(n13571), .ZN(n13575) );
  NAND2_X1 U14988 ( .A1(n12541), .A2(n13575), .ZN(n12531) );
  OAI211_X1 U14989 ( .C1(n13580), .C2(n12615), .A(n12532), .B(n12531), .ZN(
        P3_U3423) );
  INV_X1 U14990 ( .A(n12541), .ZN(n12538) );
  MUX2_X1 U14991 ( .A(n12533), .B(n12539), .S(n15597), .Z(n12537) );
  INV_X1 U14992 ( .A(n12615), .ZN(n12535) );
  INV_X1 U14993 ( .A(n12534), .ZN(n12612) );
  AOI22_X1 U14994 ( .A1(n12535), .A2(n13427), .B1(n15592), .B2(n12612), .ZN(
        n12536) );
  OAI211_X1 U14995 ( .C1(n12538), .C2(n13431), .A(n12537), .B(n12536), .ZN(
        P3_U3222) );
  INV_X1 U14996 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n12540) );
  MUX2_X1 U14997 ( .A(n12540), .B(n12539), .S(n15639), .Z(n12543) );
  INV_X1 U14998 ( .A(n13480), .ZN(n13482) );
  NAND2_X1 U14999 ( .A1(n12541), .A2(n13482), .ZN(n12542) );
  OAI211_X1 U15000 ( .C1(n13485), .C2(n12615), .A(n12543), .B(n12542), .ZN(
        P3_U3470) );
  INV_X1 U15001 ( .A(n12544), .ZN(n14782) );
  AOI22_X1 U15002 ( .A1(n15192), .A2(n14841), .B1(n14843), .B2(n15190), .ZN(
        n14779) );
  INV_X1 U15003 ( .A(n14779), .ZN(n12548) );
  XNOR2_X1 U15004 ( .A(n12545), .B(n12546), .ZN(n12547) );
  NOR2_X1 U15005 ( .A1(n12547), .A2(n15300), .ZN(n12662) );
  AOI211_X1 U15006 ( .C1(n15480), .C2(n14782), .A(n12548), .B(n12662), .ZN(
        n12556) );
  OAI21_X1 U15007 ( .B1(n12551), .B2(n12550), .A(n12549), .ZN(n12664) );
  INV_X1 U15008 ( .A(n12552), .ZN(n14785) );
  OAI211_X1 U15009 ( .C1(n14785), .C2(n6602), .A(n12653), .B(n15283), .ZN(
        n12661) );
  AOI22_X1 U15010 ( .A1(n12552), .A2(n15212), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n15484), .ZN(n12553) );
  OAI21_X1 U15011 ( .B1(n12661), .B2(n15215), .A(n12553), .ZN(n12554) );
  AOI21_X1 U15012 ( .B1(n12664), .B2(n15224), .A(n12554), .ZN(n12555) );
  OAI21_X1 U15013 ( .B1(n12556), .B2(n15484), .A(n12555), .ZN(P1_U3280) );
  XNOR2_X1 U15014 ( .A(n12632), .B(n12972), .ZN(n12578) );
  NAND2_X1 U15015 ( .A1(n12578), .A2(n13096), .ZN(n12576) );
  OAI21_X1 U15016 ( .B1(n12578), .B2(n13096), .A(n12576), .ZN(n12569) );
  XNOR2_X1 U15017 ( .A(n12955), .B(n12972), .ZN(n12565) );
  XNOR2_X1 U15018 ( .A(n12565), .B(n13098), .ZN(n12952) );
  NAND2_X1 U15019 ( .A1(n12560), .A2(n12559), .ZN(n12948) );
  OAI211_X1 U15020 ( .C1(n12562), .C2(n12561), .A(n12952), .B(n12948), .ZN(
        n12563) );
  INV_X1 U15021 ( .A(n12563), .ZN(n12564) );
  INV_X1 U15022 ( .A(n12565), .ZN(n12566) );
  NAND2_X1 U15023 ( .A1(n12566), .A2(n13098), .ZN(n12567) );
  XNOR2_X1 U15024 ( .A(n12615), .B(n12972), .ZN(n12580) );
  INV_X1 U15025 ( .A(n12580), .ZN(n12577) );
  NOR2_X1 U15026 ( .A1(n12586), .A2(n12577), .ZN(n12603) );
  NAND2_X1 U15027 ( .A1(n12586), .A2(n12577), .ZN(n12604) );
  OAI21_X1 U15028 ( .B1(n12603), .B2(n12579), .A(n12604), .ZN(n12568) );
  XOR2_X1 U15029 ( .A(n12569), .B(n12568), .Z(n12575) );
  NAND2_X1 U15030 ( .A1(n13095), .A2(n13060), .ZN(n12571) );
  NAND2_X1 U15031 ( .A1(n13059), .A2(n13097), .ZN(n12570) );
  AND2_X1 U15032 ( .A1(n12571), .A2(n12570), .ZN(n12621) );
  NAND2_X1 U15033 ( .A1(n13074), .A2(n12631), .ZN(n12572) );
  NAND2_X1 U15034 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13121)
         );
  OAI211_X1 U15035 ( .C1(n12621), .C2(n13071), .A(n12572), .B(n13121), .ZN(
        n12573) );
  AOI21_X1 U15036 ( .B1(n12632), .B2(n13063), .A(n12573), .ZN(n12574) );
  OAI21_X1 U15037 ( .B1(n12575), .B2(n13066), .A(n12574), .ZN(P3_U3164) );
  OAI21_X1 U15038 ( .B1(n12579), .B2(n12580), .A(n12576), .ZN(n12585) );
  OAI21_X1 U15039 ( .B1(n12577), .B2(n13097), .A(n13096), .ZN(n12583) );
  INV_X1 U15040 ( .A(n12578), .ZN(n12582) );
  AND2_X1 U15041 ( .A1(n12579), .A2(n12589), .ZN(n12581) );
  XNOR2_X1 U15042 ( .A(n12757), .B(n12972), .ZN(n12686) );
  XNOR2_X1 U15043 ( .A(n12686), .B(n13095), .ZN(n12587) );
  XNOR2_X1 U15044 ( .A(n12688), .B(n12587), .ZN(n12593) );
  NAND2_X1 U15045 ( .A1(n13060), .A2(n13094), .ZN(n12588) );
  OAI21_X1 U15046 ( .B1(n12589), .B2(n13048), .A(n12588), .ZN(n12745) );
  AND2_X1 U15047 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13143) );
  AOI21_X1 U15048 ( .B1(n12745), .B2(n13034), .A(n13143), .ZN(n12591) );
  NAND2_X1 U15049 ( .A1(n13074), .A2(n12758), .ZN(n12590) );
  OAI211_X1 U15050 ( .C1(n12757), .C2(n13078), .A(n12591), .B(n12590), .ZN(
        n12592) );
  AOI21_X1 U15051 ( .B1(n12593), .B2(n13044), .A(n12592), .ZN(n12594) );
  INV_X1 U15052 ( .A(n12594), .ZN(P3_U3174) );
  INV_X1 U15053 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12598) );
  AOI211_X1 U15054 ( .C1(n15314), .C2(n12597), .A(n12596), .B(n12595), .ZN(
        n12600) );
  MUX2_X1 U15055 ( .A(n12598), .B(n12600), .S(n15512), .Z(n12599) );
  OAI21_X1 U15056 ( .B1(n12708), .B2(n15389), .A(n12599), .ZN(P1_U3495) );
  MUX2_X1 U15057 ( .A(n12601), .B(n12600), .S(n15518), .Z(n12602) );
  OAI21_X1 U15058 ( .B1(n12708), .B2(n15346), .A(n12602), .ZN(P1_U3540) );
  INV_X1 U15059 ( .A(n12603), .ZN(n12605) );
  NAND2_X1 U15060 ( .A1(n12605), .A2(n12604), .ZN(n12606) );
  XNOR2_X1 U15061 ( .A(n12606), .B(n13097), .ZN(n12607) );
  NAND2_X1 U15062 ( .A1(n12607), .A2(n13044), .ZN(n12614) );
  NAND2_X1 U15063 ( .A1(n12608), .A2(n13034), .ZN(n12610) );
  NAND2_X1 U15064 ( .A1(n12610), .A2(n12609), .ZN(n12611) );
  AOI21_X1 U15065 ( .B1(n13074), .B2(n12612), .A(n12611), .ZN(n12613) );
  OAI211_X1 U15066 ( .C1(n13078), .C2(n12615), .A(n12614), .B(n12613), .ZN(
        P3_U3176) );
  XOR2_X1 U15067 ( .A(n12616), .B(n12617), .Z(n12635) );
  NAND2_X1 U15068 ( .A1(n12618), .A2(n12617), .ZN(n12619) );
  NAND3_X1 U15069 ( .A1(n12620), .A2(n13493), .A3(n12619), .ZN(n12622) );
  AND2_X1 U15070 ( .A1(n12622), .A2(n12621), .ZN(n12630) );
  MUX2_X1 U15071 ( .A(n12630), .B(n12623), .S(n15637), .Z(n12625) );
  NAND2_X1 U15072 ( .A1(n12632), .A2(n13471), .ZN(n12624) );
  OAI211_X1 U15073 ( .C1(n13480), .C2(n12635), .A(n12625), .B(n12624), .ZN(
        P3_U3471) );
  MUX2_X1 U15074 ( .A(n12626), .B(n12630), .S(n15631), .Z(n12628) );
  NAND2_X1 U15075 ( .A1(n12632), .A2(n9136), .ZN(n12627) );
  OAI211_X1 U15076 ( .C1(n12635), .C2(n13571), .A(n12628), .B(n12627), .ZN(
        P3_U3426) );
  MUX2_X1 U15077 ( .A(n12630), .B(n12629), .S(n15587), .Z(n12634) );
  AOI22_X1 U15078 ( .A1(n12632), .A2(n13427), .B1(n15592), .B2(n12631), .ZN(
        n12633) );
  OAI211_X1 U15079 ( .C1(n12635), .C2(n13431), .A(n12634), .B(n12633), .ZN(
        P3_U3221) );
  NAND2_X1 U15080 ( .A1(n12636), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n12638) );
  INV_X1 U15081 ( .A(n12636), .ZN(n12637) );
  NAND2_X1 U15082 ( .A1(n12641), .A2(n12640), .ZN(n12643) );
  NAND2_X1 U15083 ( .A1(n12643), .A2(n12642), .ZN(n15412) );
  INV_X1 U15084 ( .A(n15412), .ZN(n12645) );
  XOR2_X1 U15085 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n12644) );
  XNOR2_X1 U15086 ( .A(n12645), .B(n12644), .ZN(n15408) );
  XNOR2_X1 U15087 ( .A(n15408), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(n12646) );
  XNOR2_X1 U15088 ( .A(n15409), .B(n12646), .ZN(SUB_1596_U66) );
  OAI22_X1 U15089 ( .A1(n14746), .A2(n15168), .B1(n12701), .B2(n15166), .ZN(
        n15340) );
  XNOR2_X1 U15090 ( .A(n12647), .B(n12648), .ZN(n12649) );
  NOR2_X1 U15091 ( .A1(n12649), .A2(n15300), .ZN(n15342) );
  AOI211_X1 U15092 ( .C1(n15480), .C2(n14692), .A(n15340), .B(n15342), .ZN(
        n12660) );
  INV_X1 U15093 ( .A(n12650), .ZN(n12652) );
  NAND2_X1 U15094 ( .A1(n12652), .A2(n12651), .ZN(n15204) );
  OAI21_X1 U15095 ( .B1(n12652), .B2(n12651), .A(n15204), .ZN(n15339) );
  AOI22_X1 U15096 ( .A1(n15338), .A2(n15212), .B1(n15484), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n12657) );
  NAND2_X1 U15097 ( .A1(n15338), .A2(n12653), .ZN(n12654) );
  NAND2_X1 U15098 ( .A1(n12654), .A2(n15283), .ZN(n12655) );
  NOR2_X1 U15099 ( .A1(n15207), .A2(n12655), .ZN(n15341) );
  NAND2_X1 U15100 ( .A1(n15341), .A2(n15175), .ZN(n12656) );
  OAI211_X1 U15101 ( .C1(n15339), .C2(n15478), .A(n12657), .B(n12656), .ZN(
        n12658) );
  INV_X1 U15102 ( .A(n12658), .ZN(n12659) );
  OAI21_X1 U15103 ( .B1(n12660), .B2(n15484), .A(n12659), .ZN(P1_U3279) );
  NAND2_X1 U15104 ( .A1(n12661), .A2(n14779), .ZN(n12663) );
  AOI211_X1 U15105 ( .C1(n15494), .C2(n12664), .A(n12663), .B(n12662), .ZN(
        n12666) );
  MUX2_X1 U15106 ( .A(n15772), .B(n12666), .S(n15512), .Z(n12665) );
  OAI21_X1 U15107 ( .B1(n14785), .B2(n15389), .A(n12665), .ZN(P1_U3498) );
  MUX2_X1 U15108 ( .A(n12667), .B(n12666), .S(n15518), .Z(n12668) );
  OAI21_X1 U15109 ( .B1(n14785), .B2(n15346), .A(n12668), .ZN(P1_U3541) );
  INV_X1 U15110 ( .A(n12669), .ZN(n12673) );
  OAI222_X1 U15111 ( .A1(n12671), .A2(P2_U3088), .B1(n14685), .B2(n12673), 
        .C1(n12670), .C2(n14682), .ZN(P2_U3301) );
  OAI222_X1 U15112 ( .A1(P1_U3086), .A2(n12674), .B1(n15400), .B2(n12673), 
        .C1(n12672), .C2(n15397), .ZN(P1_U3329) );
  XNOR2_X1 U15113 ( .A(n12793), .B(n15336), .ZN(n12685) );
  NAND2_X1 U15114 ( .A1(n12680), .A2(n15210), .ZN(n12800) );
  OAI21_X1 U15115 ( .B1(n12680), .B2(n15210), .A(n12800), .ZN(n12683) );
  NOR2_X1 U15116 ( .A1(n15692), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14821) );
  AOI21_X1 U15117 ( .B1(n14945), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n14821), 
        .ZN(n12681) );
  OAI21_X1 U15118 ( .B1(n12797), .B2(n14959), .A(n12681), .ZN(n12682) );
  AOI21_X1 U15119 ( .B1(n12683), .B2(n14964), .A(n12682), .ZN(n12684) );
  OAI21_X1 U15120 ( .B1(n12685), .B2(n14940), .A(n12684), .ZN(P1_U3258) );
  XNOR2_X1 U15121 ( .A(n13579), .B(n12972), .ZN(n12901) );
  XNOR2_X1 U15122 ( .A(n12901), .B(n13094), .ZN(n12898) );
  XNOR2_X1 U15123 ( .A(n12899), .B(n12898), .ZN(n12689) );
  NAND2_X1 U15124 ( .A1(n12689), .A2(n13044), .ZN(n12696) );
  NAND2_X1 U15125 ( .A1(n13093), .A2(n13060), .ZN(n12691) );
  NAND2_X1 U15126 ( .A1(n13095), .A2(n13059), .ZN(n12690) );
  NAND2_X1 U15127 ( .A1(n12691), .A2(n12690), .ZN(n13423) );
  NAND2_X1 U15128 ( .A1(n13423), .A2(n13034), .ZN(n12693) );
  NAND2_X1 U15129 ( .A1(n12693), .A2(n12692), .ZN(n12694) );
  AOI21_X1 U15130 ( .B1(n13074), .B2(n13426), .A(n12694), .ZN(n12695) );
  OAI211_X1 U15131 ( .C1(n13078), .C2(n13579), .A(n12696), .B(n12695), .ZN(
        P3_U3155) );
  OAI211_X1 U15132 ( .C1(n12699), .C2(n12698), .A(n12697), .B(n14801), .ZN(
        n12707) );
  INV_X1 U15133 ( .A(n12700), .ZN(n12705) );
  OAI22_X1 U15134 ( .A1(n14804), .A2(n12702), .B1(n12701), .B2(n14815), .ZN(
        n12703) );
  AOI211_X1 U15135 ( .C1(n14810), .C2(n12705), .A(n12704), .B(n12703), .ZN(
        n12706) );
  OAI211_X1 U15136 ( .C1(n12708), .C2(n14808), .A(n12707), .B(n12706), .ZN(
        P1_U3224) );
  INV_X1 U15137 ( .A(n12709), .ZN(n14684) );
  AOI21_X1 U15138 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n15394), .A(n12710), 
        .ZN(n12711) );
  OAI21_X1 U15139 ( .B1(n14684), .B2(n15400), .A(n12711), .ZN(P1_U3328) );
  XNOR2_X1 U15140 ( .A(n12712), .B(n14060), .ZN(n12715) );
  OAI22_X1 U15141 ( .A1(n12713), .A2(n13734), .B1(n13882), .B2(n13732), .ZN(
        n13745) );
  INV_X1 U15142 ( .A(n13745), .ZN(n12714) );
  OAI21_X1 U15143 ( .B1(n12715), .B2(n14443), .A(n12714), .ZN(n14586) );
  INV_X1 U15144 ( .A(n14586), .ZN(n12724) );
  XNOR2_X1 U15145 ( .A(n12716), .B(n14060), .ZN(n14588) );
  INV_X1 U15146 ( .A(n14487), .ZN(n12717) );
  AOI211_X1 U15147 ( .C1(n13887), .C2(n12718), .A(n14486), .B(n12717), .ZN(
        n14587) );
  NAND2_X1 U15148 ( .A1(n14587), .A2(n14507), .ZN(n12721) );
  INV_X1 U15149 ( .A(n13749), .ZN(n12719) );
  AOI22_X1 U15150 ( .A1(n14473), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12719), 
        .B2(n14510), .ZN(n12720) );
  OAI211_X1 U15151 ( .C1(n10039), .C2(n14455), .A(n12721), .B(n12720), .ZN(
        n12722) );
  AOI21_X1 U15152 ( .B1(n14477), .B2(n14588), .A(n12722), .ZN(n12723) );
  OAI21_X1 U15153 ( .B1(n14473), .B2(n12724), .A(n12723), .ZN(P2_U3250) );
  INV_X1 U15154 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n15719) );
  INV_X1 U15155 ( .A(n13880), .ZN(n12727) );
  OAI21_X1 U15156 ( .B1(n12727), .B2(n12726), .A(n12725), .ZN(n12728) );
  AOI21_X1 U15157 ( .B1(n12729), .B2(n14589), .A(n12728), .ZN(n12730) );
  AND2_X1 U15158 ( .A1(n12731), .A2(n12730), .ZN(n12733) );
  MUX2_X1 U15159 ( .A(n15719), .B(n12733), .S(n15572), .Z(n12732) );
  INV_X1 U15160 ( .A(n12732), .ZN(P2_U3472) );
  MUX2_X1 U15161 ( .A(n12772), .B(n12733), .S(n14618), .Z(n12734) );
  INV_X1 U15162 ( .A(n12734), .ZN(P2_U3513) );
  AOI21_X1 U15163 ( .B1(n12736), .B2(n12735), .A(n6614), .ZN(n12743) );
  NAND2_X1 U15164 ( .A1(n13746), .A2(n12737), .ZN(n12738) );
  OAI211_X1 U15165 ( .C1(n13748), .C2(n12740), .A(n12739), .B(n12738), .ZN(
        n12741) );
  AOI21_X1 U15166 ( .B1(n13880), .B2(n13751), .A(n12741), .ZN(n12742) );
  OAI21_X1 U15167 ( .B1(n12743), .B2(n13753), .A(n12742), .ZN(P2_U3187) );
  XNOR2_X1 U15168 ( .A(n12744), .B(n12749), .ZN(n12746) );
  AOI21_X1 U15169 ( .B1(n12746), .B2(n13493), .A(n12745), .ZN(n12756) );
  MUX2_X1 U15170 ( .A(n12756), .B(n12747), .S(n15629), .Z(n12751) );
  XNOR2_X1 U15171 ( .A(n12748), .B(n12749), .ZN(n12754) );
  NAND2_X1 U15172 ( .A1(n12754), .A2(n13575), .ZN(n12750) );
  OAI211_X1 U15173 ( .C1(n13580), .C2(n12757), .A(n12751), .B(n12750), .ZN(
        P3_U3429) );
  MUX2_X1 U15174 ( .A(n12756), .B(n13134), .S(n15637), .Z(n12753) );
  NAND2_X1 U15175 ( .A1(n12754), .A2(n13482), .ZN(n12752) );
  OAI211_X1 U15176 ( .C1(n13485), .C2(n12757), .A(n12753), .B(n12752), .ZN(
        P3_U3472) );
  INV_X1 U15177 ( .A(n12754), .ZN(n12762) );
  MUX2_X1 U15178 ( .A(n12756), .B(n12755), .S(n15587), .Z(n12761) );
  INV_X1 U15179 ( .A(n12757), .ZN(n12759) );
  AOI22_X1 U15180 ( .A1(n12759), .A2(n13427), .B1(n15592), .B2(n12758), .ZN(
        n12760) );
  OAI211_X1 U15181 ( .C1(n12762), .C2(n13431), .A(n12761), .B(n12760), .ZN(
        P3_U3220) );
  NAND2_X1 U15182 ( .A1(n12765), .A2(n12764), .ZN(n12766) );
  NAND2_X1 U15183 ( .A1(n12767), .A2(n12766), .ZN(n14229) );
  XNOR2_X1 U15184 ( .A(n14229), .B(n7272), .ZN(n14227) );
  XNOR2_X1 U15185 ( .A(n14227), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n12777) );
  OR2_X1 U15186 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12768), .ZN(n12769) );
  OAI21_X1 U15187 ( .B1(n15543), .B2(n7272), .A(n12769), .ZN(n12775) );
  AOI211_X1 U15188 ( .C1(n12773), .C2(n14590), .A(n15529), .B(n14221), .ZN(
        n12774) );
  AOI211_X1 U15189 ( .C1(n15525), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n12775), 
        .B(n12774), .ZN(n12776) );
  OAI21_X1 U15190 ( .B1(n12777), .B2(n14269), .A(n12776), .ZN(P2_U3229) );
  XNOR2_X1 U15191 ( .A(n12778), .B(n12782), .ZN(n13572) );
  NAND2_X1 U15192 ( .A1(n13420), .A2(n12779), .ZN(n12781) );
  AND2_X1 U15193 ( .A1(n12781), .A2(n12780), .ZN(n12783) );
  XNOR2_X1 U15194 ( .A(n12783), .B(n12782), .ZN(n12784) );
  AOI22_X1 U15195 ( .A1(n13092), .A2(n13060), .B1(n13059), .B2(n13094), .ZN(
        n13072) );
  OAI21_X1 U15196 ( .B1(n12784), .B2(n13397), .A(n13072), .ZN(n13476) );
  NAND2_X1 U15197 ( .A1(n13476), .A2(n15597), .ZN(n12789) );
  INV_X1 U15198 ( .A(n13075), .ZN(n12785) );
  OAI22_X1 U15199 ( .A1(n15597), .A2(n12786), .B1(n12785), .B2(n15578), .ZN(
        n12787) );
  AOI21_X1 U15200 ( .B1(n13477), .B2(n13427), .A(n12787), .ZN(n12788) );
  OAI211_X1 U15201 ( .C1(n13572), .C2(n13431), .A(n12789), .B(n12788), .ZN(
        P3_U3218) );
  XNOR2_X1 U15202 ( .A(n14922), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12795) );
  INV_X1 U15203 ( .A(n12797), .ZN(n12792) );
  INV_X1 U15204 ( .A(n12790), .ZN(n12791) );
  NOR2_X1 U15205 ( .A1(n12794), .A2(n12795), .ZN(n14921) );
  AOI211_X1 U15206 ( .C1(n12795), .C2(n12794), .A(n14940), .B(n14921), .ZN(
        n12807) );
  INV_X1 U15207 ( .A(n12796), .ZN(n12798) );
  NAND2_X1 U15208 ( .A1(n12798), .A2(n12797), .ZN(n12799) );
  AND2_X1 U15209 ( .A1(n12800), .A2(n12799), .ZN(n12802) );
  XOR2_X1 U15210 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n14922), .Z(n12801) );
  NAND3_X1 U15211 ( .A1(n12800), .A2(n12801), .A3(n12799), .ZN(n14925) );
  OAI211_X1 U15212 ( .C1(n12802), .C2(n12801), .A(n14964), .B(n14925), .ZN(
        n12805) );
  NOR2_X1 U15213 ( .A1(n12803), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14748) );
  AOI21_X1 U15214 ( .B1(n14945), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14748), 
        .ZN(n12804) );
  OAI211_X1 U15215 ( .C1(n14959), .C2(n14927), .A(n12805), .B(n12804), .ZN(
        n12806) );
  OR2_X1 U15216 ( .A1(n12807), .A2(n12806), .ZN(P1_U3259) );
  INV_X1 U15217 ( .A(n12808), .ZN(n12809) );
  OAI222_X1 U15218 ( .A1(n13607), .A2(n12810), .B1(P3_U3151), .B2(n7509), .C1(
        n13610), .C2(n12809), .ZN(P3_U3265) );
  INV_X1 U15219 ( .A(n12811), .ZN(n12812) );
  OAI222_X1 U15220 ( .A1(n13598), .A2(n15760), .B1(P3_U3151), .B2(n12813), 
        .C1(n13610), .C2(n12812), .ZN(P3_U3267) );
  XNOR2_X1 U15221 ( .A(n12815), .B(n12814), .ZN(n12822) );
  OAI22_X1 U15222 ( .A1(n12817), .A2(n14824), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12816), .ZN(n12818) );
  AOI21_X1 U15223 ( .B1(n14834), .B2(n14812), .A(n12818), .ZN(n12819) );
  OAI21_X1 U15224 ( .B1(n15013), .B2(n14815), .A(n12819), .ZN(n12820) );
  AOI21_X1 U15225 ( .B1(n15258), .B2(n10664), .A(n12820), .ZN(n12821) );
  OAI21_X1 U15226 ( .B1(n12822), .B2(n14826), .A(n12821), .ZN(P1_U3214) );
  OAI222_X1 U15227 ( .A1(n14967), .A2(P1_U3086), .B1(n15400), .B2(n12824), 
        .C1(n12823), .C2(n15397), .ZN(P1_U3336) );
  OAI222_X1 U15228 ( .A1(n13610), .A2(n12827), .B1(n13607), .B2(n12826), .C1(
        P3_U3151), .C2(n12825), .ZN(P3_U3274) );
  OAI21_X1 U15229 ( .B1(n14288), .B2(n7043), .A(n12830), .ZN(P2_U3530) );
  INV_X1 U15230 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n12832) );
  INV_X1 U15231 ( .A(n12831), .ZN(n12835) );
  MUX2_X1 U15232 ( .A(n12832), .B(n12835), .S(n15631), .Z(n12833) );
  OAI21_X1 U15233 ( .B1(n9292), .B2(n13580), .A(n12833), .ZN(P3_U3390) );
  MUX2_X1 U15234 ( .A(n12835), .B(n12834), .S(n15637), .Z(n12836) );
  OAI21_X1 U15235 ( .B1(n9292), .B2(n13485), .A(n12836), .ZN(P3_U3459) );
  INV_X1 U15236 ( .A(n12839), .ZN(n12842) );
  AOI21_X1 U15237 ( .B1(n14584), .B2(n14622), .A(n12840), .ZN(n12841) );
  INV_X1 U15238 ( .A(n12841), .ZN(P2_U3529) );
  NOR2_X1 U15239 ( .A1(n14473), .A2(n12842), .ZN(n14285) );
  NOR2_X1 U15240 ( .A1(n14502), .A2(n12843), .ZN(n12844) );
  AOI211_X1 U15241 ( .C1(n14622), .C2(n14511), .A(n14285), .B(n12844), .ZN(
        n12845) );
  OAI21_X1 U15242 ( .B1(n12846), .B2(n14492), .A(n12845), .ZN(P2_U3235) );
  NAND2_X1 U15243 ( .A1(n14082), .A2(n7907), .ZN(n12848) );
  XNOR2_X1 U15244 ( .A(n12848), .B(n12847), .ZN(n12849) );
  XNOR2_X1 U15245 ( .A(n14293), .B(n12849), .ZN(n12852) );
  INV_X1 U15246 ( .A(n12852), .ZN(n12850) );
  NAND2_X1 U15247 ( .A1(n12850), .A2(n13714), .ZN(n12862) );
  INV_X1 U15248 ( .A(n12851), .ZN(n12856) );
  INV_X1 U15249 ( .A(n12853), .ZN(n14291) );
  AOI22_X1 U15250 ( .A1(n14291), .A2(n13700), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12854) );
  OAI21_X1 U15251 ( .B1(n12855), .B2(n13726), .A(n12854), .ZN(n12858) );
  NOR2_X1 U15252 ( .A1(n12862), .A2(n12856), .ZN(n12857) );
  AOI211_X1 U15253 ( .C1(n14293), .C2(n13751), .A(n12858), .B(n12857), .ZN(
        n12859) );
  OAI211_X1 U15254 ( .C1(n12862), .C2(n12861), .A(n12860), .B(n12859), .ZN(
        P2_U3192) );
  INV_X1 U15255 ( .A(n10274), .ZN(n15399) );
  OAI222_X1 U15256 ( .A1(P2_U3088), .A2(n7876), .B1(n14685), .B2(n15399), .C1(
        n12863), .C2(n14682), .ZN(P2_U3298) );
  NOR2_X1 U15257 ( .A1(n15027), .A2(n12865), .ZN(n12867) );
  XNOR2_X1 U15258 ( .A(n12867), .B(n12866), .ZN(n15268) );
  NOR2_X1 U15259 ( .A1(n12868), .A2(n15196), .ZN(n12881) );
  INV_X1 U15260 ( .A(n15058), .ZN(n12870) );
  NAND3_X1 U15261 ( .A1(n15031), .A2(n12873), .A3(n12872), .ZN(n12874) );
  AOI21_X1 U15262 ( .B1(n15264), .B2(n6718), .A(n12877), .ZN(n15265) );
  INV_X1 U15263 ( .A(n12878), .ZN(n12879) );
  AOI22_X1 U15264 ( .A1(n15265), .A2(n12879), .B1(n14811), .B2(n15480), .ZN(
        n12880) );
  OAI21_X1 U15265 ( .B1(n15268), .B2(n15478), .A(n12882), .ZN(P1_U3267) );
  INV_X1 U15266 ( .A(n14678), .ZN(n12884) );
  OAI222_X1 U15267 ( .A1(P1_U3086), .A2(n12885), .B1(n15400), .B2(n12884), 
        .C1(n12883), .C2(n15397), .ZN(P1_U3327) );
  INV_X1 U15268 ( .A(n12888), .ZN(n12894) );
  AOI22_X1 U15269 ( .A1(n12889), .A2(n15480), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15484), .ZN(n12890) );
  OAI21_X1 U15270 ( .B1(n14997), .B2(n15196), .A(n12890), .ZN(n12893) );
  NOR2_X1 U15271 ( .A1(n12891), .A2(n15484), .ZN(n12892) );
  OAI21_X1 U15272 ( .B1(n12896), .B2(n15478), .A(n12895), .ZN(P1_U3265) );
  OAI222_X1 U15273 ( .A1(n15400), .A2(n14676), .B1(n9487), .B2(P1_U3086), .C1(
        n12897), .C2(n15397), .ZN(P1_U3325) );
  XNOR2_X1 U15274 ( .A(n12969), .B(n13081), .ZN(n12970) );
  NAND2_X1 U15275 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  XNOR2_X1 U15276 ( .A(n13477), .B(n12972), .ZN(n12904) );
  XNOR2_X1 U15277 ( .A(n12904), .B(n13093), .ZN(n13067) );
  INV_X1 U15278 ( .A(n13067), .ZN(n12903) );
  NAND2_X1 U15279 ( .A1(n12904), .A2(n13093), .ZN(n12905) );
  NAND2_X1 U15280 ( .A1(n13069), .A2(n12905), .ZN(n12999) );
  XNOR2_X1 U15281 ( .A(n13414), .B(n12972), .ZN(n12907) );
  XNOR2_X1 U15282 ( .A(n12907), .B(n13008), .ZN(n12998) );
  NAND2_X1 U15283 ( .A1(n12907), .A2(n13092), .ZN(n12908) );
  NAND2_X1 U15284 ( .A1(n12997), .A2(n12908), .ZN(n13007) );
  XNOR2_X1 U15285 ( .A(n13559), .B(n12972), .ZN(n12909) );
  XNOR2_X1 U15286 ( .A(n12909), .B(n13049), .ZN(n13006) );
  NAND2_X1 U15287 ( .A1(n13007), .A2(n13006), .ZN(n13005) );
  NAND2_X1 U15288 ( .A1(n12909), .A2(n13091), .ZN(n12910) );
  XNOR2_X1 U15289 ( .A(n13553), .B(n12972), .ZN(n12911) );
  XNOR2_X1 U15290 ( .A(n12911), .B(n13009), .ZN(n13046) );
  NAND2_X1 U15291 ( .A1(n12911), .A2(n13090), .ZN(n12912) );
  XNOR2_X1 U15292 ( .A(n13546), .B(n12972), .ZN(n12913) );
  XNOR2_X1 U15293 ( .A(n12913), .B(n13089), .ZN(n12962) );
  INV_X1 U15294 ( .A(n12913), .ZN(n12914) );
  NAND2_X1 U15295 ( .A1(n12914), .A2(n13089), .ZN(n12915) );
  XNOR2_X1 U15296 ( .A(n13334), .B(n12972), .ZN(n12916) );
  XNOR2_X1 U15297 ( .A(n12916), .B(n13088), .ZN(n13029) );
  INV_X1 U15298 ( .A(n12916), .ZN(n12917) );
  XNOR2_X1 U15299 ( .A(n13538), .B(n12972), .ZN(n12918) );
  XNOR2_X1 U15300 ( .A(n12918), .B(n13031), .ZN(n12984) );
  XNOR2_X1 U15301 ( .A(n13026), .B(n12972), .ZN(n13022) );
  XNOR2_X1 U15302 ( .A(n13452), .B(n12972), .ZN(n13017) );
  AOI22_X1 U15303 ( .A1(n13022), .A2(n13084), .B1(n13085), .B2(n13017), .ZN(
        n12922) );
  OAI21_X1 U15304 ( .B1(n12941), .B2(n12937), .A(n12922), .ZN(n12925) );
  INV_X1 U15305 ( .A(n13022), .ZN(n12921) );
  OAI21_X1 U15306 ( .B1(n13017), .B2(n13085), .A(n13084), .ZN(n12920) );
  NOR3_X1 U15307 ( .A1(n13017), .A2(n13084), .A3(n13085), .ZN(n12919) );
  AOI21_X1 U15308 ( .B1(n12921), .B2(n12920), .A(n12919), .ZN(n12924) );
  NAND3_X1 U15309 ( .A1(n12922), .A2(n12941), .A3(n12937), .ZN(n12923) );
  XNOR2_X1 U15310 ( .A(n12926), .B(n13083), .ZN(n12991) );
  AOI22_X2 U15311 ( .A1(n12990), .A2(n12991), .B1(n12927), .B2(n12926), .ZN(
        n13057) );
  XNOR2_X1 U15312 ( .A(n12929), .B(n12928), .ZN(n13058) );
  INV_X1 U15313 ( .A(n12929), .ZN(n12930) );
  XOR2_X1 U15314 ( .A(n12970), .B(n12971), .Z(n12936) );
  AOI22_X1 U15315 ( .A1(n13258), .A2(n13074), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12931) );
  OAI21_X1 U15316 ( .B1(n12932), .B2(n13071), .A(n12931), .ZN(n12933) );
  AOI21_X1 U15317 ( .B1(n12934), .B2(n13063), .A(n12933), .ZN(n12935) );
  OAI21_X1 U15318 ( .B1(n12936), .B2(n13066), .A(n12935), .ZN(P3_U3154) );
  INV_X1 U15319 ( .A(n12937), .ZN(n12938) );
  NOR2_X1 U15320 ( .A1(n12939), .A2(n12938), .ZN(n12940) );
  XNOR2_X1 U15321 ( .A(n13021), .B(n12942), .ZN(n12947) );
  AND2_X1 U15322 ( .A1(n13086), .A2(n13059), .ZN(n12943) );
  AOI21_X1 U15323 ( .B1(n13084), .B2(n13060), .A(n12943), .ZN(n13307) );
  AOI22_X1 U15324 ( .A1(n13308), .A2(n13074), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12944) );
  OAI21_X1 U15325 ( .B1(n13307), .B2(n13071), .A(n12944), .ZN(n12945) );
  AOI21_X1 U15326 ( .B1(n13452), .B2(n13063), .A(n12945), .ZN(n12946) );
  OAI21_X1 U15327 ( .B1(n12947), .B2(n13066), .A(n12946), .ZN(P3_U3156) );
  INV_X1 U15328 ( .A(n12948), .ZN(n12949) );
  NOR2_X1 U15329 ( .A1(n12950), .A2(n12949), .ZN(n12953) );
  OAI211_X1 U15330 ( .C1(n12953), .C2(n12952), .A(n13044), .B(n12951), .ZN(
        n12960) );
  AOI22_X1 U15331 ( .A1(n12954), .A2(n13034), .B1(P3_REG3_REG_10__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12959) );
  OR2_X1 U15332 ( .A1(n12955), .A2(n13078), .ZN(n12958) );
  NAND2_X1 U15333 ( .A1(n13074), .A2(n12956), .ZN(n12957) );
  NAND4_X1 U15334 ( .A1(n12960), .A2(n12959), .A3(n12958), .A4(n12957), .ZN(
        P3_U3157) );
  OAI211_X1 U15335 ( .C1(n12963), .C2(n12962), .A(n12961), .B(n13044), .ZN(
        n12968) );
  NOR2_X1 U15336 ( .A1(n13009), .A2(n13048), .ZN(n12964) );
  AOI21_X1 U15337 ( .B1(n13088), .B2(n13060), .A(n12964), .ZN(n13368) );
  OAI21_X1 U15338 ( .B1(n13368), .B2(n13071), .A(n12965), .ZN(n12966) );
  AOI21_X1 U15339 ( .B1(n13361), .B2(n13074), .A(n12966), .ZN(n12967) );
  OAI211_X1 U15340 ( .C1(n13078), .C2(n13546), .A(n12968), .B(n12967), .ZN(
        P3_U3159) );
  AOI22_X1 U15341 ( .A1(n12971), .A2(n12970), .B1(n12976), .B2(n12969), .ZN(
        n12974) );
  XNOR2_X1 U15342 ( .A(n13250), .B(n12972), .ZN(n12973) );
  XNOR2_X1 U15343 ( .A(n12974), .B(n12973), .ZN(n12982) );
  INV_X1 U15344 ( .A(n13060), .ZN(n13050) );
  OR2_X1 U15345 ( .A1(n12975), .A2(n13050), .ZN(n12978) );
  OR2_X1 U15346 ( .A1(n12976), .A2(n13048), .ZN(n12977) );
  AND2_X1 U15347 ( .A1(n12978), .A2(n12977), .ZN(n13247) );
  AOI22_X1 U15348 ( .A1(n13252), .A2(n13074), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12979) );
  OAI21_X1 U15349 ( .B1(n13247), .B2(n13071), .A(n12979), .ZN(n12980) );
  AOI21_X1 U15350 ( .B1(n13253), .B2(n13063), .A(n12980), .ZN(n12981) );
  OAI21_X1 U15351 ( .B1(n12982), .B2(n13066), .A(n12981), .ZN(P3_U3160) );
  OAI211_X1 U15352 ( .C1(n12985), .C2(n12984), .A(n12983), .B(n13044), .ZN(
        n12989) );
  AOI22_X1 U15353 ( .A1(n13086), .A2(n13060), .B1(n13059), .B2(n13088), .ZN(
        n13340) );
  AOI22_X1 U15354 ( .A1(n13329), .A2(n13074), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12986) );
  OAI21_X1 U15355 ( .B1(n13340), .B2(n13071), .A(n12986), .ZN(n12987) );
  AOI21_X1 U15356 ( .B1(n13538), .B2(n13063), .A(n12987), .ZN(n12988) );
  NAND2_X1 U15357 ( .A1(n12989), .A2(n12988), .ZN(P3_U3163) );
  XOR2_X1 U15358 ( .A(n12991), .B(n12990), .Z(n12996) );
  AND2_X1 U15359 ( .A1(n13084), .A2(n13059), .ZN(n12992) );
  AOI21_X1 U15360 ( .B1(n13082), .B2(n13060), .A(n12992), .ZN(n13279) );
  AOI22_X1 U15361 ( .A1(n13283), .A2(n13074), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12993) );
  OAI21_X1 U15362 ( .B1(n13279), .B2(n13071), .A(n12993), .ZN(n12994) );
  AOI21_X1 U15363 ( .B1(n13520), .B2(n13063), .A(n12994), .ZN(n12995) );
  OAI21_X1 U15364 ( .B1(n12996), .B2(n13066), .A(n12995), .ZN(P3_U3165) );
  INV_X1 U15365 ( .A(n13414), .ZN(n13564) );
  OAI211_X1 U15366 ( .C1(n12999), .C2(n12998), .A(n12997), .B(n13044), .ZN(
        n13004) );
  OR2_X1 U15367 ( .A1(n13049), .A2(n13050), .ZN(n13001) );
  NAND2_X1 U15368 ( .A1(n13093), .A2(n13059), .ZN(n13000) );
  AND2_X1 U15369 ( .A1(n13001), .A2(n13000), .ZN(n13410) );
  NAND2_X1 U15370 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13180)
         );
  OAI21_X1 U15371 ( .B1(n13410), .B2(n13071), .A(n13180), .ZN(n13002) );
  AOI21_X1 U15372 ( .B1(n13413), .B2(n13074), .A(n13002), .ZN(n13003) );
  OAI211_X1 U15373 ( .C1(n13564), .C2(n13078), .A(n13004), .B(n13003), .ZN(
        P3_U3166) );
  INV_X1 U15374 ( .A(n13559), .ZN(n13015) );
  OAI211_X1 U15375 ( .C1(n13007), .C2(n13006), .A(n13005), .B(n13044), .ZN(
        n13014) );
  OAI22_X1 U15376 ( .A1(n13009), .A2(n13050), .B1(n13008), .B2(n13048), .ZN(
        n13399) );
  NOR2_X1 U15377 ( .A1(n15748), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13192) );
  INV_X1 U15378 ( .A(n13402), .ZN(n13010) );
  NOR2_X1 U15379 ( .A1(n13011), .A2(n13010), .ZN(n13012) );
  AOI211_X1 U15380 ( .C1(n13034), .C2(n13399), .A(n13192), .B(n13012), .ZN(
        n13013) );
  OAI211_X1 U15381 ( .C1(n13015), .C2(n13078), .A(n13014), .B(n13013), .ZN(
        P3_U3168) );
  INV_X1 U15382 ( .A(n13017), .ZN(n13018) );
  XNOR2_X1 U15383 ( .A(n13022), .B(n13084), .ZN(n13023) );
  AOI22_X1 U15384 ( .A1(n13083), .A2(n13060), .B1(n13059), .B2(n13085), .ZN(
        n13291) );
  AOI22_X1 U15385 ( .A1(n13294), .A2(n13074), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13024) );
  OAI21_X1 U15386 ( .B1(n13291), .B2(n13071), .A(n13024), .ZN(n13025) );
  AOI21_X1 U15387 ( .B1(n13026), .B2(n13063), .A(n13025), .ZN(n13027) );
  OAI211_X1 U15388 ( .C1(n13030), .C2(n13029), .A(n13028), .B(n13044), .ZN(
        n13038) );
  OR2_X1 U15389 ( .A1(n13031), .A2(n13050), .ZN(n13033) );
  NAND2_X1 U15390 ( .A1(n13089), .A2(n13059), .ZN(n13032) );
  NAND2_X1 U15391 ( .A1(n13033), .A2(n13032), .ZN(n13352) );
  AOI22_X1 U15392 ( .A1(n13352), .A2(n13034), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13037) );
  OR2_X1 U15393 ( .A1(n13334), .A2(n13078), .ZN(n13036) );
  NAND2_X1 U15394 ( .A1(n13348), .A2(n13074), .ZN(n13035) );
  NAND4_X1 U15395 ( .A1(n13038), .A2(n13037), .A3(n13036), .A4(n13035), .ZN(
        P3_U3173) );
  XNOR2_X1 U15396 ( .A(n13039), .B(n13086), .ZN(n13043) );
  AOI22_X1 U15397 ( .A1(n13085), .A2(n13060), .B1(n13059), .B2(n13087), .ZN(
        n13318) );
  AOI22_X1 U15398 ( .A1(n13322), .A2(n13074), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13040) );
  OAI21_X1 U15399 ( .B1(n13318), .B2(n13071), .A(n13040), .ZN(n13041) );
  AOI21_X1 U15400 ( .B1(n13532), .B2(n13063), .A(n13041), .ZN(n13042) );
  OAI21_X1 U15401 ( .B1(n13043), .B2(n13066), .A(n13042), .ZN(P3_U3175) );
  INV_X1 U15402 ( .A(n13553), .ZN(n13056) );
  OAI211_X1 U15403 ( .C1(n13047), .C2(n13046), .A(n13045), .B(n13044), .ZN(
        n13055) );
  OAI22_X1 U15404 ( .A1(n13051), .A2(n13050), .B1(n13049), .B2(n13048), .ZN(
        n13384) );
  INV_X1 U15405 ( .A(n13384), .ZN(n13052) );
  NAND2_X1 U15406 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13213)
         );
  OAI21_X1 U15407 ( .B1(n13052), .B2(n13071), .A(n13213), .ZN(n13053) );
  AOI21_X1 U15408 ( .B1(n13387), .B2(n13074), .A(n13053), .ZN(n13054) );
  OAI211_X1 U15409 ( .C1(n13056), .C2(n13078), .A(n13055), .B(n13054), .ZN(
        P3_U3178) );
  XOR2_X1 U15410 ( .A(n13058), .B(n13057), .Z(n13065) );
  AOI22_X1 U15411 ( .A1(n13081), .A2(n13060), .B1(n13059), .B2(n13083), .ZN(
        n13268) );
  AOI22_X1 U15412 ( .A1(n13271), .A2(n13074), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13061) );
  OAI21_X1 U15413 ( .B1(n13268), .B2(n13071), .A(n13061), .ZN(n13062) );
  AOI21_X1 U15414 ( .B1(n13270), .B2(n13063), .A(n13062), .ZN(n13064) );
  OAI21_X1 U15415 ( .B1(n13065), .B2(n13066), .A(n13064), .ZN(P3_U3180) );
  INV_X1 U15416 ( .A(n13477), .ZN(n13079) );
  AOI21_X1 U15417 ( .B1(n13068), .B2(n13067), .A(n13066), .ZN(n13070) );
  NAND2_X1 U15418 ( .A1(n13070), .A2(n13069), .ZN(n13077) );
  NAND2_X1 U15419 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13159)
         );
  OAI21_X1 U15420 ( .B1(n13072), .B2(n13071), .A(n13159), .ZN(n13073) );
  AOI21_X1 U15421 ( .B1(n13075), .B2(n13074), .A(n13073), .ZN(n13076) );
  OAI211_X1 U15422 ( .C1(n13079), .C2(n13078), .A(n13077), .B(n13076), .ZN(
        P3_U3181) );
  MUX2_X1 U15423 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13080), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15424 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13081), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15425 ( .A(n13082), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13107), .Z(
        P3_U3517) );
  MUX2_X1 U15426 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13083), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15427 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13084), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15428 ( .A(n13085), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13107), .Z(
        P3_U3514) );
  MUX2_X1 U15429 ( .A(n13086), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13107), .Z(
        P3_U3513) );
  MUX2_X1 U15430 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13087), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15431 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13088), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15432 ( .A(n13089), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13107), .Z(
        P3_U3510) );
  MUX2_X1 U15433 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13090), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15434 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13091), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15435 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13092), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15436 ( .A(n13093), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13107), .Z(
        P3_U3506) );
  MUX2_X1 U15437 ( .A(n13094), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13107), .Z(
        P3_U3505) );
  MUX2_X1 U15438 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13095), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15439 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13096), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15440 ( .A(n13097), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13107), .Z(
        P3_U3502) );
  MUX2_X1 U15441 ( .A(n13098), .B(P3_DATAO_REG_10__SCAN_IN), .S(n13107), .Z(
        P3_U3501) );
  MUX2_X1 U15442 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13099), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15443 ( .A(n13100), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13107), .Z(
        P3_U3499) );
  MUX2_X1 U15444 ( .A(n13101), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13107), .Z(
        P3_U3498) );
  MUX2_X1 U15445 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13102), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15446 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13103), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15447 ( .A(n13104), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13107), .Z(
        P3_U3495) );
  MUX2_X1 U15448 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13105), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15449 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13106), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15450 ( .A(n13108), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13107), .Z(
        P3_U3491) );
  INV_X1 U15451 ( .A(n13109), .ZN(n13114) );
  NOR3_X1 U15452 ( .A1(n13112), .A2(n13111), .A3(n13110), .ZN(n13113) );
  OAI21_X1 U15453 ( .B1(n13114), .B2(n13113), .A(n13217), .ZN(n13130) );
  INV_X1 U15454 ( .A(n13115), .ZN(n13117) );
  NOR3_X1 U15455 ( .A1(n6601), .A2(n13117), .A3(n13116), .ZN(n13120) );
  INV_X1 U15456 ( .A(n13118), .ZN(n13119) );
  OAI21_X1 U15457 ( .B1(n13120), .B2(n13119), .A(n13222), .ZN(n13129) );
  OAI21_X1 U15458 ( .B1(n13215), .B2(n13122), .A(n13121), .ZN(n13123) );
  AOI21_X1 U15459 ( .B1(n13124), .B2(n13212), .A(n13123), .ZN(n13128) );
  OAI211_X1 U15460 ( .C1(n13126), .C2(n13125), .A(n13139), .B(n13140), .ZN(
        n13127) );
  NAND4_X1 U15461 ( .A1(n13130), .A2(n13129), .A3(n13128), .A4(n13127), .ZN(
        P3_U3194) );
  INV_X1 U15462 ( .A(n13131), .ZN(n13132) );
  AOI21_X1 U15463 ( .B1(n13134), .B2(n13133), .A(n13132), .ZN(n13150) );
  OAI21_X1 U15464 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n13135), .A(n10688), 
        .ZN(n13148) );
  INV_X1 U15465 ( .A(n13136), .ZN(n13142) );
  AOI21_X1 U15466 ( .B1(n13139), .B2(n13138), .A(n13137), .ZN(n13141) );
  OAI21_X1 U15467 ( .B1(n13142), .B2(n13141), .A(n13140), .ZN(n13145) );
  AOI21_X1 U15468 ( .B1(n15575), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n13143), 
        .ZN(n13144) );
  OAI211_X1 U15469 ( .C1(n13195), .C2(n13146), .A(n13145), .B(n13144), .ZN(
        n13147) );
  AOI21_X1 U15470 ( .B1(n13148), .B2(n13222), .A(n13147), .ZN(n13149) );
  OAI21_X1 U15471 ( .B1(n13150), .B2(n13165), .A(n13149), .ZN(P3_U3195) );
  INV_X1 U15472 ( .A(n13170), .ZN(n13151) );
  AOI21_X1 U15473 ( .B1(n13478), .B2(n13152), .A(n13151), .ZN(n13166) );
  OAI21_X1 U15474 ( .B1(n6507), .B2(P3_REG2_REG_15__SCAN_IN), .A(n13153), .ZN(
        n13163) );
  AOI21_X1 U15475 ( .B1(n13156), .B2(n13155), .A(n13154), .ZN(n13157) );
  NOR2_X1 U15476 ( .A1(n13157), .A2(n13226), .ZN(n13162) );
  NAND2_X1 U15477 ( .A1(n15575), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n13158) );
  OAI211_X1 U15478 ( .C1(n13195), .C2(n13160), .A(n13159), .B(n13158), .ZN(
        n13161) );
  AOI211_X1 U15479 ( .C1(n13163), .C2(n13222), .A(n13162), .B(n13161), .ZN(
        n13164) );
  OAI21_X1 U15480 ( .B1(n13166), .B2(n13165), .A(n13164), .ZN(P3_U3197) );
  NOR2_X1 U15481 ( .A1(n13167), .A2(n6625), .ZN(n13168) );
  XNOR2_X1 U15482 ( .A(n6567), .B(n13168), .ZN(n13185) );
  NAND3_X1 U15483 ( .A1(n13170), .A2(n6632), .A3(n13169), .ZN(n13171) );
  NAND2_X1 U15484 ( .A1(n13172), .A2(n13171), .ZN(n13179) );
  INV_X1 U15485 ( .A(n13173), .ZN(n13175) );
  NAND3_X1 U15486 ( .A1(n13153), .A2(n13175), .A3(n13174), .ZN(n13176) );
  AOI21_X1 U15487 ( .B1(n13177), .B2(n13176), .A(n13200), .ZN(n13178) );
  AOI21_X1 U15488 ( .B1(n13217), .B2(n13179), .A(n13178), .ZN(n13184) );
  INV_X1 U15489 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15438) );
  OAI21_X1 U15490 ( .B1(n13215), .B2(n15438), .A(n13180), .ZN(n13181) );
  AOI21_X1 U15491 ( .B1(n13182), .B2(n13212), .A(n13181), .ZN(n13183) );
  OAI211_X1 U15492 ( .C1(n13226), .C2(n13185), .A(n13184), .B(n13183), .ZN(
        P3_U3198) );
  INV_X1 U15493 ( .A(n13221), .ZN(n13186) );
  AOI21_X1 U15494 ( .B1(n13401), .B2(n13187), .A(n13186), .ZN(n13201) );
  OAI21_X1 U15495 ( .B1(n13188), .B2(P3_REG1_REG_17__SCAN_IN), .A(n13208), 
        .ZN(n13198) );
  AOI211_X1 U15496 ( .C1(n13191), .C2(n13190), .A(n13226), .B(n13189), .ZN(
        n13197) );
  AOI21_X1 U15497 ( .B1(n15575), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13192), 
        .ZN(n13193) );
  OAI21_X1 U15498 ( .B1(n13195), .B2(n13194), .A(n13193), .ZN(n13196) );
  AOI211_X1 U15499 ( .C1(n13198), .C2(n13217), .A(n13197), .B(n13196), .ZN(
        n13199) );
  OAI21_X1 U15500 ( .B1(n13201), .B2(n13200), .A(n13199), .ZN(P3_U3199) );
  INV_X1 U15501 ( .A(n13205), .ZN(n13210) );
  NAND3_X1 U15502 ( .A1(n13208), .A2(n13207), .A3(n13206), .ZN(n13209) );
  NAND2_X1 U15503 ( .A1(n13210), .A2(n13209), .ZN(n13218) );
  INV_X1 U15504 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15773) );
  NAND2_X1 U15505 ( .A1(n13212), .A2(n13211), .ZN(n13214) );
  OAI211_X1 U15506 ( .C1(n13215), .C2(n15773), .A(n13214), .B(n13213), .ZN(
        n13216) );
  AND3_X1 U15507 ( .A1(n13221), .A2(n13220), .A3(n13219), .ZN(n13223) );
  OAI21_X1 U15508 ( .B1(n13224), .B2(n13223), .A(n13222), .ZN(n13225) );
  NAND2_X1 U15509 ( .A1(n13228), .A2(n13427), .ZN(n13232) );
  NOR2_X1 U15510 ( .A1(n13230), .A2(n13229), .ZN(n13503) );
  NOR2_X1 U15511 ( .A1(n13231), .A2(n15578), .ZN(n13238) );
  AOI21_X1 U15512 ( .B1(n13503), .B2(n15597), .A(n13238), .ZN(n13235) );
  OAI211_X1 U15513 ( .C1(n15597), .C2(n13233), .A(n13232), .B(n13235), .ZN(
        P3_U3202) );
  NAND2_X1 U15514 ( .A1(n13234), .A2(n13427), .ZN(n13236) );
  OAI211_X1 U15515 ( .C1(n15597), .C2(n15744), .A(n13236), .B(n13235), .ZN(
        P3_U3203) );
  INV_X1 U15516 ( .A(n13237), .ZN(n13244) );
  AOI21_X1 U15517 ( .B1(n15587), .B2(P3_REG2_REG_29__SCAN_IN), .A(n13238), 
        .ZN(n13239) );
  OAI21_X1 U15518 ( .B1(n13240), .B2(n13363), .A(n13239), .ZN(n13241) );
  AOI21_X1 U15519 ( .B1(n13242), .B2(n15597), .A(n13241), .ZN(n13243) );
  OAI21_X1 U15520 ( .B1(n13244), .B2(n13431), .A(n13243), .ZN(P3_U3204) );
  OAI211_X1 U15521 ( .C1(n13246), .C2(n13250), .A(n13245), .B(n13493), .ZN(
        n13248) );
  NAND2_X1 U15522 ( .A1(n13248), .A2(n13247), .ZN(n13509) );
  NAND2_X1 U15523 ( .A1(n9442), .A2(n13249), .ZN(n13251) );
  XNOR2_X1 U15524 ( .A(n13251), .B(n13250), .ZN(n13511) );
  AOI22_X1 U15525 ( .A1(n13253), .A2(n13427), .B1(n15592), .B2(n13252), .ZN(
        n13254) );
  OAI21_X1 U15526 ( .B1(n13511), .B2(n13431), .A(n13254), .ZN(n13255) );
  INV_X1 U15527 ( .A(n13257), .ZN(n13264) );
  AOI22_X1 U15528 ( .A1(n13258), .A2(n15592), .B1(n15587), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13259) );
  OAI21_X1 U15529 ( .B1(n13260), .B2(n13363), .A(n13259), .ZN(n13261) );
  AOI21_X1 U15530 ( .B1(n13262), .B2(n15594), .A(n13261), .ZN(n13263) );
  OAI21_X1 U15531 ( .B1(n13264), .B2(n15587), .A(n13263), .ZN(P3_U3206) );
  XNOR2_X1 U15532 ( .A(n13265), .B(n13266), .ZN(n13440) );
  INV_X1 U15533 ( .A(n13440), .ZN(n13275) );
  XOR2_X1 U15534 ( .A(n13267), .B(n13266), .Z(n13269) );
  OAI21_X1 U15535 ( .B1(n13269), .B2(n13397), .A(n13268), .ZN(n13439) );
  INV_X1 U15536 ( .A(n13270), .ZN(n13517) );
  AOI22_X1 U15537 ( .A1(n13271), .A2(n15592), .B1(n15587), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13272) );
  OAI21_X1 U15538 ( .B1(n13517), .B2(n13363), .A(n13272), .ZN(n13273) );
  AOI21_X1 U15539 ( .B1(n13439), .B2(n15597), .A(n13273), .ZN(n13274) );
  OAI21_X1 U15540 ( .B1(n13431), .B2(n13275), .A(n13274), .ZN(P3_U3207) );
  OAI211_X1 U15541 ( .C1(n13278), .C2(n13277), .A(n13276), .B(n13493), .ZN(
        n13280) );
  INV_X1 U15542 ( .A(n13520), .ZN(n13285) );
  AOI22_X1 U15543 ( .A1(n13283), .A2(n15592), .B1(n15587), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13284) );
  OAI21_X1 U15544 ( .B1(n13285), .B2(n13363), .A(n13284), .ZN(n13286) );
  AOI21_X1 U15545 ( .B1(n13443), .B2(n15594), .A(n13286), .ZN(n13287) );
  OAI21_X1 U15546 ( .B1(n13445), .B2(n15587), .A(n13287), .ZN(P3_U3208) );
  XNOR2_X1 U15547 ( .A(n13288), .B(n13289), .ZN(n13293) );
  XNOR2_X1 U15548 ( .A(n13290), .B(n13289), .ZN(n13449) );
  NAND2_X1 U15549 ( .A1(n13449), .A2(n15627), .ZN(n13292) );
  OAI211_X1 U15550 ( .C1(n13397), .C2(n13293), .A(n13292), .B(n13291), .ZN(
        n13448) );
  INV_X1 U15551 ( .A(n13448), .ZN(n13298) );
  AOI22_X1 U15552 ( .A1(n13294), .A2(n15592), .B1(n15587), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13295) );
  OAI21_X1 U15553 ( .B1(n13525), .B2(n13363), .A(n13295), .ZN(n13296) );
  AOI21_X1 U15554 ( .B1(n13449), .B2(n15594), .A(n13296), .ZN(n13297) );
  OAI21_X1 U15555 ( .B1(n13298), .B2(n15587), .A(n13297), .ZN(P3_U3209) );
  NAND2_X1 U15556 ( .A1(n13300), .A2(n13299), .ZN(n13302) );
  NAND2_X1 U15557 ( .A1(n13302), .A2(n13304), .ZN(n13301) );
  OAI21_X1 U15558 ( .B1(n13302), .B2(n13304), .A(n13301), .ZN(n13453) );
  XNOR2_X1 U15559 ( .A(n13303), .B(n13304), .ZN(n13305) );
  NAND2_X1 U15560 ( .A1(n13305), .A2(n13493), .ZN(n13306) );
  OAI211_X1 U15561 ( .C1(n13453), .C2(n15609), .A(n13307), .B(n13306), .ZN(
        n13454) );
  NAND2_X1 U15562 ( .A1(n13454), .A2(n15597), .ZN(n13313) );
  INV_X1 U15563 ( .A(n13308), .ZN(n13310) );
  OAI22_X1 U15564 ( .A1(n13310), .A2(n15578), .B1(n15597), .B2(n13309), .ZN(
        n13311) );
  AOI21_X1 U15565 ( .B1(n13452), .B2(n13427), .A(n13311), .ZN(n13312) );
  OAI211_X1 U15566 ( .C1(n13453), .C2(n13314), .A(n13313), .B(n13312), .ZN(
        P3_U3210) );
  XOR2_X1 U15567 ( .A(n13315), .B(n13316), .Z(n13535) );
  XNOR2_X1 U15568 ( .A(n13317), .B(n13316), .ZN(n13320) );
  INV_X1 U15569 ( .A(n13318), .ZN(n13319) );
  AOI21_X1 U15570 ( .B1(n13320), .B2(n13493), .A(n13319), .ZN(n13530) );
  MUX2_X1 U15571 ( .A(n13321), .B(n13530), .S(n15597), .Z(n13324) );
  AOI22_X1 U15572 ( .A1(n13532), .A2(n13427), .B1(n15592), .B2(n13322), .ZN(
        n13323) );
  OAI211_X1 U15573 ( .C1(n13535), .C2(n13431), .A(n13324), .B(n13323), .ZN(
        P3_U3211) );
  NAND2_X1 U15574 ( .A1(n13376), .A2(n13325), .ZN(n13360) );
  NOR2_X1 U15575 ( .A1(n13359), .A2(n13326), .ZN(n13347) );
  NAND2_X1 U15576 ( .A1(n13347), .A2(n7238), .ZN(n13346) );
  NAND2_X1 U15577 ( .A1(n13346), .A2(n13327), .ZN(n13328) );
  XNOR2_X1 U15578 ( .A(n13328), .B(n13338), .ZN(n13540) );
  AOI22_X1 U15579 ( .A1(n13538), .A2(n13427), .B1(n15592), .B2(n13329), .ZN(
        n13345) );
  INV_X1 U15580 ( .A(n13331), .ZN(n13332) );
  NAND2_X1 U15581 ( .A1(n13330), .A2(n13332), .ZN(n13365) );
  NAND2_X1 U15582 ( .A1(n13365), .A2(n13333), .ZN(n13351) );
  NAND2_X1 U15583 ( .A1(n13351), .A2(n13350), .ZN(n13349) );
  OAI21_X1 U15584 ( .B1(n13335), .B2(n13334), .A(n13349), .ZN(n13339) );
  INV_X1 U15585 ( .A(n13336), .ZN(n13337) );
  AOI21_X1 U15586 ( .B1(n13339), .B2(n13338), .A(n13337), .ZN(n13341) );
  OAI21_X1 U15587 ( .B1(n13341), .B2(n13397), .A(n13340), .ZN(n13536) );
  INV_X1 U15588 ( .A(n13536), .ZN(n13342) );
  MUX2_X1 U15589 ( .A(n13343), .B(n13342), .S(n15597), .Z(n13344) );
  OAI211_X1 U15590 ( .C1(n13540), .C2(n13431), .A(n13345), .B(n13344), .ZN(
        P3_U3212) );
  OAI21_X1 U15591 ( .B1(n13347), .B2(n7238), .A(n13346), .ZN(n13545) );
  AOI22_X1 U15592 ( .A1(n13543), .A2(n13427), .B1(n15592), .B2(n13348), .ZN(
        n13358) );
  OAI211_X1 U15593 ( .C1(n13351), .C2(n13350), .A(n13349), .B(n13493), .ZN(
        n13354) );
  INV_X1 U15594 ( .A(n13352), .ZN(n13353) );
  NAND2_X1 U15595 ( .A1(n13354), .A2(n13353), .ZN(n13541) );
  INV_X1 U15596 ( .A(n13541), .ZN(n13355) );
  MUX2_X1 U15597 ( .A(n13356), .B(n13355), .S(n15597), .Z(n13357) );
  OAI211_X1 U15598 ( .C1(n13545), .C2(n13431), .A(n13358), .B(n13357), .ZN(
        P3_U3213) );
  AOI21_X1 U15599 ( .B1(n13366), .B2(n13360), .A(n13359), .ZN(n13547) );
  INV_X1 U15600 ( .A(n13361), .ZN(n13362) );
  OAI22_X1 U15601 ( .A1(n13546), .A2(n13363), .B1(n13362), .B2(n15578), .ZN(
        n13364) );
  INV_X1 U15602 ( .A(n13364), .ZN(n13374) );
  NAND2_X1 U15603 ( .A1(n13365), .A2(n13493), .ZN(n13370) );
  AOI21_X1 U15604 ( .B1(n13330), .B2(n13367), .A(n13366), .ZN(n13369) );
  OAI21_X1 U15605 ( .B1(n13370), .B2(n13369), .A(n13368), .ZN(n13548) );
  INV_X1 U15606 ( .A(n13548), .ZN(n13371) );
  MUX2_X1 U15607 ( .A(n13372), .B(n13371), .S(n15597), .Z(n13373) );
  OAI211_X1 U15608 ( .C1(n13547), .C2(n13431), .A(n13374), .B(n13373), .ZN(
        P3_U3214) );
  INV_X1 U15609 ( .A(n13382), .ZN(n13377) );
  OAI21_X1 U15610 ( .B1(n7713), .B2(n13377), .A(n13376), .ZN(n13556) );
  NAND2_X1 U15611 ( .A1(n13378), .A2(n13409), .ZN(n13408) );
  AOI21_X1 U15612 ( .B1(n13408), .B2(n13393), .A(n13379), .ZN(n13396) );
  INV_X1 U15613 ( .A(n13380), .ZN(n13381) );
  NOR2_X1 U15614 ( .A1(n13396), .A2(n13381), .ZN(n13383) );
  OAI21_X1 U15615 ( .B1(n13383), .B2(n13382), .A(n13330), .ZN(n13385) );
  AOI21_X1 U15616 ( .B1(n13385), .B2(n13493), .A(n13384), .ZN(n13551) );
  MUX2_X1 U15617 ( .A(n13386), .B(n13551), .S(n15597), .Z(n13389) );
  AOI22_X1 U15618 ( .A1(n13553), .A2(n13427), .B1(n15592), .B2(n13387), .ZN(
        n13388) );
  OAI211_X1 U15619 ( .C1(n13556), .C2(n13431), .A(n13389), .B(n13388), .ZN(
        P3_U3215) );
  NAND2_X1 U15620 ( .A1(n13390), .A2(n13391), .ZN(n13392) );
  XNOR2_X1 U15621 ( .A(n13392), .B(n13395), .ZN(n13562) );
  INV_X1 U15622 ( .A(n13393), .ZN(n13394) );
  NOR2_X1 U15623 ( .A1(n13395), .A2(n13394), .ZN(n13398) );
  AOI211_X1 U15624 ( .C1(n13398), .C2(n13408), .A(n13397), .B(n13396), .ZN(
        n13400) );
  NOR2_X1 U15625 ( .A1(n13400), .A2(n13399), .ZN(n13557) );
  MUX2_X1 U15626 ( .A(n13401), .B(n13557), .S(n15597), .Z(n13404) );
  AOI22_X1 U15627 ( .A1(n13559), .A2(n13427), .B1(n15592), .B2(n13402), .ZN(
        n13403) );
  OAI211_X1 U15628 ( .C1(n13562), .C2(n13431), .A(n13404), .B(n13403), .ZN(
        P3_U3216) );
  OAI21_X1 U15629 ( .B1(n13406), .B2(n13405), .A(n13390), .ZN(n13407) );
  INV_X1 U15630 ( .A(n13407), .ZN(n13565) );
  OAI211_X1 U15631 ( .C1(n13378), .C2(n13409), .A(n13408), .B(n13493), .ZN(
        n13411) );
  NAND2_X1 U15632 ( .A1(n13411), .A2(n13410), .ZN(n13563) );
  MUX2_X1 U15633 ( .A(n13563), .B(P3_REG2_REG_16__SCAN_IN), .S(n15587), .Z(
        n13412) );
  INV_X1 U15634 ( .A(n13412), .ZN(n13416) );
  AOI22_X1 U15635 ( .A1(n13414), .A2(n13427), .B1(n15592), .B2(n13413), .ZN(
        n13415) );
  OAI211_X1 U15636 ( .C1(n13565), .C2(n13431), .A(n13416), .B(n13415), .ZN(
        P3_U3217) );
  XNOR2_X1 U15637 ( .A(n13418), .B(n13417), .ZN(n13576) );
  INV_X1 U15638 ( .A(n13576), .ZN(n13432) );
  NAND2_X1 U15639 ( .A1(n13420), .A2(n13419), .ZN(n13422) );
  XNOR2_X1 U15640 ( .A(n13422), .B(n13421), .ZN(n13424) );
  AOI21_X1 U15641 ( .B1(n13424), .B2(n13493), .A(n13423), .ZN(n13573) );
  MUX2_X1 U15642 ( .A(n13425), .B(n13573), .S(n15597), .Z(n13430) );
  INV_X1 U15643 ( .A(n13579), .ZN(n13428) );
  AOI22_X1 U15644 ( .A1(n13428), .A2(n13427), .B1(n15592), .B2(n13426), .ZN(
        n13429) );
  OAI211_X1 U15645 ( .C1(n13432), .C2(n13431), .A(n13430), .B(n13429), .ZN(
        P3_U3219) );
  NAND2_X1 U15646 ( .A1(n13228), .A2(n13471), .ZN(n13433) );
  NAND2_X1 U15647 ( .A1(n13503), .A2(n15639), .ZN(n13436) );
  OAI211_X1 U15648 ( .C1(n15639), .C2(n13434), .A(n13433), .B(n13436), .ZN(
        P3_U3490) );
  NAND2_X1 U15649 ( .A1(n15637), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13435) );
  OAI211_X1 U15650 ( .C1(n13508), .C2(n13485), .A(n13436), .B(n13435), .ZN(
        P3_U3489) );
  OAI22_X1 U15651 ( .A1(n13511), .A2(n13480), .B1(n13510), .B2(n13485), .ZN(
        n13437) );
  INV_X1 U15652 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13441) );
  AOI21_X1 U15653 ( .B1(n13440), .B2(n13486), .A(n13439), .ZN(n13514) );
  MUX2_X1 U15654 ( .A(n13441), .B(n13514), .S(n15639), .Z(n13442) );
  OAI21_X1 U15655 ( .B1(n13517), .B2(n13485), .A(n13442), .ZN(P3_U3485) );
  NAND2_X1 U15656 ( .A1(n13443), .A2(n15607), .ZN(n13444) );
  NAND2_X1 U15657 ( .A1(n13445), .A2(n13444), .ZN(n13518) );
  MUX2_X1 U15658 ( .A(n13518), .B(P3_REG1_REG_25__SCAN_IN), .S(n15637), .Z(
        n13446) );
  AOI21_X1 U15659 ( .B1(n13471), .B2(n13520), .A(n13446), .ZN(n13447) );
  INV_X1 U15660 ( .A(n13447), .ZN(P3_U3484) );
  INV_X1 U15661 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13450) );
  AOI21_X1 U15662 ( .B1(n15607), .B2(n13449), .A(n13448), .ZN(n13522) );
  MUX2_X1 U15663 ( .A(n13450), .B(n13522), .S(n15639), .Z(n13451) );
  OAI21_X1 U15664 ( .B1(n13525), .B2(n13485), .A(n13451), .ZN(P3_U3483) );
  INV_X1 U15665 ( .A(n13452), .ZN(n13529) );
  INV_X1 U15666 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13456) );
  INV_X1 U15667 ( .A(n13453), .ZN(n13455) );
  AOI21_X1 U15668 ( .B1(n15607), .B2(n13455), .A(n13454), .ZN(n13526) );
  MUX2_X1 U15669 ( .A(n13456), .B(n13526), .S(n15639), .Z(n13457) );
  OAI21_X1 U15670 ( .B1(n13529), .B2(n13485), .A(n13457), .ZN(P3_U3482) );
  INV_X1 U15671 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13458) );
  MUX2_X1 U15672 ( .A(n13458), .B(n13530), .S(n15639), .Z(n13460) );
  NAND2_X1 U15673 ( .A1(n13532), .A2(n13471), .ZN(n13459) );
  OAI211_X1 U15674 ( .C1(n13535), .C2(n13480), .A(n13460), .B(n13459), .ZN(
        P3_U3481) );
  MUX2_X1 U15675 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n13536), .S(n15639), .Z(
        n13461) );
  AOI21_X1 U15676 ( .B1(n13471), .B2(n13538), .A(n13461), .ZN(n13462) );
  OAI21_X1 U15677 ( .B1(n13540), .B2(n13480), .A(n13462), .ZN(P3_U3480) );
  MUX2_X1 U15678 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13541), .S(n15639), .Z(
        n13463) );
  AOI21_X1 U15679 ( .B1(n13471), .B2(n13543), .A(n13463), .ZN(n13464) );
  OAI21_X1 U15680 ( .B1(n13545), .B2(n13480), .A(n13464), .ZN(P3_U3479) );
  OAI22_X1 U15681 ( .A1(n13547), .A2(n13480), .B1(n13546), .B2(n13485), .ZN(
        n13466) );
  MUX2_X1 U15682 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13548), .S(n15639), .Z(
        n13465) );
  OR2_X1 U15683 ( .A1(n13466), .A2(n13465), .ZN(P3_U3478) );
  MUX2_X1 U15684 ( .A(n13467), .B(n13551), .S(n15639), .Z(n13469) );
  NAND2_X1 U15685 ( .A1(n13553), .A2(n13471), .ZN(n13468) );
  OAI211_X1 U15686 ( .C1(n13480), .C2(n13556), .A(n13469), .B(n13468), .ZN(
        P3_U3477) );
  MUX2_X1 U15687 ( .A(n13470), .B(n13557), .S(n15639), .Z(n13473) );
  NAND2_X1 U15688 ( .A1(n13559), .A2(n13471), .ZN(n13472) );
  OAI211_X1 U15689 ( .C1(n13480), .C2(n13562), .A(n13473), .B(n13472), .ZN(
        P3_U3476) );
  MUX2_X1 U15690 ( .A(n13563), .B(P3_REG1_REG_16__SCAN_IN), .S(n15637), .Z(
        n13475) );
  OAI22_X1 U15691 ( .A1(n13565), .A2(n13480), .B1(n13564), .B2(n13485), .ZN(
        n13474) );
  OR2_X1 U15692 ( .A1(n13475), .A2(n13474), .ZN(P3_U3475) );
  AOI21_X1 U15693 ( .B1(n15614), .B2(n13477), .A(n13476), .ZN(n13568) );
  MUX2_X1 U15694 ( .A(n13478), .B(n13568), .S(n15639), .Z(n13479) );
  OAI21_X1 U15695 ( .B1(n13572), .B2(n13480), .A(n13479), .ZN(P3_U3474) );
  MUX2_X1 U15696 ( .A(n13481), .B(n13573), .S(n15639), .Z(n13484) );
  NAND2_X1 U15697 ( .A1(n13576), .A2(n13482), .ZN(n13483) );
  OAI211_X1 U15698 ( .C1(n13485), .C2(n13579), .A(n13484), .B(n13483), .ZN(
        P3_U3473) );
  NAND2_X1 U15699 ( .A1(n13487), .A2(n13486), .ZN(n13488) );
  OAI211_X1 U15700 ( .C1(n13490), .C2(n15621), .A(n13489), .B(n13488), .ZN(
        n13581) );
  MUX2_X1 U15701 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n13581), .S(n15639), .Z(
        P3_U3467) );
  XNOR2_X1 U15702 ( .A(n13496), .B(n13491), .ZN(n13494) );
  AOI21_X1 U15703 ( .B1(n13494), .B2(n13493), .A(n13492), .ZN(n13498) );
  XNOR2_X1 U15704 ( .A(n13496), .B(n13495), .ZN(n13499) );
  OR2_X1 U15705 ( .A1(n13499), .A2(n15609), .ZN(n13497) );
  AND2_X1 U15706 ( .A1(n13498), .A2(n13497), .ZN(n15588) );
  INV_X1 U15707 ( .A(n13499), .ZN(n15593) );
  NOR2_X1 U15708 ( .A1(n15621), .A2(n13500), .ZN(n15591) );
  AOI21_X1 U15709 ( .B1(n15593), .B2(n15607), .A(n15591), .ZN(n13501) );
  AND2_X1 U15710 ( .A1(n15588), .A2(n13501), .ZN(n15599) );
  INV_X1 U15711 ( .A(n15599), .ZN(n13502) );
  MUX2_X1 U15712 ( .A(n13502), .B(P3_REG1_REG_1__SCAN_IN), .S(n15637), .Z(
        P3_U3460) );
  NAND2_X1 U15713 ( .A1(n15629), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13504) );
  NAND2_X1 U15714 ( .A1(n13503), .A2(n15631), .ZN(n13507) );
  OAI211_X1 U15715 ( .C1(n13505), .C2(n13580), .A(n13504), .B(n13507), .ZN(
        P3_U3458) );
  NAND2_X1 U15716 ( .A1(n15629), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13506) );
  OAI211_X1 U15717 ( .C1(n13508), .C2(n13580), .A(n13507), .B(n13506), .ZN(
        P3_U3457) );
  OAI22_X1 U15718 ( .A1(n13511), .A2(n13571), .B1(n13510), .B2(n13580), .ZN(
        n13512) );
  INV_X1 U15719 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13515) );
  MUX2_X1 U15720 ( .A(n13515), .B(n13514), .S(n15631), .Z(n13516) );
  OAI21_X1 U15721 ( .B1(n13517), .B2(n13580), .A(n13516), .ZN(P3_U3453) );
  MUX2_X1 U15722 ( .A(n13518), .B(P3_REG0_REG_25__SCAN_IN), .S(n15629), .Z(
        n13519) );
  AOI21_X1 U15723 ( .B1(n9136), .B2(n13520), .A(n13519), .ZN(n13521) );
  INV_X1 U15724 ( .A(n13521), .ZN(P3_U3452) );
  INV_X1 U15725 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13523) );
  MUX2_X1 U15726 ( .A(n13523), .B(n13522), .S(n15631), .Z(n13524) );
  OAI21_X1 U15727 ( .B1(n13525), .B2(n13580), .A(n13524), .ZN(P3_U3451) );
  INV_X1 U15728 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13527) );
  MUX2_X1 U15729 ( .A(n13527), .B(n13526), .S(n15631), .Z(n13528) );
  OAI21_X1 U15730 ( .B1(n13529), .B2(n13580), .A(n13528), .ZN(P3_U3450) );
  INV_X1 U15731 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13531) );
  MUX2_X1 U15732 ( .A(n13531), .B(n13530), .S(n15631), .Z(n13534) );
  NAND2_X1 U15733 ( .A1(n13532), .A2(n9136), .ZN(n13533) );
  OAI211_X1 U15734 ( .C1(n13535), .C2(n13571), .A(n13534), .B(n13533), .ZN(
        P3_U3449) );
  MUX2_X1 U15735 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n13536), .S(n15631), .Z(
        n13537) );
  AOI21_X1 U15736 ( .B1(n9136), .B2(n13538), .A(n13537), .ZN(n13539) );
  OAI21_X1 U15737 ( .B1(n13540), .B2(n13571), .A(n13539), .ZN(P3_U3448) );
  MUX2_X1 U15738 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13541), .S(n15631), .Z(
        n13542) );
  AOI21_X1 U15739 ( .B1(n9136), .B2(n13543), .A(n13542), .ZN(n13544) );
  OAI21_X1 U15740 ( .B1(n13545), .B2(n13571), .A(n13544), .ZN(P3_U3447) );
  OAI22_X1 U15741 ( .A1(n13547), .A2(n13571), .B1(n13546), .B2(n13580), .ZN(
        n13550) );
  MUX2_X1 U15742 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13548), .S(n15631), .Z(
        n13549) );
  OR2_X1 U15743 ( .A1(n13550), .A2(n13549), .ZN(P3_U3446) );
  INV_X1 U15744 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13552) );
  MUX2_X1 U15745 ( .A(n13552), .B(n13551), .S(n15631), .Z(n13555) );
  NAND2_X1 U15746 ( .A1(n13553), .A2(n9136), .ZN(n13554) );
  OAI211_X1 U15747 ( .C1(n13556), .C2(n13571), .A(n13555), .B(n13554), .ZN(
        P3_U3444) );
  INV_X1 U15748 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13558) );
  MUX2_X1 U15749 ( .A(n13558), .B(n13557), .S(n15631), .Z(n13561) );
  NAND2_X1 U15750 ( .A1(n13559), .A2(n9136), .ZN(n13560) );
  OAI211_X1 U15751 ( .C1(n13562), .C2(n13571), .A(n13561), .B(n13560), .ZN(
        P3_U3441) );
  MUX2_X1 U15752 ( .A(n13563), .B(P3_REG0_REG_16__SCAN_IN), .S(n15629), .Z(
        n13567) );
  OAI22_X1 U15753 ( .A1(n13565), .A2(n13571), .B1(n13564), .B2(n13580), .ZN(
        n13566) );
  OR2_X1 U15754 ( .A1(n13567), .A2(n13566), .ZN(P3_U3438) );
  INV_X1 U15755 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13569) );
  MUX2_X1 U15756 ( .A(n13569), .B(n13568), .S(n15631), .Z(n13570) );
  OAI21_X1 U15757 ( .B1(n13572), .B2(n13571), .A(n13570), .ZN(P3_U3435) );
  INV_X1 U15758 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13574) );
  MUX2_X1 U15759 ( .A(n13574), .B(n13573), .S(n15631), .Z(n13578) );
  NAND2_X1 U15760 ( .A1(n13576), .A2(n13575), .ZN(n13577) );
  OAI211_X1 U15761 ( .C1(n13580), .C2(n13579), .A(n13578), .B(n13577), .ZN(
        P3_U3432) );
  MUX2_X1 U15762 ( .A(P3_REG0_REG_8__SCAN_IN), .B(n13581), .S(n15631), .Z(
        P3_U3414) );
  MUX2_X1 U15763 ( .A(n13582), .B(P3_D_REG_1__SCAN_IN), .S(n13583), .Z(
        P3_U3377) );
  MUX2_X1 U15764 ( .A(n13584), .B(P3_D_REG_0__SCAN_IN), .S(n13583), .Z(
        P3_U3376) );
  NAND2_X1 U15765 ( .A1(n13586), .A2(n13585), .ZN(n13591) );
  INV_X1 U15766 ( .A(n13587), .ZN(n13589) );
  NAND4_X1 U15767 ( .A1(n13589), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n13588), .ZN(n13590) );
  OAI211_X1 U15768 ( .C1(n13592), .C2(n13607), .A(n13591), .B(n13590), .ZN(
        P3_U3264) );
  INV_X1 U15769 ( .A(n13593), .ZN(n13595) );
  OAI222_X1 U15770 ( .A1(n13598), .A2(n13596), .B1(n13610), .B2(n13595), .C1(
        P3_U3151), .C2(n13594), .ZN(P3_U3266) );
  INV_X1 U15771 ( .A(n13597), .ZN(n13600) );
  OAI222_X1 U15772 ( .A1(P3_U3151), .A2(n6983), .B1(n13610), .B2(n13600), .C1(
        n13599), .C2(n13598), .ZN(P3_U3268) );
  INV_X1 U15773 ( .A(n13602), .ZN(n13603) );
  OAI222_X1 U15774 ( .A1(P3_U3151), .A2(n13605), .B1(n13607), .B2(n13604), 
        .C1(n13610), .C2(n13603), .ZN(P3_U3269) );
  INV_X1 U15775 ( .A(n13606), .ZN(n13609) );
  OAI222_X1 U15776 ( .A1(P3_U3151), .A2(n13611), .B1(n13610), .B2(n13609), 
        .C1(n13608), .C2(n13607), .ZN(P3_U3270) );
  INV_X1 U15777 ( .A(n14541), .ZN(n14370) );
  NOR2_X1 U15778 ( .A1(n13721), .A2(n13614), .ZN(n13616) );
  XNOR2_X1 U15779 ( .A(n13616), .B(n13615), .ZN(n13618) );
  AOI21_X1 U15780 ( .B1(n13618), .B2(n13619), .A(n13753), .ZN(n13617) );
  OAI21_X1 U15781 ( .B1(n13619), .B2(n13618), .A(n13617), .ZN(n13626) );
  NAND2_X1 U15782 ( .A1(n14086), .A2(n13725), .ZN(n13621) );
  NAND2_X1 U15783 ( .A1(n14088), .A2(n14073), .ZN(n13620) );
  NAND2_X1 U15784 ( .A1(n13621), .A2(n13620), .ZN(n14361) );
  INV_X1 U15785 ( .A(n14367), .ZN(n13623) );
  OAI22_X1 U15786 ( .A1(n13623), .A2(n13748), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13622), .ZN(n13624) );
  AOI21_X1 U15787 ( .B1(n14361), .B2(n13746), .A(n13624), .ZN(n13625) );
  OAI211_X1 U15788 ( .C1(n14370), .C2(n13738), .A(n13626), .B(n13625), .ZN(
        P2_U3188) );
  INV_X1 U15789 ( .A(n14433), .ZN(n14644) );
  OAI21_X1 U15790 ( .B1(n13627), .B2(n13629), .A(n13628), .ZN(n13630) );
  NAND2_X1 U15791 ( .A1(n13630), .A2(n13714), .ZN(n13633) );
  AOI22_X1 U15792 ( .A1(n14090), .A2(n13725), .B1(n14073), .B2(n14092), .ZN(
        n14429) );
  NAND2_X1 U15793 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14282)
         );
  OAI21_X1 U15794 ( .B1(n14429), .B2(n13726), .A(n14282), .ZN(n13631) );
  AOI21_X1 U15795 ( .B1(n14434), .B2(n13700), .A(n13631), .ZN(n13632) );
  OAI211_X1 U15796 ( .C1(n14644), .C2(n13738), .A(n13633), .B(n13632), .ZN(
        P2_U3191) );
  OAI211_X1 U15797 ( .C1(n13636), .C2(n13635), .A(n13634), .B(n13714), .ZN(
        n13641) );
  OAI22_X1 U15798 ( .A1(n13960), .A2(n13734), .B1(n14039), .B2(n13732), .ZN(
        n14392) );
  INV_X1 U15799 ( .A(n14392), .ZN(n13638) );
  OAI22_X1 U15800 ( .A1(n13638), .A2(n13726), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13637), .ZN(n13639) );
  AOI21_X1 U15801 ( .B1(n14399), .B2(n13700), .A(n13639), .ZN(n13640) );
  OAI211_X1 U15802 ( .C1(n7763), .C2(n13738), .A(n13641), .B(n13640), .ZN(
        P2_U3195) );
  OAI211_X1 U15803 ( .C1(n13644), .C2(n13643), .A(n13642), .B(n13714), .ZN(
        n13648) );
  AOI22_X1 U15804 ( .A1(n14084), .A2(n13725), .B1(n14073), .B2(n14086), .ZN(
        n14335) );
  AOI22_X1 U15805 ( .A1(n14340), .A2(n13700), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13645) );
  OAI21_X1 U15806 ( .B1(n14335), .B2(n13726), .A(n13645), .ZN(n13646) );
  AOI21_X1 U15807 ( .B1(n14629), .B2(n13751), .A(n13646), .ZN(n13647) );
  NAND2_X1 U15808 ( .A1(n13648), .A2(n13647), .ZN(P2_U3197) );
  XNOR2_X1 U15809 ( .A(n13649), .B(n13650), .ZN(n13744) );
  INV_X1 U15810 ( .A(n13650), .ZN(n13651) );
  AOI22_X1 U15811 ( .A1(n13744), .A2(n13743), .B1(n13649), .B2(n13651), .ZN(
        n13655) );
  NAND2_X1 U15812 ( .A1(n13653), .A2(n13652), .ZN(n13654) );
  XNOR2_X1 U15813 ( .A(n13655), .B(n13654), .ZN(n13662) );
  INV_X1 U15814 ( .A(n13656), .ZN(n14484) );
  OAI22_X1 U15815 ( .A1(n13896), .A2(n13734), .B1(n13657), .B2(n13732), .ZN(
        n14483) );
  NOR2_X1 U15816 ( .A1(n13658), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14219) );
  AOI21_X1 U15817 ( .B1(n13746), .B2(n14483), .A(n14219), .ZN(n13659) );
  OAI21_X1 U15818 ( .B1(n14484), .B2(n13748), .A(n13659), .ZN(n13660) );
  AOI21_X1 U15819 ( .B1(n14655), .B2(n13751), .A(n13660), .ZN(n13661) );
  OAI21_X1 U15820 ( .B1(n13662), .B2(n13753), .A(n13661), .ZN(P2_U3198) );
  OAI21_X1 U15821 ( .B1(n13665), .B2(n13664), .A(n13663), .ZN(n13666) );
  NAND2_X1 U15822 ( .A1(n13666), .A2(n13714), .ZN(n13672) );
  NAND2_X1 U15823 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14152) );
  INV_X1 U15824 ( .A(n13667), .ZN(n13668) );
  AOI22_X1 U15825 ( .A1(n13751), .A2(n13806), .B1(n13700), .B2(n13668), .ZN(
        n13671) );
  NAND2_X1 U15826 ( .A1(n13746), .A2(n13669), .ZN(n13670) );
  NAND4_X1 U15827 ( .A1(n13672), .A2(n14152), .A3(n13671), .A4(n13670), .ZN(
        P2_U3199) );
  OAI21_X1 U15828 ( .B1(n13675), .B2(n13674), .A(n13673), .ZN(n13676) );
  NAND2_X1 U15829 ( .A1(n13676), .A2(n13714), .ZN(n13682) );
  NAND2_X1 U15830 ( .A1(n14092), .A2(n13725), .ZN(n13678) );
  NAND2_X1 U15831 ( .A1(n14094), .A2(n14073), .ZN(n13677) );
  NAND2_X1 U15832 ( .A1(n13678), .A2(n13677), .ZN(n14460) );
  INV_X1 U15833 ( .A(n14460), .ZN(n13679) );
  NAND2_X1 U15834 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14235)
         );
  OAI21_X1 U15835 ( .B1(n13679), .B2(n13726), .A(n14235), .ZN(n13680) );
  AOI21_X1 U15836 ( .B1(n14472), .B2(n13700), .A(n13680), .ZN(n13681) );
  OAI211_X1 U15837 ( .C1(n7729), .C2(n13738), .A(n13682), .B(n13681), .ZN(
        P2_U3200) );
  INV_X1 U15838 ( .A(n14536), .ZN(n13690) );
  OAI211_X1 U15839 ( .C1(n13685), .C2(n13684), .A(n13683), .B(n13714), .ZN(
        n13689) );
  OAI22_X1 U15840 ( .A1(n13733), .A2(n13734), .B1(n14064), .B2(n13732), .ZN(
        n14349) );
  OAI22_X1 U15841 ( .A1(n14353), .A2(n13748), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13686), .ZN(n13687) );
  AOI21_X1 U15842 ( .B1(n14349), .B2(n13746), .A(n13687), .ZN(n13688) );
  OAI211_X1 U15843 ( .C1(n13690), .C2(n13738), .A(n13689), .B(n13688), .ZN(
        P2_U3201) );
  AOI21_X1 U15844 ( .B1(n13693), .B2(n13692), .A(n13691), .ZN(n13697) );
  INV_X1 U15845 ( .A(n13694), .ZN(n13696) );
  OAI21_X1 U15846 ( .B1(n13697), .B2(n13696), .A(n13695), .ZN(n13698) );
  NAND2_X1 U15847 ( .A1(n13698), .A2(n13714), .ZN(n13704) );
  NAND2_X1 U15848 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14137) );
  AOI22_X1 U15849 ( .A1(n13751), .A2(n13791), .B1(n13700), .B2(n13699), .ZN(
        n13703) );
  NAND2_X1 U15850 ( .A1(n13746), .A2(n13701), .ZN(n13702) );
  NAND4_X1 U15851 ( .A1(n13704), .A2(n14137), .A3(n13703), .A4(n13702), .ZN(
        P2_U3202) );
  NAND2_X1 U15852 ( .A1(n6616), .A2(n13706), .ZN(n13707) );
  XNOR2_X1 U15853 ( .A(n13705), .B(n13707), .ZN(n13713) );
  OAI22_X1 U15854 ( .A1(n13709), .A2(n13734), .B1(n13708), .B2(n13732), .ZN(
        n14408) );
  AOI22_X1 U15855 ( .A1(n14408), .A2(n13746), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13710) );
  OAI21_X1 U15856 ( .B1(n14410), .B2(n13748), .A(n13710), .ZN(n13711) );
  AOI21_X1 U15857 ( .B1(n14557), .B2(n13751), .A(n13711), .ZN(n13712) );
  OAI21_X1 U15858 ( .B1(n13713), .B2(n13753), .A(n13712), .ZN(P2_U3205) );
  OAI21_X1 U15859 ( .B1(n13613), .B2(n13715), .A(n13714), .ZN(n13722) );
  NAND2_X1 U15860 ( .A1(n14087), .A2(n13725), .ZN(n13717) );
  NAND2_X1 U15861 ( .A1(n14089), .A2(n14073), .ZN(n13716) );
  NAND2_X1 U15862 ( .A1(n13717), .A2(n13716), .ZN(n14375) );
  AOI22_X1 U15863 ( .A1(n14375), .A2(n13746), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13718) );
  OAI21_X1 U15864 ( .B1(n14384), .B2(n13748), .A(n13718), .ZN(n13719) );
  AOI21_X1 U15865 ( .B1(n14634), .B2(n13751), .A(n13719), .ZN(n13720) );
  OAI21_X1 U15866 ( .B1(n13722), .B2(n13721), .A(n13720), .ZN(P2_U3207) );
  XNOR2_X1 U15867 ( .A(n13723), .B(n13724), .ZN(n13730) );
  NOR2_X1 U15868 ( .A1(n13748), .A2(n14451), .ZN(n13728) );
  AOI22_X1 U15869 ( .A1(n14091), .A2(n13725), .B1(n14073), .B2(n14093), .ZN(
        n14442) );
  OAI22_X1 U15870 ( .A1(n14442), .A2(n13726), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14263), .ZN(n13727) );
  AOI211_X1 U15871 ( .C1(n14450), .C2(n13751), .A(n13728), .B(n13727), .ZN(
        n13729) );
  OAI21_X1 U15872 ( .B1(n13730), .B2(n13753), .A(n13729), .ZN(P2_U3210) );
  OAI22_X1 U15873 ( .A1(n13735), .A2(n13734), .B1(n13733), .B2(n13732), .ZN(
        n14320) );
  INV_X1 U15874 ( .A(n14323), .ZN(n13737) );
  OAI22_X1 U15875 ( .A1(n13737), .A2(n13748), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13736), .ZN(n13740) );
  NOR2_X1 U15876 ( .A1(n14325), .A2(n13738), .ZN(n13739) );
  AOI211_X1 U15877 ( .C1(n13746), .C2(n14320), .A(n13740), .B(n13739), .ZN(
        n13741) );
  OAI21_X1 U15878 ( .B1(n13742), .B2(n13753), .A(n13741), .ZN(P2_U3212) );
  XNOR2_X1 U15879 ( .A(n13744), .B(n13743), .ZN(n13754) );
  AOI22_X1 U15880 ( .A1(n13746), .A2(n13745), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13747) );
  OAI21_X1 U15881 ( .B1(n13749), .B2(n13748), .A(n13747), .ZN(n13750) );
  AOI21_X1 U15882 ( .B1(n13887), .B2(n13751), .A(n13750), .ZN(n13752) );
  OAI21_X1 U15883 ( .B1(n13754), .B2(n13753), .A(n13752), .ZN(P2_U3213) );
  AND2_X1 U15884 ( .A1(n13757), .A2(n14280), .ZN(n13758) );
  NOR2_X1 U15885 ( .A1(n14033), .A2(n13758), .ZN(n13762) );
  AOI21_X1 U15886 ( .B1(n13763), .B2(n13956), .A(n13762), .ZN(n13759) );
  NAND2_X1 U15887 ( .A1(n13760), .A2(n13759), .ZN(n13766) );
  NAND2_X1 U15888 ( .A1(n13763), .A2(n13762), .ZN(n13764) );
  NAND2_X1 U15889 ( .A1(n13766), .A2(n13765), .ZN(n13777) );
  NAND2_X1 U15890 ( .A1(n14110), .A2(n13956), .ZN(n13768) );
  NAND2_X1 U15891 ( .A1(n7087), .A2(n13761), .ZN(n13767) );
  NAND2_X1 U15892 ( .A1(n13768), .A2(n13767), .ZN(n13778) );
  NAND2_X1 U15893 ( .A1(n13777), .A2(n13778), .ZN(n13771) );
  NAND2_X1 U15894 ( .A1(n14110), .A2(n13761), .ZN(n13769) );
  OAI21_X1 U15895 ( .B1(n10034), .B2(n13761), .A(n13769), .ZN(n13770) );
  NAND2_X1 U15896 ( .A1(n13771), .A2(n13770), .ZN(n13781) );
  NAND2_X1 U15897 ( .A1(n14109), .A2(n13761), .ZN(n13772) );
  NAND2_X1 U15898 ( .A1(n13773), .A2(n13772), .ZN(n13784) );
  NAND2_X1 U15899 ( .A1(n14109), .A2(n13956), .ZN(n13776) );
  OR2_X1 U15900 ( .A1(n13774), .A2(n13956), .ZN(n13775) );
  AND2_X1 U15901 ( .A1(n13776), .A2(n13775), .ZN(n13785) );
  NAND2_X1 U15902 ( .A1(n13784), .A2(n13785), .ZN(n13780) );
  NAND3_X1 U15903 ( .A1(n13781), .A2(n13780), .A3(n13779), .ZN(n13790) );
  NAND2_X1 U15904 ( .A1(n14108), .A2(n13761), .ZN(n13782) );
  OAI21_X1 U15905 ( .B1(n13783), .B2(n13761), .A(n13782), .ZN(n13794) );
  AOI22_X1 U15906 ( .A1(n15563), .A2(n13761), .B1(n14108), .B2(n13956), .ZN(
        n13795) );
  OR2_X1 U15907 ( .A1(n13794), .A2(n13795), .ZN(n13789) );
  INV_X1 U15908 ( .A(n13784), .ZN(n13787) );
  INV_X1 U15909 ( .A(n13785), .ZN(n13786) );
  NAND2_X1 U15910 ( .A1(n13787), .A2(n13786), .ZN(n13788) );
  NAND3_X1 U15911 ( .A1(n13790), .A2(n13789), .A3(n13788), .ZN(n13797) );
  AOI22_X1 U15912 ( .A1(n13791), .A2(n13761), .B1(n14107), .B2(n13956), .ZN(
        n13799) );
  NAND2_X1 U15913 ( .A1(n13791), .A2(n13956), .ZN(n13793) );
  NAND2_X1 U15914 ( .A1(n14107), .A2(n13761), .ZN(n13792) );
  NAND2_X1 U15915 ( .A1(n13793), .A2(n13792), .ZN(n13798) );
  AOI22_X1 U15916 ( .A1(n13799), .A2(n13798), .B1(n13795), .B2(n13794), .ZN(
        n13796) );
  NAND2_X1 U15917 ( .A1(n13797), .A2(n13796), .ZN(n13803) );
  INV_X1 U15918 ( .A(n13798), .ZN(n13801) );
  INV_X1 U15919 ( .A(n13799), .ZN(n13800) );
  NAND2_X1 U15920 ( .A1(n13801), .A2(n13800), .ZN(n13802) );
  NAND2_X1 U15921 ( .A1(n13803), .A2(n13802), .ZN(n13810) );
  NAND2_X1 U15922 ( .A1(n13806), .A2(n6440), .ZN(n13805) );
  OR2_X1 U15923 ( .A1(n13808), .A2(n13761), .ZN(n13804) );
  NAND2_X1 U15924 ( .A1(n13806), .A2(n13956), .ZN(n13807) );
  OAI21_X1 U15925 ( .B1(n13808), .B2(n13956), .A(n13807), .ZN(n13809) );
  NAND2_X1 U15926 ( .A1(n13813), .A2(n6433), .ZN(n13812) );
  OR2_X1 U15927 ( .A1(n13815), .A2(n13956), .ZN(n13811) );
  NAND2_X1 U15928 ( .A1(n13813), .A2(n13818), .ZN(n13814) );
  OAI21_X1 U15929 ( .B1(n13815), .B2(n6441), .A(n13814), .ZN(n13816) );
  NAND2_X1 U15930 ( .A1(n13817), .A2(n13816), .ZN(n13827) );
  NOR2_X1 U15931 ( .A1(n13820), .A2(n6433), .ZN(n13819) );
  AOI21_X1 U15932 ( .B1(n14614), .B2(n6433), .A(n13819), .ZN(n13829) );
  NAND2_X1 U15933 ( .A1(n14614), .A2(n13985), .ZN(n13822) );
  OR2_X1 U15934 ( .A1(n13820), .A2(n6440), .ZN(n13821) );
  NAND2_X1 U15935 ( .A1(n13822), .A2(n13821), .ZN(n13828) );
  NAND2_X1 U15936 ( .A1(n13829), .A2(n13828), .ZN(n13826) );
  INV_X1 U15937 ( .A(n13823), .ZN(n13824) );
  NAND2_X1 U15938 ( .A1(n13824), .A2(n6541), .ZN(n13825) );
  NAND3_X1 U15939 ( .A1(n13827), .A2(n13826), .A3(n13825), .ZN(n13833) );
  INV_X1 U15940 ( .A(n13828), .ZN(n13831) );
  INV_X1 U15941 ( .A(n13829), .ZN(n13830) );
  NAND2_X1 U15942 ( .A1(n13831), .A2(n13830), .ZN(n13832) );
  NAND2_X1 U15943 ( .A1(n13840), .A2(n6433), .ZN(n13835) );
  NAND2_X1 U15944 ( .A1(n14103), .A2(n13985), .ZN(n13834) );
  NOR2_X1 U15945 ( .A1(n13837), .A2(n6441), .ZN(n13836) );
  AOI21_X1 U15946 ( .B1(n14610), .B2(n13818), .A(n13836), .ZN(n13843) );
  NAND2_X1 U15947 ( .A1(n14610), .A2(n6433), .ZN(n13839) );
  OR2_X1 U15948 ( .A1(n13837), .A2(n6433), .ZN(n13838) );
  NAND2_X1 U15949 ( .A1(n13839), .A2(n13838), .ZN(n13842) );
  AOI22_X1 U15950 ( .A1(n13840), .A2(n6441), .B1(n14103), .B2(n13956), .ZN(
        n13841) );
  NAND2_X1 U15951 ( .A1(n13843), .A2(n13842), .ZN(n13844) );
  NAND2_X1 U15952 ( .A1(n14604), .A2(n13956), .ZN(n13846) );
  OR2_X1 U15953 ( .A1(n13848), .A2(n6433), .ZN(n13845) );
  NAND2_X1 U15954 ( .A1(n13846), .A2(n13845), .ZN(n13852) );
  NAND2_X1 U15955 ( .A1(n13851), .A2(n13852), .ZN(n13850) );
  NAND2_X1 U15956 ( .A1(n14604), .A2(n6440), .ZN(n13847) );
  OAI21_X1 U15957 ( .B1(n13848), .B2(n13818), .A(n13847), .ZN(n13849) );
  INV_X1 U15958 ( .A(n13851), .ZN(n13854) );
  INV_X1 U15959 ( .A(n13852), .ZN(n13853) );
  NAND2_X1 U15960 ( .A1(n13860), .A2(n6441), .ZN(n13856) );
  NAND2_X1 U15961 ( .A1(n14099), .A2(n6433), .ZN(n13855) );
  AND2_X1 U15962 ( .A1(n14098), .A2(n13818), .ZN(n13857) );
  AOI21_X1 U15963 ( .B1(n14599), .B2(n6433), .A(n13857), .ZN(n13863) );
  NAND2_X1 U15964 ( .A1(n14599), .A2(n13818), .ZN(n13859) );
  NAND2_X1 U15965 ( .A1(n14098), .A2(n6433), .ZN(n13858) );
  NAND2_X1 U15966 ( .A1(n13859), .A2(n13858), .ZN(n13862) );
  AOI22_X1 U15967 ( .A1(n13860), .A2(n6433), .B1(n13818), .B2(n14099), .ZN(
        n13861) );
  NAND2_X1 U15968 ( .A1(n13863), .A2(n13862), .ZN(n13864) );
  NAND2_X1 U15969 ( .A1(n13865), .A2(n13864), .ZN(n13872) );
  NAND2_X1 U15970 ( .A1(n14594), .A2(n6440), .ZN(n13867) );
  NAND2_X1 U15971 ( .A1(n14097), .A2(n13956), .ZN(n13866) );
  NAND2_X1 U15972 ( .A1(n13867), .A2(n13866), .ZN(n13873) );
  NAND2_X1 U15973 ( .A1(n13872), .A2(n13873), .ZN(n13871) );
  NAND2_X1 U15974 ( .A1(n14594), .A2(n6433), .ZN(n13868) );
  OAI21_X1 U15975 ( .B1(n13869), .B2(n13956), .A(n13868), .ZN(n13870) );
  NAND2_X1 U15976 ( .A1(n13871), .A2(n13870), .ZN(n13877) );
  INV_X1 U15977 ( .A(n13872), .ZN(n13875) );
  INV_X1 U15978 ( .A(n13873), .ZN(n13874) );
  NAND2_X1 U15979 ( .A1(n13875), .A2(n13874), .ZN(n13876) );
  NAND2_X1 U15980 ( .A1(n13877), .A2(n13876), .ZN(n13884) );
  NAND2_X1 U15981 ( .A1(n13880), .A2(n6433), .ZN(n13879) );
  NAND2_X1 U15982 ( .A1(n14096), .A2(n13818), .ZN(n13878) );
  NAND2_X1 U15983 ( .A1(n13879), .A2(n13878), .ZN(n13885) );
  NAND2_X1 U15984 ( .A1(n13880), .A2(n13985), .ZN(n13881) );
  OAI21_X1 U15985 ( .B1(n13882), .B2(n13985), .A(n13881), .ZN(n13883) );
  AND2_X1 U15986 ( .A1(n14095), .A2(n13818), .ZN(n13886) );
  AOI21_X1 U15987 ( .B1(n13887), .B2(n6433), .A(n13886), .ZN(n13904) );
  NAND2_X1 U15988 ( .A1(n13887), .A2(n6441), .ZN(n13889) );
  NAND2_X1 U15989 ( .A1(n14095), .A2(n13956), .ZN(n13888) );
  NAND2_X1 U15990 ( .A1(n13889), .A2(n13888), .ZN(n13903) );
  NAND2_X1 U15991 ( .A1(n13904), .A2(n13903), .ZN(n13902) );
  AND2_X1 U15992 ( .A1(n14094), .A2(n13985), .ZN(n13890) );
  AOI21_X1 U15993 ( .B1(n14655), .B2(n6433), .A(n13890), .ZN(n13906) );
  NAND2_X1 U15994 ( .A1(n14655), .A2(n13985), .ZN(n13892) );
  NAND2_X1 U15995 ( .A1(n14094), .A2(n6433), .ZN(n13891) );
  NAND2_X1 U15996 ( .A1(n13892), .A2(n13891), .ZN(n13905) );
  NAND2_X1 U15997 ( .A1(n13906), .A2(n13905), .ZN(n13901) );
  NAND3_X1 U15998 ( .A1(n13899), .A2(n13893), .A3(n6441), .ZN(n13898) );
  NAND2_X1 U15999 ( .A1(n13893), .A2(n6433), .ZN(n13895) );
  NAND2_X1 U16000 ( .A1(n13896), .A2(n13985), .ZN(n13894) );
  OAI21_X1 U16001 ( .B1(n13896), .B2(n13895), .A(n13894), .ZN(n13897) );
  OAI211_X1 U16002 ( .C1(n13899), .C2(n6441), .A(n13898), .B(n13897), .ZN(
        n13900) );
  AND2_X1 U16003 ( .A1(n13901), .A2(n13900), .ZN(n13911) );
  INV_X1 U16004 ( .A(n13903), .ZN(n13910) );
  INV_X1 U16005 ( .A(n13904), .ZN(n13909) );
  INV_X1 U16006 ( .A(n13905), .ZN(n13908) );
  INV_X1 U16007 ( .A(n13906), .ZN(n13907) );
  AOI22_X1 U16008 ( .A1(n13910), .A2(n13909), .B1(n13908), .B2(n13907), .ZN(
        n13913) );
  INV_X1 U16009 ( .A(n13911), .ZN(n13912) );
  NAND2_X1 U16010 ( .A1(n14651), .A2(n6440), .ZN(n13915) );
  NAND2_X1 U16011 ( .A1(n14093), .A2(n13956), .ZN(n13914) );
  OAI211_X1 U16012 ( .C1(n14651), .C2(n14093), .A(n13915), .B(n13914), .ZN(
        n13916) );
  AND2_X1 U16013 ( .A1(n13917), .A2(n13916), .ZN(n13918) );
  AND2_X1 U16014 ( .A1(n14092), .A2(n6433), .ZN(n13919) );
  AOI21_X1 U16015 ( .B1(n14450), .B2(n6441), .A(n13919), .ZN(n13929) );
  NAND2_X1 U16016 ( .A1(n14450), .A2(n13956), .ZN(n13921) );
  NAND2_X1 U16017 ( .A1(n14092), .A2(n13985), .ZN(n13920) );
  NAND2_X1 U16018 ( .A1(n13921), .A2(n13920), .ZN(n13928) );
  NAND2_X1 U16019 ( .A1(n14091), .A2(n13956), .ZN(n13922) );
  NAND2_X1 U16020 ( .A1(n13923), .A2(n13922), .ZN(n13936) );
  AND2_X1 U16021 ( .A1(n14091), .A2(n6441), .ZN(n13924) );
  AOI21_X1 U16022 ( .B1(n14433), .B2(n13956), .A(n13924), .ZN(n13937) );
  NAND2_X1 U16023 ( .A1(n13936), .A2(n13937), .ZN(n13930) );
  INV_X1 U16024 ( .A(n13925), .ZN(n13926) );
  NAND2_X1 U16025 ( .A1(n13927), .A2(n13926), .ZN(n13943) );
  NAND3_X1 U16026 ( .A1(n13930), .A2(n13929), .A3(n13928), .ZN(n13942) );
  NAND2_X1 U16027 ( .A1(n14557), .A2(n6441), .ZN(n13932) );
  NAND2_X1 U16028 ( .A1(n14090), .A2(n13956), .ZN(n13931) );
  NAND2_X1 U16029 ( .A1(n13932), .A2(n13931), .ZN(n13947) );
  INV_X1 U16030 ( .A(n13947), .ZN(n13935) );
  AND2_X1 U16031 ( .A1(n14090), .A2(n6441), .ZN(n13933) );
  AOI21_X1 U16032 ( .B1(n14557), .B2(n13956), .A(n13933), .ZN(n13948) );
  INV_X1 U16033 ( .A(n13948), .ZN(n13934) );
  NAND2_X1 U16034 ( .A1(n13935), .A2(n13934), .ZN(n13941) );
  INV_X1 U16035 ( .A(n13936), .ZN(n13939) );
  INV_X1 U16036 ( .A(n13937), .ZN(n13938) );
  NAND2_X1 U16037 ( .A1(n13939), .A2(n13938), .ZN(n13940) );
  NAND4_X1 U16038 ( .A1(n13943), .A2(n13942), .A3(n13941), .A4(n13940), .ZN(
        n13955) );
  AND2_X1 U16039 ( .A1(n14089), .A2(n13818), .ZN(n13944) );
  AOI21_X1 U16040 ( .B1(n14638), .B2(n13956), .A(n13944), .ZN(n13950) );
  NAND2_X1 U16041 ( .A1(n14638), .A2(n6441), .ZN(n13946) );
  NAND2_X1 U16042 ( .A1(n14089), .A2(n13956), .ZN(n13945) );
  NAND2_X1 U16043 ( .A1(n13946), .A2(n13945), .ZN(n13949) );
  AOI22_X1 U16044 ( .A1(n13950), .A2(n13949), .B1(n13948), .B2(n13947), .ZN(
        n13954) );
  INV_X1 U16045 ( .A(n13949), .ZN(n13952) );
  INV_X1 U16046 ( .A(n13950), .ZN(n13951) );
  AND2_X1 U16047 ( .A1(n13952), .A2(n13951), .ZN(n13953) );
  NOR2_X1 U16048 ( .A1(n13960), .A2(n13956), .ZN(n13957) );
  AOI21_X1 U16049 ( .B1(n14634), .B2(n13956), .A(n13957), .ZN(n13962) );
  INV_X1 U16050 ( .A(n13962), .ZN(n13958) );
  NAND2_X1 U16051 ( .A1(n14634), .A2(n6440), .ZN(n13959) );
  OAI21_X1 U16052 ( .B1(n13960), .B2(n13985), .A(n13959), .ZN(n13961) );
  NAND2_X1 U16053 ( .A1(n13963), .A2(n13962), .ZN(n13964) );
  NAND2_X1 U16054 ( .A1(n14541), .A2(n6440), .ZN(n13967) );
  NAND2_X1 U16055 ( .A1(n14087), .A2(n6433), .ZN(n13966) );
  NAND2_X1 U16056 ( .A1(n13967), .A2(n13966), .ZN(n13969) );
  NAND2_X1 U16057 ( .A1(n14536), .A2(n13956), .ZN(n13971) );
  NAND2_X1 U16058 ( .A1(n14086), .A2(n6440), .ZN(n13970) );
  NAND2_X1 U16059 ( .A1(n13971), .A2(n13970), .ZN(n13973) );
  AOI22_X1 U16060 ( .A1(n14536), .A2(n6440), .B1(n14086), .B2(n13956), .ZN(
        n13972) );
  NAND2_X1 U16061 ( .A1(n14629), .A2(n13985), .ZN(n13976) );
  NAND2_X1 U16062 ( .A1(n14085), .A2(n6433), .ZN(n13975) );
  NAND2_X1 U16063 ( .A1(n13976), .A2(n13975), .ZN(n13978) );
  AOI22_X1 U16064 ( .A1(n14629), .A2(n13956), .B1(n13818), .B2(n14085), .ZN(
        n13977) );
  AOI21_X1 U16065 ( .B1(n13979), .B2(n13978), .A(n13977), .ZN(n13981) );
  NAND2_X1 U16066 ( .A1(n14527), .A2(n13956), .ZN(n13983) );
  NAND2_X1 U16067 ( .A1(n14084), .A2(n13818), .ZN(n13982) );
  NAND2_X1 U16068 ( .A1(n14527), .A2(n13985), .ZN(n13984) );
  OAI21_X1 U16069 ( .B1(n13986), .B2(n13985), .A(n13984), .ZN(n13987) );
  NAND2_X1 U16070 ( .A1(n14519), .A2(n6441), .ZN(n13989) );
  NAND2_X1 U16071 ( .A1(n14083), .A2(n13956), .ZN(n13988) );
  NAND2_X1 U16072 ( .A1(n13989), .A2(n13988), .ZN(n14000) );
  AND2_X1 U16073 ( .A1(n14081), .A2(n13956), .ZN(n13990) );
  AOI21_X1 U16074 ( .B1(n14516), .B2(n6441), .A(n13990), .ZN(n14014) );
  NAND2_X1 U16075 ( .A1(n14516), .A2(n13956), .ZN(n13992) );
  NAND2_X1 U16076 ( .A1(n14081), .A2(n13985), .ZN(n13991) );
  NAND2_X1 U16077 ( .A1(n13992), .A2(n13991), .ZN(n14013) );
  NAND2_X1 U16078 ( .A1(n14014), .A2(n14013), .ZN(n14004) );
  AND2_X1 U16079 ( .A1(n14082), .A2(n13956), .ZN(n13993) );
  AOI21_X1 U16080 ( .B1(n14293), .B2(n6440), .A(n13993), .ZN(n14002) );
  NAND2_X1 U16081 ( .A1(n14293), .A2(n13956), .ZN(n13995) );
  NAND2_X1 U16082 ( .A1(n14082), .A2(n6440), .ZN(n13994) );
  NAND2_X1 U16083 ( .A1(n13995), .A2(n13994), .ZN(n14001) );
  NAND2_X1 U16084 ( .A1(n14002), .A2(n14001), .ZN(n13996) );
  AND2_X1 U16085 ( .A1(n14004), .A2(n13996), .ZN(n13998) );
  NAND2_X1 U16086 ( .A1(n14023), .A2(n14079), .ZN(n13997) );
  AOI22_X1 U16087 ( .A1(n14519), .A2(n6433), .B1(n13985), .B2(n14083), .ZN(
        n13999) );
  INV_X1 U16088 ( .A(n14001), .ZN(n14005) );
  INV_X1 U16089 ( .A(n14002), .ZN(n14003) );
  NAND4_X1 U16090 ( .A1(n14036), .A2(n14005), .A3(n14004), .A4(n14003), .ZN(
        n14018) );
  NAND2_X1 U16091 ( .A1(n14079), .A2(n13985), .ZN(n14007) );
  NAND2_X1 U16092 ( .A1(n14023), .A2(n6433), .ZN(n14006) );
  NAND3_X1 U16093 ( .A1(n14024), .A2(n14007), .A3(n14006), .ZN(n14016) );
  NOR2_X1 U16094 ( .A1(n14072), .A2(n8505), .ZN(n14008) );
  NAND2_X1 U16095 ( .A1(n14070), .A2(n14076), .ZN(n14029) );
  AND2_X1 U16096 ( .A1(n14008), .A2(n14029), .ZN(n14009) );
  NAND2_X1 U16097 ( .A1(n14079), .A2(n13956), .ZN(n14021) );
  INV_X1 U16098 ( .A(n14080), .ZN(n14037) );
  AOI21_X1 U16099 ( .B1(n14009), .B2(n14021), .A(n14037), .ZN(n14010) );
  AOI21_X1 U16100 ( .B1(n14622), .B2(n6440), .A(n14010), .ZN(n14020) );
  NAND2_X1 U16101 ( .A1(n14622), .A2(n13956), .ZN(n14012) );
  NAND2_X1 U16102 ( .A1(n14080), .A2(n6440), .ZN(n14011) );
  NAND2_X1 U16103 ( .A1(n14012), .A2(n14011), .ZN(n14019) );
  OAI22_X1 U16104 ( .A1(n14020), .A2(n14019), .B1(n14014), .B2(n14013), .ZN(
        n14015) );
  NAND2_X1 U16105 ( .A1(n14016), .A2(n14015), .ZN(n14017) );
  NAND2_X1 U16106 ( .A1(n14020), .A2(n14019), .ZN(n14027) );
  INV_X1 U16107 ( .A(n14021), .ZN(n14022) );
  AOI21_X1 U16108 ( .B1(n14023), .B2(n13985), .A(n14022), .ZN(n14025) );
  AND2_X1 U16109 ( .A1(n14025), .A2(n14024), .ZN(n14026) );
  NAND3_X1 U16110 ( .A1(n13756), .A2(n14280), .A3(n14041), .ZN(n14030) );
  AOI21_X1 U16111 ( .B1(n13756), .B2(n14031), .A(n14072), .ZN(n14032) );
  OAI21_X1 U16112 ( .B1(n14076), .B2(n14033), .A(n14032), .ZN(n14034) );
  NAND2_X1 U16113 ( .A1(n14071), .A2(n14034), .ZN(n14035) );
  XNOR2_X1 U16114 ( .A(n14622), .B(n14037), .ZN(n14069) );
  XNOR2_X1 U16115 ( .A(n14557), .B(n14039), .ZN(n14415) );
  INV_X1 U16116 ( .A(n14493), .ZN(n14480) );
  AND4_X1 U16117 ( .A1(n14042), .A2(n11429), .A3(n14041), .A4(n14040), .ZN(
        n14045) );
  NAND4_X1 U16118 ( .A1(n14046), .A2(n14045), .A3(n14044), .A4(n14043), .ZN(
        n14047) );
  NOR3_X1 U16119 ( .A1(n14049), .A2(n14048), .A3(n14047), .ZN(n14051) );
  NAND3_X1 U16120 ( .A1(n14052), .A2(n14051), .A3(n14050), .ZN(n14053) );
  NOR2_X1 U16121 ( .A1(n14054), .A2(n14053), .ZN(n14056) );
  NAND4_X1 U16122 ( .A1(n14057), .A2(n14056), .A3(n14055), .A4(n10061), .ZN(
        n14058) );
  NAND3_X1 U16123 ( .A1(n14445), .A2(n7793), .A3(n14060), .ZN(n14061) );
  NAND4_X1 U16124 ( .A1(n14347), .A2(n14378), .A3(n7810), .A4(n14394), .ZN(
        n14066) );
  NAND2_X1 U16125 ( .A1(n14063), .A2(n14062), .ZN(n14327) );
  INV_X1 U16126 ( .A(n14332), .ZN(n14065) );
  XNOR2_X1 U16127 ( .A(n14541), .B(n14064), .ZN(n14363) );
  NAND4_X1 U16128 ( .A1(n15558), .A2(n14074), .A3(n14073), .A4(n14072), .ZN(
        n14075) );
  OAI211_X1 U16129 ( .C1(n14076), .C2(n14078), .A(n14075), .B(P2_B_REG_SCAN_IN), .ZN(n14077) );
  INV_X2 U16130 ( .A(P2_U3947), .ZN(n14102) );
  MUX2_X1 U16131 ( .A(n14079), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14102), .Z(
        P2_U3562) );
  MUX2_X1 U16132 ( .A(n14080), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14102), .Z(
        P2_U3561) );
  MUX2_X1 U16133 ( .A(n14081), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14102), .Z(
        P2_U3560) );
  MUX2_X1 U16134 ( .A(n14082), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14102), .Z(
        P2_U3559) );
  MUX2_X1 U16135 ( .A(n14083), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14102), .Z(
        P2_U3558) );
  MUX2_X1 U16136 ( .A(n14084), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14102), .Z(
        P2_U3557) );
  MUX2_X1 U16137 ( .A(n14085), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14102), .Z(
        P2_U3556) );
  MUX2_X1 U16138 ( .A(n14086), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14102), .Z(
        P2_U3555) );
  MUX2_X1 U16139 ( .A(n14087), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14102), .Z(
        P2_U3554) );
  MUX2_X1 U16140 ( .A(n14088), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14102), .Z(
        P2_U3553) );
  MUX2_X1 U16141 ( .A(n14089), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14102), .Z(
        P2_U3552) );
  MUX2_X1 U16142 ( .A(n14090), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14102), .Z(
        P2_U3551) );
  MUX2_X1 U16143 ( .A(n14091), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14102), .Z(
        P2_U3550) );
  MUX2_X1 U16144 ( .A(n14092), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14102), .Z(
        P2_U3549) );
  MUX2_X1 U16145 ( .A(n14093), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14102), .Z(
        P2_U3548) );
  MUX2_X1 U16146 ( .A(n14094), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14102), .Z(
        P2_U3547) );
  MUX2_X1 U16147 ( .A(n14095), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14102), .Z(
        P2_U3546) );
  MUX2_X1 U16148 ( .A(n14096), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14102), .Z(
        P2_U3545) );
  MUX2_X1 U16149 ( .A(n14097), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14102), .Z(
        P2_U3544) );
  MUX2_X1 U16150 ( .A(n14098), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14102), .Z(
        P2_U3543) );
  MUX2_X1 U16151 ( .A(n14099), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14102), .Z(
        P2_U3542) );
  MUX2_X1 U16152 ( .A(n14100), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14102), .Z(
        P2_U3541) );
  MUX2_X1 U16153 ( .A(n14101), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14102), .Z(
        P2_U3540) );
  MUX2_X1 U16154 ( .A(n14103), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14102), .Z(
        P2_U3539) );
  MUX2_X1 U16155 ( .A(n14104), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14102), .Z(
        P2_U3538) );
  MUX2_X1 U16156 ( .A(n14105), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14102), .Z(
        P2_U3537) );
  MUX2_X1 U16157 ( .A(n14106), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14102), .Z(
        P2_U3536) );
  MUX2_X1 U16158 ( .A(n14107), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14102), .Z(
        P2_U3535) );
  MUX2_X1 U16159 ( .A(n14108), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14102), .Z(
        P2_U3534) );
  MUX2_X1 U16160 ( .A(n14109), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14102), .Z(
        P2_U3533) );
  MUX2_X1 U16161 ( .A(n14110), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14102), .Z(
        P2_U3532) );
  INV_X1 U16162 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n14111) );
  OAI22_X1 U16163 ( .A1(n15543), .A2(n14113), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14111), .ZN(n14112) );
  AOI21_X1 U16164 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n15525), .A(n14112), .ZN(
        n14122) );
  MUX2_X1 U16165 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n14504), .S(n14113), .Z(
        n14114) );
  OAI21_X1 U16166 ( .B1(n10908), .B2(n7134), .A(n14114), .ZN(n14115) );
  NAND3_X1 U16167 ( .A1(n15546), .A2(n14116), .A3(n14115), .ZN(n14121) );
  OAI211_X1 U16168 ( .C1(n14119), .C2(n14118), .A(n15537), .B(n14117), .ZN(
        n14120) );
  NAND3_X1 U16169 ( .A1(n14122), .A2(n14121), .A3(n14120), .ZN(P2_U3215) );
  NOR2_X1 U16170 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14123), .ZN(n14126) );
  NOR2_X1 U16171 ( .A1(n15543), .A2(n14124), .ZN(n14125) );
  AOI211_X1 U16172 ( .C1(n15525), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n14126), .B(
        n14125), .ZN(n14136) );
  OAI211_X1 U16173 ( .C1(n14129), .C2(n14128), .A(n15537), .B(n14127), .ZN(
        n14135) );
  MUX2_X1 U16174 ( .A(n11374), .B(P2_REG2_REG_3__SCAN_IN), .S(n14130), .Z(
        n14132) );
  NAND3_X1 U16175 ( .A1(n15531), .A2(n14132), .A3(n14131), .ZN(n14133) );
  NAND3_X1 U16176 ( .A1(n15546), .A2(n14147), .A3(n14133), .ZN(n14134) );
  NAND3_X1 U16177 ( .A1(n14136), .A2(n14135), .A3(n14134), .ZN(P2_U3217) );
  INV_X1 U16178 ( .A(n14137), .ZN(n14140) );
  NOR2_X1 U16179 ( .A1(n15543), .A2(n14138), .ZN(n14139) );
  AOI211_X1 U16180 ( .C1(n15525), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n14140), .B(
        n14139), .ZN(n14151) );
  OAI211_X1 U16181 ( .C1(n14143), .C2(n14142), .A(n15537), .B(n14141), .ZN(
        n14150) );
  MUX2_X1 U16182 ( .A(n11436), .B(P2_REG2_REG_4__SCAN_IN), .S(n14144), .Z(
        n14145) );
  NAND3_X1 U16183 ( .A1(n14147), .A2(n14146), .A3(n14145), .ZN(n14148) );
  NAND3_X1 U16184 ( .A1(n15546), .A2(n14161), .A3(n14148), .ZN(n14149) );
  NAND3_X1 U16185 ( .A1(n14151), .A2(n14150), .A3(n14149), .ZN(P2_U3218) );
  INV_X1 U16186 ( .A(n14152), .ZN(n14155) );
  NOR2_X1 U16187 ( .A1(n15543), .A2(n14153), .ZN(n14154) );
  AOI211_X1 U16188 ( .C1(n15525), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n14155), .B(
        n14154), .ZN(n14166) );
  OAI211_X1 U16189 ( .C1(n14158), .C2(n14157), .A(n15537), .B(n14156), .ZN(
        n14165) );
  MUX2_X1 U16190 ( .A(n11640), .B(P2_REG2_REG_5__SCAN_IN), .S(n14159), .Z(
        n14162) );
  NAND3_X1 U16191 ( .A1(n14162), .A2(n14161), .A3(n14160), .ZN(n14163) );
  NAND3_X1 U16192 ( .A1(n15546), .A2(n14174), .A3(n14163), .ZN(n14164) );
  NAND3_X1 U16193 ( .A1(n14166), .A2(n14165), .A3(n14164), .ZN(P2_U3219) );
  NOR2_X1 U16194 ( .A1(n15543), .A2(n14172), .ZN(n14167) );
  AOI211_X1 U16195 ( .C1(n15525), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n14168), .B(
        n14167), .ZN(n14180) );
  OAI211_X1 U16196 ( .C1(n14171), .C2(n14170), .A(n15537), .B(n14169), .ZN(
        n14179) );
  MUX2_X1 U16197 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11660), .S(n14172), .Z(
        n14175) );
  NAND3_X1 U16198 ( .A1(n14175), .A2(n14174), .A3(n14173), .ZN(n14176) );
  NAND3_X1 U16199 ( .A1(n15546), .A2(n14177), .A3(n14176), .ZN(n14178) );
  NAND3_X1 U16200 ( .A1(n14180), .A2(n14179), .A3(n14178), .ZN(P2_U3220) );
  INV_X1 U16201 ( .A(n14181), .ZN(n14183) );
  NOR2_X1 U16202 ( .A1(n15543), .A2(n14187), .ZN(n14182) );
  AOI211_X1 U16203 ( .C1(n15525), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n14183), .B(
        n14182), .ZN(n14194) );
  OAI211_X1 U16204 ( .C1(n14186), .C2(n14185), .A(n15537), .B(n14184), .ZN(
        n14193) );
  MUX2_X1 U16205 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11019), .S(n14187), .Z(
        n14188) );
  NAND3_X1 U16206 ( .A1(n15545), .A2(n14189), .A3(n14188), .ZN(n14190) );
  NAND3_X1 U16207 ( .A1(n15546), .A2(n14191), .A3(n14190), .ZN(n14192) );
  NAND3_X1 U16208 ( .A1(n14194), .A2(n14193), .A3(n14192), .ZN(P2_U3222) );
  OAI211_X1 U16209 ( .C1(n14197), .C2(n14196), .A(n14195), .B(n15537), .ZN(
        n14206) );
  NOR2_X1 U16210 ( .A1(n15543), .A2(n14198), .ZN(n14199) );
  AOI211_X1 U16211 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n15525), .A(n14200), 
        .B(n14199), .ZN(n14205) );
  OAI211_X1 U16212 ( .C1(n14203), .C2(n14202), .A(n14201), .B(n15546), .ZN(
        n14204) );
  NAND3_X1 U16213 ( .A1(n14206), .A2(n14205), .A3(n14204), .ZN(P2_U3224) );
  OAI211_X1 U16214 ( .C1(n14209), .C2(n14208), .A(n14207), .B(n15537), .ZN(
        n14218) );
  OAI21_X1 U16215 ( .B1(n15543), .B2(n14211), .A(n14210), .ZN(n14212) );
  AOI21_X1 U16216 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n15525), .A(n14212), 
        .ZN(n14217) );
  OAI211_X1 U16217 ( .C1(n14215), .C2(n14214), .A(n14213), .B(n15546), .ZN(
        n14216) );
  NAND3_X1 U16218 ( .A1(n14218), .A2(n14217), .A3(n14216), .ZN(P2_U3227) );
  INV_X1 U16219 ( .A(n14219), .ZN(n14220) );
  OAI21_X1 U16220 ( .B1(n15543), .B2(n14237), .A(n14220), .ZN(n14225) );
  XOR2_X1 U16221 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14237), .Z(n14222) );
  AOI211_X1 U16222 ( .C1(n14223), .C2(n14222), .A(n15529), .B(n14238), .ZN(
        n14224) );
  AOI211_X1 U16223 ( .C1(n15525), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n14225), 
        .B(n14224), .ZN(n14234) );
  MUX2_X1 U16224 ( .A(n14226), .B(P2_REG2_REG_16__SCAN_IN), .S(n14237), .Z(
        n14232) );
  NAND2_X1 U16225 ( .A1(n14227), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n14231) );
  NAND2_X1 U16226 ( .A1(n14229), .A2(n14228), .ZN(n14230) );
  NAND2_X1 U16227 ( .A1(n14234), .A2(n14233), .ZN(P2_U3230) );
  OAI21_X1 U16228 ( .B1(n15543), .B2(n14236), .A(n14235), .ZN(n14242) );
  INV_X1 U16229 ( .A(n14237), .ZN(n14243) );
  XNOR2_X1 U16230 ( .A(n14261), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14239) );
  AOI211_X1 U16231 ( .C1(n14240), .C2(n14239), .A(n15529), .B(n14260), .ZN(
        n14241) );
  AOI211_X1 U16232 ( .C1(n15525), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n14242), 
        .B(n14241), .ZN(n14252) );
  NAND2_X1 U16233 ( .A1(n14243), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14248) );
  NAND2_X1 U16234 ( .A1(n14249), .A2(n14248), .ZN(n14246) );
  MUX2_X1 U16235 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n14244), .S(n14261), .Z(
        n14245) );
  MUX2_X1 U16236 ( .A(n14244), .B(P2_REG2_REG_17__SCAN_IN), .S(n14261), .Z(
        n14247) );
  NAND3_X1 U16237 ( .A1(n14249), .A2(n14248), .A3(n14247), .ZN(n14250) );
  NAND3_X1 U16238 ( .A1(n14254), .A2(n15546), .A3(n14250), .ZN(n14251) );
  NAND2_X1 U16239 ( .A1(n14252), .A2(n14251), .ZN(P2_U3231) );
  NAND2_X1 U16240 ( .A1(n14261), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U16241 ( .A1(n14256), .A2(n14255), .ZN(n14257) );
  INV_X1 U16242 ( .A(n14275), .ZN(n14258) );
  AOI21_X1 U16243 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14259), .A(n14258), 
        .ZN(n14270) );
  NAND2_X1 U16244 ( .A1(n14262), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n14273) );
  OAI211_X1 U16245 ( .C1(n14262), .C2(P2_REG1_REG_18__SCAN_IN), .A(n14273), 
        .B(n15537), .ZN(n14268) );
  NOR2_X1 U16246 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14263), .ZN(n14266) );
  NOR2_X1 U16247 ( .A1(n15543), .A2(n14264), .ZN(n14265) );
  AOI211_X1 U16248 ( .C1(n15525), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n14266), 
        .B(n14265), .ZN(n14267) );
  OAI211_X1 U16249 ( .C1(n14270), .C2(n14269), .A(n14268), .B(n14267), .ZN(
        P2_U3232) );
  INV_X1 U16250 ( .A(n14271), .ZN(n14272) );
  INV_X1 U16251 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14565) );
  NAND2_X1 U16252 ( .A1(n14275), .A2(n14274), .ZN(n14276) );
  XNOR2_X1 U16253 ( .A(n14276), .B(n8281), .ZN(n14279) );
  INV_X1 U16254 ( .A(n14279), .ZN(n14277) );
  AOI22_X1 U16255 ( .A1(n14278), .A2(n15537), .B1(n15546), .B2(n14277), .ZN(
        n14281) );
  NAND2_X1 U16256 ( .A1(n14284), .A2(n14507), .ZN(n14287) );
  AOI21_X1 U16257 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n14490), .A(n14285), 
        .ZN(n14286) );
  OAI211_X1 U16258 ( .C1(n14288), .C2(n14455), .A(n14287), .B(n14286), .ZN(
        P2_U3234) );
  INV_X1 U16259 ( .A(n14292), .ZN(n14297) );
  AOI22_X1 U16260 ( .A1(n14293), .A2(n14511), .B1(n14473), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n14294) );
  OAI21_X1 U16261 ( .B1(n14295), .B2(n14492), .A(n14294), .ZN(n14296) );
  AOI21_X1 U16262 ( .B1(n14297), .B2(n14477), .A(n14296), .ZN(n14298) );
  XNOR2_X1 U16263 ( .A(n14299), .B(n14300), .ZN(n14302) );
  INV_X1 U16264 ( .A(n14303), .ZN(n14523) );
  NOR2_X1 U16265 ( .A1(n14306), .A2(n14305), .ZN(n14524) );
  OR3_X1 U16266 ( .A1(n14523), .A2(n14524), .A3(n14497), .ZN(n14315) );
  OAI22_X1 U16267 ( .A1(n14308), .A2(n14485), .B1(n14307), .B2(n14502), .ZN(
        n14309) );
  AOI21_X1 U16268 ( .B1(n14519), .B2(n14511), .A(n14309), .ZN(n14314) );
  OAI21_X1 U16269 ( .B1(n14321), .B2(n14310), .A(n14469), .ZN(n14312) );
  NOR2_X1 U16270 ( .A1(n14312), .A2(n14311), .ZN(n14521) );
  NAND2_X1 U16271 ( .A1(n14521), .A2(n14507), .ZN(n14313) );
  OAI21_X1 U16272 ( .B1(n14473), .B2(n14522), .A(n14316), .ZN(P2_U3238) );
  NAND2_X1 U16273 ( .A1(n14317), .A2(n14318), .ZN(n14319) );
  OAI21_X1 U16274 ( .B1(n14339), .B2(n14325), .A(n14469), .ZN(n14322) );
  NOR2_X1 U16275 ( .A1(n14322), .A2(n14321), .ZN(n14526) );
  AOI22_X1 U16276 ( .A1(n14323), .A2(n14510), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14490), .ZN(n14324) );
  OAI21_X1 U16277 ( .B1(n14325), .B2(n14455), .A(n14324), .ZN(n14329) );
  XNOR2_X1 U16278 ( .A(n14326), .B(n14327), .ZN(n14530) );
  NOR2_X1 U16279 ( .A1(n14530), .A2(n14497), .ZN(n14328) );
  AOI211_X1 U16280 ( .C1(n14526), .C2(n14507), .A(n14329), .B(n14328), .ZN(
        n14330) );
  OAI21_X1 U16281 ( .B1(n14473), .B2(n14529), .A(n14330), .ZN(P2_U3239) );
  XNOR2_X1 U16282 ( .A(n14332), .B(n14331), .ZN(n14531) );
  INV_X1 U16283 ( .A(n14531), .ZN(n14346) );
  OAI21_X1 U16284 ( .B1(n14333), .B2(n14332), .A(n14317), .ZN(n14334) );
  NAND2_X1 U16285 ( .A1(n14334), .A2(n14481), .ZN(n14336) );
  NAND2_X1 U16286 ( .A1(n14336), .A2(n14335), .ZN(n14533) );
  INV_X1 U16287 ( .A(n14629), .ZN(n14343) );
  NAND2_X1 U16288 ( .A1(n6561), .A2(n14629), .ZN(n14337) );
  NAND2_X1 U16289 ( .A1(n14337), .A2(n14469), .ZN(n14338) );
  NOR2_X1 U16290 ( .A1(n14339), .A2(n14338), .ZN(n14532) );
  NAND2_X1 U16291 ( .A1(n14532), .A2(n14507), .ZN(n14342) );
  AOI22_X1 U16292 ( .A1(n14340), .A2(n14510), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14490), .ZN(n14341) );
  OAI211_X1 U16293 ( .C1(n14343), .C2(n14455), .A(n14342), .B(n14341), .ZN(
        n14344) );
  AOI21_X1 U16294 ( .B1(n14533), .B2(n14502), .A(n14344), .ZN(n14345) );
  OAI21_X1 U16295 ( .B1(n14346), .B2(n14497), .A(n14345), .ZN(P2_U3240) );
  XNOR2_X1 U16296 ( .A(n14348), .B(n10081), .ZN(n14350) );
  AOI21_X1 U16297 ( .B1(n14350), .B2(n14481), .A(n14349), .ZN(n14538) );
  OAI21_X1 U16298 ( .B1(n6514), .B2(n10081), .A(n14351), .ZN(n14539) );
  OAI22_X1 U16299 ( .A1(n14353), .A2(n14485), .B1(n14352), .B2(n14502), .ZN(
        n14354) );
  AOI21_X1 U16300 ( .B1(n14536), .B2(n14511), .A(n14354), .ZN(n14357) );
  AOI21_X1 U16301 ( .B1(n14365), .B2(n14536), .A(n14486), .ZN(n14355) );
  AND2_X1 U16302 ( .A1(n6561), .A2(n14355), .ZN(n14535) );
  NAND2_X1 U16303 ( .A1(n14535), .A2(n14507), .ZN(n14356) );
  OAI211_X1 U16304 ( .C1(n14539), .C2(n14497), .A(n14357), .B(n14356), .ZN(
        n14358) );
  INV_X1 U16305 ( .A(n14358), .ZN(n14359) );
  OAI21_X1 U16306 ( .B1(n14490), .B2(n14538), .A(n14359), .ZN(P2_U3241) );
  XNOR2_X1 U16307 ( .A(n14360), .B(n14363), .ZN(n14362) );
  AOI21_X1 U16308 ( .B1(n14362), .B2(n14481), .A(n14361), .ZN(n14543) );
  XNOR2_X1 U16309 ( .A(n14364), .B(n14363), .ZN(n14544) );
  INV_X1 U16310 ( .A(n14544), .ZN(n14372) );
  AOI21_X1 U16311 ( .B1(n14382), .B2(n14541), .A(n14486), .ZN(n14366) );
  AND2_X1 U16312 ( .A1(n14366), .A2(n14365), .ZN(n14540) );
  NAND2_X1 U16313 ( .A1(n14540), .A2(n14507), .ZN(n14369) );
  AOI22_X1 U16314 ( .A1(n14367), .A2(n14510), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14490), .ZN(n14368) );
  OAI211_X1 U16315 ( .C1(n14370), .C2(n14455), .A(n14369), .B(n14368), .ZN(
        n14371) );
  AOI21_X1 U16316 ( .B1(n14372), .B2(n14477), .A(n14371), .ZN(n14373) );
  OAI21_X1 U16317 ( .B1(n14473), .B2(n14543), .A(n14373), .ZN(P2_U3242) );
  AOI21_X1 U16318 ( .B1(n14374), .B2(n10004), .A(n14443), .ZN(n14377) );
  AOI21_X1 U16319 ( .B1(n14377), .B2(n14376), .A(n14375), .ZN(n14546) );
  NAND2_X1 U16320 ( .A1(n14379), .A2(n14378), .ZN(n14380) );
  NAND2_X1 U16321 ( .A1(n14381), .A2(n14380), .ZN(n14547) );
  INV_X1 U16322 ( .A(n14547), .ZN(n14389) );
  OAI211_X1 U16323 ( .C1(n14397), .C2(n14383), .A(n14469), .B(n14382), .ZN(
        n14545) );
  INV_X1 U16324 ( .A(n14384), .ZN(n14385) );
  AOI22_X1 U16325 ( .A1(n14385), .A2(n14510), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n14490), .ZN(n14387) );
  NAND2_X1 U16326 ( .A1(n14634), .A2(n14511), .ZN(n14386) );
  OAI211_X1 U16327 ( .C1(n14545), .C2(n14492), .A(n14387), .B(n14386), .ZN(
        n14388) );
  AOI21_X1 U16328 ( .B1(n14389), .B2(n14477), .A(n14388), .ZN(n14390) );
  OAI21_X1 U16329 ( .B1(n14473), .B2(n14546), .A(n14390), .ZN(P2_U3243) );
  XNOR2_X1 U16330 ( .A(n14391), .B(n14394), .ZN(n14393) );
  AOI21_X1 U16331 ( .B1(n14393), .B2(n14481), .A(n14392), .ZN(n14552) );
  XNOR2_X1 U16332 ( .A(n14395), .B(n14394), .ZN(n14550) );
  OAI21_X1 U16333 ( .B1(n14396), .B2(n7763), .A(n14469), .ZN(n14398) );
  OR2_X1 U16334 ( .A1(n14398), .A2(n14397), .ZN(n14551) );
  AOI22_X1 U16335 ( .A1(n14473), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14399), 
        .B2(n14510), .ZN(n14401) );
  NAND2_X1 U16336 ( .A1(n14638), .A2(n14511), .ZN(n14400) );
  OAI211_X1 U16337 ( .C1(n14551), .C2(n14492), .A(n14401), .B(n14400), .ZN(
        n14402) );
  AOI21_X1 U16338 ( .B1(n14550), .B2(n14477), .A(n14402), .ZN(n14403) );
  OAI21_X1 U16339 ( .B1(n14473), .B2(n14552), .A(n14403), .ZN(P2_U3244) );
  NOR2_X1 U16340 ( .A1(n14425), .A2(n14424), .ZN(n14423) );
  NOR2_X1 U16341 ( .A1(n14423), .A2(n14404), .ZN(n14407) );
  INV_X1 U16342 ( .A(n14404), .ZN(n14405) );
  NAND2_X1 U16343 ( .A1(n14415), .A2(n14405), .ZN(n14406) );
  OAI22_X1 U16344 ( .A1(n14407), .A2(n14415), .B1(n14423), .B2(n14406), .ZN(
        n14409) );
  AOI21_X1 U16345 ( .B1(n14409), .B2(n14481), .A(n14408), .ZN(n14559) );
  AOI211_X1 U16346 ( .C1(n14557), .C2(n14432), .A(n14486), .B(n14396), .ZN(
        n14556) );
  INV_X1 U16347 ( .A(n14410), .ZN(n14411) );
  AOI22_X1 U16348 ( .A1(n14473), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14411), 
        .B2(n14510), .ZN(n14412) );
  OAI21_X1 U16349 ( .B1(n7058), .B2(n14455), .A(n14412), .ZN(n14418) );
  NAND2_X1 U16350 ( .A1(n14414), .A2(n14413), .ZN(n14416) );
  XOR2_X1 U16351 ( .A(n14416), .B(n14415), .Z(n14560) );
  NOR2_X1 U16352 ( .A1(n14560), .A2(n14497), .ZN(n14417) );
  AOI211_X1 U16353 ( .C1(n14556), .C2(n14507), .A(n14418), .B(n14417), .ZN(
        n14419) );
  OAI21_X1 U16354 ( .B1(n14473), .B2(n14559), .A(n14419), .ZN(P2_U3245) );
  NAND2_X1 U16355 ( .A1(n14446), .A2(n14421), .ZN(n14422) );
  XNOR2_X1 U16356 ( .A(n14422), .B(n14424), .ZN(n14563) );
  INV_X1 U16357 ( .A(n14563), .ZN(n14440) );
  AOI21_X1 U16358 ( .B1(n14425), .B2(n14424), .A(n14423), .ZN(n14430) );
  INV_X1 U16359 ( .A(n14426), .ZN(n14427) );
  NAND2_X1 U16360 ( .A1(n14563), .A2(n14427), .ZN(n14428) );
  OAI211_X1 U16361 ( .C1(n14430), .C2(n14443), .A(n14429), .B(n14428), .ZN(
        n14561) );
  NAND2_X1 U16362 ( .A1(n14561), .A2(n14502), .ZN(n14438) );
  AOI211_X1 U16363 ( .C1(n14433), .C2(n14431), .A(n7907), .B(n10040), .ZN(
        n14562) );
  AOI22_X1 U16364 ( .A1(n14473), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14434), 
        .B2(n14510), .ZN(n14435) );
  OAI21_X1 U16365 ( .B1(n14644), .B2(n14455), .A(n14435), .ZN(n14436) );
  AOI21_X1 U16366 ( .B1(n14562), .B2(n14507), .A(n14436), .ZN(n14437) );
  OAI211_X1 U16367 ( .C1(n14440), .C2(n14439), .A(n14438), .B(n14437), .ZN(
        P2_U3246) );
  XNOR2_X1 U16368 ( .A(n14441), .B(n14445), .ZN(n14444) );
  OAI21_X1 U16369 ( .B1(n14444), .B2(n14443), .A(n14442), .ZN(n14567) );
  INV_X1 U16370 ( .A(n14567), .ZN(n14458) );
  INV_X1 U16371 ( .A(n14420), .ZN(n14448) );
  INV_X1 U16372 ( .A(n14445), .ZN(n14447) );
  OAI21_X1 U16373 ( .B1(n14448), .B2(n14447), .A(n14446), .ZN(n14569) );
  INV_X1 U16374 ( .A(n14431), .ZN(n14449) );
  AOI211_X1 U16375 ( .C1(n14450), .C2(n7731), .A(n14486), .B(n14449), .ZN(
        n14568) );
  NAND2_X1 U16376 ( .A1(n14568), .A2(n14507), .ZN(n14454) );
  INV_X1 U16377 ( .A(n14451), .ZN(n14452) );
  AOI22_X1 U16378 ( .A1(n14473), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14452), 
        .B2(n14510), .ZN(n14453) );
  OAI211_X1 U16379 ( .C1(n14648), .C2(n14455), .A(n14454), .B(n14453), .ZN(
        n14456) );
  AOI21_X1 U16380 ( .B1(n14477), .B2(n14569), .A(n14456), .ZN(n14457) );
  OAI21_X1 U16381 ( .B1(n14473), .B2(n14458), .A(n14457), .ZN(P2_U3247) );
  XNOR2_X1 U16382 ( .A(n14459), .B(n14466), .ZN(n14461) );
  AOI21_X1 U16383 ( .B1(n14461), .B2(n14481), .A(n14460), .ZN(n14575) );
  INV_X1 U16384 ( .A(n14462), .ZN(n14463) );
  NAND2_X1 U16385 ( .A1(n14464), .A2(n14463), .ZN(n14494) );
  OR2_X1 U16386 ( .A1(n14494), .A2(n14493), .ZN(n14496) );
  NAND2_X1 U16387 ( .A1(n14496), .A2(n14465), .ZN(n14468) );
  INV_X1 U16388 ( .A(n14466), .ZN(n14467) );
  XNOR2_X1 U16389 ( .A(n14468), .B(n14467), .ZN(n14572) );
  NAND2_X1 U16390 ( .A1(n14488), .A2(n14651), .ZN(n14470) );
  NAND2_X1 U16391 ( .A1(n14470), .A2(n14469), .ZN(n14471) );
  OR2_X1 U16392 ( .A1(n14471), .A2(n7728), .ZN(n14573) );
  AOI22_X1 U16393 ( .A1(n14473), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14472), 
        .B2(n14510), .ZN(n14475) );
  NAND2_X1 U16394 ( .A1(n14651), .A2(n14511), .ZN(n14474) );
  OAI211_X1 U16395 ( .C1(n14573), .C2(n14492), .A(n14475), .B(n14474), .ZN(
        n14476) );
  AOI21_X1 U16396 ( .B1(n14572), .B2(n14477), .A(n14476), .ZN(n14478) );
  OAI21_X1 U16397 ( .B1(n14575), .B2(n14490), .A(n14478), .ZN(P2_U3248) );
  XNOR2_X1 U16398 ( .A(n14479), .B(n14480), .ZN(n14482) );
  NAND2_X1 U16399 ( .A1(n14482), .A2(n14481), .ZN(n14580) );
  INV_X1 U16400 ( .A(n14483), .ZN(n14578) );
  OAI211_X1 U16401 ( .C1(n14485), .C2(n14484), .A(n14580), .B(n14578), .ZN(
        n14500) );
  AOI21_X1 U16402 ( .B1(n14487), .B2(n14655), .A(n14486), .ZN(n14489) );
  NAND2_X1 U16403 ( .A1(n14489), .A2(n14488), .ZN(n14579) );
  AOI22_X1 U16404 ( .A1(n14655), .A2(n14511), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n14490), .ZN(n14491) );
  OAI21_X1 U16405 ( .B1(n14579), .B2(n14492), .A(n14491), .ZN(n14499) );
  NAND2_X1 U16406 ( .A1(n14494), .A2(n14493), .ZN(n14495) );
  NAND2_X1 U16407 ( .A1(n14496), .A2(n14495), .ZN(n14582) );
  NOR2_X1 U16408 ( .A1(n14582), .A2(n14497), .ZN(n14498) );
  AOI211_X1 U16409 ( .C1(n14502), .C2(n14500), .A(n14499), .B(n14498), .ZN(
        n14501) );
  INV_X1 U16410 ( .A(n14501), .ZN(P2_U3249) );
  MUX2_X1 U16411 ( .A(n14504), .B(n14503), .S(n14502), .Z(n14514) );
  INV_X1 U16412 ( .A(n14505), .ZN(n14508) );
  AOI22_X1 U16413 ( .A1(n14509), .A2(n14508), .B1(n14507), .B2(n14506), .ZN(
        n14513) );
  AOI22_X1 U16414 ( .A1(n14511), .A2(n7087), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n14510), .ZN(n14512) );
  NAND3_X1 U16415 ( .A1(n14514), .A2(n14513), .A3(n14512), .ZN(P2_U3264) );
  NOR3_X1 U16416 ( .A1(n14524), .A2(n14523), .A3(n15567), .ZN(n14525) );
  MUX2_X1 U16417 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14625), .S(n14618), .Z(
        P2_U3526) );
  AOI21_X1 U16418 ( .B1(n15564), .B2(n14527), .A(n14526), .ZN(n14528) );
  MUX2_X1 U16419 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14626), .S(n14618), .Z(
        P2_U3525) );
  MUX2_X1 U16420 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14627), .S(n14618), .Z(
        n14534) );
  AOI21_X1 U16421 ( .B1(n15564), .B2(n14536), .A(n14535), .ZN(n14537) );
  OAI211_X1 U16422 ( .C1(n14539), .C2(n15567), .A(n14538), .B(n14537), .ZN(
        n14630) );
  MUX2_X1 U16423 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14630), .S(n14618), .Z(
        P2_U3523) );
  AOI21_X1 U16424 ( .B1(n15564), .B2(n14541), .A(n14540), .ZN(n14542) );
  OAI211_X1 U16425 ( .C1(n14544), .C2(n15567), .A(n14543), .B(n14542), .ZN(
        n14631) );
  MUX2_X1 U16426 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14631), .S(n14618), .Z(
        P2_U3522) );
  OAI211_X1 U16427 ( .C1(n14547), .C2(n15567), .A(n14546), .B(n14545), .ZN(
        n14632) );
  MUX2_X1 U16428 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14632), .S(n14618), .Z(
        n14548) );
  AOI21_X1 U16429 ( .B1(n14584), .B2(n14634), .A(n14548), .ZN(n14549) );
  INV_X1 U16430 ( .A(n14549), .ZN(P2_U3521) );
  NAND2_X1 U16431 ( .A1(n14550), .A2(n14589), .ZN(n14553) );
  NAND3_X1 U16432 ( .A1(n14553), .A2(n14552), .A3(n14551), .ZN(n14636) );
  MUX2_X1 U16433 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14636), .S(n14618), .Z(
        n14554) );
  AOI21_X1 U16434 ( .B1(n14584), .B2(n14638), .A(n14554), .ZN(n14555) );
  INV_X1 U16435 ( .A(n14555), .ZN(P2_U3520) );
  AOI21_X1 U16436 ( .B1(n15564), .B2(n14557), .A(n14556), .ZN(n14558) );
  OAI211_X1 U16437 ( .C1(n15567), .C2(n14560), .A(n14559), .B(n14558), .ZN(
        n14640) );
  MUX2_X1 U16438 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14640), .S(n14618), .Z(
        P2_U3519) );
  AOI211_X1 U16439 ( .C1(n14564), .C2(n14563), .A(n14562), .B(n14561), .ZN(
        n14641) );
  MUX2_X1 U16440 ( .A(n14565), .B(n14641), .S(n14618), .Z(n14566) );
  OAI21_X1 U16441 ( .B1(n14644), .B2(n7043), .A(n14566), .ZN(P2_U3518) );
  INV_X1 U16442 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14570) );
  AOI211_X1 U16443 ( .C1(n14589), .C2(n14569), .A(n14568), .B(n14567), .ZN(
        n14645) );
  MUX2_X1 U16444 ( .A(n14570), .B(n14645), .S(n14618), .Z(n14571) );
  OAI21_X1 U16445 ( .B1(n14648), .B2(n7043), .A(n14571), .ZN(P2_U3517) );
  NAND2_X1 U16446 ( .A1(n14572), .A2(n14589), .ZN(n14574) );
  NAND3_X1 U16447 ( .A1(n14575), .A2(n14574), .A3(n14573), .ZN(n14649) );
  MUX2_X1 U16448 ( .A(n14649), .B(P2_REG1_REG_17__SCAN_IN), .S(n15573), .Z(
        n14576) );
  AOI21_X1 U16449 ( .B1(n14584), .B2(n14651), .A(n14576), .ZN(n14577) );
  INV_X1 U16450 ( .A(n14577), .ZN(P2_U3516) );
  AND2_X1 U16451 ( .A1(n14579), .A2(n14578), .ZN(n14581) );
  OAI211_X1 U16452 ( .C1(n14582), .C2(n15567), .A(n14581), .B(n14580), .ZN(
        n14653) );
  MUX2_X1 U16453 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14653), .S(n14618), .Z(
        n14583) );
  AOI21_X1 U16454 ( .B1(n14584), .B2(n14655), .A(n14583), .ZN(n14585) );
  INV_X1 U16455 ( .A(n14585), .ZN(P2_U3515) );
  AOI211_X1 U16456 ( .C1(n14589), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        n14657) );
  MUX2_X1 U16457 ( .A(n14590), .B(n14657), .S(n14618), .Z(n14591) );
  OAI21_X1 U16458 ( .B1(n10039), .B2(n7043), .A(n14591), .ZN(P2_U3514) );
  AOI211_X1 U16459 ( .C1(n15564), .C2(n14594), .A(n14593), .B(n14592), .ZN(
        n14595) );
  OAI21_X1 U16460 ( .B1(n15567), .B2(n14596), .A(n14595), .ZN(n14661) );
  MUX2_X1 U16461 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14661), .S(n14618), .Z(
        P2_U3512) );
  AOI211_X1 U16462 ( .C1(n15564), .C2(n14599), .A(n14598), .B(n14597), .ZN(
        n14601) );
  OAI211_X1 U16463 ( .C1(n15567), .C2(n14602), .A(n14601), .B(n14600), .ZN(
        n14662) );
  MUX2_X1 U16464 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14662), .S(n14618), .Z(
        P2_U3511) );
  AOI21_X1 U16465 ( .B1(n15564), .B2(n14604), .A(n14603), .ZN(n14605) );
  OAI211_X1 U16466 ( .C1(n15567), .C2(n14607), .A(n14606), .B(n14605), .ZN(
        n14663) );
  MUX2_X1 U16467 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14663), .S(n14618), .Z(
        P2_U3509) );
  AOI211_X1 U16468 ( .C1(n15564), .C2(n14610), .A(n14609), .B(n14608), .ZN(
        n14611) );
  OAI21_X1 U16469 ( .B1(n15567), .B2(n14612), .A(n14611), .ZN(n14664) );
  MUX2_X1 U16470 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14664), .S(n14618), .Z(
        P2_U3508) );
  AOI21_X1 U16471 ( .B1(n15564), .B2(n14614), .A(n14613), .ZN(n14616) );
  OAI211_X1 U16472 ( .C1(n15567), .C2(n14617), .A(n14616), .B(n14615), .ZN(
        n14665) );
  MUX2_X1 U16473 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n14665), .S(n14618), .Z(
        P2_U3506) );
  MUX2_X1 U16474 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n14619), .S(n14618), .Z(
        P2_U3499) );
  AOI21_X1 U16475 ( .B1(n10388), .B2(n14622), .A(n14621), .ZN(n14623) );
  INV_X1 U16476 ( .A(n14623), .ZN(P2_U3497) );
  MUX2_X1 U16477 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14625), .S(n15572), .Z(
        P2_U3494) );
  MUX2_X1 U16478 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14626), .S(n15572), .Z(
        P2_U3493) );
  MUX2_X1 U16479 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14627), .S(n15572), .Z(
        n14628) );
  MUX2_X1 U16480 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14630), .S(n15572), .Z(
        P2_U3491) );
  MUX2_X1 U16481 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14631), .S(n15572), .Z(
        P2_U3490) );
  MUX2_X1 U16482 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14632), .S(n15572), .Z(
        n14633) );
  AOI21_X1 U16483 ( .B1(n10388), .B2(n14634), .A(n14633), .ZN(n14635) );
  INV_X1 U16484 ( .A(n14635), .ZN(P2_U3489) );
  MUX2_X1 U16485 ( .A(n14636), .B(P2_REG0_REG_21__SCAN_IN), .S(n15570), .Z(
        n14637) );
  AOI21_X1 U16486 ( .B1(n10388), .B2(n14638), .A(n14637), .ZN(n14639) );
  INV_X1 U16487 ( .A(n14639), .ZN(P2_U3488) );
  MUX2_X1 U16488 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14640), .S(n15572), .Z(
        P2_U3487) );
  INV_X1 U16489 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14642) );
  MUX2_X1 U16490 ( .A(n14642), .B(n14641), .S(n15572), .Z(n14643) );
  OAI21_X1 U16491 ( .B1(n14644), .B2(n14660), .A(n14643), .ZN(P2_U3486) );
  INV_X1 U16492 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14646) );
  MUX2_X1 U16493 ( .A(n14646), .B(n14645), .S(n15572), .Z(n14647) );
  OAI21_X1 U16494 ( .B1(n14648), .B2(n14660), .A(n14647), .ZN(P2_U3484) );
  MUX2_X1 U16495 ( .A(n14649), .B(P2_REG0_REG_17__SCAN_IN), .S(n15570), .Z(
        n14650) );
  AOI21_X1 U16496 ( .B1(n10388), .B2(n14651), .A(n14650), .ZN(n14652) );
  INV_X1 U16497 ( .A(n14652), .ZN(P2_U3481) );
  MUX2_X1 U16498 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14653), .S(n15572), .Z(
        n14654) );
  AOI21_X1 U16499 ( .B1(n10388), .B2(n14655), .A(n14654), .ZN(n14656) );
  INV_X1 U16500 ( .A(n14656), .ZN(P2_U3478) );
  INV_X1 U16501 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14658) );
  MUX2_X1 U16502 ( .A(n14658), .B(n14657), .S(n15572), .Z(n14659) );
  OAI21_X1 U16503 ( .B1(n10039), .B2(n14660), .A(n14659), .ZN(P2_U3475) );
  MUX2_X1 U16504 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14661), .S(n15572), .Z(
        P2_U3469) );
  MUX2_X1 U16505 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14662), .S(n15572), .Z(
        P2_U3466) );
  MUX2_X1 U16506 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n14663), .S(n15572), .Z(
        P2_U3460) );
  MUX2_X1 U16507 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n14664), .S(n15572), .Z(
        P2_U3457) );
  MUX2_X1 U16508 ( .A(P2_REG0_REG_7__SCAN_IN), .B(n14665), .S(n15572), .Z(
        P2_U3451) );
  INV_X1 U16509 ( .A(n14666), .ZN(n15396) );
  NAND3_X1 U16510 ( .A1(n14668), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14670) );
  OAI22_X1 U16511 ( .A1(n14667), .A2(n14670), .B1(n14669), .B2(n14682), .ZN(
        n14671) );
  INV_X1 U16512 ( .A(n14671), .ZN(n14672) );
  OAI21_X1 U16513 ( .B1(n15396), .B2(n14673), .A(n14672), .ZN(P2_U3296) );
  OAI222_X1 U16514 ( .A1(n14685), .A2(n14676), .B1(P2_U3088), .B2(n14674), 
        .C1(n14675), .C2(n14682), .ZN(P2_U3297) );
  NAND2_X1 U16515 ( .A1(n14678), .A2(n14677), .ZN(n14680) );
  OAI211_X1 U16516 ( .C1(n14682), .C2(n14681), .A(n14680), .B(n14679), .ZN(
        P2_U3299) );
  OAI222_X1 U16517 ( .A1(n14682), .A2(n14686), .B1(n14685), .B2(n14684), .C1(
        n14683), .C2(P2_U3088), .ZN(P2_U3300) );
  MUX2_X1 U16518 ( .A(n14687), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U16519 ( .A(n14688), .ZN(n14689) );
  AOI21_X1 U16520 ( .B1(n14691), .B2(n14690), .A(n14689), .ZN(n14698) );
  INV_X1 U16521 ( .A(n14692), .ZN(n14695) );
  AOI21_X1 U16522 ( .B1(n14822), .B2(n15340), .A(n14693), .ZN(n14694) );
  OAI21_X1 U16523 ( .B1(n14695), .B2(n14824), .A(n14694), .ZN(n14696) );
  AOI21_X1 U16524 ( .B1(n15338), .B2(n10664), .A(n14696), .ZN(n14697) );
  OAI21_X1 U16525 ( .B1(n14698), .B2(n14826), .A(n14697), .ZN(P1_U3215) );
  XOR2_X1 U16526 ( .A(n14700), .B(n14699), .Z(n14705) );
  AOI22_X1 U16527 ( .A1(n14836), .A2(n15192), .B1(n15190), .B2(n14838), .ZN(
        n15061) );
  INV_X1 U16528 ( .A(n15064), .ZN(n14701) );
  AOI22_X1 U16529 ( .A1(n14701), .A2(n14810), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14702) );
  OAI21_X1 U16530 ( .B1(n15061), .B2(n14780), .A(n14702), .ZN(n14703) );
  AOI21_X1 U16531 ( .B1(n15282), .B2(n10664), .A(n14703), .ZN(n14704) );
  OAI21_X1 U16532 ( .B1(n14705), .B2(n14826), .A(n14704), .ZN(P1_U3216) );
  AOI21_X1 U16533 ( .B1(n14707), .B2(n14706), .A(n14826), .ZN(n14709) );
  NAND2_X1 U16534 ( .A1(n14709), .A2(n14708), .ZN(n14713) );
  NAND2_X1 U16535 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14970)
         );
  INV_X1 U16536 ( .A(n14970), .ZN(n14711) );
  OAI22_X1 U16537 ( .A1(n14804), .A2(n15169), .B1(n15089), .B2(n14815), .ZN(
        n14710) );
  AOI211_X1 U16538 ( .C1(n14810), .C2(n15129), .A(n14711), .B(n14710), .ZN(
        n14712) );
  OAI211_X1 U16539 ( .C1(n15132), .C2(n14808), .A(n14713), .B(n14712), .ZN(
        P1_U3219) );
  AOI22_X1 U16540 ( .A1(n14812), .A2(n10460), .B1(n9506), .B2(n10664), .ZN(
        n14722) );
  OAI21_X1 U16541 ( .B1(n14714), .B2(n14716), .A(n14715), .ZN(n14717) );
  NAND2_X1 U16542 ( .A1(n14717), .A2(n14801), .ZN(n14721) );
  AOI22_X1 U16543 ( .A1(n14719), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n14822), 
        .B2(n14718), .ZN(n14720) );
  NAND3_X1 U16544 ( .A1(n14722), .A2(n14721), .A3(n14720), .ZN(P1_U3222) );
  OR2_X1 U16545 ( .A1(n14724), .A2(n14725), .ZN(n14787) );
  INV_X1 U16546 ( .A(n14787), .ZN(n14723) );
  AOI21_X1 U16547 ( .B1(n14725), .B2(n14724), .A(n14723), .ZN(n14730) );
  OAI22_X1 U16548 ( .A1(n15097), .A2(n14824), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14726), .ZN(n14728) );
  OAI22_X1 U16549 ( .A1(n15090), .A2(n14815), .B1(n15089), .B2(n14804), .ZN(
        n14727) );
  AOI211_X1 U16550 ( .C1(n15099), .C2(n10664), .A(n14728), .B(n14727), .ZN(
        n14729) );
  OAI21_X1 U16551 ( .B1(n14730), .B2(n14826), .A(n14729), .ZN(P1_U3223) );
  XOR2_X1 U16552 ( .A(n14732), .B(n14731), .Z(n14737) );
  AOI22_X1 U16553 ( .A1(n14834), .A2(n15192), .B1(n15190), .B2(n14836), .ZN(
        n15269) );
  INV_X1 U16554 ( .A(n14733), .ZN(n15036) );
  AOI22_X1 U16555 ( .A1(n15036), .A2(n14810), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14734) );
  OAI21_X1 U16556 ( .B1(n15269), .B2(n14780), .A(n14734), .ZN(n14735) );
  AOI21_X1 U16557 ( .B1(n15035), .B2(n10664), .A(n14735), .ZN(n14736) );
  OAI21_X1 U16558 ( .B1(n14737), .B2(n14826), .A(n14736), .ZN(P1_U3225) );
  XNOR2_X1 U16559 ( .A(n14739), .B(n14738), .ZN(n14744) );
  INV_X1 U16560 ( .A(n14740), .ZN(n14742) );
  XOR2_X1 U16561 ( .A(n14741), .B(n14740), .Z(n14827) );
  NOR2_X1 U16562 ( .A1(n14827), .A2(n14828), .ZN(n14825) );
  AOI21_X1 U16563 ( .B1(n14742), .B2(n14741), .A(n14825), .ZN(n14743) );
  NAND2_X1 U16564 ( .A1(n14743), .A2(n14744), .ZN(n14755) );
  OAI21_X1 U16565 ( .B1(n14744), .B2(n14743), .A(n14755), .ZN(n14745) );
  NAND2_X1 U16566 ( .A1(n14745), .A2(n14801), .ZN(n14750) );
  OAI22_X1 U16567 ( .A1(n14804), .A2(n14746), .B1(n15142), .B2(n14815), .ZN(
        n14747) );
  AOI211_X1 U16568 ( .C1(n14810), .C2(n15194), .A(n14748), .B(n14747), .ZN(
        n14749) );
  OAI211_X1 U16569 ( .C1(n15325), .C2(n14808), .A(n14750), .B(n14749), .ZN(
        P1_U3226) );
  AOI22_X1 U16570 ( .A1(n14751), .A2(n15125), .B1(n14812), .B2(n14840), .ZN(
        n14752) );
  NAND2_X1 U16571 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14932)
         );
  OAI211_X1 U16572 ( .C1(n14824), .C2(n15160), .A(n14752), .B(n14932), .ZN(
        n14759) );
  NAND3_X1 U16573 ( .A1(n14755), .A2(n14754), .A3(n14753), .ZN(n14757) );
  AOI21_X1 U16574 ( .B1(n14757), .B2(n14756), .A(n14826), .ZN(n14758) );
  AOI211_X1 U16575 ( .C1(n15319), .C2(n10664), .A(n14759), .B(n14758), .ZN(
        n14760) );
  INV_X1 U16576 ( .A(n14760), .ZN(P1_U3228) );
  XOR2_X1 U16577 ( .A(n14762), .B(n14761), .Z(n14767) );
  AOI22_X1 U16578 ( .A1(n15050), .A2(n14810), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14764) );
  NAND2_X1 U16579 ( .A1(n14837), .A2(n14812), .ZN(n14763) );
  OAI211_X1 U16580 ( .C1(n15045), .C2(n14815), .A(n14764), .B(n14763), .ZN(
        n14765) );
  AOI21_X1 U16581 ( .B1(n15049), .B2(n10664), .A(n14765), .ZN(n14766) );
  OAI21_X1 U16582 ( .B1(n14767), .B2(n14826), .A(n14766), .ZN(P1_U3229) );
  OAI211_X1 U16583 ( .C1(n14768), .C2(n14770), .A(n14769), .B(n14801), .ZN(
        n14774) );
  AOI22_X1 U16584 ( .A1(n15069), .A2(n15192), .B1(n15190), .B2(n14839), .ZN(
        n15299) );
  OAI22_X1 U16585 ( .A1(n15299), .A2(n14780), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14771), .ZN(n14772) );
  AOI21_X1 U16586 ( .B1(n15108), .B2(n14810), .A(n14772), .ZN(n14773) );
  OAI211_X1 U16587 ( .C1(n15375), .C2(n14808), .A(n14774), .B(n14773), .ZN(
        P1_U3233) );
  OAI211_X1 U16588 ( .C1(n14777), .C2(n14776), .A(n14775), .B(n14801), .ZN(
        n14784) );
  OAI21_X1 U16589 ( .B1(n14780), .B2(n14779), .A(n14778), .ZN(n14781) );
  AOI21_X1 U16590 ( .B1(n14782), .B2(n14810), .A(n14781), .ZN(n14783) );
  OAI211_X1 U16591 ( .C1(n14785), .C2(n14808), .A(n14784), .B(n14783), .ZN(
        P1_U3234) );
  NAND2_X1 U16592 ( .A1(n14787), .A2(n14786), .ZN(n14789) );
  OAI21_X1 U16593 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n14791) );
  NAND2_X1 U16594 ( .A1(n14791), .A2(n14801), .ZN(n14798) );
  NOR2_X1 U16595 ( .A1(n14792), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14793) );
  AOI21_X1 U16596 ( .B1(n15079), .B2(n14810), .A(n14793), .ZN(n14795) );
  NAND2_X1 U16597 ( .A1(n15069), .A2(n14812), .ZN(n14794) );
  OAI211_X1 U16598 ( .C1(n15072), .C2(n14815), .A(n14795), .B(n14794), .ZN(
        n14796) );
  AOI21_X1 U16599 ( .B1(n15078), .B2(n10664), .A(n14796), .ZN(n14797) );
  NAND2_X1 U16600 ( .A1(n14798), .A2(n14797), .ZN(P1_U3235) );
  INV_X1 U16601 ( .A(n15149), .ZN(n15380) );
  XNOR2_X1 U16602 ( .A(n14800), .B(n14799), .ZN(n14802) );
  NAND2_X1 U16603 ( .A1(n14802), .A2(n14801), .ZN(n14807) );
  NOR2_X1 U16604 ( .A1(n14803), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14944) );
  OAI22_X1 U16605 ( .A1(n14804), .A2(n15142), .B1(n15143), .B2(n14815), .ZN(
        n14805) );
  AOI211_X1 U16606 ( .C1(n14810), .C2(n15150), .A(n14944), .B(n14805), .ZN(
        n14806) );
  OAI211_X1 U16607 ( .C1(n15380), .C2(n14808), .A(n14807), .B(n14806), .ZN(
        P1_U3238) );
  AOI22_X1 U16608 ( .A1(n14811), .A2(n14810), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14814) );
  NAND2_X1 U16609 ( .A1(n14835), .A2(n14812), .ZN(n14813) );
  OAI211_X1 U16610 ( .C1(n14816), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        n14817) );
  AOI21_X1 U16611 ( .B1(n15264), .B2(n10664), .A(n14817), .ZN(n14818) );
  OAI21_X1 U16612 ( .B1(n14819), .B2(n14826), .A(n14818), .ZN(P1_U3240) );
  OAI22_X1 U16613 ( .A1(n15167), .A2(n15168), .B1(n14820), .B2(n15166), .ZN(
        n15221) );
  AOI21_X1 U16614 ( .B1(n15221), .B2(n14822), .A(n14821), .ZN(n14823) );
  OAI21_X1 U16615 ( .B1(n15209), .B2(n14824), .A(n14823), .ZN(n14830) );
  AOI211_X1 U16616 ( .C1(n14828), .C2(n14827), .A(n14826), .B(n14825), .ZN(
        n14829) );
  AOI211_X1 U16617 ( .C1(n15213), .C2(n10664), .A(n14830), .B(n14829), .ZN(
        n14831) );
  INV_X1 U16618 ( .A(n14831), .ZN(P1_U3241) );
  MUX2_X1 U16619 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14832), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16620 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15242), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16621 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15243), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16622 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14833), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16623 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14834), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16624 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14835), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16625 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14836), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16626 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14837), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16627 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14838), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16628 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15069), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16629 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15126), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16630 ( .A(n14839), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14854), .Z(
        P1_U3579) );
  MUX2_X1 U16631 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15125), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16632 ( .A(n15193), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14854), .Z(
        P1_U3577) );
  MUX2_X1 U16633 ( .A(n14840), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14854), .Z(
        P1_U3576) );
  MUX2_X1 U16634 ( .A(n15191), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14854), .Z(
        P1_U3575) );
  MUX2_X1 U16635 ( .A(n14841), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14854), .Z(
        P1_U3574) );
  MUX2_X1 U16636 ( .A(n14842), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14854), .Z(
        P1_U3573) );
  MUX2_X1 U16637 ( .A(n14843), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14854), .Z(
        P1_U3572) );
  MUX2_X1 U16638 ( .A(n14844), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14854), .Z(
        P1_U3571) );
  MUX2_X1 U16639 ( .A(n14845), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14854), .Z(
        P1_U3570) );
  MUX2_X1 U16640 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14846), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16641 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14847), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16642 ( .A(n14848), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14854), .Z(
        P1_U3567) );
  MUX2_X1 U16643 ( .A(n14849), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14854), .Z(
        P1_U3566) );
  MUX2_X1 U16644 ( .A(n14850), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14854), .Z(
        P1_U3565) );
  MUX2_X1 U16645 ( .A(n14851), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14854), .Z(
        P1_U3564) );
  MUX2_X1 U16646 ( .A(n14852), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14854), .Z(
        P1_U3563) );
  MUX2_X1 U16647 ( .A(n14853), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14854), .Z(
        P1_U3562) );
  MUX2_X1 U16648 ( .A(n14855), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14854), .Z(
        P1_U3561) );
  MUX2_X1 U16649 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10460), .S(P1_U4016), .Z(
        P1_U3560) );
  INV_X1 U16650 ( .A(n14856), .ZN(n14871) );
  INV_X1 U16651 ( .A(n14883), .ZN(n14861) );
  NOR3_X1 U16652 ( .A1(n14859), .A2(n14858), .A3(n14857), .ZN(n14860) );
  NOR3_X1 U16653 ( .A1(n14960), .A2(n14861), .A3(n14860), .ZN(n14862) );
  AOI211_X1 U16654 ( .C1(n14945), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n14863), .B(
        n14862), .ZN(n14870) );
  AOI211_X1 U16655 ( .C1(n14866), .C2(n14865), .A(n14940), .B(n14864), .ZN(
        n14867) );
  AOI21_X1 U16656 ( .B1(n14902), .B2(n14868), .A(n14867), .ZN(n14869) );
  NAND3_X1 U16657 ( .A1(n14871), .A2(n14870), .A3(n14869), .ZN(P1_U3247) );
  OAI21_X1 U16658 ( .B1(n14874), .B2(n14873), .A(n14872), .ZN(n14875) );
  NAND2_X1 U16659 ( .A1(n14875), .A2(n14965), .ZN(n14888) );
  OAI21_X1 U16660 ( .B1(n14972), .B2(n14877), .A(n14876), .ZN(n14878) );
  AOI21_X1 U16661 ( .B1(n14902), .B2(n14879), .A(n14878), .ZN(n14887) );
  INV_X1 U16662 ( .A(n14880), .ZN(n14885) );
  NAND3_X1 U16663 ( .A1(n14883), .A2(n14882), .A3(n14881), .ZN(n14884) );
  NAND3_X1 U16664 ( .A1(n14964), .A2(n14885), .A3(n14884), .ZN(n14886) );
  NAND3_X1 U16665 ( .A1(n14888), .A2(n14887), .A3(n14886), .ZN(P1_U3248) );
  OAI21_X1 U16666 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n14892) );
  NAND2_X1 U16667 ( .A1(n14892), .A2(n14965), .ZN(n14906) );
  INV_X1 U16668 ( .A(n14893), .ZN(n14894) );
  AOI21_X1 U16669 ( .B1(n14945), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n14894), .ZN(
        n14905) );
  MUX2_X1 U16670 ( .A(n11960), .B(P1_REG2_REG_8__SCAN_IN), .S(n14901), .Z(
        n14897) );
  INV_X1 U16671 ( .A(n14895), .ZN(n14896) );
  NAND2_X1 U16672 ( .A1(n14897), .A2(n14896), .ZN(n14899) );
  OAI211_X1 U16673 ( .C1(n14900), .C2(n14899), .A(n14898), .B(n14964), .ZN(
        n14904) );
  NAND2_X1 U16674 ( .A1(n14902), .A2(n14901), .ZN(n14903) );
  NAND4_X1 U16675 ( .A1(n14906), .A2(n14905), .A3(n14904), .A4(n14903), .ZN(
        P1_U3251) );
  OAI211_X1 U16676 ( .C1(n14909), .C2(n14908), .A(n14907), .B(n14965), .ZN(
        n14920) );
  NOR2_X1 U16677 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9629), .ZN(n14912) );
  NOR2_X1 U16678 ( .A1(n14959), .A2(n14910), .ZN(n14911) );
  AOI211_X1 U16679 ( .C1(n14945), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n14912), 
        .B(n14911), .ZN(n14919) );
  OR3_X1 U16680 ( .A1(n14915), .A2(n14914), .A3(n14913), .ZN(n14916) );
  NAND3_X1 U16681 ( .A1(n14917), .A2(n14964), .A3(n14916), .ZN(n14918) );
  NAND3_X1 U16682 ( .A1(n14920), .A2(n14919), .A3(n14918), .ZN(P1_U3253) );
  AOI21_X1 U16683 ( .B1(n14922), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14921), 
        .ZN(n14924) );
  XNOR2_X1 U16684 ( .A(n14939), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14923) );
  NOR2_X1 U16685 ( .A1(n14924), .A2(n14923), .ZN(n14938) );
  AOI211_X1 U16686 ( .C1(n14924), .C2(n14923), .A(n14938), .B(n14940), .ZN(
        n14937) );
  INV_X1 U16687 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14926) );
  NOR2_X1 U16688 ( .A1(n14947), .A2(n14928), .ZN(n14929) );
  AOI21_X1 U16689 ( .B1(n14928), .B2(n14947), .A(n14929), .ZN(n14930) );
  OAI211_X1 U16690 ( .C1(n14931), .C2(n14930), .A(n14964), .B(n14946), .ZN(
        n14935) );
  INV_X1 U16691 ( .A(n14932), .ZN(n14933) );
  AOI21_X1 U16692 ( .B1(n14945), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14933), 
        .ZN(n14934) );
  OAI211_X1 U16693 ( .C1(n14959), .C2(n14947), .A(n14935), .B(n14934), .ZN(
        n14936) );
  OR2_X1 U16694 ( .A1(n14937), .A2(n14936), .ZN(P1_U3260) );
  AOI211_X1 U16695 ( .C1(n14941), .C2(n15316), .A(n14953), .B(n14940), .ZN(
        n14942) );
  INV_X1 U16696 ( .A(n14942), .ZN(n14951) );
  NOR2_X1 U16697 ( .A1(n14959), .A2(n14952), .ZN(n14943) );
  AOI211_X1 U16698 ( .C1(P1_ADDR_REG_18__SCAN_IN), .C2(n14945), .A(n14944), 
        .B(n14943), .ZN(n14950) );
  OAI21_X1 U16699 ( .B1(n14928), .B2(n14947), .A(n14946), .ZN(n14955) );
  OAI211_X1 U16700 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14948), .A(n14964), 
        .B(n14958), .ZN(n14949) );
  NAND3_X1 U16701 ( .A1(n14951), .A2(n14950), .A3(n14949), .ZN(P1_U3261) );
  INV_X1 U16702 ( .A(n14966), .ZN(n14962) );
  NAND2_X1 U16703 ( .A1(n14956), .A2(n14955), .ZN(n14957) );
  OAI21_X1 U16704 ( .B1(n14963), .B2(n14960), .A(n14959), .ZN(n14961) );
  AOI21_X1 U16705 ( .B1(n14962), .B2(n14965), .A(n14961), .ZN(n14969) );
  AOI22_X1 U16706 ( .A1(n14966), .A2(n14965), .B1(n14964), .B2(n14963), .ZN(
        n14968) );
  OAI211_X1 U16707 ( .C1(n7813), .C2(n14972), .A(n14971), .B(n14970), .ZN(
        P1_U3262) );
  NAND2_X1 U16708 ( .A1(n14973), .A2(n15175), .ZN(n14976) );
  INV_X1 U16709 ( .A(n14974), .ZN(n15230) );
  NOR2_X1 U16710 ( .A1(n15484), .A2(n15230), .ZN(n14979) );
  AOI21_X1 U16711 ( .B1(n15484), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14979), 
        .ZN(n14975) );
  OAI211_X1 U16712 ( .C1(n15229), .C2(n15196), .A(n14976), .B(n14975), .ZN(
        P1_U3263) );
  OAI211_X1 U16713 ( .C1(n14984), .C2(n15357), .A(n15283), .B(n14977), .ZN(
        n15231) );
  NOR2_X1 U16714 ( .A1(n15482), .A2(n14978), .ZN(n14980) );
  AOI211_X1 U16715 ( .C1(n10333), .C2(n15212), .A(n14980), .B(n14979), .ZN(
        n14981) );
  OAI21_X1 U16716 ( .B1(n15231), .B2(n15215), .A(n14981), .ZN(P1_U3264) );
  NAND2_X1 U16717 ( .A1(n15482), .A2(n15327), .ZN(n15477) );
  AOI211_X1 U16718 ( .C1(n14985), .C2(n15246), .A(n15187), .B(n14984), .ZN(
        n15251) );
  NOR2_X1 U16719 ( .A1(n14986), .A2(n15196), .ZN(n14996) );
  NAND2_X1 U16720 ( .A1(n15243), .A2(n15190), .ZN(n15238) );
  OR2_X1 U16721 ( .A1(n14988), .A2(n14987), .ZN(n15239) );
  NOR2_X1 U16722 ( .A1(n14989), .A2(n15239), .ZN(n14990) );
  AOI21_X1 U16723 ( .B1(n15484), .B2(P1_REG2_REG_29__SCAN_IN), .A(n14990), 
        .ZN(n14994) );
  INV_X1 U16724 ( .A(n14991), .ZN(n14992) );
  NAND3_X1 U16725 ( .A1(n14992), .A2(n15480), .A3(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n14993) );
  OAI211_X1 U16726 ( .C1(n15238), .C2(n15484), .A(n14994), .B(n14993), .ZN(
        n14995) );
  AOI211_X1 U16727 ( .C1(n15251), .C2(n15175), .A(n14996), .B(n14995), .ZN(
        n15002) );
  INV_X1 U16728 ( .A(n15253), .ZN(n14998) );
  NOR2_X1 U16729 ( .A1(n14997), .A2(n15013), .ZN(n15234) );
  XNOR2_X1 U16730 ( .A(n14999), .B(n15252), .ZN(n15000) );
  NAND2_X1 U16731 ( .A1(n15000), .A2(n15224), .ZN(n15001) );
  OAI211_X1 U16732 ( .C1(n15254), .C2(n15477), .A(n15002), .B(n15001), .ZN(
        P1_U3356) );
  INV_X1 U16733 ( .A(n15003), .ZN(n15007) );
  NAND3_X1 U16734 ( .A1(n15005), .A2(n15010), .A3(n15004), .ZN(n15006) );
  AOI21_X1 U16735 ( .B1(n15007), .B2(n15006), .A(n15300), .ZN(n15008) );
  OAI22_X1 U16736 ( .A1(n15013), .A2(n15168), .B1(n15012), .B2(n15166), .ZN(
        n15014) );
  INV_X1 U16737 ( .A(n12877), .ZN(n15019) );
  AOI211_X1 U16738 ( .C1(n15258), .C2(n15019), .A(n15187), .B(n15018), .ZN(
        n15257) );
  NAND2_X1 U16739 ( .A1(n15257), .A2(n15175), .ZN(n15022) );
  AOI22_X1 U16740 ( .A1(n15020), .A2(n15480), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15484), .ZN(n15021) );
  OAI211_X1 U16741 ( .C1(n15023), .C2(n15196), .A(n15022), .B(n15021), .ZN(
        n15024) );
  AOI21_X1 U16742 ( .B1(n15255), .B2(n15025), .A(n15024), .ZN(n15026) );
  OAI21_X1 U16743 ( .B1(n15263), .B2(n15484), .A(n15026), .ZN(P1_U3266) );
  INV_X1 U16744 ( .A(n12864), .ZN(n15030) );
  INV_X1 U16745 ( .A(n15027), .ZN(n15028) );
  OAI21_X1 U16746 ( .B1(n15030), .B2(n15029), .A(n15028), .ZN(n15275) );
  OAI21_X1 U16747 ( .B1(n15033), .B2(n15032), .A(n15031), .ZN(n15273) );
  INV_X1 U16748 ( .A(n15477), .ZN(n15201) );
  NAND2_X1 U16749 ( .A1(n15273), .A2(n15201), .ZN(n15041) );
  AOI211_X1 U16750 ( .C1(n15035), .C2(n15047), .A(n15187), .B(n15034), .ZN(
        n15272) );
  NOR2_X1 U16751 ( .A1(n15270), .A2(n15196), .ZN(n15039) );
  AOI22_X1 U16752 ( .A1(n15036), .A2(n15480), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15484), .ZN(n15037) );
  OAI21_X1 U16753 ( .B1(n15269), .B2(n15484), .A(n15037), .ZN(n15038) );
  AOI211_X1 U16754 ( .C1(n15272), .C2(n15175), .A(n15039), .B(n15038), .ZN(
        n15040) );
  OAI211_X1 U16755 ( .C1(n15275), .C2(n15478), .A(n15041), .B(n15040), .ZN(
        P1_U3268) );
  XNOR2_X1 U16756 ( .A(n15043), .B(n15042), .ZN(n15278) );
  INV_X1 U16757 ( .A(n15278), .ZN(n15055) );
  OAI22_X1 U16758 ( .A1(n15045), .A2(n15168), .B1(n15072), .B2(n15166), .ZN(
        n15046) );
  INV_X1 U16759 ( .A(n15047), .ZN(n15048) );
  AOI211_X1 U16760 ( .C1(n15049), .C2(n15063), .A(n15187), .B(n15048), .ZN(
        n15277) );
  NAND2_X1 U16761 ( .A1(n15277), .A2(n15175), .ZN(n15052) );
  AOI22_X1 U16762 ( .A1(n15050), .A2(n15480), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15484), .ZN(n15051) );
  OAI211_X1 U16763 ( .C1(n15365), .C2(n15196), .A(n15052), .B(n15051), .ZN(
        n15053) );
  AOI21_X1 U16764 ( .B1(n15276), .B2(n15482), .A(n15053), .ZN(n15054) );
  OAI21_X1 U16765 ( .B1(n15055), .B2(n15478), .A(n15054), .ZN(P1_U3269) );
  OAI21_X1 U16766 ( .B1(n15057), .B2(n15059), .A(n15056), .ZN(n15287) );
  AOI21_X1 U16767 ( .B1(n15060), .B2(n15059), .A(n15058), .ZN(n15062) );
  OAI21_X1 U16768 ( .B1(n15062), .B2(n15300), .A(n15061), .ZN(n15281) );
  AOI21_X1 U16769 ( .B1(n15282), .B2(n6723), .A(n7077), .ZN(n15284) );
  INV_X1 U16770 ( .A(n15284), .ZN(n15065) );
  OAI22_X1 U16771 ( .A1(n15065), .A2(n12878), .B1(n15064), .B2(n15208), .ZN(
        n15066) );
  OAI21_X1 U16772 ( .B1(n15281), .B2(n15066), .A(n15482), .ZN(n15068) );
  AOI22_X1 U16773 ( .A1(n15282), .A2(n15212), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15484), .ZN(n15067) );
  OAI211_X1 U16774 ( .C1(n15287), .C2(n15478), .A(n15068), .B(n15067), .ZN(
        P1_U3270) );
  INV_X1 U16775 ( .A(n15069), .ZN(n15073) );
  XNOR2_X1 U16776 ( .A(n15070), .B(n15075), .ZN(n15071) );
  OAI222_X1 U16777 ( .A1(n15166), .A2(n15073), .B1(n15168), .B2(n15072), .C1(
        n15300), .C2(n15071), .ZN(n15288) );
  INV_X1 U16778 ( .A(n15288), .ZN(n15084) );
  OAI21_X1 U16779 ( .B1(n15076), .B2(n15075), .A(n15074), .ZN(n15290) );
  AOI211_X1 U16780 ( .C1(n15078), .C2(n15094), .A(n15187), .B(n15077), .ZN(
        n15289) );
  NAND2_X1 U16781 ( .A1(n15289), .A2(n15175), .ZN(n15081) );
  AOI22_X1 U16782 ( .A1(n15079), .A2(n15480), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15484), .ZN(n15080) );
  OAI211_X1 U16783 ( .C1(n15196), .C2(n15370), .A(n15081), .B(n15080), .ZN(
        n15082) );
  AOI21_X1 U16784 ( .B1(n15290), .B2(n15224), .A(n15082), .ZN(n15083) );
  OAI21_X1 U16785 ( .B1(n15084), .B2(n15484), .A(n15083), .ZN(P1_U3271) );
  XNOR2_X1 U16786 ( .A(n15085), .B(n15086), .ZN(n15293) );
  INV_X1 U16787 ( .A(n15293), .ZN(n15103) );
  XNOR2_X1 U16788 ( .A(n15087), .B(n7414), .ZN(n15088) );
  NAND2_X1 U16789 ( .A1(n15088), .A2(n15327), .ZN(n15093) );
  OAI22_X1 U16790 ( .A1(n15090), .A2(n15168), .B1(n15089), .B2(n15166), .ZN(
        n15091) );
  INV_X1 U16791 ( .A(n15091), .ZN(n15092) );
  NAND2_X1 U16792 ( .A1(n15093), .A2(n15092), .ZN(n15296) );
  AOI21_X1 U16793 ( .B1(n15111), .B2(n15099), .A(n15187), .ZN(n15095) );
  NAND2_X1 U16794 ( .A1(n15095), .A2(n15094), .ZN(n15294) );
  INV_X1 U16795 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n15096) );
  OAI22_X1 U16796 ( .A1(n15097), .A2(n15208), .B1(n15096), .B2(n15482), .ZN(
        n15098) );
  AOI21_X1 U16797 ( .B1(n15099), .B2(n15212), .A(n15098), .ZN(n15100) );
  OAI21_X1 U16798 ( .B1(n15294), .B2(n15215), .A(n15100), .ZN(n15101) );
  AOI21_X1 U16799 ( .B1(n15296), .B2(n15482), .A(n15101), .ZN(n15102) );
  OAI21_X1 U16800 ( .B1(n15103), .B2(n15478), .A(n15102), .ZN(P1_U3272) );
  XNOR2_X1 U16801 ( .A(n15105), .B(n15104), .ZN(n15301) );
  AOI21_X1 U16802 ( .B1(n15107), .B2(n15106), .A(n6503), .ZN(n15303) );
  NAND2_X1 U16803 ( .A1(n15303), .A2(n15224), .ZN(n15117) );
  AOI22_X1 U16804 ( .A1(n15484), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n15108), 
        .B2(n15480), .ZN(n15109) );
  OAI21_X1 U16805 ( .B1(n15299), .B2(n15484), .A(n15109), .ZN(n15114) );
  INV_X1 U16806 ( .A(n15110), .ZN(n15112) );
  OAI211_X1 U16807 ( .C1(n15112), .C2(n15375), .A(n15283), .B(n15111), .ZN(
        n15298) );
  NOR2_X1 U16808 ( .A1(n15298), .A2(n15215), .ZN(n15113) );
  AOI211_X1 U16809 ( .C1(n15212), .C2(n15115), .A(n15114), .B(n15113), .ZN(
        n15116) );
  OAI211_X1 U16810 ( .C1(n15301), .C2(n15477), .A(n15117), .B(n15116), .ZN(
        P1_U3273) );
  XOR2_X1 U16811 ( .A(n7051), .B(n15123), .Z(n15310) );
  INV_X1 U16812 ( .A(n15119), .ZN(n15120) );
  NAND2_X1 U16813 ( .A1(n15172), .A2(n15120), .ZN(n15141) );
  AOI21_X1 U16814 ( .B1(n15141), .B2(n15138), .A(n15121), .ZN(n15124) );
  OAI21_X1 U16815 ( .B1(n15124), .B2(n15123), .A(n15122), .ZN(n15127) );
  AOI222_X1 U16816 ( .A1(n15327), .A2(n15127), .B1(n15126), .B2(n15192), .C1(
        n15125), .C2(n15190), .ZN(n15309) );
  INV_X1 U16817 ( .A(n15309), .ZN(n15134) );
  OR2_X1 U16818 ( .A1(n15132), .A2(n15148), .ZN(n15128) );
  AND3_X1 U16819 ( .A1(n15110), .A2(n15128), .A3(n15283), .ZN(n15306) );
  NAND2_X1 U16820 ( .A1(n15306), .A2(n15175), .ZN(n15131) );
  AOI22_X1 U16821 ( .A1(n15484), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n15129), 
        .B2(n15480), .ZN(n15130) );
  OAI211_X1 U16822 ( .C1(n15132), .C2(n15196), .A(n15131), .B(n15130), .ZN(
        n15133) );
  AOI21_X1 U16823 ( .B1(n15134), .B2(n15482), .A(n15133), .ZN(n15135) );
  OAI21_X1 U16824 ( .B1(n15310), .B2(n15478), .A(n15135), .ZN(P1_U3274) );
  NAND2_X1 U16825 ( .A1(n15137), .A2(n15136), .ZN(n15139) );
  XNOR2_X1 U16826 ( .A(n15139), .B(n15138), .ZN(n15311) );
  XNOR2_X1 U16827 ( .A(n15141), .B(n15140), .ZN(n15145) );
  OAI22_X1 U16828 ( .A1(n15143), .A2(n15168), .B1(n15142), .B2(n15166), .ZN(
        n15144) );
  AOI21_X1 U16829 ( .B1(n15145), .B2(n15327), .A(n15144), .ZN(n15146) );
  OAI21_X1 U16830 ( .B1(n15147), .B2(n15311), .A(n15146), .ZN(n15312) );
  NAND2_X1 U16831 ( .A1(n15312), .A2(n15482), .ZN(n15154) );
  AOI211_X1 U16832 ( .C1(n15149), .C2(n15158), .A(n15187), .B(n15148), .ZN(
        n15313) );
  AOI22_X1 U16833 ( .A1(n15484), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15150), 
        .B2(n15480), .ZN(n15151) );
  OAI21_X1 U16834 ( .B1(n15380), .B2(n15196), .A(n15151), .ZN(n15152) );
  AOI21_X1 U16835 ( .B1(n15313), .B2(n15175), .A(n15152), .ZN(n15153) );
  OAI211_X1 U16836 ( .C1(n15311), .C2(n15155), .A(n15154), .B(n15153), .ZN(
        P1_U3275) );
  XOR2_X1 U16837 ( .A(n15156), .B(n15164), .Z(n15322) );
  INV_X1 U16838 ( .A(n15158), .ZN(n15159) );
  AOI211_X1 U16839 ( .C1(n15319), .C2(n15157), .A(n15159), .B(n15187), .ZN(
        n15318) );
  INV_X1 U16840 ( .A(n15160), .ZN(n15161) );
  AOI22_X1 U16841 ( .A1(n15484), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15161), 
        .B2(n15480), .ZN(n15162) );
  OAI21_X1 U16842 ( .B1(n6724), .B2(n15196), .A(n15162), .ZN(n15174) );
  NAND2_X1 U16843 ( .A1(n15184), .A2(n15163), .ZN(n15165) );
  AOI21_X1 U16844 ( .B1(n15165), .B2(n15164), .A(n15300), .ZN(n15171) );
  OAI22_X1 U16845 ( .A1(n15169), .A2(n15168), .B1(n15167), .B2(n15166), .ZN(
        n15170) );
  AOI21_X1 U16846 ( .B1(n15172), .B2(n15171), .A(n15170), .ZN(n15321) );
  NOR2_X1 U16847 ( .A1(n15321), .A2(n15484), .ZN(n15173) );
  AOI211_X1 U16848 ( .C1(n15318), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        n15176) );
  OAI21_X1 U16849 ( .B1(n15478), .B2(n15322), .A(n15176), .ZN(P1_U3276) );
  INV_X1 U16850 ( .A(n15177), .ZN(n15181) );
  AOI211_X1 U16851 ( .C1(n12650), .C2(n15179), .A(n15183), .B(n15178), .ZN(
        n15180) );
  NOR2_X1 U16852 ( .A1(n15181), .A2(n15180), .ZN(n15330) );
  INV_X1 U16853 ( .A(n15182), .ZN(n15186) );
  INV_X1 U16854 ( .A(n15183), .ZN(n15185) );
  OAI21_X1 U16855 ( .B1(n15186), .B2(n15185), .A(n15184), .ZN(n15328) );
  AOI21_X1 U16856 ( .B1(n15206), .B2(n15188), .A(n15187), .ZN(n15189) );
  NAND2_X1 U16857 ( .A1(n15189), .A2(n15157), .ZN(n15324) );
  AOI22_X1 U16858 ( .A1(n15193), .A2(n15192), .B1(n15191), .B2(n15190), .ZN(
        n15323) );
  INV_X1 U16859 ( .A(n15194), .ZN(n15195) );
  OAI22_X1 U16860 ( .A1(n15323), .A2(n15484), .B1(n15195), .B2(n15208), .ZN(
        n15198) );
  NOR2_X1 U16861 ( .A1(n15325), .A2(n15196), .ZN(n15197) );
  AOI211_X1 U16862 ( .C1(n15484), .C2(P1_REG2_REG_16__SCAN_IN), .A(n15198), 
        .B(n15197), .ZN(n15199) );
  OAI21_X1 U16863 ( .B1(n15324), .B2(n15215), .A(n15199), .ZN(n15200) );
  AOI21_X1 U16864 ( .B1(n15328), .B2(n15201), .A(n15200), .ZN(n15202) );
  OAI21_X1 U16865 ( .B1(n15330), .B2(n15478), .A(n15202), .ZN(P1_U3277) );
  NAND2_X1 U16866 ( .A1(n15204), .A2(n15203), .ZN(n15205) );
  XNOR2_X1 U16867 ( .A(n15205), .B(n7084), .ZN(n15335) );
  OAI211_X1 U16868 ( .C1(n15386), .C2(n15207), .A(n15283), .B(n15206), .ZN(
        n15331) );
  OAI22_X1 U16869 ( .A1(n15482), .A2(n15210), .B1(n15209), .B2(n15208), .ZN(
        n15211) );
  AOI21_X1 U16870 ( .B1(n15213), .B2(n15212), .A(n15211), .ZN(n15214) );
  OAI21_X1 U16871 ( .B1(n15331), .B2(n15215), .A(n15214), .ZN(n15223) );
  NAND2_X1 U16872 ( .A1(n15217), .A2(n15216), .ZN(n15219) );
  XNOR2_X1 U16873 ( .A(n15218), .B(n15219), .ZN(n15220) );
  NAND2_X1 U16874 ( .A1(n15220), .A2(n15327), .ZN(n15333) );
  INV_X1 U16875 ( .A(n15221), .ZN(n15332) );
  AOI21_X1 U16876 ( .B1(n15333), .B2(n15332), .A(n15484), .ZN(n15222) );
  AOI211_X1 U16877 ( .C1(n15335), .C2(n15224), .A(n15223), .B(n15222), .ZN(
        n15225) );
  INV_X1 U16878 ( .A(n15225), .ZN(P1_U3278) );
  INV_X1 U16879 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15227) );
  OAI21_X1 U16880 ( .B1(n15229), .B2(n15346), .A(n15228), .ZN(P1_U3559) );
  INV_X1 U16881 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n15232) );
  MUX2_X1 U16882 ( .A(n15232), .B(n15354), .S(n15518), .Z(n15233) );
  OAI21_X1 U16883 ( .B1(n15357), .B2(n15346), .A(n15233), .ZN(P1_U3558) );
  NOR3_X1 U16884 ( .A1(n15235), .A2(n15353), .A3(n15234), .ZN(n15236) );
  NAND4_X1 U16885 ( .A1(n15244), .A2(n15237), .A3(n15243), .A4(n15494), .ZN(
        n15240) );
  OAI211_X1 U16886 ( .C1(n15246), .C2(n15240), .A(n15239), .B(n15238), .ZN(
        n15241) );
  INV_X1 U16887 ( .A(n15241), .ZN(n15249) );
  NAND4_X1 U16888 ( .A1(n15244), .A2(n15243), .A3(n15494), .A4(n15242), .ZN(
        n15245) );
  NAND2_X1 U16889 ( .A1(n15245), .A2(n15489), .ZN(n15247) );
  INV_X1 U16890 ( .A(n15255), .ZN(n15256) );
  AOI21_X1 U16891 ( .B1(n15504), .B2(n15258), .A(n15257), .ZN(n15259) );
  MUX2_X1 U16892 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15359), .S(n15518), .Z(
        P1_U3555) );
  AOI22_X1 U16893 ( .A1(n15265), .A2(n15283), .B1(n15504), .B2(n15264), .ZN(
        n15266) );
  OAI211_X1 U16894 ( .C1(n15353), .C2(n15268), .A(n15267), .B(n15266), .ZN(
        n15360) );
  MUX2_X1 U16895 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15360), .S(n15518), .Z(
        P1_U3554) );
  OAI21_X1 U16896 ( .B1(n15270), .B2(n15489), .A(n15269), .ZN(n15271) );
  AOI211_X1 U16897 ( .C1(n15273), .C2(n15327), .A(n15272), .B(n15271), .ZN(
        n15274) );
  OAI21_X1 U16898 ( .B1(n15353), .B2(n15275), .A(n15274), .ZN(n15361) );
  MUX2_X1 U16899 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15361), .S(n15518), .Z(
        P1_U3553) );
  MUX2_X1 U16900 ( .A(n15279), .B(n15362), .S(n15518), .Z(n15280) );
  OAI21_X1 U16901 ( .B1(n15365), .B2(n15346), .A(n15280), .ZN(P1_U3552) );
  INV_X1 U16902 ( .A(n15281), .ZN(n15286) );
  AOI22_X1 U16903 ( .A1(n15284), .A2(n15283), .B1(n15504), .B2(n15282), .ZN(
        n15285) );
  OAI211_X1 U16904 ( .C1(n15353), .C2(n15287), .A(n15286), .B(n15285), .ZN(
        n15366) );
  MUX2_X1 U16905 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15366), .S(n15518), .Z(
        P1_U3551) );
  AOI211_X1 U16906 ( .C1(n15494), .C2(n15290), .A(n15289), .B(n15288), .ZN(
        n15367) );
  MUX2_X1 U16907 ( .A(n15291), .B(n15367), .S(n15518), .Z(n15292) );
  OAI21_X1 U16908 ( .B1(n15346), .B2(n15370), .A(n15292), .ZN(P1_U3550) );
  AND2_X1 U16909 ( .A1(n15293), .A2(n15494), .ZN(n15297) );
  OAI21_X1 U16910 ( .B1(n7461), .B2(n15489), .A(n15294), .ZN(n15295) );
  MUX2_X1 U16911 ( .A(n15371), .B(P1_REG1_REG_21__SCAN_IN), .S(n15516), .Z(
        P1_U3549) );
  OAI211_X1 U16912 ( .C1(n15301), .C2(n15300), .A(n15299), .B(n15298), .ZN(
        n15302) );
  AOI21_X1 U16913 ( .B1(n15303), .B2(n15494), .A(n15302), .ZN(n15372) );
  MUX2_X1 U16914 ( .A(n15304), .B(n15372), .S(n15518), .Z(n15305) );
  OAI21_X1 U16915 ( .B1(n15375), .B2(n15346), .A(n15305), .ZN(P1_U3548) );
  AOI21_X1 U16916 ( .B1(n15504), .B2(n15307), .A(n15306), .ZN(n15308) );
  OAI211_X1 U16917 ( .C1(n15353), .C2(n15310), .A(n15309), .B(n15308), .ZN(
        n15376) );
  MUX2_X1 U16918 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15376), .S(n15518), .Z(
        P1_U3547) );
  INV_X1 U16919 ( .A(n15311), .ZN(n15315) );
  AOI211_X1 U16920 ( .C1(n15315), .C2(n15314), .A(n15313), .B(n15312), .ZN(
        n15377) );
  MUX2_X1 U16921 ( .A(n15316), .B(n15377), .S(n15518), .Z(n15317) );
  OAI21_X1 U16922 ( .B1(n15380), .B2(n15346), .A(n15317), .ZN(P1_U3546) );
  AOI21_X1 U16923 ( .B1(n15504), .B2(n15319), .A(n15318), .ZN(n15320) );
  OAI211_X1 U16924 ( .C1(n15353), .C2(n15322), .A(n15321), .B(n15320), .ZN(
        n15381) );
  MUX2_X1 U16925 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15381), .S(n15518), .Z(
        P1_U3545) );
  OAI211_X1 U16926 ( .C1(n15325), .C2(n15489), .A(n15324), .B(n15323), .ZN(
        n15326) );
  AOI21_X1 U16927 ( .B1(n15328), .B2(n15327), .A(n15326), .ZN(n15329) );
  OAI21_X1 U16928 ( .B1(n15353), .B2(n15330), .A(n15329), .ZN(n15382) );
  MUX2_X1 U16929 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15382), .S(n15518), .Z(
        P1_U3544) );
  NAND3_X1 U16930 ( .A1(n15333), .A2(n15332), .A3(n15331), .ZN(n15334) );
  AOI21_X1 U16931 ( .B1(n15335), .B2(n15494), .A(n15334), .ZN(n15383) );
  MUX2_X1 U16932 ( .A(n15336), .B(n15383), .S(n15518), .Z(n15337) );
  OAI21_X1 U16933 ( .B1(n15386), .B2(n15346), .A(n15337), .ZN(P1_U3543) );
  NOR2_X1 U16934 ( .A1(n15339), .A2(n15353), .ZN(n15343) );
  NOR4_X1 U16935 ( .A1(n15343), .A2(n15342), .A3(n15341), .A4(n15340), .ZN(
        n15387) );
  MUX2_X1 U16936 ( .A(n15344), .B(n15387), .S(n15518), .Z(n15345) );
  OAI21_X1 U16937 ( .B1(n7457), .B2(n15346), .A(n15345), .ZN(P1_U3542) );
  INV_X1 U16938 ( .A(n15347), .ZN(n15352) );
  AOI21_X1 U16939 ( .B1(n15504), .B2(n15349), .A(n15348), .ZN(n15350) );
  OAI211_X1 U16940 ( .C1(n15353), .C2(n15352), .A(n15351), .B(n15350), .ZN(
        n15390) );
  MUX2_X1 U16941 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15390), .S(n15518), .Z(
        P1_U3539) );
  MUX2_X1 U16942 ( .A(n15355), .B(n15354), .S(n15512), .Z(n15356) );
  OAI21_X1 U16943 ( .B1(n15357), .B2(n15389), .A(n15356), .ZN(P1_U3526) );
  MUX2_X1 U16944 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15358), .S(n15512), .Z(
        P1_U3525) );
  MUX2_X1 U16945 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15359), .S(n15512), .Z(
        P1_U3523) );
  MUX2_X1 U16946 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15360), .S(n15512), .Z(
        P1_U3522) );
  MUX2_X1 U16947 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15361), .S(n15512), .Z(
        P1_U3521) );
  INV_X1 U16948 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15363) );
  MUX2_X1 U16949 ( .A(n15363), .B(n15362), .S(n15512), .Z(n15364) );
  OAI21_X1 U16950 ( .B1(n15365), .B2(n15389), .A(n15364), .ZN(P1_U3520) );
  MUX2_X1 U16951 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15366), .S(n15512), .Z(
        P1_U3519) );
  INV_X1 U16952 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n15368) );
  MUX2_X1 U16953 ( .A(n15368), .B(n15367), .S(n15512), .Z(n15369) );
  OAI21_X1 U16954 ( .B1(n15389), .B2(n15370), .A(n15369), .ZN(P1_U3518) );
  MUX2_X1 U16955 ( .A(n15371), .B(P1_REG0_REG_21__SCAN_IN), .S(n15510), .Z(
        P1_U3517) );
  INV_X1 U16956 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15373) );
  MUX2_X1 U16957 ( .A(n15373), .B(n15372), .S(n15512), .Z(n15374) );
  OAI21_X1 U16958 ( .B1(n15375), .B2(n15389), .A(n15374), .ZN(P1_U3516) );
  MUX2_X1 U16959 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15376), .S(n15512), .Z(
        P1_U3515) );
  INV_X1 U16960 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n15378) );
  MUX2_X1 U16961 ( .A(n15378), .B(n15377), .S(n15512), .Z(n15379) );
  OAI21_X1 U16962 ( .B1(n15380), .B2(n15389), .A(n15379), .ZN(P1_U3513) );
  MUX2_X1 U16963 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15381), .S(n15512), .Z(
        P1_U3510) );
  MUX2_X1 U16964 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15382), .S(n15512), .Z(
        P1_U3507) );
  INV_X1 U16965 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15384) );
  MUX2_X1 U16966 ( .A(n15384), .B(n15383), .S(n15512), .Z(n15385) );
  OAI21_X1 U16967 ( .B1(n15386), .B2(n15389), .A(n15385), .ZN(P1_U3504) );
  MUX2_X1 U16968 ( .A(n15730), .B(n15387), .S(n15512), .Z(n15388) );
  OAI21_X1 U16969 ( .B1(n7457), .B2(n15389), .A(n15388), .ZN(P1_U3501) );
  MUX2_X1 U16970 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15390), .S(n15512), .Z(
        P1_U3492) );
  NOR4_X1 U16971 ( .A1(n15392), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n9863), .ZN(n15393) );
  AOI21_X1 U16972 ( .B1(n15394), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15393), 
        .ZN(n15395) );
  OAI21_X1 U16973 ( .B1(n15396), .B2(n15400), .A(n15395), .ZN(P1_U3324) );
  OAI222_X1 U16974 ( .A1(P1_U3086), .A2(n15401), .B1(n15400), .B2(n15399), 
        .C1(n15398), .C2(n15397), .ZN(P1_U3326) );
  MUX2_X1 U16975 ( .A(n15403), .B(n15402), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16976 ( .A(n15404), .ZN(n15405) );
  MUX2_X1 U16977 ( .A(n15405), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U16978 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15406), .Z(SUB_1596_U53) );
  XOR2_X1 U16979 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n15407), .Z(SUB_1596_U54) );
  INV_X1 U16980 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15410) );
  INV_X1 U16981 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15424) );
  NAND2_X1 U16982 ( .A1(n15424), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n15425) );
  OAI21_X1 U16983 ( .B1(n15424), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n15425), 
        .ZN(n15417) );
  NOR2_X1 U16984 ( .A1(n15413), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15411) );
  NAND2_X1 U16985 ( .A1(n15413), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15414) );
  NAND2_X1 U16986 ( .A1(n15415), .A2(n15414), .ZN(n15427) );
  INV_X1 U16987 ( .A(n15427), .ZN(n15416) );
  XOR2_X1 U16988 ( .A(n15417), .B(n15416), .Z(n15419) );
  INV_X1 U16989 ( .A(n15419), .ZN(n15420) );
  NAND2_X1 U16990 ( .A1(n15431), .A2(n15423), .ZN(n15422) );
  XNOR2_X1 U16991 ( .A(n15422), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  NOR2_X1 U16992 ( .A1(n15424), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n15426) );
  OAI21_X1 U16993 ( .B1(n15427), .B2(n15426), .A(n15425), .ZN(n15437) );
  XNOR2_X1 U16994 ( .A(n15438), .B(P1_ADDR_REG_16__SCAN_IN), .ZN(n15428) );
  XNOR2_X1 U16995 ( .A(n15437), .B(n15428), .ZN(n15429) );
  INV_X1 U16996 ( .A(n15435), .ZN(n15432) );
  NAND2_X1 U16997 ( .A1(n15432), .A2(n15434), .ZN(n15433) );
  XNOR2_X1 U16998 ( .A(n15433), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NOR2_X1 U16999 ( .A1(n15438), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15436) );
  OR2_X1 U17000 ( .A1(n15437), .A2(n15436), .ZN(n15440) );
  NAND2_X1 U17001 ( .A1(n15438), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15439) );
  XNOR2_X1 U17002 ( .A(n15449), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n15447) );
  XOR2_X1 U17003 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15447), .Z(n15441) );
  INV_X1 U17004 ( .A(n15446), .ZN(n15443) );
  NAND2_X1 U17005 ( .A1(n15442), .A2(n15441), .ZN(n15445) );
  NAND2_X1 U17006 ( .A1(n15443), .A2(n15445), .ZN(n15444) );
  XNOR2_X1 U17007 ( .A(n15444), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  NAND2_X1 U17008 ( .A1(n15447), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n15451) );
  INV_X1 U17009 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15448) );
  NAND2_X1 U17010 ( .A1(n15449), .A2(n15448), .ZN(n15450) );
  NAND2_X1 U17011 ( .A1(n15451), .A2(n15450), .ZN(n15455) );
  NAND2_X1 U17012 ( .A1(n15773), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n15463) );
  INV_X1 U17013 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15452) );
  NAND2_X1 U17014 ( .A1(n15452), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n15453) );
  NAND2_X1 U17015 ( .A1(n15463), .A2(n15453), .ZN(n15454) );
  NAND2_X1 U17016 ( .A1(n15455), .A2(n15454), .ZN(n15456) );
  INV_X1 U17017 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15459) );
  XNOR2_X1 U17018 ( .A(n15458), .B(n15459), .ZN(n15457) );
  XNOR2_X1 U17019 ( .A(n15462), .B(n15457), .ZN(SUB_1596_U62) );
  NAND2_X1 U17020 ( .A1(n15458), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15461) );
  INV_X1 U17021 ( .A(n15458), .ZN(n15460) );
  NAND2_X1 U17022 ( .A1(n15464), .A2(n15463), .ZN(n15468) );
  XNOR2_X1 U17023 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15466) );
  XNOR2_X1 U17024 ( .A(n15466), .B(n15465), .ZN(n15467) );
  XNOR2_X1 U17025 ( .A(n15468), .B(n15467), .ZN(n15469) );
  XNOR2_X1 U17026 ( .A(n15470), .B(n15469), .ZN(SUB_1596_U4) );
  AOI21_X1 U17027 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15471) );
  OAI21_X1 U17028 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15471), 
        .ZN(U28) );
  AOI21_X1 U17029 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15472) );
  OAI21_X1 U17030 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15472), 
        .ZN(U29) );
  AOI21_X1 U17031 ( .B1(n9877), .B2(n6435), .A(n15473), .ZN(n15474) );
  NOR2_X1 U17032 ( .A1(n15475), .A2(n15474), .ZN(n15483) );
  AOI21_X1 U17033 ( .B1(n15478), .B2(n15477), .A(n15476), .ZN(n15479) );
  AOI21_X1 U17034 ( .B1(n15480), .B2(P1_REG3_REG_0__SCAN_IN), .A(n15479), .ZN(
        n15481) );
  OAI221_X1 U17035 ( .B1(n15484), .B2(n15483), .C1(n15482), .C2(n10724), .A(
        n15481), .ZN(P1_U3293) );
  AND2_X1 U17036 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15487), .ZN(P1_U3294) );
  AND2_X1 U17037 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15487), .ZN(P1_U3295) );
  INV_X1 U17038 ( .A(n15487), .ZN(n15486) );
  INV_X1 U17039 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15670) );
  NOR2_X1 U17040 ( .A1(n15486), .A2(n15670), .ZN(P1_U3296) );
  INV_X1 U17041 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15679) );
  NOR2_X1 U17042 ( .A1(n15486), .A2(n15679), .ZN(P1_U3297) );
  AND2_X1 U17043 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15487), .ZN(P1_U3298) );
  AND2_X1 U17044 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15487), .ZN(P1_U3299) );
  INV_X1 U17045 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15485) );
  NOR2_X1 U17046 ( .A1(n15486), .A2(n15485), .ZN(P1_U3300) );
  AND2_X1 U17047 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15487), .ZN(P1_U3301) );
  AND2_X1 U17048 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15487), .ZN(P1_U3302) );
  AND2_X1 U17049 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15487), .ZN(P1_U3303) );
  AND2_X1 U17050 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15487), .ZN(P1_U3304) );
  AND2_X1 U17051 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15487), .ZN(P1_U3305) );
  INV_X1 U17052 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15684) );
  NOR2_X1 U17053 ( .A1(n15486), .A2(n15684), .ZN(P1_U3306) );
  AND2_X1 U17054 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15487), .ZN(P1_U3307) );
  AND2_X1 U17055 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15487), .ZN(P1_U3308) );
  AND2_X1 U17056 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15487), .ZN(P1_U3309) );
  AND2_X1 U17057 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15487), .ZN(P1_U3310) );
  AND2_X1 U17058 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15487), .ZN(P1_U3311) );
  INV_X1 U17059 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15678) );
  NOR2_X1 U17060 ( .A1(n15486), .A2(n15678), .ZN(P1_U3312) );
  AND2_X1 U17061 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15487), .ZN(P1_U3313) );
  INV_X1 U17062 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15761) );
  NOR2_X1 U17063 ( .A1(n15486), .A2(n15761), .ZN(P1_U3314) );
  AND2_X1 U17064 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15487), .ZN(P1_U3315) );
  AND2_X1 U17065 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15487), .ZN(P1_U3316) );
  AND2_X1 U17066 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15487), .ZN(P1_U3317) );
  AND2_X1 U17067 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15487), .ZN(P1_U3318) );
  AND2_X1 U17068 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15487), .ZN(P1_U3319) );
  AND2_X1 U17069 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15487), .ZN(P1_U3320) );
  AND2_X1 U17070 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15487), .ZN(P1_U3321) );
  AND2_X1 U17071 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15487), .ZN(P1_U3322) );
  AND2_X1 U17072 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15487), .ZN(P1_U3323) );
  OAI21_X1 U17073 ( .B1(n10469), .B2(n15489), .A(n15488), .ZN(n15492) );
  INV_X1 U17074 ( .A(n15490), .ZN(n15491) );
  AOI211_X1 U17075 ( .C1(n15494), .C2(n15493), .A(n15492), .B(n15491), .ZN(
        n15514) );
  AOI22_X1 U17076 ( .A1(n15512), .A2(n15514), .B1(n9529), .B2(n15510), .ZN(
        P1_U3468) );
  AOI21_X1 U17077 ( .B1(n15504), .B2(n15496), .A(n15495), .ZN(n15497) );
  OAI211_X1 U17078 ( .C1(n15499), .C2(n15507), .A(n15498), .B(n15497), .ZN(
        n15500) );
  INV_X1 U17079 ( .A(n15500), .ZN(n15515) );
  INV_X1 U17080 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15501) );
  AOI22_X1 U17081 ( .A1(n15512), .A2(n15515), .B1(n15501), .B2(n15510), .ZN(
        P1_U3474) );
  AOI21_X1 U17082 ( .B1(n15504), .B2(n15503), .A(n15502), .ZN(n15505) );
  OAI211_X1 U17083 ( .C1(n15508), .C2(n15507), .A(n15506), .B(n15505), .ZN(
        n15509) );
  INV_X1 U17084 ( .A(n15509), .ZN(n15517) );
  INV_X1 U17085 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15511) );
  AOI22_X1 U17086 ( .A1(n15512), .A2(n15517), .B1(n15511), .B2(n15510), .ZN(
        P1_U3480) );
  INV_X1 U17087 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n15513) );
  AOI22_X1 U17088 ( .A1(n15518), .A2(n15514), .B1(n15513), .B2(n15516), .ZN(
        P1_U3531) );
  AOI22_X1 U17089 ( .A1(n15518), .A2(n15515), .B1(n10926), .B2(n15516), .ZN(
        P1_U3533) );
  AOI22_X1 U17090 ( .A1(n15518), .A2(n15517), .B1(n10980), .B2(n15516), .ZN(
        P1_U3535) );
  NOR2_X1 U17091 ( .A1(n15525), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI21_X1 U17092 ( .B1(n15521), .B2(n15520), .A(n15519), .ZN(n15528) );
  OAI22_X1 U17093 ( .A1(n15543), .A2(n15523), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15522), .ZN(n15524) );
  INV_X1 U17094 ( .A(n15524), .ZN(n15527) );
  NAND2_X1 U17095 ( .A1(n15525), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n15526) );
  OAI211_X1 U17096 ( .C1(n15529), .C2(n15528), .A(n15527), .B(n15526), .ZN(
        n15530) );
  INV_X1 U17097 ( .A(n15530), .ZN(n15535) );
  OAI211_X1 U17098 ( .C1(n15533), .C2(n15532), .A(n15546), .B(n15531), .ZN(
        n15534) );
  NAND2_X1 U17099 ( .A1(n15535), .A2(n15534), .ZN(P2_U3216) );
  OAI211_X1 U17100 ( .C1(n15539), .C2(n15538), .A(n15537), .B(n15536), .ZN(
        n15541) );
  OAI211_X1 U17101 ( .C1(n15543), .C2(n15542), .A(n15541), .B(n15540), .ZN(
        n15544) );
  INV_X1 U17102 ( .A(n15544), .ZN(n15550) );
  OAI211_X1 U17103 ( .C1(n15548), .C2(n15547), .A(n15546), .B(n15545), .ZN(
        n15549) );
  OAI211_X1 U17104 ( .C1(n15552), .C2(n15551), .A(n15550), .B(n15549), .ZN(
        P2_U3221) );
  AND2_X1 U17105 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15555), .ZN(P2_U3266) );
  AND2_X1 U17106 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15555), .ZN(P2_U3267) );
  AND2_X1 U17107 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15555), .ZN(P2_U3268) );
  AND2_X1 U17108 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15555), .ZN(P2_U3269) );
  AND2_X1 U17109 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15555), .ZN(P2_U3270) );
  INV_X1 U17110 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15707) );
  NOR2_X1 U17111 ( .A1(n15554), .A2(n15707), .ZN(P2_U3271) );
  AND2_X1 U17112 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15555), .ZN(P2_U3272) );
  INV_X1 U17113 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15682) );
  NOR2_X1 U17114 ( .A1(n15554), .A2(n15682), .ZN(P2_U3273) );
  AND2_X1 U17115 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15555), .ZN(P2_U3274) );
  INV_X1 U17116 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15681) );
  NOR2_X1 U17117 ( .A1(n15554), .A2(n15681), .ZN(P2_U3275) );
  AND2_X1 U17118 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15555), .ZN(P2_U3276) );
  INV_X1 U17119 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15756) );
  NOR2_X1 U17120 ( .A1(n15554), .A2(n15756), .ZN(P2_U3277) );
  AND2_X1 U17121 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15555), .ZN(P2_U3278) );
  AND2_X1 U17122 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15555), .ZN(P2_U3279) );
  AND2_X1 U17123 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15555), .ZN(P2_U3280) );
  INV_X1 U17124 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15770) );
  NOR2_X1 U17125 ( .A1(n15554), .A2(n15770), .ZN(P2_U3281) );
  AND2_X1 U17126 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15555), .ZN(P2_U3282) );
  AND2_X1 U17127 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15555), .ZN(P2_U3283) );
  AND2_X1 U17128 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15555), .ZN(P2_U3284) );
  AND2_X1 U17129 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15555), .ZN(P2_U3285) );
  AND2_X1 U17130 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15555), .ZN(P2_U3286) );
  AND2_X1 U17131 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15555), .ZN(P2_U3287) );
  AND2_X1 U17132 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15555), .ZN(P2_U3288) );
  AND2_X1 U17133 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15555), .ZN(P2_U3289) );
  AND2_X1 U17134 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15555), .ZN(P2_U3290) );
  INV_X1 U17135 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15774) );
  NOR2_X1 U17136 ( .A1(n15554), .A2(n15774), .ZN(P2_U3291) );
  AND2_X1 U17137 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15555), .ZN(P2_U3292) );
  AND2_X1 U17138 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15555), .ZN(P2_U3293) );
  AND2_X1 U17139 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15555), .ZN(P2_U3294) );
  AND2_X1 U17140 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15555), .ZN(P2_U3295) );
  AOI22_X1 U17141 ( .A1(n15558), .A2(n15557), .B1(n15556), .B2(n15560), .ZN(
        P2_U3416) );
  AOI21_X1 U17142 ( .B1(n15561), .B2(n15560), .A(n15559), .ZN(P2_U3417) );
  AOI21_X1 U17143 ( .B1(n15564), .B2(n15563), .A(n15562), .ZN(n15565) );
  OAI21_X1 U17144 ( .B1(n15567), .B2(n15566), .A(n15565), .ZN(n15569) );
  NOR2_X1 U17145 ( .A1(n15569), .A2(n15568), .ZN(n15574) );
  INV_X1 U17146 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15571) );
  AOI22_X1 U17147 ( .A1(n15572), .A2(n15574), .B1(n15571), .B2(n15570), .ZN(
        P2_U3439) );
  AOI22_X1 U17148 ( .A1(n14618), .A2(n15574), .B1(n10995), .B2(n15573), .ZN(
        P2_U3502) );
  NOR2_X1 U17149 ( .A1(P3_U3897), .A2(n15575), .ZN(P3_U3150) );
  INV_X1 U17150 ( .A(n15576), .ZN(n15580) );
  OAI22_X1 U17151 ( .A1(n15580), .A2(n15579), .B1(n15578), .B2(n15577), .ZN(
        n15583) );
  INV_X1 U17152 ( .A(n15581), .ZN(n15582) );
  AOI211_X1 U17153 ( .C1(n15585), .C2(n15584), .A(n15583), .B(n15582), .ZN(
        n15586) );
  AOI22_X1 U17154 ( .A1(n15587), .A2(n9177), .B1(n15586), .B2(n15597), .ZN(
        P3_U3231) );
  INV_X1 U17155 ( .A(n15588), .ZN(n15589) );
  AOI21_X1 U17156 ( .B1(n15591), .B2(n15590), .A(n15589), .ZN(n15598) );
  AOI22_X1 U17157 ( .A1(n15594), .A2(n15593), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15592), .ZN(n15595) );
  OAI221_X1 U17158 ( .B1(n15587), .B2(n15598), .C1(n15597), .C2(n15596), .A(
        n15595), .ZN(P3_U3232) );
  AOI22_X1 U17159 ( .A1(n15631), .A2(n15599), .B1(n7751), .B2(n15629), .ZN(
        P3_U3393) );
  AOI22_X1 U17160 ( .A1(n15631), .A2(n15600), .B1(n8562), .B2(n15629), .ZN(
        P3_U3396) );
  NAND2_X1 U17161 ( .A1(n15605), .A2(n15607), .ZN(n15601) );
  OAI211_X1 U17162 ( .C1(n15603), .C2(n15621), .A(n15602), .B(n15601), .ZN(
        n15604) );
  AOI21_X1 U17163 ( .B1(n15605), .B2(n15627), .A(n15604), .ZN(n15633) );
  INV_X1 U17164 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15606) );
  AOI22_X1 U17165 ( .A1(n15631), .A2(n15633), .B1(n15606), .B2(n15629), .ZN(
        P3_U3399) );
  AOI21_X1 U17166 ( .B1(n15609), .B2(n9076), .A(n15608), .ZN(n15612) );
  INV_X1 U17167 ( .A(n15610), .ZN(n15611) );
  AOI211_X1 U17168 ( .C1(n15614), .C2(n15613), .A(n15612), .B(n15611), .ZN(
        n15634) );
  INV_X1 U17169 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15615) );
  AOI22_X1 U17170 ( .A1(n15631), .A2(n15634), .B1(n15615), .B2(n15629), .ZN(
        P3_U3402) );
  OAI22_X1 U17171 ( .A1(n15617), .A2(n9076), .B1(n15621), .B2(n15616), .ZN(
        n15618) );
  NOR2_X1 U17172 ( .A1(n15619), .A2(n15618), .ZN(n15636) );
  INV_X1 U17173 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15620) );
  AOI22_X1 U17174 ( .A1(n15631), .A2(n15636), .B1(n15620), .B2(n15629), .ZN(
        P3_U3405) );
  INV_X1 U17175 ( .A(n15623), .ZN(n15628) );
  OAI22_X1 U17176 ( .A1(n15623), .A2(n9076), .B1(n15622), .B2(n15621), .ZN(
        n15626) );
  INV_X1 U17177 ( .A(n15624), .ZN(n15625) );
  AOI211_X1 U17178 ( .C1(n15628), .C2(n15627), .A(n15626), .B(n15625), .ZN(
        n15638) );
  INV_X1 U17179 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15630) );
  AOI22_X1 U17180 ( .A1(n15631), .A2(n15638), .B1(n15630), .B2(n15629), .ZN(
        P3_U3408) );
  AOI22_X1 U17181 ( .A1(n15639), .A2(n15633), .B1(n15632), .B2(n15637), .ZN(
        P3_U3462) );
  AOI22_X1 U17182 ( .A1(n15639), .A2(n15634), .B1(n9144), .B2(n15637), .ZN(
        P3_U3463) );
  AOI22_X1 U17183 ( .A1(n15639), .A2(n15636), .B1(n15635), .B2(n15637), .ZN(
        P3_U3464) );
  AOI22_X1 U17184 ( .A1(n15639), .A2(n15638), .B1(n8626), .B2(n15637), .ZN(
        P3_U3465) );
  OAI22_X1 U17185 ( .A1(n15740), .A2(keyinput28), .B1(n15641), .B2(keyinput58), 
        .ZN(n15640) );
  AOI221_X1 U17186 ( .B1(n15740), .B2(keyinput28), .C1(keyinput58), .C2(n15641), .A(n15640), .ZN(n15649) );
  OAI22_X1 U17187 ( .A1(n15732), .A2(keyinput18), .B1(n15731), .B2(keyinput44), 
        .ZN(n15642) );
  AOI221_X1 U17188 ( .B1(n15732), .B2(keyinput18), .C1(keyinput44), .C2(n15731), .A(n15642), .ZN(n15648) );
  XNOR2_X1 U17189 ( .A(SI_27_), .B(keyinput53), .ZN(n15646) );
  XNOR2_X1 U17190 ( .A(P3_IR_REG_14__SCAN_IN), .B(keyinput0), .ZN(n15645) );
  XNOR2_X1 U17191 ( .A(P3_IR_REG_11__SCAN_IN), .B(keyinput45), .ZN(n15644) );
  XNOR2_X1 U17192 ( .A(keyinput19), .B(P1_D_REG_25__SCAN_IN), .ZN(n15643) );
  AND4_X1 U17193 ( .A1(n15646), .A2(n15645), .A3(n15644), .A4(n15643), .ZN(
        n15647) );
  NAND3_X1 U17194 ( .A1(n15649), .A2(n15648), .A3(n15647), .ZN(n15789) );
  XNOR2_X1 U17195 ( .A(n15733), .B(keyinput5), .ZN(n15655) );
  XNOR2_X1 U17196 ( .A(n15650), .B(keyinput21), .ZN(n15654) );
  XNOR2_X1 U17197 ( .A(n7134), .B(keyinput11), .ZN(n15653) );
  XNOR2_X1 U17198 ( .A(n15651), .B(keyinput14), .ZN(n15652) );
  NOR4_X1 U17199 ( .A1(n15655), .A2(n15654), .A3(n15653), .A4(n15652), .ZN(
        n15663) );
  OAI22_X1 U17200 ( .A1(n15734), .A2(keyinput31), .B1(n15657), .B2(keyinput22), 
        .ZN(n15656) );
  AOI221_X1 U17201 ( .B1(n15734), .B2(keyinput31), .C1(keyinput22), .C2(n15657), .A(n15656), .ZN(n15662) );
  INV_X1 U17202 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15660) );
  OAI22_X1 U17203 ( .A1(n15660), .A2(keyinput48), .B1(n15659), .B2(keyinput42), 
        .ZN(n15658) );
  AOI221_X1 U17204 ( .B1(n15660), .B2(keyinput48), .C1(keyinput42), .C2(n15659), .A(n15658), .ZN(n15661) );
  NAND3_X1 U17205 ( .A1(n15663), .A2(n15662), .A3(n15661), .ZN(n15788) );
  AOI22_X1 U17206 ( .A1(n15666), .A2(keyinput10), .B1(keyinput50), .B2(n15665), 
        .ZN(n15664) );
  OAI221_X1 U17207 ( .B1(n15666), .B2(keyinput10), .C1(n15665), .C2(keyinput50), .A(n15664), .ZN(n15676) );
  AOI22_X1 U17208 ( .A1(n15668), .A2(keyinput49), .B1(keyinput27), .B2(n9602), 
        .ZN(n15667) );
  OAI221_X1 U17209 ( .B1(n15668), .B2(keyinput49), .C1(n9602), .C2(keyinput27), 
        .A(n15667), .ZN(n15675) );
  AOI22_X1 U17210 ( .A1(n15720), .A2(keyinput39), .B1(keyinput60), .B2(n15670), 
        .ZN(n15669) );
  OAI221_X1 U17211 ( .B1(n15720), .B2(keyinput39), .C1(n15670), .C2(keyinput60), .A(n15669), .ZN(n15674) );
  XNOR2_X1 U17212 ( .A(P3_D_REG_0__SCAN_IN), .B(keyinput24), .ZN(n15672) );
  XNOR2_X1 U17213 ( .A(P2_REG0_REG_14__SCAN_IN), .B(keyinput12), .ZN(n15671)
         );
  NAND2_X1 U17214 ( .A1(n15672), .A2(n15671), .ZN(n15673) );
  NOR4_X1 U17215 ( .A1(n15676), .A2(n15675), .A3(n15674), .A4(n15673), .ZN(
        n15718) );
  AOI22_X1 U17216 ( .A1(n15679), .A2(keyinput33), .B1(keyinput26), .B2(n15678), 
        .ZN(n15677) );
  OAI221_X1 U17217 ( .B1(n15679), .B2(keyinput33), .C1(n15678), .C2(keyinput26), .A(n15677), .ZN(n15690) );
  AOI22_X1 U17218 ( .A1(n15682), .A2(keyinput9), .B1(keyinput57), .B2(n15681), 
        .ZN(n15680) );
  OAI221_X1 U17219 ( .B1(n15682), .B2(keyinput9), .C1(n15681), .C2(keyinput57), 
        .A(n15680), .ZN(n15689) );
  INV_X1 U17220 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15721) );
  AOI22_X1 U17221 ( .A1(n15721), .A2(keyinput17), .B1(keyinput16), .B2(n15684), 
        .ZN(n15683) );
  OAI221_X1 U17222 ( .B1(n15721), .B2(keyinput17), .C1(n15684), .C2(keyinput16), .A(n15683), .ZN(n15688) );
  XNOR2_X1 U17223 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput2), .ZN(n15686) );
  XNOR2_X1 U17224 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput43), .ZN(n15685)
         );
  NAND2_X1 U17225 ( .A1(n15686), .A2(n15685), .ZN(n15687) );
  NOR4_X1 U17226 ( .A1(n15690), .A2(n15689), .A3(n15688), .A4(n15687), .ZN(
        n15717) );
  AOI22_X1 U17227 ( .A1(n15693), .A2(keyinput3), .B1(keyinput62), .B2(n15692), 
        .ZN(n15691) );
  OAI221_X1 U17228 ( .B1(n15693), .B2(keyinput3), .C1(n15692), .C2(keyinput62), 
        .A(n15691), .ZN(n15702) );
  AOI22_X1 U17229 ( .A1(n15695), .A2(keyinput34), .B1(keyinput7), .B2(n15730), 
        .ZN(n15694) );
  OAI221_X1 U17230 ( .B1(n15695), .B2(keyinput34), .C1(n15730), .C2(keyinput7), 
        .A(n15694), .ZN(n15701) );
  XOR2_X1 U17231 ( .A(n7812), .B(keyinput23), .Z(n15699) );
  XNOR2_X1 U17232 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput61), .ZN(n15698) );
  XNOR2_X1 U17233 ( .A(P3_REG2_REG_30__SCAN_IN), .B(keyinput56), .ZN(n15697)
         );
  XNOR2_X1 U17234 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput15), .ZN(n15696) );
  NAND4_X1 U17235 ( .A1(n15699), .A2(n15698), .A3(n15697), .A4(n15696), .ZN(
        n15700) );
  NOR3_X1 U17236 ( .A1(n15702), .A2(n15701), .A3(n15700), .ZN(n15716) );
  INV_X1 U17237 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15705) );
  AOI22_X1 U17238 ( .A1(n15705), .A2(keyinput40), .B1(n15704), .B2(keyinput52), 
        .ZN(n15703) );
  OAI221_X1 U17239 ( .B1(n15705), .B2(keyinput40), .C1(n15704), .C2(keyinput52), .A(n15703), .ZN(n15714) );
  INV_X1 U17240 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15726) );
  AOI22_X1 U17241 ( .A1(n8281), .A2(keyinput4), .B1(keyinput51), .B2(n15726), 
        .ZN(n15706) );
  OAI221_X1 U17242 ( .B1(n8281), .B2(keyinput4), .C1(n15726), .C2(keyinput51), 
        .A(n15706), .ZN(n15713) );
  XNOR2_X1 U17243 ( .A(n15707), .B(keyinput8), .ZN(n15712) );
  XOR2_X1 U17244 ( .A(n15729), .B(keyinput29), .Z(n15710) );
  XNOR2_X1 U17245 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput32), .ZN(n15709) );
  XNOR2_X1 U17246 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput63), .ZN(n15708) );
  NAND3_X1 U17247 ( .A1(n15710), .A2(n15709), .A3(n15708), .ZN(n15711) );
  NOR4_X1 U17248 ( .A1(n15714), .A2(n15713), .A3(n15712), .A4(n15711), .ZN(
        n15715) );
  NAND4_X1 U17249 ( .A1(n15718), .A2(n15717), .A3(n15716), .A4(n15715), .ZN(
        n15787) );
  NOR4_X1 U17250 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_0__SCAN_IN), .A3(
        n15720), .A4(n15719), .ZN(n15724) );
  NOR4_X1 U17251 ( .A1(P1_REG0_REG_8__SCAN_IN), .A2(P1_REG1_REG_9__SCAN_IN), 
        .A3(P2_ADDR_REG_13__SCAN_IN), .A4(n15721), .ZN(n15722) );
  AND4_X1 U17252 ( .A1(n15681), .A2(P3_REG3_REG_16__SCAN_IN), .A3(
        P1_IR_REG_7__SCAN_IN), .A4(n15722), .ZN(n15723) );
  NAND4_X1 U17253 ( .A1(n15725), .A2(n15724), .A3(n15723), .A4(
        P2_D_REG_24__SCAN_IN), .ZN(n15785) );
  NAND4_X1 U17254 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), 
        .A3(P1_IR_REG_22__SCAN_IN), .A4(n15726), .ZN(n15743) );
  NAND4_X1 U17255 ( .A1(n15730), .A2(n15729), .A3(n15728), .A4(n15727), .ZN(
        n15742) );
  NAND4_X1 U17256 ( .A1(n15754), .A2(n15760), .A3(n15759), .A4(n10724), .ZN(
        n15738) );
  NAND4_X1 U17257 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(SI_27_), .A3(n15732), .A4(
        n15731), .ZN(n15737) );
  NAND4_X1 U17258 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(P3_REG3_REG_14__SCAN_IN), 
        .A3(P2_IR_REG_0__SCAN_IN), .A4(n15733), .ZN(n15736) );
  NAND4_X1 U17259 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(P2_REG1_REG_30__SCAN_IN), 
        .A3(P1_REG3_REG_11__SCAN_IN), .A4(n15734), .ZN(n15735) );
  NOR4_X1 U17260 ( .A1(n15738), .A2(n15737), .A3(n15736), .A4(n15735), .ZN(
        n15739) );
  NAND4_X1 U17261 ( .A1(n15740), .A2(n15757), .A3(P1_REG3_REG_5__SCAN_IN), 
        .A4(n15739), .ZN(n15741) );
  NOR3_X1 U17262 ( .A1(n15743), .A2(n15742), .A3(n15741), .ZN(n15747) );
  NOR4_X1 U17263 ( .A1(n15744), .A2(P2_REG3_REG_20__SCAN_IN), .A3(
        P2_REG0_REG_20__SCAN_IN), .A4(P3_REG1_REG_2__SCAN_IN), .ZN(n15746) );
  AND4_X1 U17264 ( .A1(n15705), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n15745) );
  NAND4_X1 U17265 ( .A1(n15747), .A2(n15746), .A3(n15745), .A4(
        P3_DATAO_REG_31__SCAN_IN), .ZN(n15752) );
  NAND4_X1 U17266 ( .A1(n15770), .A2(n15772), .A3(n15773), .A4(n15769), .ZN(
        n15751) );
  NAND4_X1 U17267 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), 
        .A3(P2_D_REG_6__SCAN_IN), .A4(n15748), .ZN(n15750) );
  NAND4_X1 U17268 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .A3(
        P1_IR_REG_24__SCAN_IN), .A4(P1_REG3_REG_15__SCAN_IN), .ZN(n15749) );
  OR4_X1 U17269 ( .A1(n15752), .A2(n15751), .A3(n15750), .A4(n15749), .ZN(
        n15784) );
  AOI22_X1 U17270 ( .A1(n15754), .A2(keyinput35), .B1(keyinput37), .B2(n10724), 
        .ZN(n15753) );
  OAI221_X1 U17271 ( .B1(n15754), .B2(keyinput35), .C1(n10724), .C2(keyinput37), .A(n15753), .ZN(n15767) );
  AOI22_X1 U17272 ( .A1(n15757), .A2(keyinput54), .B1(n15756), .B2(keyinput59), 
        .ZN(n15755) );
  OAI221_X1 U17273 ( .B1(n15757), .B2(keyinput54), .C1(n15756), .C2(keyinput59), .A(n15755), .ZN(n15766) );
  AOI22_X1 U17274 ( .A1(n15760), .A2(keyinput25), .B1(keyinput20), .B2(n15759), 
        .ZN(n15758) );
  OAI221_X1 U17275 ( .B1(n15760), .B2(keyinput25), .C1(n15759), .C2(keyinput20), .A(n15758), .ZN(n15765) );
  XOR2_X1 U17276 ( .A(n15761), .B(keyinput6), .Z(n15763) );
  XNOR2_X1 U17277 ( .A(P3_REG1_REG_2__SCAN_IN), .B(keyinput30), .ZN(n15762) );
  NAND2_X1 U17278 ( .A1(n15763), .A2(n15762), .ZN(n15764) );
  NOR4_X1 U17279 ( .A1(n15767), .A2(n15766), .A3(n15765), .A4(n15764), .ZN(
        n15783) );
  AOI22_X1 U17280 ( .A1(n15770), .A2(keyinput36), .B1(keyinput46), .B2(n15769), 
        .ZN(n15768) );
  OAI221_X1 U17281 ( .B1(n15770), .B2(keyinput36), .C1(n15769), .C2(keyinput46), .A(n15768), .ZN(n15781) );
  AOI22_X1 U17282 ( .A1(n15773), .A2(keyinput41), .B1(n15772), .B2(keyinput47), 
        .ZN(n15771) );
  OAI221_X1 U17283 ( .B1(n15773), .B2(keyinput41), .C1(n15772), .C2(keyinput47), .A(n15771), .ZN(n15780) );
  XNOR2_X1 U17284 ( .A(n15774), .B(keyinput13), .ZN(n15779) );
  XNOR2_X1 U17285 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput38), .ZN(n15777) );
  XNOR2_X1 U17286 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput55), .ZN(n15776)
         );
  XNOR2_X1 U17287 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput1), .ZN(n15775) );
  NAND3_X1 U17288 ( .A1(n15777), .A2(n15776), .A3(n15775), .ZN(n15778) );
  NOR4_X1 U17289 ( .A1(n15781), .A2(n15780), .A3(n15779), .A4(n15778), .ZN(
        n15782) );
  OAI211_X1 U17290 ( .C1(n15785), .C2(n15784), .A(n15783), .B(n15782), .ZN(
        n15786) );
  NOR4_X1 U17291 ( .A1(n15789), .A2(n15788), .A3(n15787), .A4(n15786), .ZN(
        n15794) );
  MUX2_X1 U17292 ( .A(n15792), .B(n15791), .S(n15790), .Z(n15793) );
  XNOR2_X1 U17293 ( .A(n15794), .B(n15793), .ZN(P1_U3446) );
  AOI21_X1 U7236 ( .B1(n7492), .B2(n15327), .A(n12876), .ZN(n15267) );
  INV_X1 U9823 ( .A(n12148), .ZN(n6845) );
  NAND2_X1 U7188 ( .A1(n7385), .A2(n10135), .ZN(n7392) );
  CLKBUF_X2 U7244 ( .A(n7901), .Z(n7987) );
  CLKBUF_X1 U7263 ( .A(n6448), .Z(n7072) );
  NAND2_X1 U7264 ( .A1(n6844), .A2(n6845), .ZN(n7385) );
  CLKBUF_X2 U7267 ( .A(n9071), .Z(n6432) );
  CLKBUF_X1 U9713 ( .A(n13601), .Z(n6983) );
  CLKBUF_X3 U9930 ( .A(n9909), .Z(n6435) );
  CLKBUF_X1 U10058 ( .A(n9880), .Z(n14967) );
endmodule

