

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6548, n6549, n6550, n6551, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551;

  OR3_X1 U7296 ( .A1(n13497), .A2(n13496), .A3(n13495), .ZN(n13864) );
  OAI21_X1 U7297 ( .B1(n12776), .B2(n7469), .A(n7467), .ZN(n12801) );
  INV_X2 U7298 ( .A(n11655), .ZN(n11807) );
  INV_X2 U7299 ( .A(n11795), .ZN(n11765) );
  CLKBUF_X2 U7300 ( .A(n8503), .Z(n8813) );
  BUF_X2 U7301 ( .A(n8518), .Z(n11951) );
  AND4_X1 U7302 ( .A1(n8490), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(n8837)
         );
  NAND4_X2 U7303 ( .A1(n8475), .A2(n8474), .A3(n8473), .A4(n8472), .ZN(n12180)
         );
  AND2_X2 U7304 ( .A1(n8443), .A2(n8444), .ZN(n8484) );
  NAND2_X1 U7306 ( .A1(n8442), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7062) );
  INV_X1 U7307 ( .A(n14617), .ZN(n14598) );
  XNOR2_X1 U7308 ( .A(n7755), .B(n7752), .ZN(n14746) );
  AND2_X1 U7309 ( .A1(n7549), .A2(n7704), .ZN(n8139) );
  OAI211_X1 U7310 ( .C1(n12067), .C2(n12066), .A(n12065), .B(n12064), .ZN(
        n12070) );
  INV_X2 U7311 ( .A(n14123), .ZN(n14252) );
  INV_X1 U7312 ( .A(n12961), .ZN(n12878) );
  OR2_X1 U7313 ( .A1(n8758), .A2(n8757), .ZN(n8399) );
  AND4_X1 U7314 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(P3_REG2_REG_19__SCAN_IN), 
        .A3(P3_DATAO_REG_5__SCAN_IN), .A4(n13973), .ZN(n13838) );
  OAI221_X1 U7315 ( .B1(n13973), .B2(keyinput43), .C1(n13742), .C2(keyinput116), .A(n13741), .ZN(n13746) );
  AND4_X1 U7316 ( .A1(n8470), .A2(n8469), .A3(n8468), .A4(n8467), .ZN(n10076)
         );
  INV_X1 U7317 ( .A(n13083), .ZN(n11382) );
  INV_X1 U7318 ( .A(n9783), .ZN(n11381) );
  INV_X2 U7319 ( .A(n11797), .ZN(n11787) );
  NAND2_X1 U7320 ( .A1(n10044), .A2(n14103), .ZN(n11794) );
  NAND2_X2 U7321 ( .A1(n8999), .A2(n13064), .ZN(n7896) );
  OR2_X1 U7322 ( .A1(n14979), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7453) );
  INV_X1 U7323 ( .A(n8458), .ZN(n8877) );
  NAND2_X1 U7324 ( .A1(n11112), .A2(n12057), .ZN(n11165) );
  AND2_X1 U7325 ( .A1(n6909), .A2(n14746), .ZN(n14076) );
  INV_X1 U7326 ( .A(n7896), .ZN(n14086) );
  AND2_X1 U7327 ( .A1(n7916), .A2(n7915), .ZN(n15147) );
  INV_X1 U7328 ( .A(n13064), .ZN(n9293) );
  NOR2_X1 U7329 ( .A1(n10803), .A2(n13794), .ZN(n10923) );
  OAI211_X1 U7330 ( .C1(n9535), .C2(n10172), .A(n8540), .B(n8539), .ZN(n10754)
         );
  OAI21_X1 U7331 ( .B1(n11083), .B2(n8813), .A(n8814), .ZN(n11819) );
  INV_X1 U7332 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n12619) );
  NAND2_X1 U7333 ( .A1(n12620), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7064) );
  NAND2_X1 U7334 ( .A1(n7143), .A2(n7142), .ZN(n14116) );
  AND4_X1 U7335 ( .A1(n8723), .A2(n8722), .A3(n8721), .A4(n8720), .ZN(n12407)
         );
  XNOR2_X1 U7336 ( .A(n7064), .B(n7063), .ZN(n11337) );
  INV_X2 U7337 ( .A(n9531), .ZN(n12275) );
  NAND2_X1 U7338 ( .A1(n7051), .A2(n12770), .ZN(n12776) );
  AOI211_X1 U7339 ( .C1(n14659), .C2(n9398), .A(n13986), .B(n13985), .ZN(
        n13987) );
  AND2_X1 U7340 ( .A1(n7074), .A2(n7061), .ZN(n6548) );
  INV_X1 U7341 ( .A(n6551), .ZN(n6549) );
  AND2_X2 U7342 ( .A1(n14846), .A2(n14845), .ZN(n14990) );
  OR2_X2 U7343 ( .A1(n7245), .A2(n14987), .ZN(n14846) );
  OR2_X4 U7344 ( .A1(n11794), .A2(n8988), .ZN(n11797) );
  NAND2_X2 U7345 ( .A1(n7244), .A2(n7243), .ZN(n6972) );
  AND2_X2 U7346 ( .A1(n6834), .A2(n6833), .ZN(n7445) );
  AOI21_X2 U7347 ( .B1(n6616), .B2(n7270), .A(n7268), .ZN(n8653) );
  OAI22_X2 U7348 ( .A1(n6627), .A2(n7553), .B1(n14134), .B2(n7555), .ZN(n14138) );
  XNOR2_X2 U7349 ( .A(n14813), .B(n14814), .ZN(n14876) );
  NAND2_X2 U7350 ( .A1(n6821), .A2(n14812), .ZN(n14813) );
  AND2_X2 U7351 ( .A1(n8330), .A2(n6658), .ZN(n8332) );
  NAND4_X4 U7352 ( .A1(n7890), .A2(n7889), .A3(n7888), .A4(n7887), .ZN(n14336)
         );
  OAI21_X2 U7353 ( .B1(n12399), .B2(n6738), .A(n6736), .ZN(n12369) );
  NAND2_X2 U7354 ( .A1(n6967), .A2(n12398), .ZN(n12399) );
  AND2_X1 U7355 ( .A1(n13455), .A2(n13561), .ZN(n13457) );
  NOR2_X2 U7356 ( .A1(n11007), .A2(n12973), .ZN(n13455) );
  NOR2_X4 U7357 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8461) );
  AOI21_X2 U7358 ( .B1(n7242), .B2(n7241), .A(n6668), .ZN(n14788) );
  OR2_X1 U7359 ( .A1(n9778), .A2(n13157), .ZN(n6550) );
  OR2_X1 U7360 ( .A1(n9778), .A2(n13157), .ZN(n13562) );
  XNOR2_X2 U7361 ( .A(n7728), .B(n7727), .ZN(n14617) );
  OAI22_X2 U7362 ( .A1(n11005), .A2(n11004), .B1(n13577), .B2(n13198), .ZN(
        n11006) );
  NAND2_X2 U7363 ( .A1(n6743), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8413) );
  XNOR2_X2 U7364 ( .A(n7062), .B(n7061), .ZN(n12628) );
  NAND2_X2 U7365 ( .A1(n12868), .A2(n12867), .ZN(n12961) );
  NAND2_X2 U7366 ( .A1(n6578), .A2(n9454), .ZN(n12888) );
  CLKBUF_X3 U7367 ( .A(n9305), .Z(n6551) );
  AND2_X1 U7368 ( .A1(n9285), .A2(n9286), .ZN(n9305) );
  AOI211_X1 U7369 ( .C1(n10754), .C2(n11904), .A(n10736), .B(n10735), .ZN(
        n10737) );
  INV_X1 U7370 ( .A(n10754), .ZN(n15491) );
  BUF_X4 U7371 ( .A(n9464), .Z(n11502) );
  NOR2_X2 U7372 ( .A1(n7239), .A2(n7240), .ZN(n14983) );
  AOI21_X2 U7373 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n14826), .A(n14825), .ZN(
        n14830) );
  XOR2_X2 U7374 ( .A(n14793), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15550) );
  OR2_X1 U7375 ( .A1(n12298), .A2(n15497), .ZN(n7353) );
  AND2_X1 U7376 ( .A1(n11584), .A2(n11583), .ZN(n11613) );
  NAND2_X1 U7377 ( .A1(n12331), .A2(n8859), .ZN(n12319) );
  OAI21_X1 U7378 ( .B1(n12131), .B2(n12304), .A(n12130), .ZN(n12133) );
  NAND2_X1 U7379 ( .A1(n11650), .A2(n6554), .ZN(n6555) );
  OR2_X1 U7380 ( .A1(n12957), .A2(n12956), .ZN(n12965) );
  OR2_X1 U7381 ( .A1(n11120), .A2(n11119), .ZN(n11121) );
  OAI22_X1 U7382 ( .A1(n14145), .A2(n7145), .B1(n7144), .B2(n14146), .ZN(
        n14151) );
  NAND2_X1 U7383 ( .A1(n6557), .A2(n12024), .ZN(n10782) );
  INV_X2 U7384 ( .A(n12900), .ZN(n15380) );
  NAND2_X1 U7385 ( .A1(n14624), .A2(n9923), .ZN(n14106) );
  INV_X2 U7386 ( .A(n14123), .ZN(n14155) );
  INV_X4 U7387 ( .A(n11798), .ZN(n10307) );
  AND2_X1 U7388 ( .A1(n8443), .A2(n8444), .ZN(n6566) );
  INV_X2 U7389 ( .A(n13036), .ZN(n13098) );
  AND2_X1 U7391 ( .A1(n11337), .A2(n8444), .ZN(n8486) );
  INV_X2 U7393 ( .A(n9296), .ZN(n7659) );
  OAI21_X1 U7395 ( .B1(n7352), .B2(n15538), .A(n7351), .ZN(n11347) );
  INV_X1 U7396 ( .A(n7352), .ZN(n11348) );
  AOI211_X1 U7397 ( .C1(n12438), .C2(n11819), .A(n11579), .B(n11578), .ZN(
        n11580) );
  OR2_X1 U7398 ( .A1(n13491), .A2(n15405), .ZN(n7394) );
  OAI22_X1 U7399 ( .A1(n13263), .A2(n13265), .B1(n13276), .B2(n11540), .ZN(
        n6783) );
  AOI21_X1 U7400 ( .B1(n8954), .B2(n8955), .A(n8953), .ZN(n11577) );
  INV_X1 U7401 ( .A(n11613), .ZN(n6553) );
  AND2_X1 U7402 ( .A1(n7356), .A2(n7355), .ZN(n7354) );
  OR2_X1 U7403 ( .A1(n12298), .A2(n11601), .ZN(n7356) );
  NAND2_X1 U7404 ( .A1(n11341), .A2(n7624), .ZN(n11584) );
  INV_X1 U7405 ( .A(n6918), .ZN(n11561) );
  OAI21_X1 U7406 ( .B1(n12319), .B2(n7068), .A(n6599), .ZN(n12303) );
  NAND2_X1 U7407 ( .A1(n12300), .A2(n6555), .ZN(n11339) );
  OR2_X1 U7408 ( .A1(n8869), .A2(n11593), .ZN(n8951) );
  NAND2_X1 U7409 ( .A1(n12302), .A2(n12301), .ZN(n12300) );
  NAND2_X1 U7410 ( .A1(n12314), .A2(n12120), .ZN(n12302) );
  NAND2_X1 U7411 ( .A1(n13349), .A2(n11531), .ZN(n13336) );
  NAND2_X1 U7412 ( .A1(n11729), .A2(n7657), .ZN(n13969) );
  NAND2_X1 U7413 ( .A1(n11986), .A2(n8863), .ZN(n11984) );
  NAND2_X1 U7414 ( .A1(n7427), .A2(n6607), .ZN(n13349) );
  NAND2_X1 U7415 ( .A1(n13389), .A2(n7429), .ZN(n7427) );
  OAI21_X1 U7416 ( .B1(n12366), .B2(n7614), .A(n7611), .ZN(n12330) );
  AOI21_X1 U7417 ( .B1(n6599), .B2(n7068), .A(n7359), .ZN(n7358) );
  AND2_X1 U7418 ( .A1(n14852), .A2(n14853), .ZN(n14993) );
  NAND2_X1 U7419 ( .A1(n12391), .A2(n12101), .ZN(n12368) );
  OR2_X1 U7420 ( .A1(n14566), .A2(n14565), .ZN(n14687) );
  NAND2_X1 U7421 ( .A1(n14098), .A2(n14316), .ZN(n7002) );
  NAND2_X1 U7422 ( .A1(n11466), .A2(n11465), .ZN(n13303) );
  INV_X1 U7423 ( .A(n14990), .ZN(n6832) );
  AND2_X1 U7424 ( .A1(n6934), .A2(n6932), .ZN(n14573) );
  NAND2_X1 U7425 ( .A1(n12758), .A2(n12757), .ZN(n12766) );
  NAND2_X1 U7426 ( .A1(n12444), .A2(n12075), .ZN(n12430) );
  OAI22_X1 U7427 ( .A1(n12085), .A2(n12420), .B1(n12094), .B2(n12084), .ZN(
        n12091) );
  NAND2_X1 U7428 ( .A1(n12446), .A2(n12445), .ZN(n12444) );
  INV_X1 U7429 ( .A(n12321), .ZN(n6554) );
  NAND2_X1 U7430 ( .A1(n11309), .A2(n11308), .ZN(n11673) );
  AND2_X1 U7431 ( .A1(n6820), .A2(n6819), .ZN(n14839) );
  NAND2_X1 U7432 ( .A1(n7602), .A2(n7600), .ZN(n12446) );
  OAI22_X1 U7433 ( .A1(n6639), .A2(n7524), .B1(n14154), .B2(n7526), .ZN(n14157) );
  NAND2_X1 U7434 ( .A1(n6904), .A2(n11121), .ZN(n11270) );
  NAND2_X1 U7435 ( .A1(n12477), .A2(n12476), .ZN(n12475) );
  OR2_X1 U7436 ( .A1(n14821), .A2(n14822), .ZN(n7455) );
  AND2_X1 U7437 ( .A1(n14822), .A2(n14821), .ZN(n14880) );
  OAI21_X1 U7438 ( .B1(n12914), .B2(n7663), .A(n6985), .ZN(n12920) );
  OR2_X1 U7439 ( .A1(n10711), .A2(n10712), .ZN(n10671) );
  NAND2_X1 U7440 ( .A1(n6556), .A2(n7595), .ZN(n10769) );
  AND2_X1 U7441 ( .A1(n7247), .A2(n7246), .ZN(n6830) );
  NAND2_X1 U7442 ( .A1(n10782), .A2(n7593), .ZN(n6556) );
  NAND2_X1 U7443 ( .A1(n6741), .A2(n6586), .ZN(n11108) );
  OR2_X1 U7444 ( .A1(n15085), .A2(n15095), .ZN(n15087) );
  NAND2_X1 U7445 ( .A1(n12635), .A2(n10124), .ZN(n10284) );
  AND3_X1 U7446 ( .A1(n7230), .A2(n7229), .A3(n10017), .ZN(n10651) );
  NAND2_X1 U7447 ( .A1(n7585), .A2(SI_18_), .ZN(n7819) );
  AND2_X1 U7448 ( .A1(n12041), .A2(n12040), .ZN(n12038) );
  NOR2_X1 U7449 ( .A1(n14779), .A2(n14778), .ZN(n14818) );
  OAI21_X1 U7450 ( .B1(n9758), .B2(n7922), .A(n7923), .ZN(n9929) );
  NAND2_X1 U7451 ( .A1(n13472), .A2(n10348), .ZN(n13465) );
  NAND2_X1 U7452 ( .A1(n8483), .A2(n12003), .ZN(n6558) );
  OAI21_X1 U7453 ( .B1(n8042), .B2(n6773), .A(n6770), .ZN(n8117) );
  NAND2_X1 U7454 ( .A1(n9871), .A2(n12479), .ZN(n11933) );
  NAND2_X2 U7455 ( .A1(n10345), .A2(n13397), .ZN(n13472) );
  AND2_X1 U7456 ( .A1(n12018), .A2(n12011), .ZN(n12012) );
  OAI21_X2 U7457 ( .B1(n9397), .B2(n15092), .A(n15091), .ZN(n9398) );
  INV_X2 U7458 ( .A(n15104), .ZN(n15106) );
  NAND2_X1 U7459 ( .A1(n7070), .A2(n8571), .ZN(n12175) );
  NOR2_X1 U7460 ( .A1(n12182), .A2(n11559), .ZN(n11991) );
  NAND2_X2 U7461 ( .A1(n9863), .A2(n12616), .ZN(n11655) );
  NAND2_X1 U7462 ( .A1(n7932), .A2(n7931), .ZN(n15152) );
  NAND2_X1 U7463 ( .A1(n8426), .A2(n8425), .ZN(n8634) );
  NAND2_X1 U7464 ( .A1(n6979), .A2(n7878), .ZN(n13965) );
  XNOR2_X1 U7465 ( .A(n14767), .B(n14768), .ZN(n14803) );
  AND3_X1 U7466 ( .A1(n8495), .A2(n8494), .A3(n8496), .ZN(n10244) );
  INV_X1 U7467 ( .A(n8611), .ZN(n8426) );
  INV_X1 U7468 ( .A(n8991), .ZN(n14338) );
  OR2_X1 U7469 ( .A1(n6956), .A2(n6784), .ZN(n13209) );
  AND2_X1 U7470 ( .A1(n8457), .A2(n8456), .ZN(n11559) );
  INV_X1 U7471 ( .A(n9796), .ZN(n12667) );
  AND2_X1 U7472 ( .A1(n6828), .A2(n6822), .ZN(n14767) );
  AND4_X1 U7473 ( .A1(n7921), .A2(n7920), .A3(n7919), .A4(n7918), .ZN(n14122)
         );
  NAND4_X1 U7474 ( .A1(n7901), .A2(n7900), .A3(n7899), .A4(n7898), .ZN(n14335)
         );
  AND2_X1 U7475 ( .A1(n9391), .A2(n9012), .ZN(n14554) );
  INV_X2 U7476 ( .A(n14242), .ZN(n14087) );
  BUF_X2 U7477 ( .A(n8486), .Z(n6568) );
  OR2_X1 U7478 ( .A1(n8503), .A2(n9068), .ZN(n8465) );
  AND4_X1 U7480 ( .A1(n7883), .A2(n7882), .A3(n7881), .A4(n7880), .ZN(n8991)
         );
  MUX2_X1 U7481 ( .A(n14085), .B(n14084), .S(n7523), .Z(n14123) );
  NAND2_X2 U7482 ( .A1(n8999), .A2(n9293), .ZN(n14242) );
  OAI21_X1 U7483 ( .B1(n8538), .B2(n8358), .A(n8359), .ZN(n8549) );
  INV_X2 U7484 ( .A(n14076), .ZN(n8267) );
  INV_X1 U7485 ( .A(n11502), .ZN(n11492) );
  OR2_X1 U7486 ( .A1(n6825), .A2(n14764), .ZN(n6824) );
  NAND2_X2 U7487 ( .A1(n12163), .A2(n8876), .ZN(n12129) );
  BUF_X2 U7488 ( .A(n9307), .Z(n13072) );
  OR2_X2 U7489 ( .A1(n14091), .A2(n14084), .ZN(n14589) );
  AND2_X1 U7490 ( .A1(n15314), .A2(n10346), .ZN(n12868) );
  AND2_X1 U7491 ( .A1(n7721), .A2(n7718), .ZN(n14084) );
  INV_X1 U7492 ( .A(n12628), .ZN(n8444) );
  XNOR2_X1 U7493 ( .A(n8415), .B(n8414), .ZN(n8875) );
  XNOR2_X1 U7494 ( .A(n7726), .B(n7725), .ZN(n14085) );
  NAND2_X1 U7495 ( .A1(n8408), .A2(n6548), .ZN(n12620) );
  NAND2_X1 U7496 ( .A1(n8890), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U7497 ( .A1(n7718), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U7498 ( .A1(n7724), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U7499 ( .A1(n7754), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U7500 ( .A1(n14737), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7753) );
  CLKBUF_X1 U7501 ( .A(n9264), .Z(n6561) );
  NAND2_X1 U7502 ( .A1(n13880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7660) );
  XNOR2_X1 U7503 ( .A(n7130), .B(n7844), .ZN(n15001) );
  CLKBUF_X1 U7504 ( .A(n13156), .Z(n6984) );
  NAND2_X1 U7505 ( .A1(n7131), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7130) );
  NAND2_X1 U7506 ( .A1(n8408), .A2(n7074), .ZN(n8442) );
  INV_X2 U7507 ( .A(n12617), .ZN(n12627) );
  NOR2_X1 U7508 ( .A1(n6661), .A2(n7075), .ZN(n7074) );
  OAI21_X1 U7509 ( .B1(n9656), .B2(n7480), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6841) );
  NOR2_X1 U7510 ( .A1(n9656), .A2(n7478), .ZN(n8966) );
  NAND2_X1 U7511 ( .A1(n9212), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9210) );
  NAND2_X2 U7512 ( .A1(n13064), .A2(P3_U3151), .ZN(n12623) );
  AND2_X1 U7513 ( .A1(n7362), .A2(n7627), .ZN(n7363) );
  AND2_X1 U7514 ( .A1(n8479), .A2(n6755), .ZN(n9664) );
  NAND2_X1 U7515 ( .A1(n9502), .A2(n8973), .ZN(n9656) );
  NOR2_X1 U7516 ( .A1(n8323), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7365) );
  NOR2_X1 U7517 ( .A1(n7628), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n7627) );
  AND2_X1 U7518 ( .A1(n6626), .A2(n7844), .ZN(n7658) );
  AND4_X1 U7519 ( .A1(n8973), .A2(n6630), .A3(n8972), .A4(n8971), .ZN(n8974)
         );
  AND3_X1 U7520 ( .A1(n9372), .A2(n9049), .A3(n8961), .ZN(n8975) );
  AND2_X1 U7521 ( .A1(n7631), .A2(n8414), .ZN(n7630) );
  AND3_X1 U7522 ( .A1(n8960), .A2(n8959), .A3(n9089), .ZN(n9372) );
  AND3_X1 U7523 ( .A1(n6840), .A2(n6839), .A3(n9057), .ZN(n8961) );
  AND2_X1 U7524 ( .A1(n13813), .A2(n8970), .ZN(n7489) );
  AND4_X1 U7525 ( .A1(n7712), .A2(n7711), .A3(n7710), .A4(n7709), .ZN(n7688)
         );
  AND2_X1 U7526 ( .A1(n8410), .A2(n8411), .ZN(n7631) );
  AND3_X1 U7527 ( .A1(n8327), .A2(n8328), .A3(n8326), .ZN(n8330) );
  INV_X1 U7528 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7128) );
  INV_X4 U7529 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7530 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8331) );
  NOR2_X1 U7531 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n8326) );
  NOR2_X2 U7532 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n7712) );
  NOR2_X1 U7533 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7699) );
  NOR2_X1 U7534 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n7700) );
  INV_X1 U7535 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n13831) );
  NOR2_X1 U7536 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8328) );
  INV_X1 U7537 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8414) );
  INV_X1 U7538 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7988) );
  INV_X1 U7539 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8409) );
  INV_X1 U7540 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8003) );
  INV_X1 U7541 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7709) );
  NOR2_X1 U7542 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7502) );
  NOR2_X1 U7543 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7501) );
  NOR2_X1 U7544 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7500) );
  NOR2_X1 U7545 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8327) );
  INV_X1 U7546 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n7063) );
  INV_X1 U7547 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7725) );
  NOR2_X1 U7548 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8322) );
  NOR2_X1 U7549 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n8960) );
  NOR2_X1 U7550 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8959) );
  INV_X1 U7551 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9261) );
  INV_X1 U7552 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8964) );
  NOR2_X1 U7553 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8963) );
  NOR2_X1 U7554 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8962) );
  INV_X1 U7555 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8324) );
  INV_X1 U7556 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9593) );
  INV_X1 U7557 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14760) );
  INV_X4 U7558 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7559 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9044) );
  INV_X1 U7560 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9045) );
  INV_X4 U7561 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7562 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9089) );
  OR2_X2 U7563 ( .A1(n11339), .A2(n11340), .ZN(n11341) );
  NAND2_X1 U7564 ( .A1(n12430), .A2(n12429), .ZN(n12428) );
  NAND2_X1 U7565 ( .A1(n10741), .A2(n10743), .ZN(n6557) );
  OR2_X2 U7566 ( .A1(n12368), .A2(n12370), .ZN(n12366) );
  NAND2_X1 U7567 ( .A1(n7621), .A2(n6683), .ZN(n12391) );
  NAND2_X1 U7568 ( .A1(n6558), .A2(n10224), .ZN(n8497) );
  XNOR2_X1 U7569 ( .A(n6558), .B(n6966), .ZN(n15476) );
  NAND3_X1 U7570 ( .A1(n7353), .A2(n7354), .A3(n7357), .ZN(n7352) );
  NOR2_X2 U7571 ( .A1(n7445), .A2(n14993), .ZN(n14996) );
  XNOR2_X1 U7572 ( .A(n7238), .B(n6608), .ZN(n14893) );
  NOR2_X2 U7573 ( .A1(n10834), .A2(n13582), .ZN(n7228) );
  AND4_X2 U7574 ( .A1(n9372), .A2(n9049), .A3(n7489), .A4(n8961), .ZN(n9502)
         );
  INV_X2 U7575 ( .A(n14111), .ZN(n9725) );
  INV_X4 U7576 ( .A(n9296), .ZN(n9306) );
  OAI21_X1 U7577 ( .B1(n14892), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n6615), .ZN(
        n7238) );
  XNOR2_X2 U7578 ( .A(n14862), .B(n14861), .ZN(n14892) );
  XNOR2_X1 U7579 ( .A(n6623), .B(n6759), .ZN(n9452) );
  OR2_X1 U7580 ( .A1(n13166), .A2(n13161), .ZN(n13181) );
  AOI21_X2 U7581 ( .B1(n11021), .B2(n11969), .A(n8596), .ZN(n11113) );
  NAND2_X2 U7582 ( .A1(n11996), .A2(n11995), .ZN(n9866) );
  OAI222_X1 U7583 ( .A1(n12623), .A2(n11950), .B1(P3_U3151), .B2(n11337), .C1(
        n12627), .C2(n11336), .ZN(P3_U3265) );
  XNOR2_X2 U7584 ( .A(n9209), .B(P2_IR_REG_21__SCAN_IN), .ZN(n10346) );
  XNOR2_X2 U7585 ( .A(n7753), .B(n6953), .ZN(n14743) );
  XNOR2_X2 U7586 ( .A(n7843), .B(n7842), .ZN(n11338) );
  INV_X1 U7587 ( .A(n15001), .ZN(n6559) );
  INV_X1 U7588 ( .A(n6559), .ZN(n6560) );
  NAND3_X1 U7589 ( .A1(n7156), .A2(n9466), .A3(n9467), .ZN(n13210) );
  NAND2_X1 U7590 ( .A1(n8875), .A2(n11081), .ZN(n6562) );
  NAND2_X2 U7591 ( .A1(n8875), .A2(n11081), .ZN(n6563) );
  NAND2_X1 U7592 ( .A1(n8875), .A2(n11081), .ZN(n9535) );
  AND3_X2 U7593 ( .A1(n12139), .A2(n12138), .A3(n12137), .ZN(n12140) );
  INV_X1 U7594 ( .A(n8518), .ZN(n6564) );
  NAND2_X1 U7595 ( .A1(n9783), .A2(n9293), .ZN(n6565) );
  AOI21_X1 U7596 ( .B1(n7790), .B2(n7567), .A(n6660), .ZN(n7566) );
  INV_X1 U7597 ( .A(n7788), .ZN(n7567) );
  OAI21_X1 U7598 ( .B1(n8369), .B2(n7312), .A(n7309), .ZN(n8373) );
  INV_X1 U7599 ( .A(n7313), .ZN(n7312) );
  AOI21_X1 U7600 ( .B1(n7311), .B2(n7313), .A(n7310), .ZN(n7309) );
  INV_X1 U7601 ( .A(n8372), .ZN(n7310) );
  NOR2_X1 U7602 ( .A1(n11530), .A2(n7430), .ZN(n7429) );
  INV_X1 U7603 ( .A(n11529), .ZN(n7430) );
  NOR2_X1 U7604 ( .A1(n7438), .A2(n10837), .ZN(n7437) );
  INV_X1 U7605 ( .A(n10584), .ZN(n7438) );
  NAND2_X1 U7606 ( .A1(n6878), .A2(n6877), .ZN(n15067) );
  AOI21_X1 U7607 ( .B1(n6880), .B2(n6882), .A(n6650), .ZN(n6877) );
  NAND2_X1 U7608 ( .A1(n10094), .A2(n6880), .ZN(n6878) );
  NOR2_X1 U7609 ( .A1(n14488), .A2(n7514), .ZN(n7512) );
  NAND2_X1 U7610 ( .A1(n6760), .A2(n7822), .ZN(n7823) );
  NAND2_X1 U7611 ( .A1(n8153), .A2(n6642), .ZN(n6760) );
  OR2_X1 U7612 ( .A1(n12295), .A2(n11860), .ZN(n12135) );
  AOI21_X1 U7613 ( .B1(n7167), .B2(n6576), .A(n7165), .ZN(n7164) );
  NOR2_X1 U7614 ( .A1(n13340), .A2(n13189), .ZN(n7165) );
  AOI21_X1 U7615 ( .B1(n7421), .B2(n7420), .A(n6692), .ZN(n7419) );
  INV_X1 U7616 ( .A(n11523), .ZN(n7420) );
  INV_X2 U7617 ( .A(n13082), .ZN(n13068) );
  NAND2_X1 U7618 ( .A1(n10643), .A2(n7437), .ZN(n7435) );
  NAND2_X1 U7619 ( .A1(n9783), .A2(n9293), .ZN(n13083) );
  NAND2_X1 U7620 ( .A1(n9783), .A2(n13064), .ZN(n13082) );
  NAND2_X2 U7621 ( .A1(n9220), .A2(n9215), .ZN(n9783) );
  NAND2_X1 U7622 ( .A1(n7506), .A2(n6647), .ZN(n11568) );
  NAND2_X1 U7623 ( .A1(n8153), .A2(n7819), .ZN(n8170) );
  INV_X1 U7624 ( .A(n12895), .ZN(n6958) );
  NAND2_X1 U7625 ( .A1(n12901), .A2(n12902), .ZN(n6861) );
  INV_X1 U7626 ( .A(n12901), .ZN(n6865) );
  NAND2_X1 U7627 ( .A1(n14129), .A2(n14128), .ZN(n14132) );
  NAND2_X1 U7628 ( .A1(n7000), .A2(n12964), .ZN(n6852) );
  AND2_X1 U7629 ( .A1(n13009), .A2(n13010), .ZN(n6866) );
  NAND2_X1 U7630 ( .A1(n14213), .A2(n7531), .ZN(n7528) );
  INV_X1 U7631 ( .A(n14214), .ZN(n7531) );
  NAND2_X1 U7632 ( .A1(n6674), .A2(n7676), .ZN(n7675) );
  NAND2_X1 U7633 ( .A1(n7146), .A2(n14223), .ZN(n14227) );
  AND2_X1 U7634 ( .A1(n14230), .A2(n7520), .ZN(n7519) );
  INV_X1 U7635 ( .A(n14228), .ZN(n7520) );
  NAND2_X1 U7636 ( .A1(n6910), .A2(n13965), .ZN(n14107) );
  INV_X1 U7637 ( .A(n7723), .ZN(n7722) );
  NAND2_X1 U7638 ( .A1(n7781), .A2(n6583), .ZN(n6766) );
  NAND2_X1 U7639 ( .A1(n6765), .A2(n6580), .ZN(n6764) );
  OR2_X1 U7640 ( .A1(n7956), .A2(n6767), .ZN(n6765) );
  INV_X1 U7641 ( .A(n7459), .ZN(n14763) );
  INV_X1 U7642 ( .A(n11337), .ZN(n8443) );
  OR2_X1 U7643 ( .A1(n11878), .A2(n12335), .ZN(n12119) );
  OR2_X1 U7644 ( .A1(n8856), .A2(n12372), .ZN(n11965) );
  AND2_X1 U7645 ( .A1(n7605), .A2(n6681), .ZN(n7603) );
  AND2_X1 U7646 ( .A1(n7348), .A2(n7346), .ZN(n7345) );
  AND2_X1 U7647 ( .A1(n15507), .A2(n12175), .ZN(n7350) );
  INV_X1 U7648 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U7649 ( .A1(n9084), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U7650 ( .A1(n12676), .A2(n12675), .ZN(n7465) );
  OR2_X1 U7651 ( .A1(n13490), .A2(n11540), .ZN(n11500) );
  NAND2_X1 U7652 ( .A1(n13281), .A2(n6758), .ZN(n13264) );
  AND2_X1 U7653 ( .A1(n13265), .A2(n13266), .ZN(n6758) );
  OAI21_X1 U7654 ( .B1(n6610), .B2(n7159), .A(n11390), .ZN(n7158) );
  INV_X1 U7655 ( .A(n13470), .ZN(n9459) );
  XNOR2_X1 U7656 ( .A(n13470), .B(n13212), .ZN(n13120) );
  AOI21_X1 U7657 ( .B1(n10904), .B2(n13136), .A(n10903), .ZN(n10998) );
  INV_X1 U7658 ( .A(n6903), .ZN(n6902) );
  MUX2_X1 U7659 ( .A(n14415), .B(n14247), .S(n14206), .Z(n14259) );
  NAND2_X1 U7660 ( .A1(n7523), .A2(n15140), .ZN(n14249) );
  INV_X1 U7661 ( .A(n14746), .ZN(n7756) );
  NAND2_X1 U7662 ( .A1(n14508), .A2(n7406), .ZN(n7405) );
  NOR2_X1 U7663 ( .A1(n14493), .A2(n7407), .ZN(n7406) );
  INV_X1 U7664 ( .A(n7689), .ZN(n7407) );
  NAND2_X1 U7665 ( .A1(n7396), .A2(n7256), .ZN(n6917) );
  NAND2_X1 U7666 ( .A1(n6917), .A2(n8220), .ZN(n6916) );
  INV_X1 U7667 ( .A(n14329), .ZN(n10879) );
  INV_X1 U7668 ( .A(n14295), .ZN(n11569) );
  OAI21_X1 U7669 ( .B1(n8262), .B2(n8261), .A(n8263), .ZN(n13060) );
  OR2_X1 U7670 ( .A1(n7859), .A2(n7858), .ZN(n7861) );
  NAND2_X1 U7671 ( .A1(n8196), .A2(n8195), .ZN(n8198) );
  XNOR2_X1 U7672 ( .A(n7791), .B(SI_9_), .ZN(n7986) );
  NAND2_X1 U7673 ( .A1(n7781), .A2(n7780), .ZN(n7944) );
  XNOR2_X1 U7674 ( .A(n7774), .B(SI_3_), .ZN(n7904) );
  NAND2_X1 U7675 ( .A1(n7772), .A2(n7771), .ZN(n7905) );
  AOI22_X1 U7676 ( .A1(n14850), .A2(n14849), .B1(P1_ADDR_REG_14__SCAN_IN), 
        .B2(n14848), .ZN(n14856) );
  NOR2_X1 U7677 ( .A1(n11824), .A2(n7095), .ZN(n7094) );
  INV_X1 U7678 ( .A(n7097), .ZN(n7095) );
  NAND2_X1 U7679 ( .A1(n6562), .A2(n13064), .ZN(n8518) );
  NAND2_X1 U7680 ( .A1(n9843), .A2(n12182), .ZN(n8835) );
  NAND3_X1 U7681 ( .A1(n10553), .A2(n10217), .A3(n6575), .ZN(n7078) );
  NOR2_X1 U7682 ( .A1(n7376), .A2(n6648), .ZN(n7374) );
  AOI22_X1 U7683 ( .A1(n11865), .A2(n11864), .B1(n12452), .B2(n11630), .ZN(
        n11871) );
  NAND2_X1 U7684 ( .A1(n7335), .A2(n11242), .ZN(n12184) );
  NAND2_X1 U7685 ( .A1(n6731), .A2(n6730), .ZN(n12232) );
  INV_X1 U7686 ( .A(n12211), .ZN(n6730) );
  NOR2_X1 U7687 ( .A1(n11983), .A2(n7625), .ZN(n7624) );
  INV_X1 U7688 ( .A(n12135), .ZN(n7625) );
  OAI22_X1 U7689 ( .A1(n12346), .A2(n8858), .B1(n11905), .B2(n12171), .ZN(
        n12333) );
  INV_X1 U7690 ( .A(n12372), .ZN(n12348) );
  INV_X1 U7691 ( .A(n6737), .ZN(n6736) );
  OAI21_X1 U7692 ( .B1(n7341), .B2(n6738), .A(n12370), .ZN(n6737) );
  INV_X1 U7693 ( .A(n7054), .ZN(n6738) );
  NAND2_X1 U7694 ( .A1(n12399), .A2(n7341), .ZN(n12384) );
  OR2_X1 U7695 ( .A1(n12535), .A2(n12434), .ZN(n12084) );
  NAND2_X1 U7696 ( .A1(n12419), .A2(n8854), .ZN(n12401) );
  OR2_X1 U7697 ( .A1(n12535), .A2(n12405), .ZN(n8854) );
  OR2_X1 U7698 ( .A1(n11625), .A2(n12605), .ZN(n8851) );
  XNOR2_X1 U7699 ( .A(n12177), .B(n10796), .ZN(n12027) );
  NAND3_X1 U7700 ( .A1(n7118), .A2(n7117), .A3(n9716), .ZN(n12151) );
  OR2_X1 U7701 ( .A1(n8329), .A2(n7123), .ZN(n7118) );
  NAND2_X1 U7702 ( .A1(n7124), .A2(n7127), .ZN(n7123) );
  INV_X1 U7703 ( .A(n11344), .ZN(n7355) );
  NAND2_X1 U7704 ( .A1(n8917), .A2(n8900), .ZN(n8915) );
  NAND2_X1 U7705 ( .A1(n8402), .A2(n8401), .ZN(n8405) );
  NAND2_X1 U7706 ( .A1(n7289), .A2(n7285), .ZN(n8402) );
  NAND2_X1 U7707 ( .A1(n8329), .A2(n7126), .ZN(n7119) );
  OR2_X1 U7708 ( .A1(n8329), .A2(n7127), .ZN(n7120) );
  INV_X1 U7709 ( .A(n7302), .ZN(n7301) );
  OAI21_X1 U7710 ( .B1(n8696), .B2(n7303), .A(n8711), .ZN(n7302) );
  AND2_X1 U7711 ( .A1(n8377), .A2(n8376), .ZN(n8640) );
  NAND2_X1 U7712 ( .A1(n8369), .A2(n7318), .ZN(n7315) );
  AOI21_X1 U7713 ( .B1(n8564), .B2(n7282), .A(n7280), .ZN(n7279) );
  OR2_X1 U7714 ( .A1(n8565), .A2(n7281), .ZN(n7278) );
  INV_X1 U7715 ( .A(n8366), .ZN(n7280) );
  NAND2_X1 U7716 ( .A1(n8565), .A2(n8363), .ZN(n7284) );
  INV_X1 U7717 ( .A(n12667), .ZN(n12732) );
  OAI211_X1 U7718 ( .C1(n6613), .C2(n7030), .A(n7028), .B(n7041), .ZN(n7027)
         );
  OR2_X1 U7719 ( .A1(n12680), .A2(n12679), .ZN(n7041) );
  NAND2_X1 U7720 ( .A1(n7466), .A2(n7465), .ZN(n7030) );
  NAND2_X1 U7721 ( .A1(n7032), .A2(n7029), .ZN(n7028) );
  NAND2_X1 U7722 ( .A1(n12776), .A2(n7470), .ZN(n12715) );
  NAND2_X1 U7723 ( .A1(n6991), .A2(n6988), .ZN(n9220) );
  NAND2_X1 U7724 ( .A1(n9211), .A2(n6978), .ZN(n6991) );
  NOR2_X1 U7725 ( .A1(n6990), .A2(n6989), .ZN(n6988) );
  NOR2_X1 U7726 ( .A1(n6992), .A2(n13881), .ZN(n6978) );
  NAND2_X1 U7727 ( .A1(n13071), .A2(n13070), .ZN(n13253) );
  INV_X1 U7728 ( .A(n13148), .ZN(n13265) );
  NAND2_X1 U7729 ( .A1(n7167), .A2(n6602), .ZN(n7166) );
  INV_X1 U7730 ( .A(n11417), .ZN(n7170) );
  NAND2_X1 U7731 ( .A1(n13370), .A2(n13361), .ZN(n13355) );
  AOI21_X1 U7732 ( .B1(n7429), .B2(n11528), .A(n6588), .ZN(n7428) );
  INV_X1 U7733 ( .A(n13364), .ZN(n7172) );
  NAND2_X1 U7734 ( .A1(n11527), .A2(n11526), .ZN(n13389) );
  OAI21_X1 U7735 ( .B1(n11353), .B2(n7387), .A(n7389), .ZN(n11368) );
  OR2_X1 U7736 ( .A1(n11352), .A2(n7388), .ZN(n7387) );
  AOI21_X1 U7737 ( .B1(n6573), .B2(n11357), .A(n6653), .ZN(n7389) );
  INV_X1 U7738 ( .A(n11357), .ZN(n7388) );
  NAND2_X1 U7739 ( .A1(n11356), .A2(n11355), .ZN(n13460) );
  NAND2_X1 U7740 ( .A1(n11522), .A2(n11521), .ZN(n13445) );
  AOI21_X1 U7741 ( .B1(n7437), .B2(n10583), .A(n6663), .ZN(n7436) );
  NAND2_X1 U7742 ( .A1(n10578), .A2(n10577), .ZN(n10643) );
  NOR2_X2 U7743 ( .A1(n10471), .A2(n15370), .ZN(n10470) );
  INV_X1 U7744 ( .A(n13332), .ZN(n13513) );
  NAND2_X1 U7745 ( .A1(n15314), .A2(n12867), .ZN(n15423) );
  NAND2_X1 U7746 ( .A1(n7202), .A2(n10034), .ZN(n7201) );
  INV_X1 U7747 ( .A(n7213), .ZN(n7212) );
  NAND2_X1 U7748 ( .A1(n11792), .A2(n7216), .ZN(n7214) );
  NAND2_X1 U7749 ( .A1(n14022), .A2(n14021), .ZN(n11729) );
  AND2_X1 U7750 ( .A1(n7636), .A2(n14014), .ZN(n7635) );
  NAND2_X1 U7751 ( .A1(n7638), .A2(n7641), .ZN(n7636) );
  NAND2_X1 U7752 ( .A1(n10039), .A2(n10040), .ZN(n7653) );
  OAI21_X1 U7753 ( .B1(n10537), .B2(n7220), .A(n7217), .ZN(n11120) );
  AOI21_X1 U7754 ( .B1(n7218), .B2(n7219), .A(n6676), .ZN(n7217) );
  INV_X1 U7755 ( .A(n10536), .ZN(n7218) );
  NAND2_X1 U7756 ( .A1(n7650), .A2(n7649), .ZN(n7652) );
  NAND2_X1 U7757 ( .A1(n13980), .A2(n13982), .ZN(n11773) );
  AND2_X1 U7758 ( .A1(n14051), .A2(n7645), .ZN(n7644) );
  NAND2_X1 U7759 ( .A1(n7646), .A2(n11774), .ZN(n7645) );
  INV_X1 U7760 ( .A(n11774), .ZN(n7647) );
  AND3_X1 U7761 ( .A1(n7937), .A2(n6889), .A3(n7940), .ZN(n10189) );
  AND2_X1 U7762 ( .A1(n7939), .A2(n7938), .ZN(n6889) );
  NOR2_X1 U7763 ( .A1(n14450), .A2(n7505), .ZN(n7504) );
  INV_X1 U7764 ( .A(n7507), .ZN(n7505) );
  XNOR2_X1 U7765 ( .A(n14644), .B(n14317), .ZN(n14450) );
  NAND2_X1 U7766 ( .A1(n14467), .A2(n6640), .ZN(n14454) );
  NAND2_X1 U7767 ( .A1(n14454), .A2(n14453), .ZN(n14452) );
  NAND2_X1 U7768 ( .A1(n7405), .A2(n7403), .ZN(n14470) );
  AND2_X1 U7769 ( .A1(n14471), .A2(n7404), .ZN(n7403) );
  INV_X1 U7770 ( .A(n7408), .ZN(n7404) );
  AND2_X1 U7771 ( .A1(n14497), .A2(n14476), .ZN(n8301) );
  XNOR2_X1 U7772 ( .A(n14664), .B(n14476), .ZN(n14493) );
  INV_X1 U7773 ( .A(n7405), .ZN(n14491) );
  NAND2_X1 U7774 ( .A1(n8299), .A2(n8298), .ZN(n14505) );
  OAI21_X1 U7775 ( .B1(n14687), .B2(n7253), .A(n7251), .ZN(n8299) );
  INV_X1 U7776 ( .A(n7252), .ZN(n7251) );
  OR2_X1 U7777 ( .A1(n14505), .A2(n14509), .ZN(n14507) );
  OR2_X1 U7778 ( .A1(n14944), .A2(n11690), .ZN(n14173) );
  AND2_X1 U7779 ( .A1(n14165), .A2(n8072), .ZN(n7409) );
  NAND2_X1 U7780 ( .A1(n6871), .A2(n6868), .ZN(n8289) );
  AOI21_X1 U7781 ( .B1(n7490), .B2(n6870), .A(n6869), .ZN(n6868) );
  NOR2_X2 U7782 ( .A1(n11030), .A2(n14961), .ZN(n11029) );
  NAND2_X1 U7783 ( .A1(n15087), .A2(n7385), .ZN(n15064) );
  NOR2_X1 U7784 ( .A1(n14280), .A2(n7386), .ZN(n7385) );
  INV_X1 U7785 ( .A(n7985), .ZN(n7386) );
  OR2_X2 U7786 ( .A1(n15098), .A2(n15076), .ZN(n15078) );
  NAND2_X1 U7787 ( .A1(n8281), .A2(n8280), .ZN(n10094) );
  INV_X1 U7788 ( .A(n14554), .ZN(n14606) );
  NAND2_X1 U7789 ( .A1(n6926), .A2(n7907), .ZN(n9758) );
  INV_X1 U7790 ( .A(n14608), .ZN(n15059) );
  NAND2_X1 U7791 ( .A1(n6763), .A2(n6762), .ZN(n8153) );
  INV_X1 U7792 ( .A(n8150), .ZN(n6762) );
  NAND2_X1 U7793 ( .A1(n7815), .A2(n7814), .ZN(n8136) );
  XNOR2_X1 U7794 ( .A(n8027), .B(n8026), .ZN(n10579) );
  INV_X1 U7795 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7246) );
  INV_X1 U7796 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7243) );
  NAND2_X1 U7797 ( .A1(n13894), .A2(n13068), .ZN(n6768) );
  NAND2_X1 U7798 ( .A1(n12870), .A2(n12869), .ZN(n6976) );
  NAND2_X1 U7799 ( .A1(n12877), .A2(n6960), .ZN(n12882) );
  OR2_X1 U7800 ( .A1(n12878), .A2(n12876), .ZN(n12874) );
  INV_X1 U7801 ( .A(n12890), .ZN(n6968) );
  NAND2_X1 U7802 ( .A1(n6864), .A2(n6862), .ZN(n12907) );
  NAND2_X1 U7803 ( .A1(n6865), .A2(n6863), .ZN(n6862) );
  INV_X1 U7804 ( .A(n12902), .ZN(n6863) );
  INV_X1 U7805 ( .A(n12912), .ZN(n6986) );
  INV_X1 U7806 ( .A(n12913), .ZN(n6987) );
  NAND2_X1 U7807 ( .A1(n6844), .A2(n6843), .ZN(n12934) );
  AOI21_X1 U7808 ( .B1(n6609), .B2(n6847), .A(n6590), .ZN(n6843) );
  NAND2_X1 U7809 ( .A1(n12920), .A2(n6609), .ZN(n6844) );
  AND2_X1 U7810 ( .A1(n12921), .A2(n6848), .ZN(n6847) );
  NAND2_X1 U7811 ( .A1(n14154), .A2(n7526), .ZN(n7525) );
  NAND2_X1 U7812 ( .A1(n7679), .A2(n12938), .ZN(n7678) );
  INV_X1 U7813 ( .A(n6697), .ZN(n7679) );
  NAND2_X1 U7814 ( .A1(n6858), .A2(n6857), .ZN(n12955) );
  AOI21_X1 U7815 ( .B1(n6577), .B2(n6860), .A(n6571), .ZN(n6857) );
  NAND2_X1 U7816 ( .A1(n12944), .A2(n6577), .ZN(n6858) );
  NOR2_X1 U7817 ( .A1(n6612), .A2(n12943), .ZN(n6860) );
  INV_X1 U7818 ( .A(n12963), .ZN(n7000) );
  NAND2_X1 U7819 ( .A1(n7139), .A2(n7138), .ZN(n7137) );
  INV_X1 U7820 ( .A(n14199), .ZN(n7139) );
  INV_X1 U7821 ( .A(n14201), .ZN(n7138) );
  NAND2_X1 U7822 ( .A1(n13031), .A2(n7670), .ZN(n7669) );
  NAND2_X1 U7823 ( .A1(n7672), .A2(n7671), .ZN(n7670) );
  INV_X1 U7824 ( .A(n14220), .ZN(n7148) );
  INV_X1 U7825 ( .A(n14221), .ZN(n7552) );
  INV_X1 U7826 ( .A(n7692), .ZN(n7573) );
  AOI21_X1 U7827 ( .B1(n7692), .B2(n7572), .A(n7571), .ZN(n7570) );
  INV_X1 U7828 ( .A(n7806), .ZN(n7571) );
  INV_X1 U7829 ( .A(n7802), .ZN(n7572) );
  OR2_X1 U7830 ( .A1(n8864), .A2(n11586), .ZN(n11592) );
  NAND2_X1 U7831 ( .A1(n7545), .A2(n14239), .ZN(n7544) );
  AND2_X1 U7832 ( .A1(n14238), .A2(n7547), .ZN(n7546) );
  INV_X1 U7833 ( .A(n14239), .ZN(n7547) );
  INV_X1 U7834 ( .A(n7836), .ZN(n7588) );
  NAND2_X1 U7835 ( .A1(n7816), .A2(n9512), .ZN(n7584) );
  AOI21_X1 U7836 ( .B1(n7809), .B2(n8097), .A(n8095), .ZN(n7810) );
  INV_X1 U7837 ( .A(n7570), .ZN(n6772) );
  OAI21_X1 U7838 ( .B1(n13064), .B2(n13630), .A(n6974), .ZN(n7783) );
  NAND2_X1 U7839 ( .A1(n13064), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6974) );
  INV_X1 U7840 ( .A(n7412), .ZN(n6776) );
  OAI21_X1 U7841 ( .B1(n14788), .B2(n14787), .A(n7460), .ZN(n7459) );
  NAND2_X1 U7842 ( .A1(n14761), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7460) );
  NAND2_X1 U7843 ( .A1(n11633), .A2(n12422), .ZN(n7116) );
  NAND2_X1 U7844 ( .A1(n11654), .A2(n7369), .ZN(n7368) );
  INV_X1 U7845 ( .A(n7109), .ZN(n7108) );
  NAND2_X1 U7846 ( .A1(n7340), .A2(n7339), .ZN(n6729) );
  NAND2_X1 U7847 ( .A1(n9670), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7339) );
  NOR2_X1 U7848 ( .A1(n9668), .A2(n6646), .ZN(n9701) );
  NAND2_X1 U7849 ( .A1(n9824), .A2(n9823), .ZN(n6733) );
  INV_X1 U7850 ( .A(n9889), .ZN(n7325) );
  OR2_X1 U7851 ( .A1(n6733), .A2(n9895), .ZN(n7324) );
  NAND2_X1 U7852 ( .A1(n12186), .A2(n12192), .ZN(n12221) );
  AND2_X1 U7853 ( .A1(n8931), .A2(n11814), .ZN(n11956) );
  AOI21_X1 U7854 ( .B1(n12318), .B2(n7069), .A(n7068), .ZN(n7067) );
  INV_X1 U7855 ( .A(n8859), .ZN(n7069) );
  NOR2_X1 U7856 ( .A1(n12109), .A2(n7616), .ZN(n7615) );
  INV_X1 U7857 ( .A(n12117), .ZN(n7616) );
  INV_X1 U7858 ( .A(n12589), .ZN(n8856) );
  NOR2_X1 U7859 ( .A1(n12392), .A2(n7343), .ZN(n7341) );
  AND2_X1 U7860 ( .A1(n12068), .A2(n6681), .ZN(n12065) );
  OR2_X1 U7861 ( .A1(n8584), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8597) );
  NOR2_X1 U7862 ( .A1(n7597), .A2(n7594), .ZN(n7593) );
  INV_X1 U7863 ( .A(n12027), .ZN(n7597) );
  INV_X1 U7864 ( .A(n12030), .ZN(n7598) );
  NAND2_X1 U7865 ( .A1(n10244), .A2(n8837), .ZN(n12002) );
  NAND2_X1 U7866 ( .A1(n9866), .A2(n8835), .ZN(n10293) );
  INV_X1 U7867 ( .A(n11990), .ZN(n8876) );
  NAND2_X1 U7868 ( .A1(n7274), .A2(n7277), .ZN(n7273) );
  NOR2_X1 U7869 ( .A1(n8370), .A2(n7319), .ZN(n7318) );
  AND2_X1 U7870 ( .A1(n9498), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8370) );
  INV_X1 U7871 ( .A(n8368), .ZN(n7319) );
  NAND2_X1 U7872 ( .A1(n9134), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8366) );
  NAND4_X1 U7873 ( .A1(n7767), .A2(n14897), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7412) );
  INV_X1 U7874 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7767) );
  NAND4_X1 U7875 ( .A1(n7766), .A2(n7765), .A3(n10971), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7413) );
  INV_X1 U7876 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7765) );
  INV_X1 U7877 ( .A(n7465), .ZN(n7029) );
  OR2_X1 U7878 ( .A1(n12777), .A2(n7038), .ZN(n7036) );
  NAND2_X1 U7879 ( .A1(n7037), .A2(n7038), .ZN(n7034) );
  INV_X1 U7880 ( .A(n10724), .ZN(n7477) );
  NOR2_X1 U7881 ( .A1(n12827), .A2(n7471), .ZN(n7470) );
  INV_X1 U7882 ( .A(n12657), .ZN(n7471) );
  INV_X1 U7883 ( .A(n12634), .ZN(n10115) );
  INV_X1 U7884 ( .A(n13099), .ZN(n7666) );
  INV_X1 U7885 ( .A(n13100), .ZN(n7667) );
  INV_X1 U7886 ( .A(n11379), .ZN(n7159) );
  NAND2_X1 U7887 ( .A1(n13444), .A2(n11523), .ZN(n7423) );
  INV_X1 U7888 ( .A(n13138), .ZN(n7178) );
  INV_X1 U7889 ( .A(n10024), .ZN(n7384) );
  NAND2_X1 U7890 ( .A1(n12867), .A2(n13155), .ZN(n9778) );
  NAND2_X1 U7891 ( .A1(n6939), .A2(n6938), .ZN(n9476) );
  INV_X1 U7892 ( .A(n13120), .ZN(n6939) );
  NAND2_X1 U7893 ( .A1(n7479), .A2(n9261), .ZN(n7478) );
  INV_X1 U7894 ( .A(n7480), .ZN(n7479) );
  OAI21_X1 U7895 ( .B1(n6901), .B2(n6900), .A(n6899), .ZN(n7655) );
  NAND2_X1 U7896 ( .A1(n11700), .A2(n11688), .ZN(n6900) );
  NAND2_X1 U7897 ( .A1(n6594), .A2(n11700), .ZN(n6899) );
  INV_X1 U7898 ( .A(n10698), .ZN(n7221) );
  NAND2_X1 U7899 ( .A1(n8992), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6897) );
  OR2_X1 U7900 ( .A1(n7190), .A2(n10185), .ZN(n7189) );
  AND2_X1 U7901 ( .A1(n10186), .A2(n10041), .ZN(n7190) );
  AND2_X1 U7902 ( .A1(n7544), .A2(n14241), .ZN(n7539) );
  NAND2_X1 U7903 ( .A1(n7517), .A2(n7515), .ZN(n14233) );
  AOI21_X1 U7904 ( .B1(n7519), .B2(n7518), .A(n7516), .ZN(n7515) );
  OAI21_X1 U7905 ( .B1(n14229), .B2(n7519), .A(n7153), .ZN(n14235) );
  AND2_X1 U7906 ( .A1(n7516), .A2(n7518), .ZN(n7153) );
  INV_X1 U7907 ( .A(n7546), .ZN(n7543) );
  NAND2_X1 U7908 ( .A1(n7539), .A2(n7546), .ZN(n7538) );
  NOR2_X1 U7909 ( .A1(n14545), .A2(n7255), .ZN(n7254) );
  INV_X1 U7910 ( .A(n8296), .ZN(n7255) );
  AND2_X1 U7911 ( .A1(n14285), .A2(n14173), .ZN(n6936) );
  NAND2_X1 U7912 ( .A1(n6617), .A2(n11210), .ZN(n6935) );
  INV_X1 U7913 ( .A(n7400), .ZN(n7399) );
  AOI21_X1 U7914 ( .B1(n8168), .B2(n7401), .A(n8167), .ZN(n7400) );
  INV_X1 U7915 ( .A(n8149), .ZN(n7401) );
  AND2_X1 U7916 ( .A1(n14602), .A2(n8132), .ZN(n7402) );
  NOR2_X1 U7917 ( .A1(n7259), .A2(n6884), .ZN(n6883) );
  INV_X1 U7918 ( .A(n8292), .ZN(n6884) );
  INV_X1 U7919 ( .A(n7260), .ZN(n7259) );
  AOI21_X1 U7920 ( .B1(n11210), .B2(n8293), .A(n14285), .ZN(n7260) );
  INV_X1 U7921 ( .A(n8293), .ZN(n7258) );
  NAND2_X1 U7922 ( .A1(n14106), .A2(n14107), .ZN(n7509) );
  NOR2_X1 U7923 ( .A1(n14613), .A2(n14710), .ZN(n14616) );
  OAI22_X1 U7924 ( .A1(n8223), .A2(n7831), .B1(SI_23_), .B2(n8221), .ZN(n7859)
         );
  OR2_X1 U7925 ( .A1(n6595), .A2(n11155), .ZN(n7577) );
  NAND2_X1 U7926 ( .A1(n7722), .A2(n7712), .ZN(n7719) );
  NAND2_X1 U7927 ( .A1(n7722), .A2(n6637), .ZN(n7718) );
  INV_X1 U7928 ( .A(n8180), .ZN(n7825) );
  NAND2_X1 U7929 ( .A1(n8117), .A2(n8116), .ZN(n7815) );
  NAND2_X1 U7930 ( .A1(n7808), .A2(SI_15_), .ZN(n8097) );
  AOI21_X1 U7931 ( .B1(n6574), .B2(n7986), .A(n7564), .ZN(n7563) );
  AND2_X1 U7932 ( .A1(n7802), .A2(n7801), .ZN(n8039) );
  XNOR2_X1 U7933 ( .A(n8021), .B(SI_10_), .ZN(n8018) );
  INV_X1 U7934 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U7935 ( .A1(n6829), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n6828) );
  OAI22_X1 U7936 ( .A1(n14807), .A2(n14771), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14806), .ZN(n14772) );
  OAI22_X1 U7937 ( .A1(n14836), .A2(n14835), .B1(P1_ADDR_REG_12__SCAN_IN), 
        .B2(n14834), .ZN(n14842) );
  NOR2_X1 U7938 ( .A1(n7099), .A2(n11623), .ZN(n7098) );
  INV_X1 U7939 ( .A(n11097), .ZN(n7099) );
  NAND2_X1 U7940 ( .A1(n7100), .A2(n6713), .ZN(n7097) );
  NAND2_X1 U7941 ( .A1(n8428), .A2(n8427), .ZN(n8646) );
  INV_X1 U7942 ( .A(n8634), .ZN(n8428) );
  AND2_X1 U7943 ( .A1(n7116), .A2(n7114), .ZN(n7111) );
  OR2_X1 U7944 ( .A1(n7112), .A2(n7110), .ZN(n7109) );
  INV_X1 U7945 ( .A(n7116), .ZN(n7110) );
  AND2_X1 U7946 ( .A1(n11908), .A2(n7113), .ZN(n7112) );
  NAND2_X1 U7947 ( .A1(n11872), .A2(n7114), .ZN(n7113) );
  NAND2_X1 U7948 ( .A1(n6564), .A2(SI_1_), .ZN(n8466) );
  NAND2_X1 U7949 ( .A1(n9865), .A2(n7088), .ZN(n10079) );
  NAND2_X1 U7950 ( .A1(n7085), .A2(n7084), .ZN(n7088) );
  NAND2_X1 U7951 ( .A1(n9866), .A2(n11655), .ZN(n7085) );
  CLKBUF_X1 U7952 ( .A(n9866), .Z(n11967) );
  NAND2_X1 U7953 ( .A1(n8436), .A2(n8435), .ZN(n8753) );
  INV_X1 U7954 ( .A(n8743), .ZN(n8436) );
  NAND2_X1 U7955 ( .A1(n8438), .A2(n8437), .ZN(n8770) );
  INV_X1 U7956 ( .A(n8768), .ZN(n8438) );
  NAND4_X1 U7957 ( .A1(n7370), .A2(n10557), .A3(n10848), .A4(n7078), .ZN(
        n10859) );
  NAND2_X1 U7958 ( .A1(n7105), .A2(n7108), .ZN(n7103) );
  AOI21_X1 U7959 ( .B1(n7109), .B2(n7107), .A(n7106), .ZN(n7105) );
  INV_X1 U7960 ( .A(n7111), .ZN(n7107) );
  INV_X1 U7961 ( .A(n11841), .ZN(n7106) );
  OAI21_X1 U7962 ( .B1(n11871), .B2(n7108), .A(n7105), .ZN(n11889) );
  AND2_X1 U7963 ( .A1(n11640), .A2(n12360), .ZN(n7378) );
  XNOR2_X1 U7964 ( .A(n10213), .B(n12180), .ZN(n10081) );
  NAND2_X1 U7965 ( .A1(n10080), .A2(n10081), .ZN(n10215) );
  OR2_X1 U7966 ( .A1(n11631), .A2(n12405), .ZN(n7114) );
  NAND2_X1 U7967 ( .A1(n8432), .A2(n8431), .ZN(n8704) );
  INV_X1 U7968 ( .A(n8690), .ZN(n8432) );
  OR2_X1 U7969 ( .A1(n8931), .A2(n11814), .ZN(n11954) );
  AND4_X1 U7970 ( .A1(n8639), .A2(n8638), .A3(n8637), .A4(n8636), .ZN(n11099)
         );
  NAND2_X1 U7971 ( .A1(n6950), .A2(n6948), .ZN(n9547) );
  NAND2_X1 U7972 ( .A1(n6949), .A2(P3_IR_REG_1__SCAN_IN), .ZN(n6948) );
  NAND2_X1 U7973 ( .A1(n9546), .A2(n9582), .ZN(n6950) );
  OR2_X1 U7974 ( .A1(n9580), .A2(n9579), .ZN(n7340) );
  XNOR2_X1 U7975 ( .A(n9701), .B(n7338), .ZN(n9703) );
  OR2_X1 U7976 ( .A1(n8479), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8521) );
  AOI22_X1 U7977 ( .A1(n9896), .A2(P3_REG1_REG_5__SCAN_IN), .B1(n9895), .B2(
        n9894), .ZN(n9897) );
  NOR2_X1 U7978 ( .A1(n9897), .A2(n9898), .ZN(n10171) );
  AOI21_X1 U7979 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10631), .A(n10630), .ZN(
        n10633) );
  NAND2_X1 U7980 ( .A1(n15460), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U7981 ( .A1(n6723), .A2(n6706), .ZN(n7336) );
  INV_X1 U7982 ( .A(n10801), .ZN(n6723) );
  NAND2_X1 U7983 ( .A1(n10924), .A2(n6722), .ZN(n6721) );
  NAND2_X1 U7984 ( .A1(n10923), .A2(n6722), .ZN(n6720) );
  OR2_X1 U7985 ( .A1(n11251), .A2(n11252), .ZN(n6995) );
  NAND2_X1 U7986 ( .A1(n11254), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n11253) );
  XNOR2_X1 U7987 ( .A(n12221), .B(n12196), .ZN(n12187) );
  NAND2_X1 U7988 ( .A1(n6732), .A2(n6606), .ZN(n6731) );
  NAND2_X1 U7989 ( .A1(n12187), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12223) );
  NAND2_X1 U7990 ( .A1(n14905), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14904) );
  OR2_X1 U7991 ( .A1(n14902), .A2(n14903), .ZN(n6997) );
  INV_X1 U7992 ( .A(n8826), .ZN(n11615) );
  INV_X1 U7993 ( .A(n11340), .ZN(n12132) );
  XNOR2_X1 U7994 ( .A(n12338), .B(n12320), .ZN(n12334) );
  NOR2_X1 U7995 ( .A1(n6678), .A2(n7619), .ZN(n7618) );
  INV_X1 U7996 ( .A(n8736), .ZN(n7619) );
  NAND2_X1 U7997 ( .A1(n12593), .A2(n12172), .ZN(n8736) );
  OR2_X1 U7998 ( .A1(n12527), .A2(n12407), .ZN(n7054) );
  NOR2_X1 U7999 ( .A1(n12398), .A2(n7623), .ZN(n7622) );
  INV_X1 U8000 ( .A(n12401), .ZN(n6967) );
  INV_X1 U8001 ( .A(n12415), .ZN(n12420) );
  NAND2_X1 U8002 ( .A1(n12431), .A2(n8853), .ZN(n12421) );
  NAND2_X1 U8003 ( .A1(n12421), .A2(n12420), .ZN(n12419) );
  AND2_X1 U8004 ( .A1(n12084), .A2(n12093), .ZN(n12415) );
  AND2_X1 U8005 ( .A1(n12078), .A2(n12074), .ZN(n12429) );
  INV_X1 U8006 ( .A(n12445), .ZN(n12450) );
  AND2_X1 U8007 ( .A1(n12075), .A2(n12071), .ZN(n12445) );
  AOI21_X1 U8008 ( .B1(n7607), .B2(n7608), .A(n7606), .ZN(n7605) );
  INV_X1 U8009 ( .A(n12063), .ZN(n7606) );
  NAND2_X1 U8010 ( .A1(n12462), .A2(n12461), .ZN(n12460) );
  NAND2_X1 U8011 ( .A1(n11165), .A2(n11164), .ZN(n11163) );
  NAND2_X1 U8012 ( .A1(n10987), .A2(n7345), .ZN(n6741) );
  OR2_X1 U8013 ( .A1(n8848), .A2(n7350), .ZN(n7348) );
  NAND2_X1 U8014 ( .A1(n8424), .A2(n8423), .ZN(n8584) );
  INV_X1 U8015 ( .A(n8568), .ZN(n8424) );
  INV_X1 U8016 ( .A(n10225), .ZN(n6965) );
  INV_X1 U8017 ( .A(n10083), .ZN(n11997) );
  INV_X1 U8018 ( .A(n12480), .ZN(n12406) );
  OR2_X1 U8019 ( .A1(n8883), .A2(n12129), .ZN(n12408) );
  NAND2_X1 U8020 ( .A1(n8934), .A2(n8874), .ZN(n12474) );
  NAND2_X1 U8021 ( .A1(n8767), .A2(n8766), .ZN(n11878) );
  OR2_X1 U8022 ( .A1(n11951), .A2(n10545), .ZN(n8766) );
  OR2_X1 U8023 ( .A1(n11951), .A2(n9717), .ZN(n8728) );
  OR2_X1 U8024 ( .A1(n9718), .A2(n8813), .ZN(n8729) );
  INV_X1 U8025 ( .A(n10244), .ZN(n15475) );
  NAND2_X1 U8026 ( .A1(n8925), .A2(n11990), .ZN(n15515) );
  INV_X1 U8027 ( .A(n12408), .ZN(n12479) );
  AND3_X1 U8028 ( .A1(n9108), .A2(n12616), .A3(n8936), .ZN(n9752) );
  AND2_X1 U8029 ( .A1(n8891), .A2(n8890), .ZN(n8917) );
  OR2_X1 U8030 ( .A1(n8405), .A2(n8404), .ZN(n8775) );
  NAND2_X1 U8031 ( .A1(n8399), .A2(n6702), .ZN(n7289) );
  INV_X1 U8032 ( .A(n7075), .ZN(n7073) );
  AOI21_X1 U8033 ( .B1(n7295), .B2(n7297), .A(n7294), .ZN(n7293) );
  INV_X1 U8034 ( .A(n8397), .ZN(n7294) );
  NAND2_X1 U8035 ( .A1(n8738), .A2(n8737), .ZN(n8740) );
  INV_X1 U8036 ( .A(n7628), .ZN(n7626) );
  AND2_X1 U8037 ( .A1(n8389), .A2(n8388), .ZN(n8711) );
  INV_X1 U8038 ( .A(n8387), .ZN(n7303) );
  AND2_X1 U8039 ( .A1(n8387), .A2(n8386), .ZN(n8696) );
  NAND2_X1 U8040 ( .A1(n8685), .A2(n8385), .ZN(n8697) );
  NAND2_X1 U8041 ( .A1(n8697), .A2(n8696), .ZN(n8699) );
  NAND2_X1 U8042 ( .A1(n8329), .A2(n8331), .ZN(n8700) );
  NAND2_X1 U8043 ( .A1(n8683), .A2(n8682), .ZN(n8685) );
  NAND2_X1 U8044 ( .A1(n8654), .A2(n8381), .ZN(n8669) );
  NAND2_X1 U8045 ( .A1(n8669), .A2(n8668), .ZN(n8671) );
  NAND2_X1 U8046 ( .A1(n7080), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8672) );
  OAI21_X1 U8047 ( .B1(n8375), .B2(n7269), .A(n8377), .ZN(n7268) );
  AND2_X1 U8048 ( .A1(n8374), .A2(n8640), .ZN(n7270) );
  INV_X1 U8049 ( .A(n8640), .ZN(n7269) );
  NAND2_X1 U8050 ( .A1(n8373), .A2(n9501), .ZN(n8375) );
  OR2_X1 U8051 ( .A1(n8373), .A2(n9501), .ZN(n8374) );
  NAND2_X1 U8052 ( .A1(n6616), .A2(n8374), .ZN(n8629) );
  NOR2_X1 U8053 ( .A1(n7314), .A2(n8622), .ZN(n7313) );
  INV_X1 U8054 ( .A(n7316), .ZN(n7314) );
  NAND2_X1 U8055 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n7317), .ZN(n7316) );
  NAND2_X1 U8056 ( .A1(n8591), .A2(n8367), .ZN(n8369) );
  NOR2_X1 U8057 ( .A1(n8578), .A2(n7283), .ZN(n7282) );
  INV_X1 U8058 ( .A(n8364), .ZN(n7283) );
  NAND2_X1 U8059 ( .A1(n8362), .A2(n8361), .ZN(n8565) );
  NAND2_X1 U8060 ( .A1(n8549), .A2(n8360), .ZN(n8362) );
  XNOR2_X1 U8061 ( .A(n9074), .B(P1_DATAO_REG_5__SCAN_IN), .ZN(n8519) );
  OAI21_X1 U8062 ( .B1(n8492), .B2(n7306), .A(n7304), .ZN(n8520) );
  INV_X1 U8063 ( .A(n7307), .ZN(n7306) );
  AOI21_X1 U8064 ( .B1(n7307), .B2(n7305), .A(n6669), .ZN(n7304) );
  AND2_X1 U8065 ( .A1(n8353), .A2(n7308), .ZN(n7307) );
  INV_X1 U8066 ( .A(n7472), .ZN(n7047) );
  AND2_X1 U8067 ( .A1(n7044), .A2(n12643), .ZN(n7046) );
  INV_X1 U8068 ( .A(n10118), .ZN(n7483) );
  NOR2_X1 U8069 ( .A1(n6613), .A2(n7029), .ZN(n7025) );
  AND2_X1 U8070 ( .A1(n6677), .A2(n7033), .ZN(n7032) );
  INV_X1 U8071 ( .A(n13209), .ZN(n10065) );
  OAI21_X1 U8072 ( .B1(n7464), .B2(n7466), .A(n7465), .ZN(n7043) );
  OR2_X1 U8073 ( .A1(n11386), .A2(n11385), .ZN(n11398) );
  INV_X1 U8074 ( .A(n7470), .ZN(n7468) );
  AND2_X1 U8075 ( .A1(n10675), .A2(n10666), .ZN(n7050) );
  NOR2_X1 U8076 ( .A1(n7018), .A2(n7487), .ZN(n7486) );
  INV_X1 U8077 ( .A(n10112), .ZN(n7487) );
  NAND2_X1 U8078 ( .A1(n10823), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n10906) );
  INV_X1 U8079 ( .A(n10825), .ZN(n10823) );
  INV_X1 U8080 ( .A(n13072), .ZN(n11513) );
  NOR2_X1 U8081 ( .A1(n9285), .A2(n13887), .ZN(n9464) );
  AOI21_X1 U8082 ( .B1(n15212), .B2(n9246), .A(n9247), .ZN(n9249) );
  OR2_X1 U8083 ( .A1(n9249), .A2(n6788), .ZN(n6787) );
  NOR2_X1 U8084 ( .A1(n9456), .A2(n10500), .ZN(n6788) );
  AND2_X1 U8085 ( .A1(n6787), .A2(n6786), .ZN(n15229) );
  INV_X1 U8086 ( .A(n15230), .ZN(n6786) );
  AOI21_X1 U8087 ( .B1(n13214), .B2(n13215), .A(n6794), .ZN(n6793) );
  INV_X1 U8088 ( .A(n9204), .ZN(n6794) );
  NOR2_X1 U8089 ( .A1(n9322), .A2(n6795), .ZN(n9325) );
  AND2_X1 U8090 ( .A1(n9998), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6795) );
  NOR2_X1 U8091 ( .A1(n9379), .A2(n9378), .ZN(n9487) );
  OR2_X1 U8092 ( .A1(n9487), .A2(n6800), .ZN(n6799) );
  AND2_X1 U8093 ( .A1(n10377), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6800) );
  INV_X1 U8094 ( .A(n11042), .ZN(n15286) );
  NAND2_X1 U8095 ( .A1(n15286), .A2(n15285), .ZN(n15284) );
  NAND2_X1 U8096 ( .A1(n15298), .A2(n15297), .ZN(n15295) );
  NAND2_X1 U8097 ( .A1(n13264), .A2(n11500), .ZN(n11510) );
  INV_X1 U8098 ( .A(n13149), .ZN(n11509) );
  NOR3_X2 U8099 ( .A1(n13311), .A2(n13493), .A3(n7232), .ZN(n13257) );
  OR2_X1 U8100 ( .A1(n7233), .A2(n13484), .ZN(n7232) );
  XNOR2_X1 U8101 ( .A(n13484), .B(n13183), .ZN(n13149) );
  AOI21_X1 U8102 ( .B1(n7169), .B2(n11416), .A(n6582), .ZN(n7167) );
  INV_X1 U8103 ( .A(n13352), .ZN(n7432) );
  XNOR2_X1 U8104 ( .A(n13526), .B(n13190), .ZN(n13352) );
  NAND2_X1 U8105 ( .A1(n11406), .A2(n11405), .ZN(n13364) );
  NAND2_X1 U8106 ( .A1(n11368), .A2(n6610), .ZN(n13412) );
  OR2_X1 U8107 ( .A1(n13445), .A2(n13444), .ZN(n13447) );
  OR2_X1 U8108 ( .A1(n7391), .A2(n6573), .ZN(n13451) );
  NAND2_X1 U8109 ( .A1(n11003), .A2(n11002), .ZN(n12973) );
  NAND2_X1 U8110 ( .A1(n10998), .A2(n10997), .ZN(n11000) );
  NAND2_X1 U8111 ( .A1(n10599), .A2(n6611), .ZN(n10644) );
  NAND2_X1 U8112 ( .A1(n6778), .A2(n6994), .ZN(n10578) );
  INV_X1 U8113 ( .A(n13134), .ZN(n6994) );
  AOI21_X1 U8114 ( .B1(n10024), .B2(n7383), .A(n6624), .ZN(n7382) );
  INV_X1 U8115 ( .A(n10023), .ZN(n7383) );
  OR2_X1 U8116 ( .A1(n10404), .A2(n7384), .ZN(n7381) );
  NAND2_X1 U8117 ( .A1(n10446), .A2(n9995), .ZN(n6781) );
  INV_X1 U8118 ( .A(n9471), .ZN(n7226) );
  NAND2_X1 U8119 ( .A1(n11436), .A2(n11435), .ZN(n13520) );
  AND2_X1 U8120 ( .A1(n10347), .A2(n15423), .ZN(n15405) );
  AND2_X1 U8121 ( .A1(n7661), .A2(n9279), .ZN(n7179) );
  NAND2_X1 U8122 ( .A1(n7574), .A2(SI_22_), .ZN(n7581) );
  XNOR2_X1 U8123 ( .A(n9047), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9224) );
  INV_X1 U8124 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9301) );
  NAND2_X1 U8125 ( .A1(n11793), .A2(n11801), .ZN(n7215) );
  NAND2_X1 U8126 ( .A1(n11276), .A2(n6644), .ZN(n11297) );
  NAND2_X1 U8127 ( .A1(n11270), .A2(n11269), .ZN(n11276) );
  INV_X1 U8128 ( .A(n6712), .ZN(n7184) );
  NOR2_X1 U8129 ( .A1(n7653), .A2(n7189), .ZN(n7187) );
  NAND2_X1 U8130 ( .A1(n13940), .A2(n6638), .ZN(n7185) );
  NAND2_X1 U8131 ( .A1(n10186), .A2(n10185), .ZN(n7191) );
  NAND2_X1 U8132 ( .A1(n6908), .A2(n7652), .ZN(n7186) );
  AND2_X1 U8133 ( .A1(n7648), .A2(n7188), .ZN(n6908) );
  INV_X1 U8134 ( .A(n7189), .ZN(n7188) );
  NAND2_X1 U8135 ( .A1(n13919), .A2(n6635), .ZN(n6903) );
  INV_X1 U8136 ( .A(n6898), .ZN(n11692) );
  AOI21_X1 U8137 ( .B1(n13919), .B2(n11688), .A(n6594), .ZN(n6898) );
  AND4_X1 U8138 ( .A1(n8115), .A2(n8114), .A3(n8113), .A4(n8112), .ZN(n11690)
         );
  AND4_X1 U8139 ( .A1(n8087), .A2(n8086), .A3(n8085), .A4(n8084), .ZN(n11683)
         );
  OR2_X1 U8140 ( .A1(n8255), .A2(n14352), .ZN(n7887) );
  NAND2_X1 U8141 ( .A1(n14076), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7872) );
  OR2_X1 U8142 ( .A1(n8255), .A2(n7870), .ZN(n6957) );
  NAND2_X1 U8143 ( .A1(n14076), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U8144 ( .A1(n14244), .A2(n14243), .ZN(n14415) );
  NAND2_X1 U8145 ( .A1(n14652), .A2(n14318), .ZN(n7507) );
  AND2_X1 U8146 ( .A1(n14497), .A2(n14512), .ZN(n7408) );
  NAND2_X1 U8147 ( .A1(n6876), .A2(n6875), .ZN(n14467) );
  NOR2_X1 U8148 ( .A1(n7510), .A2(n14471), .ZN(n6875) );
  OR2_X1 U8149 ( .A1(n8300), .A2(n14320), .ZN(n7689) );
  AOI21_X1 U8150 ( .B1(n6917), .B2(n6914), .A(n6913), .ZN(n6912) );
  INV_X1 U8151 ( .A(n14533), .ZN(n6915) );
  INV_X1 U8152 ( .A(n14509), .ZN(n6913) );
  XNOR2_X1 U8153 ( .A(n14676), .B(n6940), .ZN(n14522) );
  INV_X1 U8154 ( .A(n14522), .ZN(n14520) );
  NAND2_X1 U8155 ( .A1(n14687), .A2(n7254), .ZN(n14542) );
  NAND2_X1 U8156 ( .A1(n14616), .A2(n14198), .ZN(n14587) );
  NOR2_X2 U8157 ( .A1(n14587), .A2(n14581), .ZN(n14575) );
  OAI21_X1 U8158 ( .B1(n14603), .B2(n14195), .A(n14196), .ZN(n14586) );
  NAND2_X1 U8159 ( .A1(n8133), .A2(n7402), .ZN(n14611) );
  OR2_X1 U8160 ( .A1(n11211), .A2(n14288), .ZN(n6937) );
  NAND2_X1 U8161 ( .A1(n7261), .A2(n14288), .ZN(n11199) );
  INV_X1 U8162 ( .A(n11201), .ZN(n7261) );
  NOR2_X1 U8163 ( .A1(n14284), .A2(n6874), .ZN(n6873) );
  INV_X1 U8164 ( .A(n7491), .ZN(n7490) );
  NAND2_X1 U8165 ( .A1(n15064), .A2(n8002), .ZN(n15049) );
  NAND2_X1 U8166 ( .A1(n7493), .A2(n7492), .ZN(n9852) );
  AOI21_X1 U8167 ( .B1(n6579), .B2(n7496), .A(n6654), .ZN(n7492) );
  INV_X1 U8168 ( .A(n7497), .ZN(n7496) );
  NAND2_X1 U8169 ( .A1(n7494), .A2(n7497), .ZN(n9928) );
  NAND2_X1 U8170 ( .A1(n9764), .A2(n7498), .ZN(n7494) );
  NAND2_X1 U8171 ( .A1(n6925), .A2(n6927), .ZN(n9682) );
  NAND2_X1 U8172 ( .A1(n14111), .A2(n14110), .ZN(n6927) );
  NAND2_X1 U8173 ( .A1(n14253), .A2(n15159), .ZN(n6808) );
  NAND2_X1 U8174 ( .A1(n6809), .A2(n6693), .ZN(n14426) );
  NAND2_X1 U8175 ( .A1(n6811), .A2(n6810), .ZN(n6809) );
  INV_X1 U8176 ( .A(n8317), .ZN(n6810) );
  AOI21_X1 U8177 ( .B1(n11565), .B2(n15139), .A(n11564), .ZN(n14641) );
  NAND2_X1 U8178 ( .A1(n11563), .A2(n11562), .ZN(n11564) );
  AND2_X1 U8179 ( .A1(n7506), .A2(n6618), .ZN(n11570) );
  NAND2_X1 U8180 ( .A1(n8252), .A2(n8251), .ZN(n14644) );
  NAND2_X1 U8181 ( .A1(n14507), .A2(n7513), .ZN(n14487) );
  AND2_X1 U8182 ( .A1(n14507), .A2(n7512), .ZN(n14486) );
  NAND2_X1 U8183 ( .A1(n8107), .A2(n8106), .ZN(n14944) );
  AOI21_X1 U8184 ( .B1(n8171), .B2(n9113), .A(n6815), .ZN(n7915) );
  NOR2_X1 U8185 ( .A1(n8171), .A2(n6814), .ZN(n6815) );
  NAND2_X1 U8186 ( .A1(n15092), .A2(n8308), .ZN(n15159) );
  NAND2_X1 U8187 ( .A1(n8274), .A2(n14245), .ZN(n15139) );
  AND2_X1 U8188 ( .A1(n7717), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9102) );
  AOI21_X1 U8189 ( .B1(n13060), .B2(n13059), .A(n13058), .ZN(n13077) );
  INV_X1 U8190 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7844) );
  INV_X1 U8191 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U8192 ( .A1(n8139), .A2(n7688), .ZN(n7750) );
  INV_X1 U8193 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7749) );
  NOR2_X1 U8194 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n7224) );
  INV_X1 U8195 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n7223) );
  INV_X1 U8196 ( .A(n7719), .ZN(n7707) );
  NAND2_X1 U8197 ( .A1(n7823), .A2(n9717), .ZN(n7824) );
  OR2_X1 U8198 ( .A1(n7823), .A2(n9717), .ZN(n7826) );
  INV_X1 U8199 ( .A(n7592), .ZN(n7591) );
  NAND2_X1 U8200 ( .A1(n7789), .A2(n7788), .ZN(n7987) );
  AND2_X1 U8201 ( .A1(n7503), .A2(n7875), .ZN(n7891) );
  NAND3_X1 U8202 ( .A1(n7249), .A2(n7416), .A3(n6604), .ZN(n6759) );
  NAND2_X1 U8203 ( .A1(n7250), .A2(n7877), .ZN(n7249) );
  XNOR2_X1 U8204 ( .A(n7769), .B(SI_1_), .ZN(n7877) );
  INV_X1 U8205 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n14791) );
  NAND2_X1 U8206 ( .A1(n14875), .A2(n14874), .ZN(n7457) );
  NOR2_X1 U8207 ( .A1(n14815), .A2(n14816), .ZN(n14819) );
  NOR2_X1 U8208 ( .A1(n14876), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n14815) );
  NAND2_X1 U8209 ( .A1(n9492), .A2(n7450), .ZN(n7449) );
  INV_X1 U8210 ( .A(n14982), .ZN(n6820) );
  NAND2_X1 U8211 ( .A1(n14833), .A2(n9519), .ZN(n6819) );
  NOR2_X1 U8212 ( .A1(n14986), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7245) );
  AND3_X1 U8213 ( .A1(n8556), .A2(n8555), .A3(n8554), .ZN(n10796) );
  AND3_X1 U8214 ( .A1(n11890), .A2(n11847), .A3(n11848), .ZN(n11850) );
  OAI21_X1 U8215 ( .B1(n7372), .B2(n12463), .A(n11928), .ZN(n11628) );
  NAND2_X1 U8216 ( .A1(n8752), .A2(n8751), .ZN(n11905) );
  NAND2_X1 U8217 ( .A1(n8449), .A2(n8448), .ZN(n12321) );
  NAND4_X1 U8218 ( .A1(n8748), .A2(n8747), .A3(n8746), .A4(n8745), .ZN(n12372)
         );
  NAND4_X1 U8219 ( .A1(n8602), .A2(n8601), .A3(n8600), .A4(n8599), .ZN(n12173)
         );
  INV_X1 U8220 ( .A(n7071), .ZN(n7070) );
  OAI211_X1 U8221 ( .C1(n8458), .C2(n7072), .A(n8570), .B(n8572), .ZN(n7071)
         );
  AOI21_X1 U8222 ( .B1(n8478), .B2(P3_IR_REG_2__SCAN_IN), .A(n6756), .ZN(n6755) );
  AND2_X1 U8223 ( .A1(n12619), .A2(n6757), .ZN(n6756) );
  OR2_X1 U8224 ( .A1(n10620), .A2(n10621), .ZN(n10811) );
  NAND2_X1 U8225 ( .A1(n12282), .A2(n6747), .ZN(n6746) );
  AND2_X1 U8226 ( .A1(n6597), .A2(n6708), .ZN(n6747) );
  XNOR2_X1 U8227 ( .A(n6749), .B(n12276), .ZN(n6748) );
  NAND2_X1 U8228 ( .A1(n12266), .A2(n7015), .ZN(n6749) );
  OR2_X1 U8229 ( .A1(n12267), .A2(n12530), .ZN(n7015) );
  AND2_X1 U8230 ( .A1(n6997), .A2(n6996), .ZN(n12235) );
  NAND2_X1 U8231 ( .A1(n12233), .A2(n12252), .ZN(n6996) );
  XNOR2_X1 U8232 ( .A(n8946), .B(n11984), .ZN(n11581) );
  NAND2_X1 U8233 ( .A1(n8793), .A2(n8792), .ZN(n11622) );
  OR2_X1 U8234 ( .A1(n11951), .A2(n11161), .ZN(n8792) );
  NAND2_X1 U8235 ( .A1(n8781), .A2(n8780), .ZN(n12295) );
  OR2_X1 U8236 ( .A1(n10873), .A2(n8813), .ZN(n8781) );
  NAND2_X1 U8237 ( .A1(n8717), .A2(n8716), .ZN(n12390) );
  OR2_X1 U8238 ( .A1(n9679), .A2(n8813), .ZN(n8717) );
  INV_X1 U8239 ( .A(n12488), .ZN(n12438) );
  NAND2_X1 U8240 ( .A1(n6553), .A2(n15509), .ZN(n7058) );
  NAND2_X1 U8241 ( .A1(n8645), .A2(n8644), .ZN(n12605) );
  OR2_X1 U8242 ( .A1(n7586), .A2(n7411), .ZN(n9302) );
  NAND2_X1 U8243 ( .A1(n10210), .A2(n9800), .ZN(n9809) );
  NAND2_X1 U8244 ( .A1(n11384), .A2(n11383), .ZN(n13543) );
  NAND2_X1 U8245 ( .A1(n11486), .A2(n11485), .ZN(n13490) );
  OAI21_X1 U8246 ( .B1(n12801), .B2(n12797), .A(n12798), .ZN(n12744) );
  NAND2_X1 U8247 ( .A1(n11410), .A2(n11409), .ZN(n13367) );
  NAND2_X1 U8248 ( .A1(n10569), .A2(n10568), .ZN(n13855) );
  NAND2_X1 U8249 ( .A1(n10063), .A2(n10066), .ZN(n10113) );
  NAND2_X1 U8250 ( .A1(n12766), .A2(n12653), .ZN(n7051) );
  NAND2_X1 U8251 ( .A1(n11396), .A2(n11395), .ZN(n13537) );
  NAND2_X1 U8252 ( .A1(n10820), .A2(n10819), .ZN(n13582) );
  NAND2_X1 U8253 ( .A1(n10671), .A2(n7050), .ZN(n10722) );
  NAND2_X1 U8254 ( .A1(n10582), .A2(n10581), .ZN(n12941) );
  NAND2_X1 U8255 ( .A1(n11371), .A2(n11370), .ZN(n13549) );
  NAND2_X1 U8256 ( .A1(n7052), .A2(n9973), .ZN(n15393) );
  NAND2_X1 U8257 ( .A1(n9971), .A2(n13068), .ZN(n7052) );
  AOI21_X1 U8258 ( .B1(n6854), .B2(n13115), .A(n13114), .ZN(n13166) );
  OAI21_X1 U8259 ( .B1(n6856), .B2(n6855), .A(n7664), .ZN(n6854) );
  NAND2_X1 U8260 ( .A1(n13179), .A2(n13180), .ZN(n6946) );
  XNOR2_X1 U8261 ( .A(n13230), .B(n13234), .ZN(n11044) );
  NOR2_X1 U8262 ( .A1(n11044), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13232) );
  NAND2_X1 U8263 ( .A1(n13085), .A2(n13084), .ZN(n13261) );
  OR2_X1 U8264 ( .A1(n14744), .A2(n13082), .ZN(n13085) );
  OR2_X1 U8265 ( .A1(n13269), .A2(n13270), .ZN(n7395) );
  NAND2_X1 U8266 ( .A1(n11446), .A2(n11445), .ZN(n13332) );
  NAND2_X1 U8267 ( .A1(n11360), .A2(n11359), .ZN(n13438) );
  NAND2_X1 U8268 ( .A1(n15358), .A2(n9779), .ZN(n13397) );
  INV_X1 U8269 ( .A(n9224), .ZN(n6805) );
  OAI21_X1 U8270 ( .B1(n10532), .B2(n10531), .A(n10530), .ZN(n10537) );
  INV_X1 U8271 ( .A(n14644), .ZN(n14447) );
  AND2_X1 U8272 ( .A1(n7906), .A2(n6625), .ZN(n7143) );
  NAND2_X1 U8273 ( .A1(n9781), .A2(n14087), .ZN(n7142) );
  AND2_X1 U8274 ( .A1(n8166), .A2(n8165), .ZN(n14609) );
  NOR2_X1 U8275 ( .A1(n7210), .A2(n14074), .ZN(n7208) );
  AND2_X1 U8276 ( .A1(n6686), .A2(n7212), .ZN(n7210) );
  NAND2_X1 U8277 ( .A1(n7212), .A2(n7215), .ZN(n7211) );
  AOI21_X1 U8278 ( .B1(n7644), .B2(n7647), .A(n11782), .ZN(n7643) );
  NAND2_X1 U8279 ( .A1(n7976), .A2(n7975), .ZN(n15089) );
  NAND2_X1 U8280 ( .A1(n8200), .A2(n8199), .ZN(n14682) );
  INV_X1 U8281 ( .A(n14326), .ZN(n13926) );
  NAND2_X1 U8282 ( .A1(n11773), .A2(n13981), .ZN(n13984) );
  NAND2_X1 U8283 ( .A1(n7863), .A2(n7862), .ZN(n14664) );
  INV_X1 U8284 ( .A(n7638), .ZN(n6907) );
  NAND2_X1 U8285 ( .A1(n7638), .A2(n6906), .ZN(n6905) );
  NAND2_X1 U8286 ( .A1(n13950), .A2(n11721), .ZN(n14022) );
  NAND2_X1 U8287 ( .A1(n8064), .A2(n8063), .ZN(n14961) );
  NAND2_X1 U8288 ( .A1(n14757), .A2(n8999), .ZN(n14676) );
  XNOR2_X1 U8289 ( .A(n6888), .B(n6887), .ZN(n6999) );
  INV_X1 U8290 ( .A(n14299), .ZN(n6887) );
  NAND2_X1 U8291 ( .A1(n11568), .A2(n8304), .ZN(n6888) );
  NAND2_X1 U8292 ( .A1(n8185), .A2(n8184), .ZN(n14688) );
  INV_X1 U8293 ( .A(n14198), .ZN(n14705) );
  NAND2_X1 U8294 ( .A1(n8079), .A2(n8078), .ZN(n14952) );
  OR2_X1 U8295 ( .A1(n9396), .A2(n9395), .ZN(n15091) );
  NOR2_X1 U8296 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n7654) );
  NAND2_X1 U8297 ( .A1(n14819), .A2(n14820), .ZN(n7247) );
  NOR2_X1 U8298 ( .A1(n14819), .A2(n14820), .ZN(n14878) );
  OR2_X1 U8299 ( .A1(n14880), .A2(n7453), .ZN(n7447) );
  INV_X1 U8300 ( .A(n14853), .ZN(n6831) );
  NAND2_X1 U8301 ( .A1(n6832), .A2(n6972), .ZN(n14852) );
  NAND2_X1 U8302 ( .A1(n12872), .A2(n15312), .ZN(n6961) );
  NAND2_X1 U8303 ( .A1(n12886), .A2(n12887), .ZN(n12890) );
  INV_X1 U8304 ( .A(n12891), .ZN(n6969) );
  NAND2_X1 U8305 ( .A1(n6943), .A2(n6942), .ZN(n6941) );
  INV_X1 U8306 ( .A(n12896), .ZN(n6942) );
  NAND2_X1 U8307 ( .A1(n7555), .A2(n14134), .ZN(n7554) );
  INV_X1 U8308 ( .A(n12919), .ZN(n6848) );
  AND2_X1 U8309 ( .A1(n12913), .A2(n12912), .ZN(n7663) );
  NAND2_X1 U8310 ( .A1(n6987), .A2(n6986), .ZN(n6985) );
  NAND2_X1 U8311 ( .A1(n12919), .A2(n6846), .ZN(n6845) );
  NAND2_X1 U8312 ( .A1(n12926), .A2(n12925), .ZN(n7682) );
  INV_X1 U8313 ( .A(n14144), .ZN(n7144) );
  NOR2_X1 U8314 ( .A1(n14147), .A2(n14144), .ZN(n7145) );
  NAND2_X1 U8315 ( .A1(n6697), .A2(n7681), .ZN(n7680) );
  NAND2_X1 U8316 ( .A1(n6612), .A2(n12943), .ZN(n6859) );
  INV_X1 U8317 ( .A(n14196), .ZN(n7141) );
  NAND2_X1 U8318 ( .A1(n14200), .A2(n14199), .ZN(n7135) );
  NAND2_X1 U8319 ( .A1(n7137), .A2(n7134), .ZN(n7133) );
  NOR2_X1 U8320 ( .A1(n14194), .A2(n14195), .ZN(n7134) );
  AOI21_X1 U8321 ( .B1(n6850), .B2(n6853), .A(n6670), .ZN(n6849) );
  NOR2_X1 U8322 ( .A1(n12964), .A2(n7000), .ZN(n6853) );
  INV_X1 U8323 ( .A(n13006), .ZN(n7687) );
  NAND2_X1 U8324 ( .A1(n6641), .A2(n7687), .ZN(n7686) );
  NAND2_X1 U8325 ( .A1(n7530), .A2(n14214), .ZN(n7529) );
  AOI21_X1 U8326 ( .B1(n13016), .B2(n13015), .A(n13014), .ZN(n13018) );
  OR2_X1 U8327 ( .A1(n13022), .A2(n13021), .ZN(n7671) );
  AND2_X1 U8328 ( .A1(n13021), .A2(n13022), .ZN(n7672) );
  NAND2_X1 U8329 ( .A1(n7674), .A2(n13039), .ZN(n7673) );
  INV_X1 U8330 ( .A(n6674), .ZN(n7674) );
  NAND2_X1 U8331 ( .A1(n7147), .A2(n7550), .ZN(n14225) );
  NAND2_X1 U8332 ( .A1(n7551), .A2(n14221), .ZN(n7550) );
  INV_X1 U8333 ( .A(n14222), .ZN(n7551) );
  NAND2_X1 U8334 ( .A1(n14225), .A2(n14224), .ZN(n7146) );
  AOI21_X1 U8335 ( .B1(n12224), .B2(n6753), .A(n6752), .ZN(n6750) );
  INV_X1 U8336 ( .A(n12247), .ZN(n6752) );
  INV_X1 U8337 ( .A(n7318), .ZN(n7311) );
  NAND2_X1 U8338 ( .A1(n14228), .A2(n14231), .ZN(n7518) );
  NAND2_X1 U8339 ( .A1(n14082), .A2(n14083), .ZN(n7523) );
  INV_X1 U8340 ( .A(n6881), .ZN(n6880) );
  OAI21_X1 U8341 ( .B1(n10093), .B2(n6882), .A(n15095), .ZN(n6881) );
  INV_X1 U8342 ( .A(n8282), .ZN(n6882) );
  INV_X1 U8343 ( .A(n8169), .ZN(n6761) );
  NOR2_X2 U8344 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8102) );
  OAI21_X1 U8345 ( .B1(n8042), .B2(n7573), .A(n7570), .ZN(n8091) );
  INV_X1 U8346 ( .A(n7798), .ZN(n7565) );
  INV_X1 U8347 ( .A(n7797), .ZN(n7564) );
  AND2_X1 U8348 ( .A1(n7022), .A2(n7020), .ZN(n7004) );
  INV_X1 U8349 ( .A(n7775), .ZN(n7020) );
  NAND2_X1 U8350 ( .A1(n7904), .A2(n7775), .ZN(n7022) );
  NAND2_X1 U8351 ( .A1(n11807), .A2(n11996), .ZN(n7084) );
  INV_X1 U8352 ( .A(n8835), .ZN(n10291) );
  AND2_X1 U8353 ( .A1(n7090), .A2(n7089), .ZN(n11638) );
  NAND2_X1 U8354 ( .A1(n11637), .A2(n12348), .ZN(n7089) );
  INV_X1 U8355 ( .A(n11850), .ZN(n7090) );
  INV_X1 U8356 ( .A(n7094), .ZN(n7093) );
  NAND2_X1 U8357 ( .A1(n10804), .A2(n6703), .ZN(n10928) );
  INV_X1 U8358 ( .A(n10926), .ZN(n6722) );
  INV_X1 U8359 ( .A(n8863), .ZN(n8862) );
  INV_X1 U8360 ( .A(n11954), .ZN(n12141) );
  OR2_X1 U8361 ( .A1(n8815), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8826) );
  OR2_X1 U8362 ( .A1(n12543), .A2(n12463), .ZN(n12075) );
  INV_X1 U8363 ( .A(n7349), .ZN(n7344) );
  NOR2_X1 U8364 ( .A1(n10860), .A2(n12175), .ZN(n8847) );
  NAND2_X1 U8365 ( .A1(n8846), .A2(n7594), .ZN(n10985) );
  NAND2_X1 U8366 ( .A1(n15475), .A2(n9508), .ZN(n12010) );
  AND2_X1 U8367 ( .A1(n7122), .A2(n7124), .ZN(n7121) );
  INV_X1 U8368 ( .A(n7126), .ZN(n7122) );
  AOI21_X1 U8369 ( .B1(n12331), .B2(n7067), .A(n7065), .ZN(n11590) );
  NAND2_X1 U8370 ( .A1(n11585), .A2(n7066), .ZN(n7065) );
  NAND2_X1 U8371 ( .A1(n7067), .A2(n12315), .ZN(n7066) );
  NAND2_X1 U8372 ( .A1(n12315), .A2(n8860), .ZN(n7361) );
  INV_X1 U8373 ( .A(n12127), .ZN(n7359) );
  OR2_X1 U8374 ( .A1(n8915), .A2(n8914), .ZN(n8936) );
  NAND2_X1 U8375 ( .A1(n8894), .A2(n7631), .ZN(n8890) );
  NOR2_X1 U8376 ( .A1(n8399), .A2(n7291), .ZN(n7286) );
  NAND2_X1 U8377 ( .A1(n6675), .A2(n8407), .ZN(n7075) );
  INV_X1 U8378 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7076) );
  INV_X1 U8379 ( .A(n7296), .ZN(n7295) );
  OAI21_X1 U8380 ( .B1(n8737), .B2(n7297), .A(n8396), .ZN(n7296) );
  INV_X1 U8381 ( .A(n8393), .ZN(n7297) );
  AND2_X1 U8382 ( .A1(n8408), .A2(n8407), .ZN(n8918) );
  NAND2_X1 U8383 ( .A1(n7629), .A2(n8324), .ZN(n7628) );
  INV_X1 U8384 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7629) );
  AND2_X1 U8385 ( .A1(n6621), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n7126) );
  INV_X1 U8386 ( .A(n7125), .ZN(n7124) );
  OAI22_X1 U8387 ( .A1(n6621), .A2(n7127), .B1(P3_IR_REG_31__SCAN_IN), .B2(
        n7128), .ZN(n7125) );
  NAND2_X1 U8388 ( .A1(n7128), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7127) );
  INV_X1 U8389 ( .A(n7282), .ZN(n7281) );
  INV_X1 U8390 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8321) );
  INV_X1 U8391 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U8392 ( .A1(n8351), .A2(n8352), .ZN(n7308) );
  INV_X1 U8393 ( .A(n8352), .ZN(n7305) );
  NOR2_X1 U8394 ( .A1(n12777), .A2(n7040), .ZN(n7037) );
  INV_X1 U8395 ( .A(n12706), .ZN(n7040) );
  NOR2_X1 U8396 ( .A1(n7049), .A2(n7477), .ZN(n7048) );
  INV_X1 U8397 ( .A(n7050), .ZN(n7049) );
  AND2_X1 U8398 ( .A1(n13152), .A2(n13151), .ZN(n13153) );
  AND2_X1 U8399 ( .A1(n13150), .A2(n13149), .ZN(n13151) );
  OR2_X1 U8400 ( .A1(n13046), .A2(n13045), .ZN(n7690) );
  AND2_X1 U8401 ( .A1(n13046), .A2(n13045), .ZN(n13048) );
  INV_X1 U8402 ( .A(n9212), .ZN(n6990) );
  NOR2_X1 U8403 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6989) );
  NAND2_X1 U8404 ( .A1(n15262), .A2(n11040), .ZN(n11041) );
  NAND2_X1 U8405 ( .A1(n13276), .A2(n7234), .ZN(n7233) );
  AOI21_X1 U8406 ( .B1(n7164), .B2(n7166), .A(n13320), .ZN(n7162) );
  OR2_X1 U8407 ( .A1(n10586), .A2(n13591), .ZN(n10825) );
  OR2_X1 U8408 ( .A1(n10571), .A2(n10570), .ZN(n10586) );
  NAND2_X1 U8409 ( .A1(n10390), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10571) );
  INV_X1 U8410 ( .A(n10392), .ZN(n10390) );
  OR2_X1 U8411 ( .A1(n10134), .A2(n10133), .ZN(n10392) );
  INV_X1 U8412 ( .A(n9996), .ZN(n6780) );
  AND2_X1 U8413 ( .A1(n10449), .A2(n10453), .ZN(n10017) );
  NAND2_X1 U8414 ( .A1(n9457), .A2(n10474), .ZN(n9944) );
  AND2_X1 U8415 ( .A1(n7662), .A2(n6992), .ZN(n7661) );
  INV_X1 U8416 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9279) );
  NOR2_X1 U8417 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7662) );
  NAND2_X1 U8418 ( .A1(n10034), .A2(n7205), .ZN(n7204) );
  NAND2_X1 U8419 ( .A1(n7206), .A2(n11765), .ZN(n7205) );
  INV_X1 U8420 ( .A(n10034), .ZN(n7198) );
  OR2_X1 U8421 ( .A1(n14639), .A2(n14316), .ZN(n8303) );
  OR2_X1 U8422 ( .A1(n8028), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8100) );
  NOR2_X1 U8423 ( .A1(n14442), .A2(n14639), .ZN(n8316) );
  INV_X1 U8424 ( .A(n8240), .ZN(n8254) );
  INV_X1 U8425 ( .A(n8297), .ZN(n7253) );
  OAI21_X1 U8426 ( .B1(n7254), .B2(n7253), .A(n14522), .ZN(n7252) );
  AND2_X1 U8427 ( .A1(n7397), .A2(n8220), .ZN(n6914) );
  OR2_X1 U8428 ( .A1(n8158), .A2(n8157), .ZN(n8174) );
  INV_X1 U8429 ( .A(n6873), .ZN(n6870) );
  NAND2_X1 U8430 ( .A1(n7499), .A2(n7497), .ZN(n7495) );
  NAND2_X1 U8431 ( .A1(n15147), .A2(n14122), .ZN(n7497) );
  INV_X1 U8432 ( .A(n14422), .ZN(n6811) );
  OAI21_X1 U8433 ( .B1(n14470), .B2(n6920), .A(n6919), .ZN(n6918) );
  NAND2_X1 U8434 ( .A1(n14450), .A2(n7694), .ZN(n6920) );
  AOI21_X1 U8435 ( .B1(n6922), .B2(n14450), .A(n6923), .ZN(n6919) );
  INV_X1 U8436 ( .A(n14493), .ZN(n14488) );
  NAND2_X1 U8437 ( .A1(n13064), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6814) );
  AOI21_X1 U8438 ( .B1(n7590), .B2(n7588), .A(n6707), .ZN(n7587) );
  INV_X1 U8439 ( .A(n7590), .ZN(n7589) );
  INV_X1 U8440 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7705) );
  NAND2_X1 U8441 ( .A1(n7582), .A2(n6695), .ZN(n7585) );
  AND2_X1 U8442 ( .A1(n7584), .A2(n7814), .ZN(n7583) );
  AOI21_X1 U8443 ( .B1(n7569), .B2(n6772), .A(n6771), .ZN(n6770) );
  INV_X1 U8444 ( .A(n7569), .ZN(n6773) );
  INV_X1 U8445 ( .A(n7810), .ZN(n6771) );
  AND2_X1 U8446 ( .A1(n7814), .A2(n7813), .ZN(n8116) );
  NAND2_X1 U8447 ( .A1(n7793), .A2(SI_11_), .ZN(n8025) );
  NAND2_X1 U8448 ( .A1(n7262), .A2(n7566), .ZN(n8021) );
  NOR2_X1 U8449 ( .A1(n7986), .A2(n7972), .ZN(n7263) );
  AND2_X1 U8450 ( .A1(n6766), .A2(n6764), .ZN(n7973) );
  INV_X1 U8451 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7928) );
  INV_X1 U8452 ( .A(n7417), .ZN(n7415) );
  NAND2_X1 U8453 ( .A1(n6774), .A2(n6775), .ZN(n7769) );
  OAI21_X1 U8454 ( .B1(n6777), .B2(n6776), .A(n9038), .ZN(n6774) );
  INV_X1 U8455 ( .A(n7413), .ZN(n6777) );
  AND2_X1 U8456 ( .A1(n7586), .A2(n7768), .ZN(n7250) );
  XNOR2_X1 U8457 ( .A(n7459), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14797) );
  NOR2_X1 U8458 ( .A1(n14775), .A2(n14774), .ZN(n14784) );
  OAI21_X1 U8459 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14782), .A(n14781), .ZN(
        n14824) );
  AOI22_X1 U8460 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14843), .B1(n14842), 
        .B2(n14841), .ZN(n14850) );
  NOR2_X1 U8461 ( .A1(n14860), .A2(n14859), .ZN(n14863) );
  AND2_X1 U8462 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14858), .ZN(n14859) );
  OAI22_X1 U8463 ( .A1(n11879), .A2(n7366), .B1(n11660), .B2(n7367), .ZN(
        n11662) );
  AND2_X1 U8464 ( .A1(n11661), .A2(n7368), .ZN(n7367) );
  NAND2_X1 U8465 ( .A1(n11659), .A2(n11654), .ZN(n7366) );
  INV_X1 U8466 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U8467 ( .A1(n7371), .A2(n10553), .ZN(n7370) );
  AND2_X1 U8468 ( .A1(n10216), .A2(n6575), .ZN(n7371) );
  NAND2_X1 U8469 ( .A1(n8434), .A2(n8433), .ZN(n8730) );
  INV_X1 U8470 ( .A(n8718), .ZN(n8434) );
  NAND2_X1 U8471 ( .A1(n11638), .A2(n11639), .ZN(n11640) );
  AND2_X1 U8472 ( .A1(n7375), .A2(n11091), .ZN(n11141) );
  AND2_X1 U8473 ( .A1(n7082), .A2(n7081), .ZN(n11916) );
  NAND2_X1 U8474 ( .A1(n11654), .A2(n7369), .ZN(n7081) );
  NAND2_X1 U8475 ( .A1(n8440), .A2(n8439), .ZN(n8782) );
  OAI21_X1 U8476 ( .B1(n11098), .B2(n7093), .A(n7091), .ZN(n7372) );
  INV_X1 U8477 ( .A(n7092), .ZN(n7091) );
  OAI21_X1 U8478 ( .B1(n7098), .B2(n7093), .A(n7373), .ZN(n7092) );
  NAND2_X1 U8479 ( .A1(n11627), .A2(n12478), .ZN(n7373) );
  NAND2_X1 U8480 ( .A1(n8430), .A2(n8429), .ZN(n8676) );
  INV_X1 U8481 ( .A(n8662), .ZN(n8430) );
  AND2_X1 U8482 ( .A1(n12145), .A2(n11959), .ZN(n12144) );
  AND4_X1 U8483 ( .A1(n8589), .A2(n8588), .A3(n8587), .A4(n8586), .ZN(n11086)
         );
  AND2_X1 U8484 ( .A1(n9547), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9583) );
  OAI21_X1 U8485 ( .B1(n9664), .B2(n15522), .A(n6754), .ZN(n9586) );
  NAND2_X1 U8486 ( .A1(n9664), .A2(n15522), .ZN(n6754) );
  AOI21_X1 U8487 ( .B1(n6949), .B2(n9584), .A(n9583), .ZN(n9585) );
  AND2_X1 U8488 ( .A1(n6727), .A2(n6726), .ZN(n9671) );
  NAND2_X1 U8489 ( .A1(n6728), .A2(n9697), .ZN(n6727) );
  NAND2_X1 U8490 ( .A1(n9671), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U8491 ( .A1(n9707), .A2(n9708), .ZN(n9824) );
  AND2_X1 U8492 ( .A1(n6745), .A2(n6744), .ZN(n9704) );
  NAND2_X1 U8493 ( .A1(n9702), .A2(n7338), .ZN(n6744) );
  NAND2_X1 U8494 ( .A1(n9703), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n6745) );
  NOR2_X1 U8495 ( .A1(n9704), .A2(n9705), .ZN(n9820) );
  NAND2_X1 U8496 ( .A1(n7324), .A2(n9886), .ZN(n9825) );
  AND2_X1 U8497 ( .A1(n7321), .A2(n7324), .ZN(n9888) );
  NOR2_X1 U8498 ( .A1(n9887), .A2(n10525), .ZN(n7321) );
  INV_X1 U8499 ( .A(n9888), .ZN(n7320) );
  NAND2_X1 U8500 ( .A1(n9887), .A2(n7325), .ZN(n7323) );
  OR2_X1 U8501 ( .A1(n10171), .A2(n6699), .ZN(n10258) );
  OR2_X1 U8502 ( .A1(n15444), .A2(n10634), .ZN(n6725) );
  AND2_X1 U8503 ( .A1(n6725), .A2(n6724), .ZN(n10801) );
  INV_X1 U8504 ( .A(n10635), .ZN(n6724) );
  NAND2_X1 U8505 ( .A1(n15459), .A2(n10625), .ZN(n10626) );
  NAND2_X1 U8506 ( .A1(n10626), .A2(n10627), .ZN(n10804) );
  INV_X1 U8507 ( .A(n7336), .ZN(n10922) );
  NAND2_X1 U8508 ( .A1(n6995), .A2(n6632), .ZN(n7335) );
  INV_X1 U8509 ( .A(n6970), .ZN(n11215) );
  NAND2_X1 U8510 ( .A1(n11253), .A2(n11222), .ZN(n11224) );
  OR2_X1 U8511 ( .A1(n11259), .A2(n11258), .ZN(n11261) );
  NAND2_X1 U8512 ( .A1(n12184), .A2(n12193), .ZN(n12207) );
  OR2_X1 U8513 ( .A1(n12185), .A2(n12197), .ZN(n6732) );
  OR2_X1 U8514 ( .A1(n14914), .A2(n14915), .ZN(n14912) );
  NAND2_X1 U8515 ( .A1(n7332), .A2(n7331), .ZN(n7330) );
  NAND2_X1 U8516 ( .A1(n12234), .A2(n12264), .ZN(n7332) );
  NAND2_X1 U8517 ( .A1(n14904), .A2(n12257), .ZN(n12254) );
  NAND2_X1 U8518 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  NOR2_X1 U8519 ( .A1(n12141), .A2(n11956), .ZN(n8872) );
  XNOR2_X1 U8520 ( .A(n11650), .B(n12321), .ZN(n12301) );
  INV_X1 U8521 ( .A(n12301), .ZN(n12304) );
  AOI21_X1 U8522 ( .B1(n7615), .B2(n7613), .A(n7612), .ZN(n7611) );
  INV_X1 U8523 ( .A(n7615), .ZN(n7614) );
  INV_X1 U8524 ( .A(n7618), .ZN(n7613) );
  NAND2_X1 U8525 ( .A1(n8857), .A2(n11964), .ZN(n12346) );
  NAND2_X1 U8526 ( .A1(n12369), .A2(n7053), .ZN(n12358) );
  NAND2_X1 U8527 ( .A1(n12104), .A2(n12172), .ZN(n7053) );
  INV_X1 U8528 ( .A(n12434), .ZN(n12405) );
  AOI21_X1 U8529 ( .B1(n7603), .B2(n7609), .A(n7601), .ZN(n7600) );
  INV_X1 U8530 ( .A(n12068), .ZN(n7601) );
  NAND2_X1 U8531 ( .A1(n12475), .A2(n6636), .ZN(n12462) );
  AOI22_X1 U8532 ( .A1(n8849), .A2(n11149), .B1(n6740), .B2(n6739), .ZN(n11167) );
  NAND2_X1 U8533 ( .A1(n11108), .A2(n12173), .ZN(n6740) );
  NOR2_X1 U8534 ( .A1(n7596), .A2(n6619), .ZN(n7595) );
  INV_X1 U8535 ( .A(n12035), .ZN(n7596) );
  AND2_X1 U8536 ( .A1(n10985), .A2(n8848), .ZN(n10774) );
  NAND2_X1 U8537 ( .A1(n8422), .A2(n8421), .ZN(n8557) );
  INV_X1 U8538 ( .A(n8541), .ZN(n8422) );
  AND4_X1 U8539 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n10844)
         );
  AND4_X1 U8540 ( .A1(n8517), .A2(n8516), .A3(n8515), .A4(n8514), .ZN(n10734)
         );
  NAND2_X1 U8541 ( .A1(n10293), .A2(n8836), .ZN(n11546) );
  NAND2_X1 U8542 ( .A1(n11546), .A2(n11542), .ZN(n11545) );
  NAND2_X1 U8543 ( .A1(n8417), .A2(n8416), .ZN(n11650) );
  OR2_X1 U8544 ( .A1(n11951), .A2(n10680), .ZN(n8416) );
  OR2_X1 U8545 ( .A1(n10681), .A2(n8813), .ZN(n8417) );
  AOI21_X1 U8546 ( .B1(n8775), .B2(n7274), .A(n7272), .ZN(n7271) );
  NAND2_X1 U8547 ( .A1(n7273), .A2(n8805), .ZN(n7272) );
  INV_X1 U8548 ( .A(n8777), .ZN(n7277) );
  AOI21_X1 U8549 ( .B1(n8777), .B2(n7276), .A(n7275), .ZN(n7274) );
  INV_X1 U8550 ( .A(n8789), .ZN(n7275) );
  INV_X1 U8551 ( .A(n8774), .ZN(n7276) );
  AOI21_X1 U8552 ( .B1(n7301), .B2(n7303), .A(n7300), .ZN(n7299) );
  INV_X1 U8553 ( .A(n8389), .ZN(n7300) );
  NAND2_X1 U8554 ( .A1(n8725), .A2(n8724), .ZN(n8727) );
  AND2_X1 U8555 ( .A1(n8385), .A2(n8384), .ZN(n8682) );
  NAND2_X1 U8556 ( .A1(n8380), .A2(n8379), .ZN(n8654) );
  OR2_X1 U8557 ( .A1(n8631), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8656) );
  AND2_X1 U8558 ( .A1(n8573), .A2(n8324), .ZN(n8325) );
  OR2_X1 U8559 ( .A1(n8535), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8550) );
  AND2_X1 U8560 ( .A1(n8359), .A2(n8357), .ZN(n8537) );
  NAND2_X1 U8561 ( .A1(n8356), .A2(n8355), .ZN(n8538) );
  XNOR2_X1 U8562 ( .A(n9063), .B(P1_DATAO_REG_4__SCAN_IN), .ZN(n8504) );
  AND2_X1 U8563 ( .A1(n9782), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8351) );
  XNOR2_X1 U8564 ( .A(n15393), .B(n12667), .ZN(n12634) );
  AND2_X1 U8565 ( .A1(n12856), .A2(n12650), .ZN(n12758) );
  OR2_X1 U8566 ( .A1(n10002), .A2(n10001), .ZN(n10009) );
  OR2_X1 U8567 ( .A1(n10719), .A2(n7477), .ZN(n7476) );
  AND2_X1 U8568 ( .A1(n6620), .A2(n7473), .ZN(n7472) );
  INV_X1 U8569 ( .A(n11195), .ZN(n7473) );
  NAND2_X1 U8570 ( .A1(n10671), .A2(n7048), .ZN(n7474) );
  NAND2_X1 U8571 ( .A1(n11372), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n11386) );
  NOR2_X1 U8572 ( .A1(n9785), .A2(n15355), .ZN(n9807) );
  INV_X1 U8573 ( .A(n10906), .ZN(n10905) );
  XNOR2_X1 U8574 ( .A(n12649), .B(n12648), .ZN(n12855) );
  AND2_X1 U8575 ( .A1(n7556), .A2(n13244), .ZN(n13174) );
  AND2_X1 U8576 ( .A1(n13111), .A2(n6685), .ZN(n7664) );
  NAND2_X1 U8577 ( .A1(n7667), .A2(n7666), .ZN(n7665) );
  NAND2_X1 U8578 ( .A1(n13154), .A2(n7558), .ZN(n13111) );
  NAND2_X1 U8579 ( .A1(n7560), .A2(n7559), .ZN(n7558) );
  NAND2_X1 U8580 ( .A1(n13103), .A2(n13104), .ZN(n7559) );
  NAND2_X1 U8581 ( .A1(n13106), .A2(n13107), .ZN(n7560) );
  XNOR2_X1 U8582 ( .A(n9224), .B(n6802), .ZN(n15217) );
  INV_X1 U8583 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6802) );
  NOR2_X1 U8584 ( .A1(n15229), .A2(n6785), .ZN(n15245) );
  NOR2_X1 U8585 ( .A1(n15224), .A2(n9198), .ZN(n6785) );
  NAND2_X1 U8586 ( .A1(n9325), .A2(n9324), .ZN(n9376) );
  OR2_X1 U8587 ( .A1(n9059), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9374) );
  INV_X1 U8588 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6840) );
  INV_X1 U8589 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6839) );
  OR2_X1 U8590 ( .A1(n6799), .A2(n6797), .ZN(n9524) );
  NAND2_X1 U8591 ( .A1(n9488), .A2(n6798), .ZN(n6797) );
  OR2_X1 U8592 ( .A1(n10580), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6798) );
  AOI21_X1 U8593 ( .B1(n9524), .B2(n9522), .A(n9523), .ZN(n11036) );
  XNOR2_X1 U8594 ( .A(n11039), .B(n15272), .ZN(n15263) );
  NAND2_X1 U8595 ( .A1(n15263), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n15262) );
  XNOR2_X1 U8596 ( .A(n11041), .B(n11054), .ZN(n15275) );
  NAND2_X1 U8597 ( .A1(n15284), .A2(n6714), .ZN(n15298) );
  NOR3_X1 U8598 ( .A1(n13311), .A2(n13493), .A3(n13303), .ZN(n13288) );
  NAND2_X1 U8599 ( .A1(n11475), .A2(n13117), .ZN(n13283) );
  INV_X1 U8600 ( .A(n13147), .ZN(n13282) );
  NAND2_X1 U8601 ( .A1(n13283), .A2(n13282), .ZN(n13281) );
  AND2_X1 U8602 ( .A1(n13118), .A2(n13117), .ZN(n13297) );
  OAI21_X1 U8603 ( .B1(n11368), .B2(n7159), .A(n7157), .ZN(n11392) );
  INV_X1 U8604 ( .A(n7158), .ZN(n7157) );
  INV_X1 U8605 ( .A(n13424), .ZN(n7016) );
  NAND2_X1 U8606 ( .A1(n7228), .A2(n7227), .ZN(n11007) );
  INV_X1 U8607 ( .A(n7177), .ZN(n7176) );
  OAI21_X1 U8608 ( .B1(n6611), .B2(n6587), .A(n10822), .ZN(n7177) );
  NAND2_X1 U8609 ( .A1(n10017), .A2(n7230), .ZN(n10384) );
  NAND2_X1 U8610 ( .A1(n7175), .A2(n7174), .ZN(n10354) );
  AOI21_X1 U8611 ( .B1(n7379), .B2(n7384), .A(n6652), .ZN(n7174) );
  NAND2_X1 U8612 ( .A1(n10354), .A2(n10353), .ZN(n10388) );
  NOR2_X1 U8613 ( .A1(n10025), .A2(n7380), .ZN(n7379) );
  INV_X1 U8614 ( .A(n7382), .ZN(n7380) );
  NAND2_X1 U8615 ( .A1(n10017), .A2(n10438), .ZN(n10358) );
  NOR2_X2 U8616 ( .A1(n10426), .A2(n15393), .ZN(n10449) );
  NAND2_X1 U8617 ( .A1(n10065), .A2(n12900), .ZN(n10418) );
  NAND2_X1 U8618 ( .A1(n12888), .A2(n7410), .ZN(n10474) );
  CLKBUF_X1 U8619 ( .A(n13120), .Z(n6954) );
  XNOR2_X1 U8620 ( .A(n6842), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13156) );
  OAI21_X1 U8621 ( .B1(n9656), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6842) );
  INV_X1 U8622 ( .A(n13261), .ZN(n13482) );
  NAND2_X1 U8623 ( .A1(n7557), .A2(n11501), .ZN(n13484) );
  NAND2_X1 U8624 ( .A1(n13885), .A2(n13068), .ZN(n7557) );
  INV_X1 U8625 ( .A(n15421), .ZN(n15379) );
  NOR2_X1 U8626 ( .A1(n6633), .A2(n7425), .ZN(n7424) );
  NAND2_X1 U8627 ( .A1(n9781), .A2(n13068), .ZN(n7426) );
  NOR2_X1 U8628 ( .A1(n9783), .A2(n15224), .ZN(n7425) );
  INV_X1 U8629 ( .A(n15405), .ZN(n13571) );
  AND2_X1 U8630 ( .A1(n15313), .A2(n13163), .ZN(n15421) );
  AND2_X1 U8631 ( .A1(n8975), .A2(n8974), .ZN(n8977) );
  NAND2_X1 U8632 ( .A1(n8967), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U8633 ( .A1(n8964), .A2(n7481), .ZN(n7480) );
  OR2_X1 U8634 ( .A1(n9095), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U8635 ( .A1(n11673), .A2(n11672), .ZN(n11679) );
  INV_X1 U8636 ( .A(n7691), .ZN(n7651) );
  OR2_X1 U8637 ( .A1(n7963), .A2(n10538), .ZN(n7977) );
  AND2_X1 U8638 ( .A1(n11736), .A2(n11728), .ZN(n7657) );
  INV_X1 U8639 ( .A(n7864), .ZN(n7853) );
  NAND2_X1 U8640 ( .A1(n13989), .A2(n13990), .ZN(n13988) );
  INV_X1 U8641 ( .A(n7656), .ZN(n7195) );
  NAND2_X1 U8642 ( .A1(n7655), .A2(n14063), .ZN(n7194) );
  NAND2_X1 U8643 ( .A1(n7655), .A2(n6902), .ZN(n7193) );
  AOI21_X1 U8644 ( .B1(n13934), .B2(n7640), .A(n7639), .ZN(n7638) );
  INV_X1 U8645 ( .A(n14016), .ZN(n7639) );
  INV_X1 U8646 ( .A(n13935), .ZN(n7640) );
  INV_X1 U8647 ( .A(n14031), .ZN(n6906) );
  AND2_X1 U8648 ( .A1(n13982), .A2(n11762), .ZN(n14014) );
  OR2_X1 U8649 ( .A1(n7977), .A2(n9154), .ZN(n7995) );
  INV_X1 U8650 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U8651 ( .A1(n11787), .A2(n14338), .ZN(n6894) );
  NAND2_X1 U8652 ( .A1(n8993), .A2(n6895), .ZN(n9605) );
  INV_X1 U8653 ( .A(n6896), .ZN(n6895) );
  OAI21_X1 U8654 ( .B1(n11794), .B2(n14099), .A(n6897), .ZN(n6896) );
  AND2_X1 U8655 ( .A1(n8992), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n8989) );
  NOR2_X1 U8656 ( .A1(n8174), .A2(n13810), .ZN(n8186) );
  NOR2_X1 U8657 ( .A1(n8049), .A2(n8048), .ZN(n8065) );
  AND2_X1 U8658 ( .A1(n8065), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8080) );
  INV_X1 U8659 ( .A(n7852), .ZN(n8241) );
  NAND2_X1 U8660 ( .A1(n7196), .A2(n11691), .ZN(n14060) );
  INV_X1 U8661 ( .A(n14062), .ZN(n7196) );
  OR2_X1 U8662 ( .A1(n8109), .A2(n8108), .ZN(n8128) );
  NAND2_X1 U8663 ( .A1(n7541), .A2(n7534), .ZN(n7533) );
  INV_X1 U8664 ( .A(n7539), .ZN(n7534) );
  AND2_X1 U8665 ( .A1(n7537), .A2(n7536), .ZN(n7535) );
  NAND2_X1 U8666 ( .A1(n7542), .A2(n7540), .ZN(n7536) );
  NAND2_X1 U8667 ( .A1(n7543), .A2(n7548), .ZN(n7542) );
  INV_X1 U8668 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14761) );
  INV_X1 U8669 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9154) );
  AND2_X1 U8670 ( .A1(n8316), .A2(n14432), .ZN(n14422) );
  XNOR2_X1 U8671 ( .A(n14253), .B(n8272), .ZN(n14299) );
  NAND2_X1 U8672 ( .A1(n14459), .A2(n14447), .ZN(n14442) );
  AND2_X1 U8673 ( .A1(n14496), .A2(n6816), .ZN(n14459) );
  NOR2_X1 U8674 ( .A1(n14652), .A2(n14659), .ZN(n6816) );
  NAND2_X1 U8675 ( .A1(n14496), .A2(n14481), .ZN(n14473) );
  INV_X1 U8676 ( .A(n8227), .ZN(n7865) );
  NAND2_X1 U8677 ( .A1(n7865), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U8678 ( .A1(n8228), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U8679 ( .A1(n6911), .A2(n6634), .ZN(n14510) );
  INV_X1 U8680 ( .A(n6916), .ZN(n6911) );
  NAND2_X1 U8681 ( .A1(n6813), .A2(n6585), .ZN(n14524) );
  INV_X1 U8682 ( .A(n14562), .ZN(n6813) );
  NOR2_X1 U8683 ( .A1(n14562), .A2(n14682), .ZN(n14537) );
  AOI21_X1 U8684 ( .B1(n6617), .B2(n6933), .A(n7399), .ZN(n6932) );
  INV_X1 U8685 ( .A(n6936), .ZN(n6933) );
  OAI21_X1 U8686 ( .B1(n14586), .B2(n14201), .A(n14200), .ZN(n14570) );
  NAND2_X1 U8687 ( .A1(n8133), .A2(n8132), .ZN(n14605) );
  NAND2_X1 U8688 ( .A1(n6886), .A2(n7257), .ZN(n14603) );
  AOI21_X1 U8689 ( .B1(n7260), .B2(n7258), .A(n6651), .ZN(n7257) );
  NAND2_X1 U8690 ( .A1(n14950), .A2(n6883), .ZN(n6886) );
  NAND2_X1 U8691 ( .A1(n14950), .A2(n8292), .ZN(n11201) );
  NAND2_X1 U8692 ( .A1(n14938), .A2(n6629), .ZN(n11030) );
  NAND2_X1 U8693 ( .A1(n14938), .A2(n14969), .ZN(n14937) );
  NOR2_X1 U8694 ( .A1(n7995), .A2(n7994), .ZN(n8009) );
  OR2_X1 U8695 ( .A1(n15097), .A2(n15089), .ZN(n15098) );
  NAND2_X1 U8696 ( .A1(n10095), .A2(n15171), .ZN(n15097) );
  AND2_X1 U8697 ( .A1(n10317), .A2(n9936), .ZN(n10095) );
  OR2_X1 U8698 ( .A1(n7941), .A2(n6930), .ZN(n6928) );
  AND2_X1 U8699 ( .A1(n6817), .A2(n15147), .ZN(n9936) );
  NOR2_X1 U8700 ( .A1(n9767), .A2(n15152), .ZN(n6817) );
  INV_X1 U8701 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7934) );
  NOR2_X1 U8702 ( .A1(n7935), .A2(n7934), .ZN(n7949) );
  OAI21_X1 U8703 ( .B1(n10189), .B2(n15152), .A(n7942), .ZN(n14272) );
  NAND2_X1 U8704 ( .A1(n6931), .A2(n7941), .ZN(n9931) );
  INV_X1 U8705 ( .A(n9929), .ZN(n6931) );
  NAND2_X1 U8706 ( .A1(n6818), .A2(n15147), .ZN(n9937) );
  NAND2_X1 U8707 ( .A1(n9683), .A2(n8278), .ZN(n9764) );
  NAND2_X1 U8708 ( .A1(n9719), .A2(n8277), .ZN(n9685) );
  NAND2_X1 U8709 ( .A1(n9685), .A2(n9684), .ZN(n9683) );
  INV_X1 U8710 ( .A(n14269), .ZN(n9684) );
  NAND2_X1 U8711 ( .A1(n9621), .A2(n8276), .ZN(n9721) );
  NAND2_X1 U8712 ( .A1(n9720), .A2(n9721), .ZN(n9719) );
  AND2_X1 U8713 ( .A1(n9722), .A2(n9725), .ZN(n9723) );
  NAND2_X1 U8714 ( .A1(n7509), .A2(n7508), .ZN(n9621) );
  INV_X1 U8715 ( .A(n9619), .ZN(n7508) );
  INV_X1 U8716 ( .A(n7509), .ZN(n14271) );
  NAND2_X1 U8717 ( .A1(n8991), .A2(n15141), .ZN(n14101) );
  INV_X1 U8718 ( .A(n14116), .ZN(n14117) );
  INV_X1 U8719 ( .A(n15159), .ZN(n15191) );
  NAND2_X1 U8720 ( .A1(n10044), .A2(n9102), .ZN(n9395) );
  XNOR2_X1 U8721 ( .A(n13067), .B(n13066), .ZN(n14088) );
  XNOR2_X1 U8722 ( .A(n13060), .B(n13059), .ZN(n13885) );
  XNOR2_X1 U8723 ( .A(n8262), .B(n8261), .ZN(n11483) );
  AND2_X1 U8724 ( .A1(n8237), .A2(n8236), .ZN(n13898) );
  AND2_X1 U8725 ( .A1(n7861), .A2(n7860), .ZN(n11444) );
  OAI21_X1 U8726 ( .B1(n8198), .B2(n6698), .A(n7575), .ZN(n8223) );
  AND2_X1 U8727 ( .A1(n7577), .A2(n7576), .ZN(n7575) );
  OR2_X1 U8728 ( .A1(n7829), .A2(n7579), .ZN(n7576) );
  NAND2_X1 U8729 ( .A1(n7707), .A2(n7224), .ZN(n7715) );
  NAND2_X1 U8730 ( .A1(n7723), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7728) );
  INV_X1 U8731 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7727) );
  OR2_X1 U8732 ( .A1(n8118), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n8120) );
  XNOR2_X1 U8733 ( .A(n8099), .B(n8098), .ZN(n11001) );
  NAND2_X1 U8734 ( .A1(n8042), .A2(n7802), .ZN(n8058) );
  NAND2_X1 U8735 ( .A1(n7568), .A2(n7784), .ZN(n7957) );
  NAND2_X1 U8736 ( .A1(n7944), .A2(n7782), .ZN(n7568) );
  INV_X1 U8737 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7912) );
  NAND2_X1 U8738 ( .A1(n7561), .A2(n7775), .ZN(n7909) );
  NAND2_X1 U8739 ( .A1(n7905), .A2(n7773), .ZN(n7561) );
  OR2_X1 U8740 ( .A1(n9302), .A2(n9301), .ZN(n7417) );
  INV_X1 U8741 ( .A(n7250), .ZN(n7885) );
  INV_X1 U8742 ( .A(n14790), .ZN(n7241) );
  XNOR2_X1 U8743 ( .A(n14785), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14786) );
  NAND2_X1 U8744 ( .A1(n6836), .A2(n6835), .ZN(n14804) );
  NAND2_X1 U8745 ( .A1(n6837), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6835) );
  OAI21_X1 U8746 ( .B1(n6837), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6838), .ZN(
        n6836) );
  NOR2_X1 U8747 ( .A1(n14770), .A2(n14769), .ZN(n14807) );
  NOR2_X1 U8748 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14803), .ZN(n14769) );
  INV_X1 U8749 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14806) );
  NAND2_X1 U8750 ( .A1(n15545), .A2(n15546), .ZN(n6821) );
  AOI22_X1 U8751 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n14831), .B1(n14830), 
        .B2(n14829), .ZN(n14835) );
  NAND2_X1 U8752 ( .A1(n7096), .A2(n7097), .ZN(n11825) );
  NAND2_X1 U8753 ( .A1(n11098), .A2(n7098), .ZN(n7096) );
  OAI21_X1 U8754 ( .B1(n11646), .B2(n11645), .A(n11644), .ZN(n11834) );
  NOR2_X1 U8755 ( .A1(n11834), .A2(n12320), .ZN(n11833) );
  NAND2_X1 U8756 ( .A1(n8760), .A2(n8759), .ZN(n12338) );
  OR2_X1 U8757 ( .A1(n11951), .A2(n10156), .ZN(n8759) );
  AND3_X1 U8758 ( .A1(n8595), .A2(n8594), .A3(n8593), .ZN(n10869) );
  NAND2_X1 U8759 ( .A1(n10215), .A2(n10214), .ZN(n10217) );
  OR2_X1 U8760 ( .A1(n8503), .A2(n9033), .ZN(n8495) );
  NAND2_X1 U8761 ( .A1(n7104), .A2(n7109), .ZN(n11840) );
  NAND2_X1 U8762 ( .A1(n11871), .A2(n7111), .ZN(n7104) );
  NAND2_X1 U8763 ( .A1(n7087), .A2(n7086), .ZN(n9869) );
  AND2_X1 U8764 ( .A1(n8788), .A2(n8787), .ZN(n11860) );
  AND2_X1 U8765 ( .A1(n8675), .A2(n8674), .ZN(n12539) );
  AND3_X1 U8766 ( .A1(n8525), .A2(n8524), .A3(n8523), .ZN(n10562) );
  NAND2_X1 U8767 ( .A1(n10859), .A2(n10858), .ZN(n11088) );
  AOI21_X1 U8768 ( .B1(n11871), .B2(n7105), .A(n7102), .ZN(n7101) );
  NAND2_X1 U8769 ( .A1(n7103), .A2(n7115), .ZN(n7102) );
  AND2_X1 U8770 ( .A1(n11891), .A2(n11888), .ZN(n7115) );
  NAND2_X1 U8771 ( .A1(n11098), .A2(n11097), .ZN(n11624) );
  AND2_X1 U8772 ( .A1(n7378), .A2(n7377), .ZN(n11899) );
  INV_X1 U8773 ( .A(n12173), .ZN(n11149) );
  OAI21_X1 U8774 ( .B1(n11871), .B2(n11872), .A(n7114), .ZN(n11909) );
  AND3_X1 U8775 ( .A1(n10849), .A2(n10732), .A3(n10846), .ZN(n10793) );
  AND2_X1 U8776 ( .A1(n9748), .A2(n12159), .ZN(n11920) );
  INV_X1 U8777 ( .A(n7372), .ZN(n11930) );
  OR2_X1 U8778 ( .A1(n10212), .A2(n10211), .ZN(n11938) );
  AND2_X1 U8779 ( .A1(n10340), .A2(n8833), .ZN(n11814) );
  INV_X1 U8780 ( .A(n11860), .ZN(n12306) );
  INV_X1 U8781 ( .A(n11099), .ZN(n12464) );
  INV_X1 U8782 ( .A(n11086), .ZN(n12174) );
  NAND4_X2 U8783 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), .ZN(n12182)
         );
  OR2_X1 U8784 ( .A1(n9735), .A2(n12615), .ZN(n12181) );
  INV_X1 U8785 ( .A(n7340), .ZN(n9669) );
  XNOR2_X1 U8786 ( .A(n8506), .B(P3_IR_REG_4__SCAN_IN), .ZN(n9816) );
  XNOR2_X1 U8787 ( .A(n10258), .B(n10254), .ZN(n10173) );
  OR2_X1 U8788 ( .A1(n15451), .A2(n15447), .ZN(n10618) );
  XNOR2_X1 U8789 ( .A(n7336), .B(n10929), .ZN(n10803) );
  NOR2_X1 U8790 ( .A1(n10924), .A2(n10923), .ZN(n10927) );
  XNOR2_X1 U8791 ( .A(n6970), .B(n11257), .ZN(n11251) );
  INV_X1 U8792 ( .A(n6995), .ZN(n11250) );
  INV_X1 U8793 ( .A(n12184), .ZN(n12183) );
  INV_X1 U8794 ( .A(n7335), .ZN(n11217) );
  INV_X1 U8795 ( .A(n6731), .ZN(n12210) );
  NAND2_X1 U8796 ( .A1(n12223), .A2(n12224), .ZN(n12248) );
  XNOR2_X1 U8797 ( .A(n12233), .B(n12252), .ZN(n14902) );
  INV_X1 U8798 ( .A(n6997), .ZN(n14901) );
  AND2_X1 U8799 ( .A1(n12235), .A2(n12234), .ZN(n7014) );
  INV_X1 U8800 ( .A(n12234), .ZN(n7333) );
  OAI21_X1 U8801 ( .B1(n11342), .B2(n12132), .A(n11341), .ZN(n12298) );
  NAND2_X1 U8802 ( .A1(n12319), .A2(n12318), .ZN(n12317) );
  AND2_X1 U8803 ( .A1(n7617), .A2(n7620), .ZN(n12344) );
  NAND2_X1 U8804 ( .A1(n12366), .A2(n7618), .ZN(n7617) );
  AND2_X1 U8805 ( .A1(n12366), .A2(n8736), .ZN(n12356) );
  NAND2_X1 U8806 ( .A1(n12384), .A2(n7054), .ZN(n12371) );
  AND2_X1 U8807 ( .A1(n7621), .A2(n8710), .ZN(n12393) );
  NAND2_X1 U8808 ( .A1(n12399), .A2(n7342), .ZN(n12380) );
  INV_X1 U8809 ( .A(n7621), .ZN(n12396) );
  AND2_X1 U8810 ( .A1(n12424), .A2(n12423), .ZN(n12534) );
  NAND2_X1 U8811 ( .A1(n8689), .A2(n8688), .ZN(n12535) );
  AND2_X1 U8812 ( .A1(n12436), .A2(n12435), .ZN(n12538) );
  AND2_X1 U8813 ( .A1(n12454), .A2(n12453), .ZN(n12542) );
  NAND2_X1 U8814 ( .A1(n7604), .A2(n7605), .ZN(n12459) );
  OR2_X1 U8815 ( .A1(n11165), .A2(n7609), .ZN(n7604) );
  NAND2_X1 U8816 ( .A1(n11163), .A2(n12058), .ZN(n12473) );
  INV_X1 U8817 ( .A(n10869), .ZN(n15514) );
  NAND2_X1 U8818 ( .A1(n7347), .A2(n7348), .ZN(n11017) );
  NAND2_X1 U8819 ( .A1(n8846), .A2(n7349), .ZN(n7347) );
  NAND2_X1 U8820 ( .A1(n10782), .A2(n12027), .ZN(n7599) );
  NAND2_X1 U8821 ( .A1(n12159), .A2(n9753), .ZN(n12387) );
  INV_X1 U8822 ( .A(n12151), .ZN(n11544) );
  NAND2_X1 U8823 ( .A1(n10243), .A2(n10242), .ZN(n12488) );
  INV_X1 U8824 ( .A(n12387), .ZN(n12485) );
  NAND2_X1 U8825 ( .A1(n15538), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7007) );
  NAND2_X1 U8826 ( .A1(n11947), .A2(n11946), .ZN(n12563) );
  INV_X1 U8827 ( .A(n11957), .ZN(n12569) );
  INV_X1 U8828 ( .A(n12295), .ZN(n11927) );
  INV_X1 U8829 ( .A(n11650), .ZN(n12573) );
  AND2_X1 U8830 ( .A1(n8742), .A2(n8741), .ZN(n12589) );
  OR2_X1 U8831 ( .A1(n11951), .A2(n9833), .ZN(n8741) );
  OR2_X1 U8832 ( .A1(n9834), .A2(n8813), .ZN(n8742) );
  AND2_X1 U8833 ( .A1(n8703), .A2(n8702), .ZN(n12598) );
  OR2_X1 U8834 ( .A1(n9618), .A2(n8813), .ZN(n8703) );
  AND2_X1 U8835 ( .A1(n8902), .A2(n8901), .ZN(n12616) );
  OR2_X1 U8836 ( .A1(n8915), .A2(P3_D_REG_0__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U8837 ( .A1(n9536), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12615) );
  NAND2_X1 U8838 ( .A1(n8894), .A2(n7630), .ZN(n6743) );
  INV_X1 U8839 ( .A(n8917), .ZN(n10875) );
  NAND2_X1 U8840 ( .A1(n8778), .A2(n8777), .ZN(n8790) );
  NAND2_X1 U8841 ( .A1(n8775), .A2(n8774), .ZN(n8778) );
  NAND2_X1 U8842 ( .A1(n7290), .A2(n7289), .ZN(n8765) );
  INV_X1 U8843 ( .A(n7287), .ZN(n7290) );
  AOI21_X1 U8844 ( .B1(n8399), .B2(n8398), .A(n7291), .ZN(n7287) );
  NAND2_X1 U8845 ( .A1(n8740), .A2(n8393), .ZN(n8750) );
  XNOR2_X1 U8846 ( .A(n8333), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12163) );
  NAND2_X1 U8847 ( .A1(n8340), .A2(n8339), .ZN(n11990) );
  INV_X1 U8848 ( .A(SI_20_), .ZN(n9717) );
  OAI21_X1 U8849 ( .B1(n8697), .B2(n7303), .A(n7301), .ZN(n8714) );
  NAND2_X1 U8850 ( .A1(n8699), .A2(n8387), .ZN(n8712) );
  INV_X1 U8851 ( .A(SI_17_), .ZN(n9512) );
  INV_X1 U8852 ( .A(SI_16_), .ZN(n13778) );
  NAND2_X1 U8853 ( .A1(n8629), .A2(n8375), .ZN(n8641) );
  INV_X1 U8854 ( .A(SI_13_), .ZN(n9128) );
  NAND2_X1 U8855 ( .A1(n7315), .A2(n7313), .ZN(n8625) );
  NAND2_X1 U8856 ( .A1(n7315), .A2(n7316), .ZN(n8623) );
  INV_X1 U8857 ( .A(SI_12_), .ZN(n13820) );
  NAND2_X1 U8858 ( .A1(n8369), .A2(n8368), .ZN(n8604) );
  INV_X1 U8859 ( .A(SI_10_), .ZN(n13829) );
  NAND2_X1 U8860 ( .A1(n7284), .A2(n7282), .ZN(n8581) );
  NAND2_X1 U8861 ( .A1(n7284), .A2(n8364), .ZN(n8579) );
  NAND2_X1 U8862 ( .A1(n8462), .A2(n8463), .ZN(n9546) );
  INV_X1 U8863 ( .A(n6734), .ZN(n8463) );
  OAI21_X1 U8864 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(P3_IR_REG_31__SCAN_IN), .A(
        n6735), .ZN(n6734) );
  NAND2_X1 U8865 ( .A1(n7462), .A2(n7461), .ZN(n12785) );
  INV_X1 U8866 ( .A(n9808), .ZN(n7461) );
  INV_X1 U8867 ( .A(n9809), .ZN(n7462) );
  OR2_X1 U8868 ( .A1(n12854), .A2(n12677), .ZN(n12852) );
  NAND2_X1 U8869 ( .A1(n12715), .A2(n12663), .ZN(n12721) );
  OAI21_X1 U8870 ( .B1(n10063), .B2(n7485), .A(n7482), .ZN(n7017) );
  AOI21_X1 U8871 ( .B1(n7486), .B2(n7484), .A(n7483), .ZN(n7482) );
  INV_X1 U8872 ( .A(n7486), .ZN(n7485) );
  INV_X1 U8873 ( .A(n7032), .ZN(n7031) );
  INV_X1 U8874 ( .A(n7027), .ZN(n7026) );
  NAND2_X1 U8875 ( .A1(n7464), .A2(n7025), .ZN(n7024) );
  NAND2_X1 U8876 ( .A1(n11455), .A2(n11454), .ZN(n13314) );
  NAND2_X1 U8877 ( .A1(n7035), .A2(n12678), .ZN(n7042) );
  NAND2_X1 U8878 ( .A1(n12707), .A2(n12706), .ZN(n7039) );
  NAND2_X1 U8879 ( .A1(n9783), .A2(n13910), .ZN(n6993) );
  AOI21_X1 U8880 ( .B1(n12663), .B2(n7468), .A(n6664), .ZN(n7467) );
  INV_X1 U8881 ( .A(n12663), .ZN(n7469) );
  NAND2_X1 U8882 ( .A1(n7474), .A2(n6620), .ZN(n11194) );
  NAND2_X1 U8883 ( .A1(n7463), .A2(n10204), .ZN(n10210) );
  NAND2_X1 U8884 ( .A1(n9908), .A2(n9795), .ZN(n7463) );
  NAND2_X1 U8885 ( .A1(n12776), .A2(n12657), .ZN(n12828) );
  NAND2_X1 U8886 ( .A1(n10113), .A2(n7486), .ZN(n12834) );
  NAND2_X1 U8887 ( .A1(n10113), .A2(n10112), .ZN(n12833) );
  AND2_X1 U8888 ( .A1(n9807), .A2(n13168), .ZN(n12838) );
  AND2_X1 U8889 ( .A1(n11489), .A2(n11468), .ZN(n13300) );
  NAND2_X1 U8890 ( .A1(n7023), .A2(n7488), .ZN(n12856) );
  NOR2_X1 U8891 ( .A1(n12853), .A2(n12677), .ZN(n7488) );
  INV_X1 U8892 ( .A(n12855), .ZN(n7023) );
  NOR2_X1 U8893 ( .A1(n11492), .A2(n12788), .ZN(n6784) );
  NAND2_X1 U8894 ( .A1(n9464), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9298) );
  OAI21_X1 U8895 ( .B1(n9224), .B2(n13474), .A(n6801), .ZN(n15213) );
  NAND2_X1 U8896 ( .A1(n9224), .A2(n13474), .ZN(n6801) );
  OAI21_X1 U8897 ( .B1(n15237), .B2(n6805), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15210) );
  INV_X1 U8898 ( .A(n6787), .ZN(n15231) );
  NAND2_X1 U8899 ( .A1(n6792), .A2(n6790), .ZN(n9322) );
  NAND2_X1 U8900 ( .A1(n6796), .A2(n6791), .ZN(n6790) );
  INV_X1 U8901 ( .A(n6793), .ZN(n6791) );
  INV_X1 U8902 ( .A(n6799), .ZN(n9489) );
  INV_X1 U8903 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7766) );
  XNOR2_X1 U8904 ( .A(n6789), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13243) );
  OR2_X1 U8905 ( .A1(n13232), .A2(n13231), .ZN(n6789) );
  AOI21_X1 U8906 ( .B1(n11517), .B2(n15409), .A(n11516), .ZN(n13486) );
  NAND2_X1 U8907 ( .A1(n11515), .A2(n11514), .ZN(n11516) );
  XNOR2_X1 U8908 ( .A(n11510), .B(n11509), .ZN(n11517) );
  INV_X1 U8909 ( .A(n13337), .ZN(n13324) );
  OAI21_X1 U8910 ( .B1(n13364), .B2(n7166), .A(n7164), .ZN(n13323) );
  NAND2_X1 U8911 ( .A1(n7163), .A2(n7167), .ZN(n13343) );
  NAND2_X1 U8912 ( .A1(n13364), .A2(n7169), .ZN(n7163) );
  NAND2_X1 U8913 ( .A1(n7427), .A2(n7428), .ZN(n13351) );
  NAND2_X1 U8914 ( .A1(n7171), .A2(n11417), .ZN(n13348) );
  NAND2_X1 U8915 ( .A1(n7172), .A2(n7173), .ZN(n7171) );
  NAND2_X1 U8916 ( .A1(n7431), .A2(n11529), .ZN(n13366) );
  OR2_X1 U8917 ( .A1(n13389), .A2(n11528), .ZN(n7431) );
  NAND2_X1 U8918 ( .A1(n13412), .A2(n11379), .ZN(n13405) );
  NAND2_X1 U8919 ( .A1(n11368), .A2(n11367), .ZN(n13410) );
  NAND2_X1 U8920 ( .A1(n13447), .A2(n11523), .ZN(n13429) );
  NAND2_X1 U8921 ( .A1(n13451), .A2(n11357), .ZN(n13428) );
  NAND2_X1 U8922 ( .A1(n7435), .A2(n7436), .ZN(n10896) );
  NAND2_X1 U8923 ( .A1(n10644), .A2(n10601), .ZN(n10821) );
  NAND2_X1 U8924 ( .A1(n7439), .A2(n10584), .ZN(n10838) );
  OR2_X1 U8925 ( .A1(n10643), .A2(n10583), .ZN(n7439) );
  NAND2_X1 U8926 ( .A1(n10599), .A2(n10598), .ZN(n10646) );
  NAND2_X1 U8927 ( .A1(n7381), .A2(n7382), .ZN(n10026) );
  NAND2_X1 U8928 ( .A1(n7381), .A2(n7379), .ZN(n10442) );
  NAND2_X1 U8929 ( .A1(n6781), .A2(n9996), .ZN(n10349) );
  NAND2_X1 U8930 ( .A1(n10404), .A2(n10023), .ZN(n10447) );
  INV_X1 U8931 ( .A(n15370), .ZN(n10472) );
  NAND2_X1 U8932 ( .A1(n13472), .A2(n13459), .ZN(n13420) );
  INV_X1 U8933 ( .A(n13467), .ZN(n13440) );
  AND2_X1 U8934 ( .A1(n13472), .A2(n13244), .ZN(n13467) );
  OR2_X1 U8935 ( .A1(n13082), .A2(n9292), .ZN(n9295) );
  INV_X1 U8936 ( .A(n13420), .ZN(n13471) );
  INV_X2 U8937 ( .A(n15441), .ZN(n15443) );
  NAND2_X1 U8938 ( .A1(n7394), .A2(n6955), .ZN(n13863) );
  NOR2_X1 U8939 ( .A1(n13488), .A2(n6589), .ZN(n6955) );
  AND2_X1 U8940 ( .A1(n9787), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15358) );
  CLKBUF_X1 U8941 ( .A(n15336), .Z(n15353) );
  INV_X1 U8942 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9280) );
  XNOR2_X1 U8943 ( .A(n8969), .B(P2_IR_REG_24__SCAN_IN), .ZN(n13904) );
  NAND2_X1 U8944 ( .A1(n8968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U8945 ( .A1(n8986), .A2(n8985), .ZN(n8968) );
  INV_X1 U8946 ( .A(n10346), .ZN(n13155) );
  INV_X1 U8947 ( .A(n6984), .ZN(n13244) );
  INV_X1 U8948 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9837) );
  INV_X1 U8949 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13792) );
  INV_X1 U8950 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9600) );
  INV_X1 U8951 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9615) );
  INV_X1 U8952 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9444) );
  INV_X1 U8953 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9450) );
  INV_X1 U8954 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9131) );
  INV_X1 U8955 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n13821) );
  INV_X1 U8956 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9094) );
  INV_X1 U8957 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9084) );
  INV_X1 U8958 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U8960 ( .A1(n10537), .A2(n10536), .ZN(n10696) );
  NAND2_X1 U8961 ( .A1(n11679), .A2(n11678), .ZN(n13920) );
  NAND2_X1 U8962 ( .A1(n13933), .A2(n13935), .ZN(n7637) );
  OAI21_X1 U8963 ( .B1(n11118), .B2(n11117), .A(n11116), .ZN(n6904) );
  NOR2_X1 U8964 ( .A1(n10038), .A2(n7691), .ZN(n13942) );
  NAND2_X1 U8965 ( .A1(n13948), .A2(n6628), .ZN(n13950) );
  NAND2_X1 U8966 ( .A1(n10696), .A2(n10695), .ZN(n10697) );
  OR2_X1 U8967 ( .A1(n7896), .A2(n9038), .ZN(n7878) );
  INV_X1 U8968 ( .A(n6980), .ZN(n6979) );
  NAND2_X1 U8969 ( .A1(n11729), .A2(n11728), .ZN(n13971) );
  INV_X1 U8970 ( .A(n7187), .ZN(n7181) );
  XNOR2_X1 U8971 ( .A(n7192), .B(n10041), .ZN(n10187) );
  NAND2_X1 U8972 ( .A1(n13940), .A2(n7653), .ZN(n7192) );
  NAND2_X1 U8973 ( .A1(n11276), .A2(n11275), .ZN(n11278) );
  INV_X1 U8974 ( .A(n7652), .ZN(n10038) );
  OR2_X1 U8975 ( .A1(n7896), .A2(n9054), .ZN(n7897) );
  INV_X1 U8976 ( .A(n6952), .ZN(n6951) );
  OAI21_X1 U8977 ( .B1(n14242), .B2(n9452), .A(n6614), .ZN(n6952) );
  AND2_X1 U8978 ( .A1(n8156), .A2(n8155), .ZN(n14198) );
  INV_X1 U8979 ( .A(n7186), .ZN(n7180) );
  NAND2_X1 U8980 ( .A1(n7185), .A2(n7183), .ZN(n7182) );
  OAI21_X1 U8981 ( .B1(n11773), .B2(n7647), .A(n7644), .ZN(n14049) );
  NAND2_X1 U8982 ( .A1(n13984), .A2(n11774), .ZN(n14050) );
  NAND2_X1 U8983 ( .A1(n11692), .A2(n6903), .ZN(n14062) );
  INV_X1 U8984 ( .A(n10189), .ZN(n14333) );
  NAND2_X1 U8985 ( .A1(n14076), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7899) );
  OR2_X1 U8986 ( .A1(n14081), .A2(n9017), .ZN(n7889) );
  INV_X1 U8987 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U8988 ( .A1(n14088), .A2(n14087), .B1(n14086), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n14633) );
  INV_X1 U8989 ( .A(n14415), .ZN(n14636) );
  OAI21_X1 U8990 ( .B1(n14470), .B2(n6924), .A(n6921), .ZN(n14438) );
  NOR2_X1 U8991 ( .A1(n14448), .A2(n7267), .ZN(n14647) );
  AND2_X1 U8992 ( .A1(n14449), .A2(n14450), .ZN(n7267) );
  NAND2_X1 U8993 ( .A1(n14452), .A2(n7507), .ZN(n14449) );
  NAND2_X1 U8994 ( .A1(n14470), .A2(n6603), .ZN(n14456) );
  NOR2_X1 U8995 ( .A1(n14491), .A2(n7408), .ZN(n14472) );
  AND2_X1 U8996 ( .A1(n6876), .A2(n7511), .ZN(n14469) );
  NAND2_X1 U8997 ( .A1(n14508), .A2(n7689), .ZN(n14492) );
  NAND2_X1 U8998 ( .A1(n14542), .A2(n8297), .ZN(n14523) );
  NAND2_X1 U8999 ( .A1(n7398), .A2(n8210), .ZN(n14521) );
  NAND2_X1 U9000 ( .A1(n14533), .A2(n14545), .ZN(n7398) );
  NAND2_X1 U9001 ( .A1(n14687), .A2(n8296), .ZN(n14544) );
  NAND2_X1 U9002 ( .A1(n8173), .A2(n8172), .ZN(n14581) );
  NAND2_X1 U9003 ( .A1(n14611), .A2(n8149), .ZN(n14592) );
  NAND2_X1 U9004 ( .A1(n8143), .A2(n8142), .ZN(n14710) );
  NAND2_X1 U9005 ( .A1(n11199), .A2(n8293), .ZN(n11324) );
  NAND2_X1 U9006 ( .A1(n6937), .A2(n14173), .ZN(n11319) );
  NAND2_X1 U9007 ( .A1(n8291), .A2(n6885), .ZN(n14950) );
  AND2_X1 U9008 ( .A1(n14289), .A2(n8290), .ZN(n6885) );
  NAND2_X1 U9009 ( .A1(n8291), .A2(n8290), .ZN(n10980) );
  NAND2_X1 U9010 ( .A1(n11025), .A2(n8072), .ZN(n10972) );
  NAND2_X1 U9011 ( .A1(n15057), .A2(n6873), .ZN(n6872) );
  NAND2_X1 U9012 ( .A1(n7248), .A2(n8029), .ZN(n14934) );
  NAND2_X1 U9013 ( .A1(n10579), .A2(n14087), .ZN(n7248) );
  NAND2_X1 U9014 ( .A1(n8286), .A2(n8285), .ZN(n14936) );
  NAND2_X1 U9015 ( .A1(n15057), .A2(n15056), .ZN(n8286) );
  NAND2_X1 U9016 ( .A1(n8007), .A2(n8006), .ZN(n15188) );
  AND2_X1 U9017 ( .A1(n15087), .A2(n7985), .ZN(n15065) );
  NAND2_X1 U9018 ( .A1(n7992), .A2(n7991), .ZN(n15076) );
  NAND2_X1 U9019 ( .A1(n6879), .A2(n8282), .ZN(n15096) );
  NAND2_X1 U9020 ( .A1(n10094), .A2(n10093), .ZN(n6879) );
  OR2_X1 U9021 ( .A1(n14431), .A2(n14598), .ZN(n14583) );
  AND2_X1 U9022 ( .A1(n15104), .A2(n15139), .ZN(n14627) );
  NOR2_X1 U9023 ( .A1(n14426), .A2(n6807), .ZN(n6806) );
  NAND2_X1 U9024 ( .A1(n6999), .A2(n15195), .ZN(n6998) );
  NAND2_X1 U9025 ( .A1(n6808), .A2(n6716), .ZN(n6807) );
  INV_X1 U9026 ( .A(n6982), .ZN(n6981) );
  OR2_X1 U9027 ( .A1(n14673), .A2(n14672), .ZN(n14726) );
  NAND2_X1 U9028 ( .A1(n13081), .A2(n13080), .ZN(n14744) );
  INV_X1 U9029 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6953) );
  XNOR2_X1 U9030 ( .A(n6769), .B(n8250), .ZN(n13894) );
  NAND2_X1 U9031 ( .A1(n8237), .A2(n7836), .ZN(n6769) );
  AND2_X1 U9032 ( .A1(n7688), .A2(n6626), .ZN(n7132) );
  XNOR2_X1 U9033 ( .A(n7713), .B(n7748), .ZN(n14748) );
  NAND2_X1 U9034 ( .A1(n7225), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7708) );
  AND2_X1 U9035 ( .A1(n7224), .A2(n7223), .ZN(n7222) );
  XNOR2_X1 U9036 ( .A(n8211), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14757) );
  INV_X1 U9037 ( .A(n8306), .ZN(n14756) );
  INV_X1 U9038 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10498) );
  NAND2_X1 U9039 ( .A1(n7591), .A2(n7826), .ZN(n8183) );
  NAND2_X1 U9040 ( .A1(n7826), .A2(n7824), .ZN(n8181) );
  INV_X1 U9041 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9835) );
  INV_X1 U9042 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n13776) );
  INV_X1 U9043 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9653) );
  INV_X1 U9044 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9617) );
  INV_X1 U9045 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9501) );
  INV_X1 U9046 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9448) );
  INV_X1 U9047 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9134) );
  INV_X1 U9048 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9087) );
  INV_X1 U9049 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9074) );
  INV_X1 U9050 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9063) );
  INV_X1 U9051 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9056) );
  INV_X1 U9052 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7902) );
  INV_X1 U9053 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9054) );
  NAND2_X1 U9054 ( .A1(n14794), .A2(n14795), .ZN(n14871) );
  NOR2_X1 U9055 ( .A1(n15548), .A2(n14800), .ZN(n15541) );
  XNOR2_X1 U9056 ( .A(n14786), .B(n7236), .ZN(n15542) );
  INV_X1 U9057 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7236) );
  XNOR2_X1 U9058 ( .A(n14804), .B(n7458), .ZN(n14875) );
  INV_X1 U9059 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7458) );
  XNOR2_X1 U9060 ( .A(n14811), .B(n7456), .ZN(n15545) );
  INV_X1 U9061 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7456) );
  NOR2_X1 U9062 ( .A1(n7455), .A2(n7451), .ZN(n7240) );
  AND2_X1 U9063 ( .A1(n14979), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7451) );
  NOR2_X1 U9064 ( .A1(n14983), .A2(n14984), .ZN(n14982) );
  AND2_X1 U9065 ( .A1(n14839), .A2(n14838), .ZN(n14986) );
  NAND2_X1 U9066 ( .A1(n7334), .A2(n6711), .ZN(n7328) );
  AOI21_X1 U9067 ( .B1(n6748), .B2(n15461), .A(n6746), .ZN(n7327) );
  NAND2_X1 U9068 ( .A1(n7008), .A2(n7005), .ZN(P3_U3487) );
  INV_X1 U9069 ( .A(n7006), .ZN(n7005) );
  NAND2_X1 U9070 ( .A1(n8957), .A2(n15540), .ZN(n7008) );
  OAI21_X1 U9071 ( .B1(n8956), .B2(n12556), .A(n7007), .ZN(n7006) );
  OAI21_X1 U9072 ( .B1(n7057), .B2(n15538), .A(n7056), .ZN(n11603) );
  NAND2_X1 U9073 ( .A1(n15538), .A2(n11602), .ZN(n7056) );
  OAI21_X1 U9074 ( .B1(n8957), .B2(n15521), .A(n6983), .ZN(n8958) );
  OR2_X1 U9075 ( .A1(n15519), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U9076 ( .A1(n7475), .A2(n10724), .ZN(n11193) );
  NAND2_X1 U9077 ( .A1(n10722), .A2(n10719), .ZN(n7475) );
  AND2_X1 U9078 ( .A1(n13165), .A2(n13177), .ZN(n6947) );
  OAI211_X1 U9079 ( .C1(n13487), .C2(n13465), .A(n7442), .B(n7440), .ZN(
        P2_U3236) );
  NAND2_X1 U9080 ( .A1(n7441), .A2(n13472), .ZN(n7440) );
  AOI21_X1 U9081 ( .B1(n13483), .B2(n13467), .A(n11541), .ZN(n7442) );
  INV_X1 U9082 ( .A(n13486), .ZN(n7441) );
  NAND2_X1 U9083 ( .A1(n7393), .A2(n7392), .ZN(P2_U3495) );
  NAND2_X1 U9084 ( .A1(n15429), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7392) );
  NAND2_X1 U9085 ( .A1(n13863), .A2(n15431), .ZN(n7393) );
  NAND2_X1 U9086 ( .A1(n6803), .A2(n6719), .ZN(P2_U3326) );
  INV_X1 U9087 ( .A(n6804), .ZN(n6803) );
  OAI22_X1 U9088 ( .A1(n13905), .A2(n9048), .B1(P2_U3088), .B2(n6805), .ZN(
        n6804) );
  INV_X1 U9089 ( .A(n6891), .ZN(n6890) );
  OAI21_X1 U9090 ( .B1(n14447), .B2(n14067), .A(n13918), .ZN(n6891) );
  NAND2_X1 U9091 ( .A1(n7211), .A2(n14052), .ZN(n7209) );
  INV_X1 U9092 ( .A(n6999), .ZN(n14437) );
  OAI21_X1 U9093 ( .B1(n14647), .B2(n14623), .A(n7264), .ZN(P1_U3266) );
  INV_X1 U9094 ( .A(n7265), .ZN(n7264) );
  OAI21_X1 U9095 ( .B1(n14646), .B2(n15106), .A(n7266), .ZN(n7265) );
  AOI21_X1 U9096 ( .B1(n14643), .B2(n15101), .A(n14451), .ZN(n7266) );
  XNOR2_X1 U9097 ( .A(n6838), .B(n6837), .ZN(n15543) );
  INV_X1 U9098 ( .A(n7247), .ZN(n14877) );
  INV_X1 U9099 ( .A(n7455), .ZN(n14881) );
  AND2_X1 U9100 ( .A1(n7452), .A2(n7455), .ZN(n14980) );
  OAI21_X1 U9101 ( .B1(n7455), .B2(n14979), .A(n7447), .ZN(n14978) );
  INV_X1 U9102 ( .A(n7244), .ZN(n14989) );
  OAI21_X1 U9103 ( .B1(n14893), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n7237), .ZN(
        n7444) );
  OR2_X1 U9104 ( .A1(n11881), .A2(n12349), .ZN(n6569) );
  AND2_X1 U9105 ( .A1(n9306), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6570) );
  AND2_X1 U9106 ( .A1(n6662), .A2(n12950), .ZN(n6571) );
  OR2_X1 U9107 ( .A1(n14524), .A2(n14668), .ZN(n6572) );
  NAND2_X1 U9108 ( .A1(n11351), .A2(n13444), .ZN(n6573) );
  AND2_X1 U9109 ( .A1(n7566), .A2(n7565), .ZN(n6574) );
  INV_X1 U9110 ( .A(n14335), .ZN(n7206) );
  OR2_X1 U9111 ( .A1(n8837), .A2(n10509), .ZN(n6575) );
  NAND2_X1 U9112 ( .A1(n14452), .A2(n7504), .ZN(n7506) );
  NAND2_X1 U9113 ( .A1(n7362), .A2(n7364), .ZN(n8552) );
  AND2_X1 U9114 ( .A1(n7168), .A2(n6602), .ZN(n6576) );
  AND2_X1 U9115 ( .A1(n6649), .A2(n6859), .ZN(n6577) );
  NAND2_X1 U9116 ( .A1(n8239), .A2(n8238), .ZN(n14652) );
  AND2_X1 U9117 ( .A1(n9455), .A2(n6622), .ZN(n6578) );
  INV_X1 U9118 ( .A(n15056), .ZN(n6874) );
  AND2_X1 U9119 ( .A1(n14272), .A2(n7495), .ZN(n6579) );
  NAND2_X1 U9120 ( .A1(n7785), .A2(SI_7_), .ZN(n6580) );
  OAI21_X1 U9121 ( .B1(n9783), .B2(P2_IR_REG_0__SCAN_IN), .A(n6993), .ZN(
        n12876) );
  AND2_X1 U9122 ( .A1(n9305), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6581) );
  AND2_X1 U9123 ( .A1(n13361), .A2(n13190), .ZN(n6582) );
  AND3_X1 U9124 ( .A1(n6580), .A2(n7780), .A3(n7784), .ZN(n6583) );
  AND3_X1 U9125 ( .A1(n14572), .A2(n7135), .A3(n7133), .ZN(n6584) );
  AND2_X1 U9126 ( .A1(n14676), .A2(n6812), .ZN(n6585) );
  INV_X1 U9127 ( .A(n12925), .ZN(n7684) );
  INV_X1 U9128 ( .A(n13039), .ZN(n7676) );
  AND2_X1 U9129 ( .A1(n7055), .A2(n6657), .ZN(n6586) );
  NAND2_X1 U9130 ( .A1(n10601), .A2(n6643), .ZN(n6587) );
  AND2_X1 U9131 ( .A1(n12082), .A2(n12101), .ZN(n12392) );
  INV_X1 U9132 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7706) );
  INV_X1 U9133 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8976) );
  INV_X1 U9134 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7842) );
  AND2_X1 U9135 ( .A1(n7433), .A2(n12807), .ZN(n6588) );
  OR2_X1 U9136 ( .A1(n13489), .A2(n6680), .ZN(n6589) );
  INV_X1 U9137 ( .A(n14098), .ZN(n14639) );
  AND2_X1 U9138 ( .A1(n7846), .A2(n7845), .ZN(n14098) );
  AND2_X1 U9139 ( .A1(n7683), .A2(n7684), .ZN(n6590) );
  INV_X1 U9140 ( .A(n14885), .ZN(n7632) );
  NAND2_X1 U9141 ( .A1(n8265), .A2(n8264), .ZN(n14253) );
  OR2_X1 U9142 ( .A1(n14219), .A2(n14218), .ZN(n6591) );
  AND2_X1 U9143 ( .A1(n11654), .A2(n11880), .ZN(n6592) );
  NOR2_X1 U9144 ( .A1(n15412), .A2(n12924), .ZN(n7230) );
  INV_X1 U9145 ( .A(n14238), .ZN(n7545) );
  AND2_X1 U9146 ( .A1(n7325), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6593) );
  XOR2_X1 U9147 ( .A(n11689), .B(n11795), .Z(n6594) );
  AND2_X1 U9148 ( .A1(n7829), .A2(n7579), .ZN(n6595) );
  AND4_X1 U9149 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n12381)
         );
  INV_X1 U9150 ( .A(n13409), .ZN(n7160) );
  AND2_X1 U9151 ( .A1(n6704), .A2(n6575), .ZN(n6596) );
  NAND2_X1 U9152 ( .A1(n7334), .A2(n6701), .ZN(n6597) );
  NAND2_X1 U9153 ( .A1(n7186), .A2(n6710), .ZN(n6598) );
  INV_X1 U9154 ( .A(n15465), .ZN(n7334) );
  XNOR2_X1 U9155 ( .A(n6841), .B(n9261), .ZN(n9264) );
  INV_X1 U9156 ( .A(n6567), .ZN(n8831) );
  INV_X1 U9157 ( .A(n8458), .ZN(n8543) );
  NAND2_X1 U9158 ( .A1(n11337), .A2(n12628), .ZN(n8458) );
  INV_X1 U9159 ( .A(n9866), .ZN(n11987) );
  NAND2_X2 U9160 ( .A1(n14743), .A2(n14746), .ZN(n8312) );
  AND2_X1 U9161 ( .A1(n12304), .A2(n7361), .ZN(n6599) );
  INV_X1 U9162 ( .A(n11164), .ZN(n7607) );
  OAI21_X1 U9163 ( .B1(n12676), .B2(n12675), .A(n12811), .ZN(n7466) );
  NAND2_X1 U9164 ( .A1(n7637), .A2(n13934), .ZN(n13932) );
  OR2_X1 U9165 ( .A1(n13311), .A2(n13303), .ZN(n6600) );
  AND3_X1 U9166 ( .A1(n8963), .A2(n8962), .A3(n9593), .ZN(n8973) );
  NAND3_X1 U9167 ( .A1(n8573), .A2(n8332), .A3(n7626), .ZN(n6601) );
  OR2_X1 U9168 ( .A1(n13520), .A2(n12809), .ZN(n6602) );
  OR2_X1 U9169 ( .A1(n14481), .A2(n14319), .ZN(n6603) );
  OR2_X1 U9170 ( .A1(n7769), .A2(n9067), .ZN(n6604) );
  OR2_X1 U9171 ( .A1(n9783), .A2(n6805), .ZN(n6605) );
  NAND2_X1 U9172 ( .A1(n12222), .A2(n12207), .ZN(n6606) );
  AND2_X1 U9173 ( .A1(n7432), .A2(n7428), .ZN(n6607) );
  XOR2_X1 U9174 ( .A(n14895), .B(n14894), .Z(n6608) );
  AND2_X1 U9175 ( .A1(n7682), .A2(n6845), .ZN(n6609) );
  AND2_X1 U9176 ( .A1(n7160), .A2(n11367), .ZN(n6610) );
  AND2_X1 U9177 ( .A1(n7178), .A2(n10598), .ZN(n6611) );
  AND2_X1 U9178 ( .A1(n12940), .A2(n12939), .ZN(n6612) );
  AND2_X1 U9179 ( .A1(n7034), .A2(n7036), .ZN(n6613) );
  OR2_X1 U9180 ( .A1(n8999), .A2(n14351), .ZN(n6614) );
  OR2_X1 U9181 ( .A1(n14862), .A2(n14861), .ZN(n6615) );
  INV_X1 U9182 ( .A(n6742), .ZN(n8894) );
  AND2_X1 U9183 ( .A1(n8375), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6616) );
  AND2_X1 U9184 ( .A1(n8168), .A2(n7402), .ZN(n6617) );
  AND2_X1 U9185 ( .A1(n9044), .A2(n9045), .ZN(n9049) );
  INV_X1 U9186 ( .A(n14281), .ZN(n6869) );
  AND3_X2 U9187 ( .A1(n8466), .A2(n8465), .A3(n8464), .ZN(n10290) );
  OR2_X1 U9188 ( .A1(n14644), .A2(n14317), .ZN(n6618) );
  XNOR2_X1 U9189 ( .A(n7522), .B(n7521), .ZN(n8306) );
  INV_X1 U9190 ( .A(n9697), .ZN(n7338) );
  AND2_X1 U9191 ( .A1(n12032), .A2(n7598), .ZN(n6619) );
  INV_X1 U9192 ( .A(n7609), .ZN(n7608) );
  NAND2_X1 U9193 ( .A1(n12058), .A2(n7610), .ZN(n7609) );
  INV_X1 U9194 ( .A(n14284), .ZN(n14935) );
  XNOR2_X1 U9195 ( .A(n14934), .B(n15058), .ZN(n14284) );
  INV_X1 U9196 ( .A(n11641), .ZN(n7377) );
  AND2_X1 U9197 ( .A1(n7476), .A2(n11192), .ZN(n6620) );
  INV_X1 U9198 ( .A(n14545), .ZN(n7256) );
  NAND2_X1 U9199 ( .A1(n7891), .A2(n7697), .ZN(n7894) );
  INV_X1 U9200 ( .A(n13303), .ZN(n7234) );
  AND2_X1 U9201 ( .A1(n8331), .A2(n7129), .ZN(n6621) );
  OR2_X1 U9202 ( .A1(n9783), .A2(n9456), .ZN(n6622) );
  INV_X1 U9203 ( .A(n12888), .ZN(n9473) );
  XOR2_X1 U9204 ( .A(n7770), .B(SI_2_), .Z(n6623) );
  AND2_X1 U9205 ( .A1(n15402), .A2(n12918), .ZN(n6624) );
  INV_X1 U9206 ( .A(n7362), .ZN(n8479) );
  OR2_X1 U9207 ( .A1(n8999), .A2(n14368), .ZN(n6625) );
  INV_X1 U9208 ( .A(n8860), .ZN(n7068) );
  AND2_X1 U9209 ( .A1(n7749), .A2(n7748), .ZN(n6626) );
  INV_X1 U9210 ( .A(n9582), .ZN(n6949) );
  NOR2_X1 U9211 ( .A1(n14132), .A2(n14131), .ZN(n6627) );
  NAND2_X2 U9212 ( .A1(n6768), .A2(n11476), .ZN(n13493) );
  INV_X1 U9213 ( .A(n13493), .ZN(n7235) );
  AND2_X1 U9214 ( .A1(n13951), .A2(n13949), .ZN(n6628) );
  AND2_X1 U9215 ( .A1(n14969), .A2(n7632), .ZN(n6629) );
  AND4_X1 U9216 ( .A1(n9261), .A2(n8964), .A3(n7481), .A4(n8970), .ZN(n6630)
         );
  NOR2_X1 U9217 ( .A1(n11087), .A2(n11090), .ZN(n6631) );
  INV_X1 U9218 ( .A(n12938), .ZN(n7681) );
  OR2_X1 U9219 ( .A1(n11235), .A2(n11215), .ZN(n6632) );
  NOR2_X1 U9220 ( .A1(n13083), .A2(n9782), .ZN(n6633) );
  INV_X1 U9221 ( .A(n7231), .ZN(n13273) );
  NOR3_X1 U9222 ( .A1(n13311), .A2(n13493), .A3(n7233), .ZN(n7231) );
  OR2_X1 U9223 ( .A1(n14533), .A2(n7397), .ZN(n6634) );
  NOR2_X1 U9224 ( .A1(n11432), .A2(n7170), .ZN(n7169) );
  INV_X1 U9225 ( .A(n14659), .ZN(n14481) );
  NAND2_X1 U9226 ( .A1(n7850), .A2(n7849), .ZN(n14659) );
  AND2_X1 U9227 ( .A1(n6594), .A2(n11688), .ZN(n6635) );
  INV_X1 U9228 ( .A(n14234), .ZN(n7516) );
  INV_X1 U9229 ( .A(n11623), .ZN(n7100) );
  OR2_X1 U9230 ( .A1(n12609), .A2(n11099), .ZN(n6636) );
  AND2_X1 U9231 ( .A1(n7712), .A2(n7706), .ZN(n6637) );
  INV_X1 U9232 ( .A(n12315), .ZN(n12318) );
  AND2_X1 U9233 ( .A1(n12119), .A2(n12120), .ZN(n12315) );
  AND2_X1 U9234 ( .A1(n7653), .A2(n7191), .ZN(n6638) );
  XNOR2_X1 U9235 ( .A(n9284), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9286) );
  NOR2_X1 U9236 ( .A1(n14151), .A2(n14150), .ZN(n6639) );
  OR2_X1 U9237 ( .A1(n14481), .A2(n14489), .ZN(n6640) );
  AND2_X1 U9238 ( .A1(n13005), .A2(n13004), .ZN(n6641) );
  AND2_X1 U9239 ( .A1(n7819), .A2(n6761), .ZN(n6642) );
  NAND2_X1 U9240 ( .A1(n13855), .A2(n12949), .ZN(n6643) );
  AND2_X1 U9241 ( .A1(n11277), .A2(n11275), .ZN(n6644) );
  AND2_X1 U9242 ( .A1(n11687), .A2(n11678), .ZN(n6645) );
  INV_X1 U9243 ( .A(n12059), .ZN(n7610) );
  AND2_X1 U9244 ( .A1(n9670), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U9245 ( .A1(n8225), .A2(n8224), .ZN(n14668) );
  INV_X1 U9246 ( .A(n7514), .ZN(n7513) );
  AND2_X1 U9247 ( .A1(n11569), .A2(n6618), .ZN(n6647) );
  INV_X1 U9248 ( .A(n7694), .ZN(n6924) );
  OR2_X1 U9249 ( .A1(n7693), .A2(n11092), .ZN(n6648) );
  INV_X1 U9250 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8412) );
  OR2_X1 U9251 ( .A1(n6662), .A2(n12950), .ZN(n6649) );
  NOR2_X1 U9252 ( .A1(n15089), .A2(n14330), .ZN(n6650) );
  NOR2_X1 U9253 ( .A1(n14714), .A2(n14323), .ZN(n6651) );
  INV_X1 U9254 ( .A(n7343), .ZN(n7342) );
  NOR2_X1 U9255 ( .A1(n8855), .A2(n12422), .ZN(n7343) );
  NOR2_X1 U9256 ( .A1(n12924), .A2(n10352), .ZN(n6652) );
  NOR2_X1 U9257 ( .A1(n13438), .A2(n12986), .ZN(n6653) );
  NOR2_X1 U9258 ( .A1(n14333), .A2(n15152), .ZN(n6654) );
  XOR2_X1 U9259 ( .A(n14900), .B(n14899), .Z(n6655) );
  INV_X1 U9260 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7481) );
  OR2_X1 U9261 ( .A1(n11905), .A2(n12360), .ZN(n12113) );
  INV_X1 U9262 ( .A(n12113), .ZN(n7612) );
  AND2_X1 U9263 ( .A1(n13493), .A2(n13185), .ZN(n6656) );
  OR2_X1 U9264 ( .A1(n15514), .A2(n11086), .ZN(n6657) );
  AND4_X1 U9265 ( .A1(n8331), .A2(n7079), .A3(n7129), .A4(n7128), .ZN(n6658)
         );
  OR2_X1 U9266 ( .A1(n12934), .A2(n12933), .ZN(n6659) );
  NAND2_X1 U9267 ( .A1(n7395), .A2(n13268), .ZN(n13488) );
  AND2_X1 U9268 ( .A1(n7791), .A2(SI_9_), .ZN(n6660) );
  NAND2_X1 U9269 ( .A1(n7630), .A2(n8412), .ZN(n6661) );
  AND2_X1 U9270 ( .A1(n12946), .A2(n12945), .ZN(n6662) );
  NOR2_X1 U9271 ( .A1(n13855), .A2(n13200), .ZN(n6663) );
  INV_X1 U9272 ( .A(n6922), .ZN(n6921) );
  OAI21_X1 U9273 ( .B1(n6924), .B2(n6603), .A(n8248), .ZN(n6922) );
  AND2_X1 U9274 ( .A1(n12666), .A2(n12665), .ZN(n6664) );
  NAND2_X1 U9275 ( .A1(n6951), .A2(n7897), .ZN(n14111) );
  INV_X1 U9276 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n13630) );
  NAND2_X1 U9277 ( .A1(n13100), .A2(n13099), .ZN(n6665) );
  INV_X1 U9278 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7752) );
  INV_X1 U9279 ( .A(n7220), .ZN(n7219) );
  NAND2_X1 U9280 ( .A1(n10695), .A2(n7221), .ZN(n7220) );
  AND2_X1 U9281 ( .A1(n7635), .A2(n6905), .ZN(n6666) );
  NAND2_X1 U9282 ( .A1(n8374), .A2(n8375), .ZN(n6667) );
  AND2_X1 U9283 ( .A1(n14760), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6668) );
  AND2_X1 U9284 ( .A1(n9063), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U9285 ( .A1(n12995), .A2(n12994), .ZN(n6670) );
  OR2_X1 U9286 ( .A1(n13582), .A2(n13199), .ZN(n6671) );
  INV_X1 U9287 ( .A(n7422), .ZN(n7421) );
  NAND2_X1 U9288 ( .A1(n13430), .A2(n7423), .ZN(n7422) );
  INV_X1 U9289 ( .A(n6851), .ZN(n6850) );
  NAND2_X1 U9290 ( .A1(n12977), .A2(n6852), .ZN(n6851) );
  INV_X1 U9291 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13881) );
  AND2_X1 U9292 ( .A1(n11774), .A2(n11772), .ZN(n13981) );
  INV_X1 U9293 ( .A(n13981), .ZN(n7646) );
  INV_X1 U9294 ( .A(n14285), .ZN(n11318) );
  INV_X1 U9295 ( .A(n7541), .ZN(n7540) );
  OAI21_X1 U9296 ( .B1(n7544), .B2(n14241), .A(n14240), .ZN(n7541) );
  OR2_X1 U9297 ( .A1(n14304), .A2(n14095), .ZN(n6672) );
  AND2_X1 U9298 ( .A1(n10858), .A2(n6631), .ZN(n6673) );
  AND2_X1 U9299 ( .A1(n13038), .A2(n13037), .ZN(n6674) );
  INV_X1 U9300 ( .A(n12926), .ZN(n7683) );
  INV_X1 U9301 ( .A(n7499), .ZN(n7498) );
  NOR2_X1 U9302 ( .A1(n15147), .A2(n14122), .ZN(n7499) );
  NAND2_X1 U9303 ( .A1(n8918), .A2(n8409), .ZN(n8892) );
  AND2_X1 U9304 ( .A1(n8409), .A2(n7076), .ZN(n6675) );
  INV_X1 U9305 ( .A(n12872), .ZN(n13164) );
  AND2_X1 U9306 ( .A1(n10346), .A2(n6561), .ZN(n12872) );
  INV_X1 U9307 ( .A(n14213), .ZN(n7530) );
  AND2_X1 U9308 ( .A1(n10876), .A2(n10877), .ZN(n6676) );
  INV_X1 U9309 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9498) );
  AND2_X1 U9310 ( .A1(n7037), .A2(n12678), .ZN(n6677) );
  AND2_X1 U9311 ( .A1(n12589), .A2(n12372), .ZN(n6678) );
  INV_X1 U9312 ( .A(n7397), .ZN(n7396) );
  NAND2_X1 U9313 ( .A1(n14520), .A2(n8210), .ZN(n7397) );
  AND2_X1 U9314 ( .A1(n13486), .A2(n13485), .ZN(n6679) );
  AND2_X1 U9315 ( .A1(n13490), .A2(n15421), .ZN(n6680) );
  NAND2_X1 U9316 ( .A1(n12605), .A2(n12478), .ZN(n6681) );
  OR2_X1 U9317 ( .A1(n14098), .A2(n14316), .ZN(n6682) );
  AND2_X1 U9318 ( .A1(n12044), .A2(n12049), .ZN(n11969) );
  INV_X1 U9319 ( .A(n11969), .ZN(n7346) );
  AND2_X1 U9320 ( .A1(n12392), .A2(n8710), .ZN(n6683) );
  AND2_X1 U9321 ( .A1(n8330), .A2(n7079), .ZN(n6684) );
  AND2_X1 U9322 ( .A1(n13097), .A2(n7665), .ZN(n6685) );
  NAND2_X1 U9323 ( .A1(n13914), .A2(n7216), .ZN(n6686) );
  INV_X1 U9324 ( .A(n14241), .ZN(n7548) );
  INV_X1 U9325 ( .A(n12921), .ZN(n6846) );
  AND2_X1 U9326 ( .A1(n7578), .A2(n7580), .ZN(n6687) );
  INV_X1 U9327 ( .A(n7942), .ZN(n6930) );
  NAND2_X1 U9328 ( .A1(n10189), .A2(n15152), .ZN(n7942) );
  INV_X1 U9329 ( .A(n11644), .ZN(n11881) );
  OR2_X1 U9330 ( .A1(n11642), .A2(n11643), .ZN(n11644) );
  NAND2_X1 U9331 ( .A1(n7552), .A2(n14222), .ZN(n6688) );
  INV_X1 U9332 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n6757) );
  INV_X1 U9333 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6992) );
  OR2_X1 U9334 ( .A1(n7687), .A2(n6641), .ZN(n6689) );
  INV_X1 U9335 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14766) );
  INV_X1 U9336 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U9337 ( .A1(n7777), .A2(SI_4_), .ZN(n6690) );
  INV_X1 U9338 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7061) );
  OAI21_X1 U9339 ( .B1(n13990), .B2(n14000), .A(n13999), .ZN(n7656) );
  INV_X1 U9340 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7521) );
  INV_X1 U9341 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7129) );
  INV_X1 U9342 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7079) );
  OAI211_X1 U9343 ( .C1(n8458), .C2(n12579), .A(n8764), .B(n8763), .ZN(n12320)
         );
  INV_X1 U9344 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7317) );
  INV_X1 U9345 ( .A(n13367), .ZN(n7433) );
  NOR2_X1 U9346 ( .A1(n11353), .A2(n11352), .ZN(n7391) );
  NAND4_X1 U9347 ( .A1(n7502), .A2(n7501), .A3(n7500), .A4(n7503), .ZN(n7958)
         );
  INV_X1 U9348 ( .A(n7958), .ZN(n7549) );
  AND2_X1 U9349 ( .A1(n7474), .A2(n7472), .ZN(n6691) );
  NAND2_X1 U9350 ( .A1(n6937), .A2(n6936), .ZN(n8133) );
  AND2_X1 U9351 ( .A1(n11856), .A2(n11649), .ZN(n11880) );
  INV_X1 U9352 ( .A(n14682), .ZN(n6812) );
  INV_X1 U9353 ( .A(n11856), .ZN(n7369) );
  AND2_X1 U9354 ( .A1(n13438), .A2(n13195), .ZN(n6692) );
  INV_X1 U9355 ( .A(n14288), .ZN(n11210) );
  NAND2_X1 U9356 ( .A1(n11679), .A2(n6645), .ZN(n13919) );
  INV_X1 U9357 ( .A(n13919), .ZN(n6901) );
  AND4_X1 U9358 ( .A1(n7764), .A2(n7763), .A3(n7762), .A4(n7761), .ZN(n14097)
         );
  INV_X1 U9359 ( .A(n7228), .ZN(n10917) );
  AND3_X1 U9360 ( .A1(n8610), .A2(n8609), .A3(n8608), .ZN(n11133) );
  INV_X1 U9361 ( .A(n11133), .ZN(n6739) );
  AND2_X1 U9362 ( .A1(n14016), .A2(n11753), .ZN(n13934) );
  INV_X1 U9363 ( .A(n13934), .ZN(n7641) );
  INV_X1 U9364 ( .A(n7634), .ZN(n11321) );
  NOR2_X1 U9365 ( .A1(n11202), .A2(n14944), .ZN(n7634) );
  OR2_X1 U9366 ( .A1(n14097), .A2(n14606), .ZN(n6693) );
  NOR2_X1 U9367 ( .A1(n10927), .A2(n10926), .ZN(n6694) );
  OR2_X1 U9368 ( .A1(n7816), .A2(n9512), .ZN(n6695) );
  AND4_X1 U9369 ( .A1(n8616), .A2(n8615), .A3(n8614), .A4(n8613), .ZN(n11144)
         );
  INV_X1 U9370 ( .A(n11144), .ZN(n12481) );
  INV_X1 U9371 ( .A(n14194), .ZN(n7140) );
  OR2_X1 U9372 ( .A1(n7140), .A2(n7141), .ZN(n6696) );
  AND2_X1 U9373 ( .A1(n12937), .A2(n12936), .ZN(n6697) );
  INV_X1 U9374 ( .A(SI_0_), .ZN(n7411) );
  NOR2_X1 U9375 ( .A1(n7580), .A2(SI_22_), .ZN(n6698) );
  INV_X1 U9376 ( .A(n12104), .ZN(n12593) );
  NAND2_X1 U9377 ( .A1(n8729), .A2(n8728), .ZN(n12104) );
  AND2_X1 U9378 ( .A1(n10172), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n6699) );
  INV_X1 U9379 ( .A(n12360), .ZN(n12171) );
  AND2_X1 U9380 ( .A1(n8756), .A2(n8755), .ZN(n12360) );
  INV_X1 U9381 ( .A(n11155), .ZN(n7580) );
  AND2_X1 U9382 ( .A1(n7096), .A2(n7094), .ZN(n6700) );
  INV_X1 U9383 ( .A(n12109), .ZN(n7620) );
  AND2_X1 U9384 ( .A1(n13156), .A2(n9264), .ZN(n15314) );
  NAND2_X2 U9385 ( .A1(n14431), .A2(n15091), .ZN(n15104) );
  NAND2_X1 U9386 ( .A1(n8126), .A2(n8125), .ZN(n14714) );
  INV_X1 U9387 ( .A(n14714), .ZN(n7633) );
  INV_X1 U9388 ( .A(n14216), .ZN(n6940) );
  NAND2_X1 U9389 ( .A1(n8977), .A2(n8976), .ZN(n8979) );
  INV_X2 U9390 ( .A(n15429), .ZN(n15431) );
  AND2_X1 U9391 ( .A1(n7330), .A2(n7329), .ZN(n6701) );
  XNOR2_X1 U9392 ( .A(n7708), .B(n7709), .ZN(n7730) );
  NAND2_X1 U9393 ( .A1(n10901), .A2(n10900), .ZN(n13577) );
  INV_X1 U9394 ( .A(n13577), .ZN(n7227) );
  NAND2_X1 U9395 ( .A1(n7599), .A2(n12030), .ZN(n10984) );
  NAND2_X1 U9396 ( .A1(n9931), .A2(n7942), .ZN(n9853) );
  AND2_X1 U9397 ( .A1(n8398), .A2(n7291), .ZN(n6702) );
  OR2_X1 U9398 ( .A1(n10805), .A2(n10604), .ZN(n6703) );
  INV_X1 U9399 ( .A(n8977), .ZN(n8981) );
  OR2_X1 U9400 ( .A1(n10217), .A2(n10216), .ZN(n6704) );
  AND2_X1 U9401 ( .A1(n10696), .A2(n7219), .ZN(n6705) );
  NAND2_X1 U9402 ( .A1(n10802), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6706) );
  INV_X1 U9403 ( .A(n8813), .ZN(n11948) );
  AND2_X1 U9404 ( .A1(n8249), .A2(SI_27_), .ZN(n6707) );
  INV_X1 U9405 ( .A(n7077), .ZN(n10849) );
  AND2_X1 U9406 ( .A1(n12271), .A2(n12270), .ZN(n6708) );
  AND2_X1 U9407 ( .A1(n7837), .A2(n11161), .ZN(n6709) );
  AND2_X1 U9408 ( .A1(n7185), .A2(n7181), .ZN(n6710) );
  OAI21_X1 U9409 ( .B1(n8398), .B2(n7291), .A(n13906), .ZN(n7288) );
  INV_X1 U9410 ( .A(n11091), .ZN(n7376) );
  INV_X1 U9411 ( .A(n13211), .ZN(n7410) );
  INV_X1 U9412 ( .A(n6910), .ZN(n14624) );
  INV_X1 U9413 ( .A(n14074), .ZN(n14052) );
  INV_X1 U9414 ( .A(n10066), .ZN(n7484) );
  NAND2_X1 U9415 ( .A1(n10131), .A2(n10130), .ZN(n15412) );
  AND2_X2 U9416 ( .A1(n10239), .A2(n8929), .ZN(n15540) );
  INV_X1 U9417 ( .A(n9886), .ZN(n9887) );
  NAND2_X1 U9418 ( .A1(n6733), .A2(n9895), .ZN(n9886) );
  AND2_X1 U9419 ( .A1(n7333), .A2(n12277), .ZN(n6711) );
  INV_X1 U9420 ( .A(n13210), .ZN(n7155) );
  NAND2_X1 U9421 ( .A1(n10379), .A2(n10378), .ZN(n15420) );
  INV_X1 U9422 ( .A(n15420), .ZN(n7229) );
  NAND2_X1 U9423 ( .A1(n8047), .A2(n8046), .ZN(n14885) );
  OR2_X1 U9424 ( .A1(n10192), .A2(n10191), .ZN(n6712) );
  AND2_X1 U9425 ( .A1(n11100), .A2(n11099), .ZN(n6713) );
  INV_X1 U9426 ( .A(n9767), .ZN(n6818) );
  NAND2_X1 U9427 ( .A1(n9393), .A2(n9392), .ZN(n14074) );
  INV_X1 U9428 ( .A(n9911), .ZN(n6938) );
  OR2_X1 U9429 ( .A1(n11058), .A2(n11035), .ZN(n6714) );
  AND2_X1 U9430 ( .A1(n9886), .A2(n7320), .ZN(n6715) );
  NAND2_X1 U9431 ( .A1(n14314), .A2(n14417), .ZN(n6716) );
  AND2_X1 U9432 ( .A1(n8990), .A2(n6894), .ZN(n6717) );
  INV_X1 U9433 ( .A(SI_22_), .ZN(n7579) );
  AND2_X1 U9434 ( .A1(n7331), .A2(n12264), .ZN(n6718) );
  INV_X1 U9435 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9584) );
  OR2_X1 U9436 ( .A1(n13908), .A2(n9292), .ZN(n6719) );
  INV_X1 U9437 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n6753) );
  INV_X1 U9438 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7503) );
  INV_X1 U9439 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n7072) );
  INV_X1 U9440 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6823) );
  INV_X1 U9441 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7450) );
  XNOR2_X1 U9442 ( .A(n7043), .B(n12678), .ZN(n12707) );
  INV_X1 U9443 ( .A(n12678), .ZN(n7038) );
  NAND3_X1 U9444 ( .A1(n6721), .A2(n6720), .A3(n11214), .ZN(n6970) );
  INV_X1 U9445 ( .A(n6725), .ZN(n10636) );
  NOR2_X1 U9446 ( .A1(n15445), .A2(n15446), .ZN(n15444) );
  NAND2_X1 U9447 ( .A1(n6729), .A2(n7338), .ZN(n6726) );
  INV_X1 U9448 ( .A(n6729), .ZN(n6728) );
  XNOR2_X1 U9449 ( .A(n12207), .B(n12222), .ZN(n12185) );
  INV_X1 U9450 ( .A(n6732), .ZN(n12208) );
  NAND3_X1 U9451 ( .A1(n7324), .A2(n9886), .A3(n6593), .ZN(n7322) );
  NAND3_X1 U9452 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        P3_IR_REG_1__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U9453 ( .A1(n11166), .A2(n8850), .ZN(n12477) );
  OR2_X2 U9454 ( .A1(n12333), .A2(n12334), .ZN(n12331) );
  INV_X1 U9455 ( .A(n11542), .ZN(n11971) );
  NAND3_X1 U9456 ( .A1(n6966), .A2(n11545), .A3(n6965), .ZN(n10227) );
  XNOR2_X2 U9457 ( .A(n12180), .B(n10083), .ZN(n11542) );
  AND3_X2 U9458 ( .A1(n7363), .A2(n8332), .A3(n7365), .ZN(n8408) );
  NAND4_X1 U9459 ( .A1(n7363), .A2(n8332), .A3(n7365), .A4(n7073), .ZN(n6742)
         );
  INV_X1 U9460 ( .A(n11220), .ZN(n11221) );
  XNOR2_X1 U9461 ( .A(n11220), .B(n11257), .ZN(n11254) );
  OAI21_X1 U9462 ( .B1(n12187), .B2(n6751), .A(n6750), .ZN(n12251) );
  INV_X1 U9463 ( .A(n12224), .ZN(n6751) );
  NAND2_X1 U9464 ( .A1(n6623), .A2(n6759), .ZN(n7772) );
  INV_X1 U9465 ( .A(n8151), .ZN(n6763) );
  NAND3_X1 U9466 ( .A1(n6766), .A2(n6764), .A3(n7786), .ZN(n7789) );
  AND2_X1 U9467 ( .A1(n7943), .A2(n7784), .ZN(n6767) );
  NAND2_X2 U9468 ( .A1(n7413), .A2(n7412), .ZN(n7586) );
  NAND3_X1 U9469 ( .A1(n7413), .A2(n7412), .A3(n9048), .ZN(n6775) );
  INV_X1 U9470 ( .A(n10383), .ZN(n6778) );
  NAND2_X1 U9471 ( .A1(n6781), .A2(n6779), .ZN(n6782) );
  NOR2_X1 U9472 ( .A1(n13130), .A2(n6780), .ZN(n6779) );
  NAND2_X1 U9473 ( .A1(n10351), .A2(n13132), .ZN(n10381) );
  NAND2_X1 U9474 ( .A1(n6782), .A2(n10350), .ZN(n10351) );
  AOI21_X2 U9475 ( .B1(n13280), .B2(n13147), .A(n6656), .ZN(n13263) );
  OAI22_X2 U9476 ( .A1(n13296), .A2(n11539), .B1(n11538), .B2(n7234), .ZN(
        n13280) );
  INV_X1 U9477 ( .A(n6783), .ZN(n7443) );
  OAI21_X2 U9478 ( .B1(n13445), .B2(n7422), .A(n7419), .ZN(n13424) );
  NAND3_X1 U9479 ( .A1(n13216), .A2(n6796), .A3(n13214), .ZN(n6792) );
  OAI21_X1 U9480 ( .B1(n13216), .B2(n13215), .A(n13214), .ZN(n13213) );
  INV_X1 U9481 ( .A(n9203), .ZN(n6796) );
  NAND2_X1 U9482 ( .A1(n7634), .A2(n7633), .ZN(n14613) );
  NAND3_X1 U9483 ( .A1(n14427), .A2(n6998), .A3(n6806), .ZN(n14637) );
  NAND2_X2 U9484 ( .A1(n15001), .A2(n11338), .ZN(n8999) );
  NAND3_X1 U9485 ( .A1(n6824), .A2(n6823), .A3(n6827), .ZN(n6822) );
  NAND2_X1 U9486 ( .A1(n6827), .A2(n6824), .ZN(n14785) );
  OR2_X1 U9487 ( .A1(n14764), .A2(n14765), .ZN(n6829) );
  NAND2_X1 U9488 ( .A1(n6826), .A2(n14766), .ZN(n6825) );
  INV_X1 U9489 ( .A(n14765), .ZN(n6826) );
  OAI21_X1 U9490 ( .B1(n14764), .B2(n14765), .A(P3_ADDR_REG_4__SCAN_IN), .ZN(
        n6827) );
  NOR2_X2 U9491 ( .A1(n6830), .A2(n14878), .ZN(n14821) );
  NAND3_X1 U9492 ( .A1(n6832), .A2(n6972), .A3(n6831), .ZN(n6834) );
  INV_X1 U9493 ( .A(n6834), .ZN(n14992) );
  INV_X1 U9494 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6833) );
  XNOR2_X1 U9495 ( .A(n14803), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U9496 ( .A1(n14801), .A2(n14802), .ZN(n6838) );
  OAI21_X1 U9497 ( .B1(n12965), .B2(n6851), .A(n6849), .ZN(n13001) );
  OAI21_X1 U9498 ( .B1(n13001), .B2(n13000), .A(n12999), .ZN(n13003) );
  OAI21_X1 U9499 ( .B1(n13053), .B2(n13052), .A(n6665), .ZN(n6855) );
  AOI21_X1 U9500 ( .B1(n13053), .B2(n13052), .A(n13051), .ZN(n6856) );
  NAND3_X1 U9501 ( .A1(n6944), .A2(n6941), .A3(n6861), .ZN(n6864) );
  OAI22_X2 U9502 ( .A1(n13011), .A2(n6866), .B1(n13009), .B2(n13010), .ZN(
        n13016) );
  NAND2_X1 U9503 ( .A1(n8284), .A2(n8283), .ZN(n15057) );
  INV_X1 U9504 ( .A(n15057), .ZN(n6867) );
  NAND2_X1 U9505 ( .A1(n6867), .A2(n7490), .ZN(n6871) );
  NAND2_X1 U9506 ( .A1(n6872), .A2(n7490), .ZN(n10757) );
  NAND2_X1 U9507 ( .A1(n14505), .A2(n7512), .ZN(n6876) );
  NAND2_X1 U9508 ( .A1(n14076), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7888) );
  NAND2_X1 U9509 ( .A1(n6892), .A2(n6890), .ZN(P1_U3214) );
  NAND2_X1 U9510 ( .A1(n6893), .A2(n14052), .ZN(n6892) );
  XNOR2_X1 U9511 ( .A(n13913), .B(n13914), .ZN(n6893) );
  NAND3_X1 U9512 ( .A1(n8990), .A2(n6894), .A3(n9605), .ZN(n9604) );
  INV_X2 U9513 ( .A(n11794), .ZN(n11783) );
  NAND2_X1 U9514 ( .A1(n11744), .A2(n14031), .ZN(n13933) );
  OAI21_X2 U9515 ( .B1(n11744), .B2(n6907), .A(n6666), .ZN(n13980) );
  NAND2_X1 U9516 ( .A1(n7652), .A2(n7648), .ZN(n13940) );
  NAND2_X2 U9517 ( .A1(n7756), .A2(n6909), .ZN(n8255) );
  INV_X1 U9518 ( .A(n14743), .ZN(n6909) );
  AND4_X2 U9519 ( .A1(n7872), .A2(n7871), .A3(n6957), .A4(n7873), .ZN(n6910)
         );
  NAND2_X1 U9520 ( .A1(n9923), .A2(n6910), .ZN(n8276) );
  OAI22_X1 U9521 ( .A1(n9923), .A2(n11794), .B1(n6910), .B2(n11798), .ZN(n9601) );
  OAI22_X1 U9522 ( .A1(n11797), .A2(n6910), .B1(n9923), .B2(n11798), .ZN(n9602) );
  XNOR2_X1 U9523 ( .A(n9628), .B(n6910), .ZN(n9623) );
  OAI21_X2 U9524 ( .B1(n6916), .B2(n6915), .A(n6912), .ZN(n14508) );
  AND2_X1 U9525 ( .A1(n14644), .A2(n8302), .ZN(n6923) );
  INV_X1 U9526 ( .A(n14268), .ZN(n9720) );
  NAND2_X1 U9527 ( .A1(n7886), .A2(n14106), .ZN(n9726) );
  NAND2_X1 U9528 ( .A1(n9682), .A2(n14269), .ZN(n6926) );
  NAND3_X1 U9529 ( .A1(n7886), .A2(n14268), .A3(n14106), .ZN(n6925) );
  NAND2_X1 U9530 ( .A1(n9929), .A2(n7942), .ZN(n6929) );
  NAND3_X1 U9531 ( .A1(n6929), .A2(n6928), .A3(n14275), .ZN(n9854) );
  OR2_X2 U9532 ( .A1(n6935), .A2(n11211), .ZN(n6934) );
  NAND2_X1 U9533 ( .A1(n9854), .A2(n7955), .ZN(n10089) );
  NAND2_X1 U9534 ( .A1(n8193), .A2(n14565), .ZN(n14552) );
  NAND2_X1 U9535 ( .A1(n7001), .A2(n6874), .ZN(n15052) );
  NAND2_X1 U9536 ( .A1(n10759), .A2(n6869), .ZN(n10758) );
  XNOR2_X1 U9537 ( .A(n14336), .B(n14111), .ZN(n14268) );
  NAND3_X1 U9538 ( .A1(n7179), .A2(n8975), .A3(n8974), .ZN(n9283) );
  NAND2_X1 U9539 ( .A1(n7016), .A2(n13409), .ZN(n13422) );
  OAI21_X2 U9540 ( .B1(n13307), .B2(n11536), .A(n11537), .ZN(n13296) );
  NAND2_X1 U9541 ( .A1(n14552), .A2(n8194), .ZN(n14533) );
  INV_X1 U9542 ( .A(n8975), .ZN(n9483) );
  NAND2_X1 U9543 ( .A1(n7818), .A2(n7819), .ZN(n8151) );
  NAND2_X1 U9544 ( .A1(n7581), .A2(n7578), .ZN(n11156) );
  NAND2_X1 U9545 ( .A1(n12416), .A2(n12415), .ZN(n12414) );
  NAND2_X1 U9546 ( .A1(n11341), .A2(n12135), .ZN(n11582) );
  AOI21_X2 U9547 ( .B1(n12330), .B2(n12334), .A(n12121), .ZN(n12316) );
  OAI21_X1 U9548 ( .B1(n10769), .B2(n8847), .A(n12040), .ZN(n11021) );
  NAND3_X1 U9549 ( .A1(n7059), .A2(n7058), .A3(n7060), .ZN(n7057) );
  NAND2_X1 U9550 ( .A1(n10806), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n10930) );
  XNOR2_X1 U9551 ( .A(n9893), .B(n9895), .ZN(n9896) );
  INV_X1 U9552 ( .A(n12897), .ZN(n6943) );
  NAND2_X1 U9553 ( .A1(n6959), .A2(n6958), .ZN(n6944) );
  NAND2_X1 U9554 ( .A1(n13181), .A2(n6945), .ZN(P2_U3328) );
  AOI21_X1 U9555 ( .B1(n13166), .B2(n6947), .A(n6946), .ZN(n6945) );
  NAND2_X1 U9556 ( .A1(n10622), .A2(n10623), .ZN(n10624) );
  AOI21_X1 U9557 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n9821), .A(n9820), .ZN(
        n9893) );
  NAND2_X2 U9558 ( .A1(n14743), .A2(n7756), .ZN(n14081) );
  NAND2_X1 U9559 ( .A1(n15052), .A2(n8017), .ZN(n14927) );
  NOR2_X1 U9560 ( .A1(n13962), .A2(n9606), .ZN(n9609) );
  NAND3_X1 U9561 ( .A1(n7549), .A2(n7705), .A3(n7704), .ZN(n7723) );
  NAND2_X1 U9562 ( .A1(n7418), .A2(n11535), .ZN(n13307) );
  MUX2_X2 U9563 ( .A(n12053), .B(n12052), .S(n12129), .Z(n12067) );
  MUX2_X2 U9564 ( .A(n12126), .B(n12125), .S(n12129), .Z(n12131) );
  NOR3_X2 U9565 ( .A1(n12048), .A2(n12046), .A3(n12045), .ZN(n12047) );
  AOI211_X2 U9566 ( .C1(n12143), .C2(n12142), .A(n12141), .B(n12140), .ZN(
        n12149) );
  INV_X1 U9567 ( .A(n7057), .ZN(n11604) );
  AOI211_X2 U9568 ( .C1(n12112), .C2(n12111), .A(n12110), .B(n12345), .ZN(
        n12116) );
  NAND3_X1 U9569 ( .A1(n9775), .A2(n9776), .A3(n9777), .ZN(n6956) );
  NAND2_X1 U9570 ( .A1(n9956), .A2(n9955), .ZN(n10417) );
  NAND2_X1 U9571 ( .A1(n7414), .A2(n9983), .ZN(n10446) );
  NAND2_X1 U9572 ( .A1(n13321), .A2(n13320), .ZN(n7418) );
  OAI21_X1 U9573 ( .B1(n13048), .B2(n13047), .A(n7690), .ZN(n13053) );
  OR2_X1 U9574 ( .A1(n13018), .A2(n13017), .ZN(n13023) );
  NAND2_X1 U9575 ( .A1(n12897), .A2(n12896), .ZN(n6959) );
  NAND3_X1 U9576 ( .A1(n9847), .A2(n12961), .A3(n6961), .ZN(n6960) );
  NAND2_X1 U9577 ( .A1(n7677), .A2(n7680), .ZN(n12944) );
  NAND2_X1 U9578 ( .A1(n6969), .A2(n6968), .ZN(n12892) );
  INV_X1 U9579 ( .A(n12889), .ZN(n7011) );
  AOI21_X1 U9580 ( .B1(n7570), .B2(n7573), .A(n7807), .ZN(n7569) );
  AND2_X1 U9581 ( .A1(n14255), .A2(n7538), .ZN(n7537) );
  NAND2_X1 U9582 ( .A1(n7815), .A2(n7583), .ZN(n7582) );
  NAND2_X1 U9583 ( .A1(n6962), .A2(n14312), .ZN(P1_U3242) );
  OAI211_X1 U9584 ( .C1(n14267), .C2(n6672), .A(n6964), .B(n6963), .ZN(n6962)
         );
  INV_X1 U9585 ( .A(n14313), .ZN(n6963) );
  NAND2_X1 U9586 ( .A1(n14267), .A2(n14303), .ZN(n6964) );
  NAND2_X1 U9587 ( .A1(n7861), .A2(n7833), .ZN(n7848) );
  NAND2_X1 U9588 ( .A1(n7592), .A2(n7826), .ZN(n8196) );
  NAND2_X1 U9589 ( .A1(n7776), .A2(n7004), .ZN(n7019) );
  NAND2_X1 U9590 ( .A1(n10262), .A2(n10263), .ZN(n10622) );
  NAND2_X1 U9591 ( .A1(n11224), .A2(n11241), .ZN(n12186) );
  NAND2_X1 U9592 ( .A1(n12251), .A2(n12250), .ZN(n12253) );
  NOR2_X1 U9593 ( .A1(n9585), .A2(n9586), .ZN(n9668) );
  OR2_X1 U9594 ( .A1(n10743), .A2(n10744), .ZN(n10742) );
  NAND2_X1 U9595 ( .A1(n12451), .A2(n12450), .ZN(n12449) );
  OAI21_X1 U9596 ( .B1(n10519), .B2(n8843), .A(n8842), .ZN(n8845) );
  INV_X1 U9597 ( .A(n10224), .ZN(n6966) );
  NAND2_X1 U9598 ( .A1(n11027), .A2(n11026), .ZN(n11025) );
  AND2_X1 U9599 ( .A1(n10178), .A2(n10254), .ZN(n7337) );
  NOR2_X1 U9600 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  NAND2_X1 U9601 ( .A1(n12433), .A2(n12432), .ZN(n12431) );
  NAND2_X1 U9602 ( .A1(n7344), .A2(n7345), .ZN(n7055) );
  NAND2_X1 U9603 ( .A1(n6971), .A2(n14995), .ZN(n14862) );
  NAND2_X1 U9604 ( .A1(n14996), .A2(n14997), .ZN(n14995) );
  OAI21_X1 U9605 ( .B1(n14996), .B2(n14997), .A(P2_ADDR_REG_16__SCAN_IN), .ZN(
        n6971) );
  NOR2_X1 U9606 ( .A1(n14784), .A2(n14783), .ZN(n14778) );
  NAND2_X1 U9607 ( .A1(n12449), .A2(n8852), .ZN(n12433) );
  NAND2_X1 U9608 ( .A1(n8840), .A2(n8839), .ZN(n10519) );
  NAND2_X1 U9609 ( .A1(n6973), .A2(n11453), .ZN(n13309) );
  NAND2_X1 U9610 ( .A1(n7162), .A2(n7161), .ZN(n6973) );
  NAND2_X1 U9611 ( .A1(n6687), .A2(n7581), .ZN(n11158) );
  INV_X1 U9612 ( .A(n7169), .ZN(n7168) );
  OAI21_X1 U9613 ( .B1(n13487), .B2(n15405), .A(n6679), .ZN(n13862) );
  NAND2_X1 U9614 ( .A1(n8040), .A2(n8039), .ZN(n8042) );
  NAND2_X1 U9615 ( .A1(n12254), .A2(n12255), .ZN(n12266) );
  NAND2_X1 U9616 ( .A1(n12885), .A2(n12884), .ZN(n12891) );
  NAND3_X1 U9617 ( .A1(n8975), .A2(n8974), .A3(n7661), .ZN(n9212) );
  NAND2_X1 U9618 ( .A1(n7010), .A2(n12892), .ZN(n12897) );
  OR2_X1 U9619 ( .A1(n12909), .A2(n12908), .ZN(n12914) );
  INV_X1 U9620 ( .A(n12882), .ZN(n6977) );
  INV_X1 U9621 ( .A(n8966), .ZN(n9208) );
  INV_X1 U9622 ( .A(n6976), .ZN(n12883) );
  NAND2_X1 U9623 ( .A1(n6975), .A2(n12881), .ZN(n12885) );
  NAND2_X1 U9624 ( .A1(n6977), .A2(n6976), .ZN(n6975) );
  AOI21_X1 U9625 ( .B1(n12955), .B2(n12954), .A(n12953), .ZN(n12957) );
  AOI21_X1 U9626 ( .B1(n12907), .B2(n12906), .A(n12905), .ZN(n12909) );
  NAND2_X1 U9627 ( .A1(n12891), .A2(n12890), .ZN(n7012) );
  OAI22_X1 U9628 ( .A1(n14242), .A2(n9292), .B1(n8999), .B2(n14342), .ZN(n6980) );
  NOR2_X2 U9629 ( .A1(n6572), .A2(n14664), .ZN(n14496) );
  INV_X1 U9630 ( .A(n7585), .ZN(n7817) );
  NAND2_X1 U9631 ( .A1(n14641), .A2(n6981), .ZN(n14721) );
  OAI21_X1 U9632 ( .B1(n14642), .B2(n14964), .A(n14640), .ZN(n6982) );
  AOI21_X1 U9633 ( .B1(n7512), .B2(n14509), .A(n8301), .ZN(n7511) );
  INV_X1 U9634 ( .A(n7511), .ZN(n7510) );
  NAND2_X1 U9635 ( .A1(n14760), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n14759) );
  AOI21_X1 U9636 ( .B1(n14872), .B2(n14796), .A(n14869), .ZN(n14798) );
  AND2_X1 U9637 ( .A1(n14799), .A2(n14798), .ZN(n15547) );
  OAI21_X2 U9638 ( .B1(n12331), .B2(n12315), .A(n7067), .ZN(n12305) );
  NAND2_X1 U9639 ( .A1(n10758), .A2(n8057), .ZN(n11027) );
  NAND2_X1 U9640 ( .A1(n8275), .A2(n15139), .ZN(n14427) );
  NAND3_X1 U9641 ( .A1(n12935), .A2(n6659), .A3(n7678), .ZN(n7677) );
  AOI21_X1 U9642 ( .B1(n13023), .B2(n7671), .A(n7669), .ZN(n7668) );
  NAND2_X1 U9643 ( .A1(n11006), .A2(n13141), .ZN(n11522) );
  NAND2_X1 U9644 ( .A1(n10898), .A2(n10897), .ZN(n11005) );
  NAND2_X1 U9645 ( .A1(n7323), .A2(n7322), .ZN(n10177) );
  AOI21_X1 U9646 ( .B1(n10266), .B2(P3_REG2_REG_7__SCAN_IN), .A(n10268), .ZN(
        n10271) );
  NAND2_X1 U9647 ( .A1(n7885), .A2(n7417), .ZN(n7876) );
  NAND2_X1 U9648 ( .A1(n9970), .A2(n9969), .ZN(n10403) );
  NAND2_X1 U9649 ( .A1(n7435), .A2(n7434), .ZN(n10898) );
  NAND2_X1 U9650 ( .A1(n14930), .A2(n8038), .ZN(n10759) );
  NAND3_X2 U9651 ( .A1(n9295), .A2(n9294), .A3(n6605), .ZN(n13470) );
  NAND2_X1 U9652 ( .A1(n7562), .A2(n7563), .ZN(n8040) );
  INV_X1 U9653 ( .A(n15049), .ZN(n7001) );
  NAND2_X1 U9654 ( .A1(n7003), .A2(n7002), .ZN(n8273) );
  NAND2_X1 U9655 ( .A1(n11561), .A2(n6682), .ZN(n7003) );
  INV_X4 U9656 ( .A(n7586), .ZN(n13064) );
  MUX2_X1 U9657 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7586), .Z(n7777) );
  INV_X1 U9658 ( .A(n14272), .ZN(n7941) );
  XNOR2_X2 U9659 ( .A(n8413), .B(n8412), .ZN(n11081) );
  NAND2_X1 U9660 ( .A1(n12460), .A2(n8851), .ZN(n12451) );
  XNOR2_X1 U9661 ( .A(n10928), .B(n10936), .ZN(n10806) );
  NAND2_X1 U9662 ( .A1(n7009), .A2(n7675), .ZN(n13046) );
  NAND3_X1 U9663 ( .A1(n13034), .A2(n13035), .A3(n7673), .ZN(n7009) );
  NAND2_X1 U9664 ( .A1(n7012), .A2(n7011), .ZN(n7010) );
  MUX2_X1 U9665 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n7586), .Z(n7770) );
  NOR2_X1 U9666 ( .A1(n14797), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n14764) );
  NAND2_X1 U9667 ( .A1(n7446), .A2(n7454), .ZN(n7239) );
  XNOR2_X1 U9668 ( .A(n7444), .B(n6655), .ZN(SUB_1596_U4) );
  NAND2_X1 U9669 ( .A1(n7013), .A2(n12263), .ZN(P3_U3200) );
  OAI21_X1 U9670 ( .B1(n12265), .B2(n7014), .A(n7334), .ZN(n7013) );
  NOR2_X1 U9671 ( .A1(n10268), .A2(n7337), .ZN(n10266) );
  NAND2_X1 U9672 ( .A1(n7132), .A2(n8139), .ZN(n7131) );
  NOR2_X2 U9673 ( .A1(n13965), .A2(n15141), .ZN(n9722) );
  NAND2_X1 U9674 ( .A1(n10284), .A2(n10127), .ZN(n10132) );
  NAND2_X1 U9675 ( .A1(n7017), .A2(n12631), .ZN(n12635) );
  AOI21_X1 U9676 ( .B1(n12833), .B2(n7018), .A(n12854), .ZN(n12835) );
  NAND2_X1 U9677 ( .A1(n10117), .A2(n10118), .ZN(n7018) );
  NAND3_X1 U9678 ( .A1(n7905), .A2(n7776), .A3(n7022), .ZN(n7021) );
  NAND3_X1 U9679 ( .A1(n7021), .A2(n6690), .A3(n7019), .ZN(n7925) );
  OAI211_X1 U9680 ( .C1(n7464), .C2(n7031), .A(n7026), .B(n7024), .ZN(n12751)
         );
  NAND2_X1 U9681 ( .A1(n7466), .A2(n7465), .ZN(n7033) );
  INV_X1 U9682 ( .A(n7043), .ZN(n7035) );
  AND2_X1 U9683 ( .A1(n7039), .A2(n7042), .ZN(n12778) );
  NAND2_X1 U9684 ( .A1(n7472), .A2(n7045), .ZN(n7044) );
  INV_X1 U9685 ( .A(n7048), .ZN(n7045) );
  OAI21_X2 U9686 ( .B1(n10671), .B2(n7047), .A(n7046), .ZN(n12700) );
  MUX2_X1 U9687 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7586), .Z(n7774) );
  NAND2_X1 U9688 ( .A1(n11600), .A2(n12474), .ZN(n7060) );
  NAND2_X1 U9689 ( .A1(n7060), .A2(n7059), .ZN(n11607) );
  AOI21_X1 U9690 ( .B1(n6553), .B2(n10988), .A(n11599), .ZN(n7059) );
  AND2_X1 U9691 ( .A1(n7365), .A2(n7362), .ZN(n8573) );
  AND2_X2 U9692 ( .A1(n8461), .A2(n6757), .ZN(n7362) );
  NAND3_X1 U9693 ( .A1(n7370), .A2(n10557), .A3(n7078), .ZN(n7077) );
  NAND2_X1 U9694 ( .A1(n8325), .A2(n6684), .ZN(n8686) );
  NAND2_X1 U9695 ( .A1(n8325), .A2(n8330), .ZN(n7080) );
  NAND2_X1 U9696 ( .A1(n11834), .A2(n11644), .ZN(n7083) );
  NAND3_X1 U9697 ( .A1(n6569), .A2(n7083), .A3(n11880), .ZN(n11879) );
  NAND3_X1 U9698 ( .A1(n6569), .A2(n7083), .A3(n6592), .ZN(n7082) );
  NAND2_X1 U9699 ( .A1(n11807), .A2(n11996), .ZN(n7086) );
  NAND2_X1 U9700 ( .A1(n9866), .A2(n11655), .ZN(n7087) );
  INV_X1 U9701 ( .A(n7101), .ZN(n11890) );
  NAND2_X1 U9702 ( .A1(n8329), .A2(n7121), .ZN(n7117) );
  NAND3_X1 U9703 ( .A1(n7120), .A2(n7119), .A3(n7124), .ZN(n12268) );
  OAI21_X1 U9704 ( .B1(n14197), .B2(n7136), .A(n6584), .ZN(n14205) );
  NAND2_X1 U9705 ( .A1(n7137), .A2(n6696), .ZN(n7136) );
  NAND2_X1 U9706 ( .A1(n14252), .A2(n14117), .ZN(n14118) );
  NAND2_X1 U9707 ( .A1(n14151), .A2(n14150), .ZN(n14149) );
  NAND3_X1 U9708 ( .A1(n7148), .A2(n6591), .A3(n6688), .ZN(n7147) );
  NAND2_X1 U9709 ( .A1(n7149), .A2(n7554), .ZN(n7553) );
  NAND2_X1 U9710 ( .A1(n7150), .A2(n14130), .ZN(n7149) );
  NAND2_X1 U9711 ( .A1(n14132), .A2(n14131), .ZN(n7150) );
  OAI22_X1 U9712 ( .A1(n14157), .A2(n7152), .B1(n14158), .B2(n7151), .ZN(
        n14163) );
  NAND2_X1 U9713 ( .A1(n14163), .A2(n14164), .ZN(n14161) );
  INV_X1 U9714 ( .A(n14156), .ZN(n7151) );
  NOR2_X1 U9715 ( .A1(n14159), .A2(n14156), .ZN(n7152) );
  NAND2_X1 U9716 ( .A1(n10370), .A2(n7154), .ZN(n10475) );
  NAND2_X1 U9717 ( .A1(n10472), .A2(n13210), .ZN(n7154) );
  NAND2_X1 U9718 ( .A1(n7155), .A2(n15370), .ZN(n10370) );
  NOR2_X1 U9719 ( .A1(n6570), .A2(n6581), .ZN(n7156) );
  NAND2_X1 U9720 ( .A1(n13364), .A2(n7164), .ZN(n7161) );
  INV_X1 U9721 ( .A(n11416), .ZN(n7173) );
  NAND2_X1 U9722 ( .A1(n10404), .A2(n7379), .ZN(n7175) );
  OAI21_X1 U9723 ( .B1(n10599), .B2(n6587), .A(n7176), .ZN(n10904) );
  INV_X1 U9724 ( .A(n9283), .ZN(n9281) );
  OAI21_X2 U9725 ( .B1(n7182), .B2(n7180), .A(n10304), .ZN(n10310) );
  NOR2_X1 U9726 ( .A1(n7187), .A2(n7184), .ZN(n7183) );
  NAND3_X1 U9727 ( .A1(n7194), .A2(n7193), .A3(n7195), .ZN(n14002) );
  NAND2_X1 U9728 ( .A1(n7204), .A2(n7197), .ZN(n7200) );
  NAND2_X1 U9729 ( .A1(n7198), .A2(n11765), .ZN(n7197) );
  INV_X1 U9730 ( .A(n10040), .ZN(n7199) );
  XNOR2_X1 U9731 ( .A(n10039), .B(n7199), .ZN(n13941) );
  NAND3_X1 U9732 ( .A1(n7201), .A2(n7200), .A3(n7203), .ZN(n10039) );
  NOR2_X1 U9733 ( .A1(n10307), .A2(n11795), .ZN(n7202) );
  NAND3_X1 U9734 ( .A1(n10307), .A2(n14335), .A3(n11795), .ZN(n7203) );
  NAND2_X1 U9735 ( .A1(n13913), .A2(n7208), .ZN(n7207) );
  OAI211_X1 U9736 ( .C1(n13913), .C2(n7209), .A(n7207), .B(n11806), .ZN(
        P1_U3220) );
  OAI21_X1 U9737 ( .B1(n13914), .B2(n7215), .A(n7214), .ZN(n7213) );
  INV_X1 U9738 ( .A(n11801), .ZN(n7216) );
  NAND2_X1 U9739 ( .A1(n7707), .A2(n7222), .ZN(n7225) );
  NAND2_X1 U9740 ( .A1(n7226), .A2(n9473), .ZN(n10471) );
  NAND2_X1 U9741 ( .A1(n9459), .A2(n12876), .ZN(n9471) );
  NAND2_X1 U9742 ( .A1(n8977), .A2(n7662), .ZN(n9211) );
  NAND2_X1 U9743 ( .A1(n10651), .A2(n10684), .ZN(n10650) );
  NOR2_X2 U9744 ( .A1(n13355), .A2(n13520), .ZN(n13337) );
  NOR2_X2 U9745 ( .A1(n13381), .A2(n13367), .ZN(n13370) );
  NAND2_X1 U9746 ( .A1(n7238), .A2(n6608), .ZN(n7237) );
  INV_X1 U9747 ( .A(n14789), .ZN(n7242) );
  OR3_X2 U9748 ( .A1(n7245), .A2(n14987), .A3(n14845), .ZN(n7244) );
  NAND2_X1 U9749 ( .A1(n7973), .A2(n7263), .ZN(n7262) );
  NAND2_X1 U9750 ( .A1(n11819), .A2(n11666), .ZN(n8863) );
  OAI21_X1 U9751 ( .B1(n8775), .B2(n7277), .A(n7274), .ZN(n8806) );
  INV_X1 U9752 ( .A(n7271), .ZN(n8808) );
  NAND2_X1 U9753 ( .A1(n7278), .A2(n7279), .ZN(n8591) );
  NOR2_X1 U9754 ( .A1(n7286), .A2(n7288), .ZN(n7285) );
  NAND2_X1 U9755 ( .A1(n8399), .A2(n8398), .ZN(n8400) );
  INV_X1 U9756 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7291) );
  NAND2_X1 U9757 ( .A1(n8738), .A2(n7295), .ZN(n7292) );
  NAND2_X1 U9758 ( .A1(n7292), .A2(n7293), .ZN(n8758) );
  NAND2_X1 U9759 ( .A1(n8697), .A2(n7301), .ZN(n7298) );
  NAND2_X1 U9760 ( .A1(n7298), .A2(n7299), .ZN(n8725) );
  OAI21_X1 U9761 ( .B1(n8492), .B2(n8351), .A(n8352), .ZN(n8505) );
  OAI211_X1 U9762 ( .C1(n12235), .C2(n7328), .A(n7327), .B(n7326), .ZN(
        P3_U3201) );
  NAND3_X1 U9763 ( .A1(n12235), .A2(n6718), .A3(n7334), .ZN(n7326) );
  NOR2_X1 U9764 ( .A1(n12235), .A2(n12234), .ZN(n12265) );
  NAND2_X1 U9765 ( .A1(n12277), .A2(n12264), .ZN(n7329) );
  INV_X1 U9766 ( .A(n12277), .ZN(n7331) );
  NOR2_X1 U9767 ( .A1(n12032), .A2(n7350), .ZN(n7349) );
  NAND2_X1 U9768 ( .A1(n11345), .A2(n12474), .ZN(n7357) );
  NAND2_X1 U9769 ( .A1(n7357), .A2(n7354), .ZN(n12290) );
  NAND2_X1 U9770 ( .A1(n15538), .A2(n11346), .ZN(n7351) );
  NAND2_X1 U9771 ( .A1(n7360), .A2(n7358), .ZN(n11343) );
  NAND2_X1 U9772 ( .A1(n12319), .A2(n6599), .ZN(n7360) );
  INV_X1 U9773 ( .A(n8323), .ZN(n7364) );
  NOR2_X2 U9774 ( .A1(n13543), .A2(n13414), .ZN(n13396) );
  NAND2_X1 U9775 ( .A1(n11662), .A2(n11663), .ZN(n11822) );
  NAND2_X1 U9776 ( .A1(n7375), .A2(n7374), .ZN(n11098) );
  NAND2_X1 U9777 ( .A1(n10859), .A2(n6673), .ZN(n7375) );
  NOR2_X1 U9778 ( .A1(n7378), .A2(n11641), .ZN(n11642) );
  NAND2_X1 U9779 ( .A1(n7377), .A2(n11640), .ZN(n11900) );
  XNOR2_X1 U9780 ( .A(n11997), .B(n11807), .ZN(n10213) );
  INV_X1 U9781 ( .A(n7391), .ZN(n7390) );
  NAND2_X1 U9782 ( .A1(n7390), .A2(n11351), .ZN(n13449) );
  NAND2_X1 U9783 ( .A1(n11025), .A2(n7409), .ZN(n8088) );
  NAND2_X1 U9784 ( .A1(n10403), .A2(n9982), .ZN(n7414) );
  NAND2_X1 U9785 ( .A1(n7877), .A2(n7415), .ZN(n7416) );
  INV_X2 U9786 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14897) );
  NAND2_X2 U9787 ( .A1(n7426), .A2(n7424), .ZN(n15370) );
  AND2_X1 U9788 ( .A1(n7436), .A2(n6671), .ZN(n7434) );
  XNOR2_X2 U9789 ( .A(n7443), .B(n13149), .ZN(n13487) );
  OR2_X1 U9790 ( .A1(n14880), .A2(n7448), .ZN(n7446) );
  AND2_X1 U9791 ( .A1(n7453), .A2(n7449), .ZN(n7448) );
  OR2_X1 U9792 ( .A1(n14880), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7452) );
  OR2_X1 U9793 ( .A1(n14979), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7454) );
  NAND2_X1 U9794 ( .A1(n7457), .A2(n14809), .ZN(n14811) );
  INV_X1 U9795 ( .A(n12812), .ZN(n7464) );
  NAND4_X1 U9796 ( .A1(n9372), .A2(n9049), .A3(n8961), .A4(n13813), .ZN(n9442)
         );
  OAI21_X1 U9797 ( .B1(n14284), .B2(n8285), .A(n8287), .ZN(n7491) );
  NAND2_X1 U9798 ( .A1(n9764), .A2(n6579), .ZN(n7493) );
  INV_X1 U9799 ( .A(n7506), .ZN(n14448) );
  NOR2_X1 U9800 ( .A1(n8300), .A2(n14490), .ZN(n7514) );
  NAND2_X1 U9801 ( .A1(n14229), .A2(n7518), .ZN(n7517) );
  NAND2_X1 U9802 ( .A1(n14152), .A2(n7525), .ZN(n7524) );
  INV_X1 U9803 ( .A(n14153), .ZN(n7526) );
  NAND3_X1 U9804 ( .A1(n14212), .A2(n14211), .A3(n7529), .ZN(n7527) );
  NAND2_X1 U9805 ( .A1(n7527), .A2(n7528), .ZN(n14219) );
  NAND2_X1 U9806 ( .A1(n7532), .A2(n7535), .ZN(n14266) );
  NAND2_X1 U9807 ( .A1(n14237), .A2(n7533), .ZN(n7532) );
  NOR2_X2 U9808 ( .A1(n7702), .A2(n7703), .ZN(n7704) );
  INV_X1 U9809 ( .A(n14133), .ZN(n7555) );
  OAI21_X1 U9810 ( .B1(n7556), .B2(n13244), .A(n13155), .ZN(n13173) );
  NAND2_X1 U9811 ( .A1(n13154), .A2(n13153), .ZN(n7556) );
  NAND2_X1 U9812 ( .A1(n13076), .A2(n13113), .ZN(n13116) );
  NAND2_X1 U9813 ( .A1(n7789), .A2(n6574), .ZN(n7562) );
  NAND2_X1 U9814 ( .A1(n8198), .A2(n7829), .ZN(n7574) );
  NAND2_X1 U9815 ( .A1(n8198), .A2(n6595), .ZN(n7578) );
  OAI21_X1 U9816 ( .B1(n8235), .B2(n7589), .A(n7587), .ZN(n8262) );
  AOI21_X1 U9817 ( .B1(n8234), .B2(n7836), .A(n6709), .ZN(n7590) );
  OR2_X1 U9818 ( .A1(n8235), .A2(n8234), .ZN(n8237) );
  NAND2_X1 U9819 ( .A1(n7824), .A2(n7825), .ZN(n7592) );
  INV_X1 U9820 ( .A(n12032), .ZN(n7594) );
  NAND2_X1 U9821 ( .A1(n11165), .A2(n7603), .ZN(n7602) );
  NAND2_X1 U9822 ( .A1(n12414), .A2(n7622), .ZN(n7621) );
  NAND2_X1 U9823 ( .A1(n12414), .A2(n12084), .ZN(n12397) );
  INV_X1 U9824 ( .A(n12084), .ZN(n7623) );
  NAND3_X1 U9825 ( .A1(n8573), .A2(n8332), .A3(n8324), .ZN(n8334) );
  AND2_X1 U9826 ( .A1(n8894), .A2(n8410), .ZN(n8888) );
  NOR2_X2 U9827 ( .A1(n15078), .A2(n15188), .ZN(n14938) );
  NAND2_X1 U9828 ( .A1(n11773), .A2(n7644), .ZN(n7642) );
  NAND2_X1 U9829 ( .A1(n7642), .A2(n7643), .ZN(n13913) );
  AND2_X1 U9830 ( .A1(n13941), .A2(n7651), .ZN(n7648) );
  INV_X1 U9831 ( .A(n9609), .ZN(n7650) );
  INV_X1 U9832 ( .A(n9608), .ZN(n7649) );
  INV_X1 U9833 ( .A(n11120), .ZN(n11118) );
  NAND2_X1 U9834 ( .A1(n7751), .A2(n7842), .ZN(n7754) );
  NAND2_X1 U9835 ( .A1(n7751), .A2(n7654), .ZN(n14737) );
  NAND2_X1 U9836 ( .A1(n14060), .A2(n11692), .ZN(n13989) );
  NAND2_X1 U9837 ( .A1(n11297), .A2(n11296), .ZN(n11309) );
  NAND2_X1 U9838 ( .A1(n13969), .A2(n14030), .ZN(n11744) );
  NAND4_X1 U9839 ( .A1(n7704), .A2(n7688), .A3(n7549), .A4(n7658), .ZN(n7841)
         );
  NAND2_X1 U9840 ( .A1(n7659), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9300) );
  NAND2_X2 U9841 ( .A1(n9285), .A2(n13887), .ZN(n9296) );
  XNOR2_X2 U9842 ( .A(n7660), .B(n9282), .ZN(n9285) );
  OAI21_X1 U9843 ( .B1(n13023), .B2(n7672), .A(n7671), .ZN(n13030) );
  INV_X1 U9844 ( .A(n7668), .ZN(n13029) );
  NAND3_X1 U9845 ( .A1(n13003), .A2(n13002), .A3(n6689), .ZN(n7685) );
  NAND2_X1 U9846 ( .A1(n7685), .A2(n7686), .ZN(n13011) );
  INV_X1 U9847 ( .A(n12366), .ZN(n12367) );
  XNOR2_X1 U9848 ( .A(n12179), .B(n12015), .ZN(n12008) );
  NAND2_X1 U9849 ( .A1(n11167), .A2(n7607), .ZN(n11166) );
  XNOR2_X1 U9850 ( .A(n11561), .B(n11569), .ZN(n11565) );
  XNOR2_X1 U9851 ( .A(n11955), .B(n8834), .ZN(n11621) );
  NAND2_X1 U9852 ( .A1(n7841), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7843) );
  OR2_X1 U9853 ( .A1(n8255), .A2(n13915), .ZN(n8258) );
  AOI21_X2 U9854 ( .B1(n11584), .B2(n11982), .A(n8861), .ZN(n11955) );
  INV_X1 U9855 ( .A(n9286), .ZN(n13887) );
  INV_X1 U9856 ( .A(n14081), .ZN(n8309) );
  NAND2_X1 U9857 ( .A1(n9283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9284) );
  INV_X1 U9858 ( .A(n13965), .ZN(n9923) );
  INV_X1 U9859 ( .A(n8827), .ZN(n10337) );
  INV_X1 U9860 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8423) );
  INV_X1 U9861 ( .A(n8139), .ZN(n8140) );
  NAND4_X1 U9862 ( .A1(n8260), .A2(n8259), .A3(n8258), .A4(n8257), .ZN(n14317)
         );
  INV_X1 U9863 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8048) );
  INV_X1 U9864 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8419) );
  NAND4_X1 U9865 ( .A1(n8246), .A2(n8245), .A3(n8244), .A4(n8243), .ZN(n14318)
         );
  AND2_X1 U9866 ( .A1(n10037), .A2(n10036), .ZN(n7691) );
  AND2_X1 U9867 ( .A1(n7806), .A2(n7805), .ZN(n7692) );
  AND2_X1 U9868 ( .A1(n11130), .A2(n11149), .ZN(n7693) );
  INV_X1 U9869 ( .A(n14278), .ZN(n15095) );
  OR2_X1 U9870 ( .A1(n14652), .A2(n8247), .ZN(n7694) );
  INV_X1 U9871 ( .A(n14652), .ZN(n14463) );
  NAND2_X1 U9872 ( .A1(n9780), .A2(n13397), .ZN(n12831) );
  OR2_X1 U9873 ( .A1(n11617), .A2(n12613), .ZN(n7695) );
  OR2_X1 U9874 ( .A1(n11617), .A2(n12556), .ZN(n7696) );
  NAND2_X2 U9875 ( .A1(n10241), .A2(n12387), .ZN(n12490) );
  NAND2_X1 U9876 ( .A1(n13212), .A2(n13036), .ZN(n12869) );
  AND2_X1 U9877 ( .A1(n12978), .A2(n12976), .ZN(n12977) );
  INV_X2 U9878 ( .A(n12961), .ZN(n13036) );
  OAI21_X1 U9879 ( .B1(n13043), .B2(n13036), .A(n13042), .ZN(n13044) );
  INV_X1 U9880 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7698) );
  NOR2_X1 U9881 ( .A1(n12481), .A2(n11093), .ZN(n11092) );
  INV_X1 U9882 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8407) );
  INV_X1 U9883 ( .A(n7986), .ZN(n7790) );
  OR2_X1 U9884 ( .A1(n11094), .A2(n11145), .ZN(n11096) );
  OR2_X1 U9885 ( .A1(n12539), .A2(n11934), .ZN(n8853) );
  OR2_X1 U9886 ( .A1(n11829), .A2(n12543), .ZN(n8852) );
  INV_X1 U9887 ( .A(n13116), .ZN(n13154) );
  INV_X1 U9888 ( .A(n11374), .ZN(n11372) );
  OR2_X1 U9889 ( .A1(n9205), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8967) );
  INV_X1 U9890 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8965) );
  INV_X1 U9891 ( .A(n14318), .ZN(n8247) );
  INV_X1 U9892 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8030) );
  INV_X1 U9893 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8421) );
  INV_X1 U9894 ( .A(n8770), .ZN(n8440) );
  AND2_X1 U9895 ( .A1(n11096), .A2(n11095), .ZN(n11097) );
  INV_X1 U9896 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n8418) );
  AND2_X1 U9897 ( .A1(n10237), .A2(n10236), .ZN(n10238) );
  INV_X1 U9898 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8410) );
  AND2_X1 U9899 ( .A1(n8383), .A2(n8382), .ZN(n8668) );
  INV_X1 U9900 ( .A(n11398), .ZN(n11397) );
  OR3_X1 U9901 ( .A1(n15357), .A2(n9942), .A3(n9774), .ZN(n9785) );
  OR2_X1 U9902 ( .A1(n11423), .A2(n11422), .ZN(n11437) );
  OR2_X1 U9903 ( .A1(n11363), .A2(n11362), .ZN(n11374) );
  AND2_X1 U9904 ( .A1(n13172), .A2(n10346), .ZN(n9805) );
  OR2_X1 U9905 ( .A1(n15423), .A2(n10346), .ZN(n9784) );
  INV_X1 U9906 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8985) );
  INV_X1 U9907 ( .A(n13921), .ZN(n11687) );
  NAND2_X1 U9908 ( .A1(n14084), .A2(n14085), .ZN(n14103) );
  AOI21_X1 U9909 ( .B1(n10307), .B2(n15141), .A(n8989), .ZN(n8990) );
  NOR2_X1 U9910 ( .A1(n13973), .A2(n8201), .ZN(n8214) );
  NAND2_X1 U9911 ( .A1(n8080), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U9912 ( .A1(n8241), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8240) );
  AND2_X1 U9913 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n8254), .ZN(n7757) );
  NAND2_X1 U9914 ( .A1(n7853), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7852) );
  INV_X1 U9915 ( .A(n8213), .ZN(n8228) );
  NAND2_X1 U9916 ( .A1(n8186), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8201) );
  OR2_X1 U9917 ( .A1(n8031), .A2(n8030), .ZN(n8049) );
  AND2_X1 U9918 ( .A1(n9391), .A2(n7729), .ZN(n10043) );
  NAND2_X1 U9919 ( .A1(n7811), .A2(n13778), .ZN(n7814) );
  NOR2_X1 U9920 ( .A1(n14810), .A2(n14773), .ZN(n14774) );
  AND2_X1 U9921 ( .A1(n10340), .A2(n10339), .ZN(n12284) );
  INV_X1 U9922 ( .A(n10259), .ZN(n10254) );
  INV_X1 U9923 ( .A(n12065), .ZN(n12461) );
  OR2_X1 U9924 ( .A1(n8527), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8541) );
  OR2_X1 U9925 ( .A1(n12284), .A2(n12283), .ZN(n12495) );
  OR2_X1 U9926 ( .A1(n11951), .A2(n10874), .ZN(n8780) );
  OR2_X1 U9927 ( .A1(n11951), .A2(n7579), .ZN(n8751) );
  INV_X1 U9928 ( .A(n12163), .ZN(n8925) );
  INV_X1 U9929 ( .A(n12474), .ZN(n12404) );
  AND2_X1 U9930 ( .A1(n8344), .A2(n8924), .ZN(n11601) );
  NAND2_X1 U9931 ( .A1(n8904), .A2(n8903), .ZN(n10235) );
  NAND2_X1 U9932 ( .A1(n8727), .A2(n8391), .ZN(n8738) );
  NAND2_X1 U9933 ( .A1(n8671), .A2(n8383), .ZN(n8683) );
  NAND2_X1 U9934 ( .A1(n11397), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n11423) );
  OR3_X1 U9935 ( .A1(n11456), .A2(n12779), .A3(n12752), .ZN(n11467) );
  NAND2_X1 U9936 ( .A1(n10905), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n11363) );
  INV_X1 U9937 ( .A(n12808), .ZN(n12848) );
  OR2_X1 U9938 ( .A1(n11467), .A2(n13662), .ZN(n11489) );
  INV_X1 U9939 ( .A(n12838), .ZN(n12860) );
  OR2_X1 U9940 ( .A1(n11437), .A2(n12711), .ZN(n11456) );
  OR2_X1 U9941 ( .A1(n13457), .A2(n13456), .ZN(n13563) );
  NAND2_X1 U9942 ( .A1(n10692), .A2(n10694), .ZN(n10695) );
  OR2_X1 U9943 ( .A1(n9400), .A2(n9399), .ZN(n14055) );
  OR2_X1 U9944 ( .A1(n8255), .A2(n11804), .ZN(n7762) );
  NAND2_X1 U9945 ( .A1(n8144), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8158) );
  NOR2_X1 U9946 ( .A1(n8128), .A2(n8127), .ZN(n8144) );
  INV_X1 U9947 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10538) );
  XNOR2_X1 U9948 ( .A(n14335), .B(n14116), .ZN(n14269) );
  NAND2_X1 U9949 ( .A1(n15104), .A2(n9768), .ZN(n14541) );
  INV_X1 U9950 ( .A(n14934), .ZN(n14969) );
  OR2_X1 U9951 ( .A1(n7730), .A2(P1_B_REG_SCAN_IN), .ZN(n7733) );
  INV_X1 U9952 ( .A(n11916), .ZN(n11858) );
  AND2_X1 U9953 ( .A1(n9871), .A2(n12480), .ZN(n11931) );
  INV_X1 U9954 ( .A(n11935), .ZN(n11904) );
  AOI21_X1 U9955 ( .B1(n11811), .B2(n8484), .A(n8819), .ZN(n11666) );
  AND3_X1 U9956 ( .A1(n8773), .A2(n8772), .A3(n8771), .ZN(n12335) );
  NAND2_X1 U9957 ( .A1(n8917), .A2(n8916), .ZN(n9735) );
  AND2_X1 U9958 ( .A1(n9548), .A2(n12275), .ZN(n15461) );
  AND2_X1 U9959 ( .A1(n9543), .A2(n9544), .ZN(n9548) );
  AND2_X1 U9960 ( .A1(n8883), .A2(n12103), .ZN(n12480) );
  AND2_X1 U9961 ( .A1(n8923), .A2(n8922), .ZN(n10239) );
  INV_X1 U9962 ( .A(n15515), .ZN(n15508) );
  INV_X1 U9963 ( .A(n12500), .ZN(n15518) );
  AND2_X1 U9964 ( .A1(n9735), .A2(n9110), .ZN(n12159) );
  AND2_X1 U9965 ( .A1(n9807), .A2(n9806), .ZN(n12846) );
  INV_X1 U9966 ( .A(n12867), .ZN(n13172) );
  INV_X1 U9967 ( .A(n13239), .ZN(n15302) );
  AND2_X1 U9968 ( .A1(n9222), .A2(n9216), .ZN(n15296) );
  NOR2_X1 U9969 ( .A1(n15320), .A2(n13575), .ZN(n13406) );
  INV_X1 U9970 ( .A(n13562), .ZN(n13431) );
  NAND2_X1 U9971 ( .A1(n9278), .A2(n15354), .ZN(n9942) );
  INV_X1 U9972 ( .A(n15409), .ZN(n13575) );
  NAND2_X1 U9973 ( .A1(n9304), .A2(n9303), .ZN(n15409) );
  INV_X1 U9974 ( .A(n9942), .ZN(n10344) );
  AND2_X1 U9975 ( .A1(n9258), .A2(n9277), .ZN(n15321) );
  AND2_X1 U9976 ( .A1(n9263), .A2(n9262), .ZN(n9787) );
  INV_X1 U9977 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9057) );
  AND4_X1 U9978 ( .A1(n8219), .A2(n8218), .A3(n8217), .A4(n8216), .ZN(n14216)
         );
  INV_X1 U9979 ( .A(n15027), .ZN(n15035) );
  INV_X1 U9980 ( .A(n15025), .ZN(n15040) );
  INV_X1 U9981 ( .A(n14583), .ZN(n15101) );
  INV_X1 U9982 ( .A(n14541), .ZN(n15075) );
  NAND2_X1 U9983 ( .A1(n7747), .A2(n7746), .ZN(n9761) );
  INV_X1 U9984 ( .A(n15139), .ZN(n15084) );
  AND2_X1 U9985 ( .A1(n15068), .A2(n15163), .ZN(n14964) );
  INV_X1 U9986 ( .A(n14964), .ZN(n15195) );
  NAND3_X1 U9987 ( .A1(n7733), .A2(n7732), .A3(n7731), .ZN(n9100) );
  AND2_X1 U9988 ( .A1(n9545), .A2(n9544), .ZN(n15458) );
  INV_X1 U9989 ( .A(n11938), .ZN(n10872) );
  AND2_X1 U9990 ( .A1(n9754), .A2(n12387), .ZN(n11935) );
  INV_X1 U9991 ( .A(n11923), .ZN(n12169) );
  INV_X1 U9992 ( .A(n12381), .ZN(n12172) );
  INV_X1 U9993 ( .A(n12280), .ZN(n15454) );
  NAND2_X1 U9994 ( .A1(n9548), .A2(n9542), .ZN(n15465) );
  NAND2_X1 U9995 ( .A1(n12490), .A2(n10301), .ZN(n12493) );
  NAND2_X1 U9996 ( .A1(n15540), .A2(n15508), .ZN(n12556) );
  INV_X1 U9997 ( .A(n15540), .ZN(n15538) );
  INV_X1 U9998 ( .A(n11622), .ZN(n11671) );
  AND2_X2 U9999 ( .A1(n8941), .A2(n12159), .ZN(n15519) );
  INV_X1 U10000 ( .A(n15519), .ZN(n15521) );
  INV_X1 U10001 ( .A(SI_18_), .ZN(n13597) );
  INV_X1 U10002 ( .A(SI_14_), .ZN(n9183) );
  INV_X1 U10003 ( .A(n10612), .ZN(n10631) );
  INV_X1 U10004 ( .A(n9882), .ZN(n9895) );
  INV_X1 U10005 ( .A(n13460), .ZN(n13561) );
  INV_X2 U10006 ( .A(n12846), .ZN(n12854) );
  INV_X1 U10007 ( .A(n12831), .ZN(n12866) );
  OR2_X1 U10008 ( .A1(n15237), .A2(P2_U3088), .ZN(n15273) );
  INV_X1 U10009 ( .A(n15296), .ZN(n15242) );
  OR2_X1 U10010 ( .A1(n9943), .A2(n9942), .ZN(n15441) );
  OR3_X1 U10011 ( .A1(n13566), .A2(n13565), .A3(n13564), .ZN(n13875) );
  OR2_X1 U10012 ( .A1(n9943), .A2(n10344), .ZN(n15429) );
  NOR2_X1 U10013 ( .A1(n15321), .A2(n15355), .ZN(n15336) );
  INV_X1 U10014 ( .A(n15358), .ZN(n15355) );
  NAND2_X1 U10015 ( .A1(n9260), .A2(n9259), .ZN(n15357) );
  INV_X1 U10016 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11434) );
  INV_X1 U10017 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9505) );
  INV_X1 U10018 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9782) );
  AND2_X1 U10019 ( .A1(n9003), .A2(n9001), .ZN(n15006) );
  INV_X1 U10020 ( .A(n14097), .ZN(n14316) );
  INV_X1 U10021 ( .A(n11690), .ZN(n14324) );
  OR2_X1 U10022 ( .A1(n15004), .A2(n6559), .ZN(n15027) );
  INV_X1 U10023 ( .A(n15006), .ZN(n15047) );
  NAND2_X1 U10024 ( .A1(n15104), .A2(n9766), .ZN(n14623) );
  OR2_X1 U10025 ( .A1(n9633), .A2(n9761), .ZN(n15206) );
  NAND2_X1 U10026 ( .A1(n15196), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8319) );
  OR2_X1 U10027 ( .A1(n9633), .A2(n9390), .ZN(n15196) );
  INV_X2 U10028 ( .A(n15196), .ZN(n15197) );
  INV_X1 U10029 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9655) );
  INV_X1 U10030 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9446) );
  INV_X1 U10031 ( .A(n12181), .ZN(P3_U3897) );
  OAI21_X1 U10032 ( .B1(n12613), .B2(n8956), .A(n8958), .ZN(P3_U3455) );
  AND2_X1 U10033 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9214), .ZN(P2_U3947) );
  INV_X1 U10034 ( .A(n14337), .ZN(P1_U4016) );
  NAND3_X1 U10035 ( .A1(n8102), .A2(n8003), .A3(n7988), .ZN(n7703) );
  NOR2_X1 U10036 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .ZN(n7701) );
  NAND4_X1 U10037 ( .A1(n7701), .A2(n7700), .A3(n7699), .A4(n7698), .ZN(n7702)
         );
  NOR2_X1 U10038 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n7711) );
  NOR2_X1 U10039 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n7710) );
  OAI21_X1 U10040 ( .B1(n7750), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U10041 ( .A1(n7750), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7714) );
  XNOR2_X1 U10042 ( .A(n7714), .B(n7749), .ZN(n14751) );
  OR3_X2 U10043 ( .A1(n7730), .A2(n14748), .A3(n14751), .ZN(n10044) );
  NAND2_X1 U10044 ( .A1(n7715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7716) );
  XNOR2_X1 U10045 ( .A(n7716), .B(P1_IR_REG_23__SCAN_IN), .ZN(n8998) );
  INV_X1 U10046 ( .A(n8998), .ZN(n7717) );
  NAND2_X1 U10047 ( .A1(n7719), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7720) );
  MUX2_X1 U10048 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7720), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n7721) );
  NAND2_X1 U10049 ( .A1(n14756), .A2(n14084), .ZN(n14092) );
  INV_X1 U10050 ( .A(n14092), .ZN(n9391) );
  NAND2_X1 U10051 ( .A1(n7728), .A2(n7727), .ZN(n7724) );
  NAND2_X1 U10052 ( .A1(n14085), .A2(n14617), .ZN(n7729) );
  NOR2_X1 U10053 ( .A1(n9395), .A2(n10043), .ZN(n14309) );
  NAND3_X1 U10054 ( .A1(n7730), .A2(P1_B_REG_SCAN_IN), .A3(n14751), .ZN(n7732)
         );
  INV_X1 U10055 ( .A(n14748), .ZN(n7731) );
  OR2_X1 U10056 ( .A1(n9100), .A2(P1_D_REG_1__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U10057 ( .A1(n14748), .A2(n14751), .ZN(n7734) );
  NAND2_X1 U10058 ( .A1(n7735), .A2(n7734), .ZN(n9389) );
  NOR2_X1 U10059 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .ZN(
        n13843) );
  NOR4_X1 U10060 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n7738) );
  NOR4_X1 U10061 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n7737) );
  NOR4_X1 U10062 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n7736) );
  AND4_X1 U10063 ( .A1(n13843), .A2(n7738), .A3(n7737), .A4(n7736), .ZN(n7744)
         );
  NOR4_X1 U10064 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n7742) );
  NOR4_X1 U10065 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n7741) );
  NOR4_X1 U10066 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n7740) );
  NOR4_X1 U10067 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n7739) );
  AND4_X1 U10068 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .ZN(n7743)
         );
  AND2_X1 U10069 ( .A1(n7744), .A2(n7743), .ZN(n7745) );
  OR2_X1 U10070 ( .A1(n9100), .A2(n7745), .ZN(n9760) );
  NAND2_X1 U10071 ( .A1(n8306), .A2(n14085), .ZN(n14091) );
  NAND2_X1 U10072 ( .A1(n8988), .A2(n14598), .ZN(n9396) );
  NAND4_X1 U10073 ( .A1(n14309), .A2(n9389), .A3(n9760), .A4(n9396), .ZN(n9633) );
  OR2_X1 U10074 ( .A1(n9100), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7747) );
  NAND2_X1 U10075 ( .A1(n7730), .A2(n14748), .ZN(n7746) );
  INV_X1 U10076 ( .A(n9761), .ZN(n9390) );
  INV_X1 U10077 ( .A(n7841), .ZN(n7751) );
  NAND2_X1 U10078 ( .A1(n14077), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7764) );
  INV_X1 U10079 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n13782) );
  OR2_X1 U10080 ( .A1(n14081), .A2(n13782), .ZN(n7763) );
  INV_X1 U10081 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13973) );
  NAND2_X1 U10082 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7935) );
  NAND2_X1 U10083 ( .A1(n7949), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U10084 ( .A1(n8009), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8031) );
  INV_X1 U10085 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8108) );
  INV_X1 U10086 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8127) );
  INV_X1 U10087 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8157) );
  INV_X1 U10088 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U10089 ( .A1(n8214), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U10090 ( .A1(n7757), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14430) );
  INV_X1 U10091 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7759) );
  INV_X1 U10092 ( .A(n7757), .ZN(n7758) );
  NAND2_X1 U10093 ( .A1(n7759), .A2(n7758), .ZN(n7760) );
  NAND2_X1 U10094 ( .A1(n14430), .A2(n7760), .ZN(n11804) );
  INV_X1 U10095 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n11567) );
  OR2_X1 U10096 ( .A1(n8267), .A2(n11567), .ZN(n7761) );
  INV_X1 U10097 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9038) );
  AND2_X1 U10098 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7768) );
  INV_X1 U10099 ( .A(SI_1_), .ZN(n9067) );
  NAND2_X1 U10100 ( .A1(n7770), .A2(SI_2_), .ZN(n7771) );
  INV_X1 U10101 ( .A(n7904), .ZN(n7773) );
  NAND2_X1 U10102 ( .A1(n7774), .A2(SI_3_), .ZN(n7775) );
  XNOR2_X1 U10103 ( .A(n7777), .B(SI_4_), .ZN(n7908) );
  INV_X1 U10104 ( .A(n7908), .ZN(n7776) );
  MUX2_X1 U10105 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n13064), .Z(n7779) );
  XNOR2_X1 U10106 ( .A(n7779), .B(SI_5_), .ZN(n7924) );
  INV_X1 U10107 ( .A(n7924), .ZN(n7778) );
  NAND2_X1 U10108 ( .A1(n7925), .A2(n7778), .ZN(n7781) );
  NAND2_X1 U10109 ( .A1(n7779), .A2(SI_5_), .ZN(n7780) );
  XNOR2_X1 U10110 ( .A(n7783), .B(SI_6_), .ZN(n7943) );
  INV_X1 U10111 ( .A(n7943), .ZN(n7782) );
  NAND2_X1 U10112 ( .A1(n7783), .A2(SI_6_), .ZN(n7784) );
  MUX2_X1 U10113 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n13064), .Z(n7785) );
  XNOR2_X1 U10114 ( .A(n7785), .B(SI_7_), .ZN(n7956) );
  MUX2_X1 U10115 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n13064), .Z(n7787) );
  XNOR2_X1 U10116 ( .A(n7787), .B(SI_8_), .ZN(n7972) );
  INV_X1 U10117 ( .A(n7972), .ZN(n7786) );
  NAND2_X1 U10118 ( .A1(n7787), .A2(SI_8_), .ZN(n7788) );
  MUX2_X1 U10119 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n13064), .Z(n7791) );
  MUX2_X1 U10120 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n13064), .Z(n8019) );
  INV_X1 U10121 ( .A(n8019), .ZN(n7792) );
  MUX2_X1 U10122 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n13064), .Z(n7793) );
  OAI21_X1 U10123 ( .B1(n7792), .B2(n13829), .A(n8025), .ZN(n7798) );
  NOR2_X1 U10124 ( .A1(n8019), .A2(SI_10_), .ZN(n7796) );
  INV_X1 U10125 ( .A(n7793), .ZN(n7794) );
  INV_X1 U10126 ( .A(SI_11_), .ZN(n9080) );
  NAND2_X1 U10127 ( .A1(n7794), .A2(n9080), .ZN(n8024) );
  INV_X1 U10128 ( .A(n8024), .ZN(n7795) );
  AOI21_X1 U10129 ( .B1(n7796), .B2(n8025), .A(n7795), .ZN(n7797) );
  MUX2_X1 U10130 ( .A(n9446), .B(n9444), .S(n13064), .Z(n7799) );
  NAND2_X1 U10131 ( .A1(n7799), .A2(n13820), .ZN(n7802) );
  INV_X1 U10132 ( .A(n7799), .ZN(n7800) );
  NAND2_X1 U10133 ( .A1(n7800), .A2(SI_12_), .ZN(n7801) );
  MUX2_X1 U10134 ( .A(n9501), .B(n9505), .S(n13064), .Z(n7803) );
  NAND2_X1 U10135 ( .A1(n7803), .A2(n9128), .ZN(n7806) );
  INV_X1 U10136 ( .A(n7803), .ZN(n7804) );
  NAND2_X1 U10137 ( .A1(n7804), .A2(SI_13_), .ZN(n7805) );
  MUX2_X1 U10138 ( .A(n9617), .B(n9615), .S(n13064), .Z(n8073) );
  MUX2_X1 U10139 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n13064), .Z(n7808) );
  OAI21_X1 U10140 ( .B1(n8073), .B2(n9183), .A(n8097), .ZN(n7807) );
  INV_X1 U10141 ( .A(n8073), .ZN(n8089) );
  NOR2_X1 U10142 ( .A1(n8089), .A2(SI_14_), .ZN(n7809) );
  NOR2_X1 U10143 ( .A1(n7808), .A2(SI_15_), .ZN(n8095) );
  MUX2_X1 U10144 ( .A(n13776), .B(n9600), .S(n13064), .Z(n7811) );
  INV_X1 U10145 ( .A(n7811), .ZN(n7812) );
  NAND2_X1 U10146 ( .A1(n7812), .A2(SI_16_), .ZN(n7813) );
  MUX2_X1 U10147 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n13064), .Z(n8134) );
  INV_X1 U10148 ( .A(n8134), .ZN(n7816) );
  NAND2_X1 U10149 ( .A1(n7817), .A2(n13597), .ZN(n7818) );
  MUX2_X1 U10150 ( .A(n9835), .B(n9837), .S(n13064), .Z(n8150) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n13064), .Z(n7820) );
  XNOR2_X1 U10152 ( .A(n7820), .B(SI_19_), .ZN(n8169) );
  INV_X1 U10153 ( .A(n7820), .ZN(n7821) );
  INV_X1 U10154 ( .A(SI_19_), .ZN(n9681) );
  NAND2_X1 U10155 ( .A1(n7821), .A2(n9681), .ZN(n7822) );
  INV_X1 U10156 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11394) );
  MUX2_X1 U10157 ( .A(n10498), .B(n11394), .S(n13064), .Z(n8180) );
  MUX2_X1 U10158 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n13064), .Z(n7827) );
  NAND2_X1 U10159 ( .A1(n7827), .A2(SI_21_), .ZN(n7829) );
  OAI21_X1 U10160 ( .B1(SI_21_), .B2(n7827), .A(n7829), .ZN(n7828) );
  INV_X1 U10161 ( .A(n7828), .ZN(n8195) );
  INV_X1 U10162 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8394) );
  INV_X1 U10163 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13738) );
  MUX2_X1 U10164 ( .A(n8394), .B(n13738), .S(n13064), .Z(n11155) );
  MUX2_X1 U10165 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n13064), .Z(n8221) );
  INV_X1 U10166 ( .A(n8221), .ZN(n7830) );
  INV_X1 U10167 ( .A(SI_23_), .ZN(n10156) );
  NOR2_X1 U10168 ( .A1(n7830), .A2(n10156), .ZN(n7831) );
  MUX2_X1 U10169 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n13064), .Z(n7832) );
  NAND2_X1 U10170 ( .A1(n7832), .A2(SI_24_), .ZN(n7833) );
  OAI21_X1 U10171 ( .B1(SI_24_), .B2(n7832), .A(n7833), .ZN(n7858) );
  MUX2_X1 U10172 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n13064), .Z(n7834) );
  XNOR2_X1 U10173 ( .A(n7834), .B(SI_25_), .ZN(n7847) );
  OAI22_X1 U10174 ( .A1(n7848), .A2(n7847), .B1(SI_25_), .B2(n7834), .ZN(n8235) );
  MUX2_X1 U10175 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n13064), .Z(n7835) );
  NAND2_X1 U10176 ( .A1(n7835), .A2(SI_26_), .ZN(n7836) );
  OAI21_X1 U10177 ( .B1(SI_26_), .B2(n7835), .A(n7836), .ZN(n8234) );
  INV_X1 U10178 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11329) );
  INV_X1 U10179 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13897) );
  MUX2_X1 U10180 ( .A(n11329), .B(n13897), .S(n13064), .Z(n7837) );
  INV_X1 U10181 ( .A(SI_27_), .ZN(n11161) );
  INV_X1 U10182 ( .A(n7837), .ZN(n8249) );
  INV_X1 U10183 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13588) );
  INV_X1 U10184 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n11484) );
  MUX2_X1 U10185 ( .A(n13588), .B(n11484), .S(n13064), .Z(n7838) );
  INV_X1 U10186 ( .A(SI_28_), .ZN(n11082) );
  NAND2_X1 U10187 ( .A1(n7838), .A2(n11082), .ZN(n8263) );
  INV_X1 U10188 ( .A(n7838), .ZN(n7839) );
  NAND2_X1 U10189 ( .A1(n7839), .A2(SI_28_), .ZN(n7840) );
  NAND2_X1 U10190 ( .A1(n8263), .A2(n7840), .ZN(n8261) );
  NAND2_X1 U10191 ( .A1(n11483), .A2(n14087), .ZN(n7846) );
  OR2_X1 U10192 ( .A1(n7896), .A2(n13588), .ZN(n7845) );
  XNOR2_X1 U10193 ( .A(n7848), .B(n7847), .ZN(n13901) );
  NAND2_X1 U10194 ( .A1(n13901), .A2(n14087), .ZN(n7850) );
  INV_X1 U10195 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14754) );
  OR2_X1 U10196 ( .A1(n7896), .A2(n14754), .ZN(n7849) );
  NAND2_X1 U10197 ( .A1(n8309), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7857) );
  INV_X1 U10198 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n7851) );
  OR2_X1 U10199 ( .A1(n8312), .A2(n7851), .ZN(n7856) );
  OAI21_X1 U10200 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n7853), .A(n7852), .ZN(
        n14479) );
  OR2_X1 U10201 ( .A1(n8255), .A2(n14479), .ZN(n7855) );
  INV_X1 U10202 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14480) );
  OR2_X1 U10203 ( .A1(n8267), .A2(n14480), .ZN(n7854) );
  NAND4_X1 U10204 ( .A1(n7857), .A2(n7856), .A3(n7855), .A4(n7854), .ZN(n14319) );
  NAND2_X1 U10205 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  NAND2_X1 U10206 ( .A1(n11444), .A2(n14087), .ZN(n7863) );
  OR2_X1 U10207 ( .A1(n7896), .A2(n7291), .ZN(n7862) );
  INV_X1 U10208 ( .A(n14664), .ZN(n14497) );
  NAND2_X1 U10209 ( .A1(n14077), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7869) );
  INV_X1 U10210 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n13730) );
  OR2_X1 U10211 ( .A1(n14081), .A2(n13730), .ZN(n7868) );
  OAI21_X1 U10212 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n7865), .A(n7864), .ZN(
        n14498) );
  OR2_X1 U10213 ( .A1(n8255), .A2(n14498), .ZN(n7867) );
  INV_X1 U10214 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14499) );
  OR2_X1 U10215 ( .A1(n8267), .A2(n14499), .ZN(n7866) );
  NAND4_X1 U10216 ( .A1(n7869), .A2(n7868), .A3(n7867), .A4(n7866), .ZN(n14512) );
  NAND2_X1 U10217 ( .A1(n14077), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7873) );
  INV_X1 U10218 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7870) );
  INV_X1 U10219 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9013) );
  OR2_X1 U10220 ( .A1(n14081), .A2(n9013), .ZN(n7871) );
  INV_X1 U10221 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10222 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n7874) );
  XNOR2_X1 U10223 ( .A(n7875), .B(n7874), .ZN(n14342) );
  XNOR2_X1 U10224 ( .A(n7877), .B(n7876), .ZN(n9292) );
  INV_X1 U10225 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n14625) );
  OR2_X1 U10226 ( .A1(n8255), .A2(n14625), .ZN(n7882) );
  INV_X1 U10227 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7879) );
  OR2_X1 U10228 ( .A1(n8312), .A2(n7879), .ZN(n7881) );
  INV_X1 U10229 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15000) );
  OR2_X1 U10230 ( .A1(n14081), .A2(n15000), .ZN(n7880) );
  INV_X1 U10231 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8454) );
  OAI21_X1 U10232 ( .B1(n13064), .B2(n7411), .A(n8454), .ZN(n7884) );
  AND2_X1 U10233 ( .A1(n7885), .A2(n7884), .ZN(n14758) );
  MUX2_X1 U10234 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14758), .S(n8999), .Z(n15141)
         );
  NAND2_X1 U10235 ( .A1(n14107), .A2(n14101), .ZN(n7886) );
  NAND2_X1 U10236 ( .A1(n14077), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7890) );
  INV_X1 U10237 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9017) );
  INV_X1 U10238 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9006) );
  INV_X1 U10239 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14352) );
  INV_X1 U10240 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14736) );
  NOR2_X1 U10241 ( .A1(n7891), .A2(n14736), .ZN(n7892) );
  MUX2_X1 U10242 ( .A(n14736), .B(n7892), .S(P1_IR_REG_2__SCAN_IN), .Z(n7893)
         );
  INV_X1 U10243 ( .A(n7893), .ZN(n7895) );
  NAND2_X1 U10244 ( .A1(n7895), .A2(n7894), .ZN(n14351) );
  NAND2_X1 U10245 ( .A1(n14077), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7901) );
  OR2_X1 U10246 ( .A1(n8255), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7900) );
  INV_X1 U10247 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10100) );
  INV_X1 U10248 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9020) );
  OR2_X1 U10249 ( .A1(n14081), .A2(n9020), .ZN(n7898) );
  NAND2_X1 U10250 ( .A1(n7894), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7903) );
  XNOR2_X1 U10251 ( .A(n7903), .B(n7902), .ZN(n14368) );
  XNOR2_X1 U10252 ( .A(n7905), .B(n7904), .ZN(n9781) );
  OR2_X1 U10253 ( .A1(n7896), .A2(n9056), .ZN(n7906) );
  NAND2_X1 U10254 ( .A1(n7206), .A2(n14116), .ZN(n7907) );
  XNOR2_X1 U10255 ( .A(n7909), .B(n7908), .ZN(n9950) );
  NAND2_X1 U10256 ( .A1(n9950), .A2(n14087), .ZN(n7916) );
  INV_X2 U10257 ( .A(n8999), .ZN(n8171) );
  OR2_X1 U10258 ( .A1(n7894), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U10259 ( .A1(n7911), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7910) );
  MUX2_X1 U10260 ( .A(n7910), .B(P1_IR_REG_31__SCAN_IN), .S(n7912), .Z(n7914)
         );
  INV_X1 U10261 ( .A(n7911), .ZN(n7913) );
  NAND2_X1 U10262 ( .A1(n7913), .A2(n7912), .ZN(n7927) );
  NAND2_X1 U10263 ( .A1(n7914), .A2(n7927), .ZN(n9116) );
  INV_X1 U10264 ( .A(n9116), .ZN(n9113) );
  INV_X1 U10265 ( .A(n15147), .ZN(n14124) );
  NAND2_X1 U10266 ( .A1(n14077), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7921) );
  INV_X1 U10267 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7917) );
  OR2_X1 U10268 ( .A1(n14081), .A2(n7917), .ZN(n7920) );
  OAI21_X1 U10269 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n7935), .ZN(n10054) );
  OR2_X1 U10270 ( .A1(n8255), .A2(n10054), .ZN(n7919) );
  INV_X1 U10271 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9763) );
  OR2_X1 U10272 ( .A1(n8267), .A2(n9763), .ZN(n7918) );
  AND2_X1 U10273 ( .A1(n14124), .A2(n14122), .ZN(n7922) );
  OR2_X1 U10274 ( .A1(n14122), .A2(n14124), .ZN(n7923) );
  XNOR2_X1 U10275 ( .A(n7925), .B(n7924), .ZN(n9957) );
  NAND2_X1 U10276 ( .A1(n9957), .A2(n14087), .ZN(n7932) );
  NAND2_X1 U10277 ( .A1(n7927), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7926) );
  MUX2_X1 U10278 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7926), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7930) );
  INV_X1 U10279 ( .A(n7927), .ZN(n7929) );
  NAND2_X1 U10280 ( .A1(n7929), .A2(n7928), .ZN(n7945) );
  AND2_X1 U10281 ( .A1(n7930), .A2(n7945), .ZN(n9138) );
  AOI22_X1 U10282 ( .A1(n14086), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8171), 
        .B2(n9138), .ZN(n7931) );
  NAND2_X1 U10283 ( .A1(n14077), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7940) );
  INV_X1 U10284 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7933) );
  OR2_X1 U10285 ( .A1(n14081), .A2(n7933), .ZN(n7939) );
  AND2_X1 U10286 ( .A1(n7935), .A2(n7934), .ZN(n7936) );
  OR2_X1 U10287 ( .A1(n7936), .A2(n7949), .ZN(n10197) );
  OR2_X1 U10288 ( .A1(n8255), .A2(n10197), .ZN(n7938) );
  INV_X1 U10289 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9935) );
  OR2_X1 U10290 ( .A1(n8267), .A2(n9935), .ZN(n7937) );
  XNOR2_X1 U10291 ( .A(n7944), .B(n7943), .ZN(n9971) );
  NAND2_X1 U10292 ( .A1(n9971), .A2(n14087), .ZN(n7948) );
  NAND2_X1 U10293 ( .A1(n7945), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7946) );
  XNOR2_X1 U10294 ( .A(n7946), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9139) );
  AOI22_X1 U10295 ( .A1(n14086), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8171), 
        .B2(n9139), .ZN(n7947) );
  NAND2_X1 U10296 ( .A1(n7948), .A2(n7947), .ZN(n15160) );
  NAND2_X1 U10297 ( .A1(n14077), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7954) );
  INV_X1 U10298 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9149) );
  OR2_X1 U10299 ( .A1(n14081), .A2(n9149), .ZN(n7953) );
  OR2_X1 U10300 ( .A1(n7949), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10301 ( .A1(n7963), .A2(n7950), .ZN(n10311) );
  OR2_X1 U10302 ( .A1(n8255), .A2(n10311), .ZN(n7952) );
  INV_X1 U10303 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9858) );
  OR2_X1 U10304 ( .A1(n8267), .A2(n9858), .ZN(n7951) );
  NAND4_X1 U10305 ( .A1(n7954), .A2(n7953), .A3(n7952), .A4(n7951), .ZN(n14332) );
  XNOR2_X1 U10306 ( .A(n15160), .B(n14332), .ZN(n14275) );
  INV_X1 U10307 ( .A(n14332), .ZN(n10305) );
  NAND2_X1 U10308 ( .A1(n15160), .A2(n10305), .ZN(n7955) );
  XNOR2_X1 U10309 ( .A(n7957), .B(n7956), .ZN(n9984) );
  NAND2_X1 U10310 ( .A1(n9984), .A2(n14087), .ZN(n7961) );
  NAND2_X1 U10311 ( .A1(n7958), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7959) );
  XNOR2_X1 U10312 ( .A(n7959), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14391) );
  AOI22_X1 U10313 ( .A1(n14086), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8171), 
        .B2(n14391), .ZN(n7960) );
  NAND2_X1 U10314 ( .A1(n7961), .A2(n7960), .ZN(n14135) );
  NAND2_X1 U10315 ( .A1(n8309), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7968) );
  INV_X1 U10316 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7962) );
  OR2_X1 U10317 ( .A1(n8312), .A2(n7962), .ZN(n7967) );
  NAND2_X1 U10318 ( .A1(n7963), .A2(n10538), .ZN(n7964) );
  NAND2_X1 U10319 ( .A1(n7977), .A2(n7964), .ZN(n10539) );
  OR2_X1 U10320 ( .A1(n8255), .A2(n10539), .ZN(n7966) );
  INV_X1 U10321 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9157) );
  OR2_X1 U10322 ( .A1(n8267), .A2(n9157), .ZN(n7965) );
  NAND4_X1 U10323 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n14331) );
  INV_X1 U10324 ( .A(n14331), .ZN(n10533) );
  OR2_X1 U10325 ( .A1(n14135), .A2(n10533), .ZN(n7969) );
  NAND2_X1 U10326 ( .A1(n10089), .A2(n7969), .ZN(n7971) );
  NAND2_X1 U10327 ( .A1(n14135), .A2(n10533), .ZN(n7970) );
  NAND2_X1 U10328 ( .A1(n7971), .A2(n7970), .ZN(n15085) );
  XNOR2_X1 U10329 ( .A(n7973), .B(n7972), .ZN(n9997) );
  NAND2_X1 U10330 ( .A1(n9997), .A2(n14087), .ZN(n7976) );
  NOR2_X1 U10331 ( .A1(n7958), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n7989) );
  OR2_X1 U10332 ( .A1(n7989), .A2(n14736), .ZN(n7974) );
  XNOR2_X1 U10333 ( .A(n7974), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9175) );
  AOI22_X1 U10334 ( .A1(n14086), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8171), 
        .B2(n9175), .ZN(n7975) );
  NAND2_X1 U10335 ( .A1(n14077), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7983) );
  INV_X1 U10336 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9148) );
  OR2_X1 U10337 ( .A1(n14081), .A2(n9148), .ZN(n7982) );
  NAND2_X1 U10338 ( .A1(n7977), .A2(n9154), .ZN(n7978) );
  NAND2_X1 U10339 ( .A1(n7995), .A2(n7978), .ZN(n15090) );
  OR2_X1 U10340 ( .A1(n8255), .A2(n15090), .ZN(n7981) );
  INV_X1 U10341 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7979) );
  OR2_X1 U10342 ( .A1(n8267), .A2(n7979), .ZN(n7980) );
  NAND4_X1 U10343 ( .A1(n7983), .A2(n7982), .A3(n7981), .A4(n7980), .ZN(n14330) );
  XNOR2_X1 U10344 ( .A(n15089), .B(n14330), .ZN(n14278) );
  INV_X1 U10345 ( .A(n14330), .ZN(n7984) );
  OR2_X1 U10346 ( .A1(n15089), .A2(n7984), .ZN(n7985) );
  XNOR2_X1 U10347 ( .A(n7987), .B(n7986), .ZN(n10128) );
  NAND2_X1 U10348 ( .A1(n10128), .A2(n14087), .ZN(n7992) );
  AND2_X1 U10349 ( .A1(n7989), .A2(n7988), .ZN(n8004) );
  OR2_X1 U10350 ( .A1(n8004), .A2(n14736), .ZN(n7990) );
  XNOR2_X1 U10351 ( .A(n7990), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9188) );
  AOI22_X1 U10352 ( .A1(n14086), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8171), 
        .B2(n9188), .ZN(n7991) );
  NAND2_X1 U10353 ( .A1(n14077), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8001) );
  INV_X1 U10354 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7993) );
  OR2_X1 U10355 ( .A1(n14081), .A2(n7993), .ZN(n8000) );
  INV_X1 U10356 ( .A(n8009), .ZN(n7997) );
  NAND2_X1 U10357 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  NAND2_X1 U10358 ( .A1(n7997), .A2(n7996), .ZN(n15072) );
  OR2_X1 U10359 ( .A1(n8255), .A2(n15072), .ZN(n7999) );
  INV_X1 U10360 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9167) );
  OR2_X1 U10361 ( .A1(n8267), .A2(n9167), .ZN(n7998) );
  NAND4_X1 U10362 ( .A1(n8001), .A2(n8000), .A3(n7999), .A4(n7998), .ZN(n14329) );
  XNOR2_X1 U10363 ( .A(n15076), .B(n10879), .ZN(n14280) );
  INV_X1 U10364 ( .A(n14280), .ZN(n15066) );
  NAND2_X1 U10365 ( .A1(n15076), .A2(n10879), .ZN(n8002) );
  XNOR2_X1 U10366 ( .A(n8018), .B(n8019), .ZN(n10376) );
  NAND2_X1 U10367 ( .A1(n10376), .A2(n14087), .ZN(n8007) );
  NAND2_X1 U10368 ( .A1(n8004), .A2(n8003), .ZN(n8028) );
  NAND2_X1 U10369 ( .A1(n8028), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8005) );
  XNOR2_X1 U10370 ( .A(n8005), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9408) );
  AOI22_X1 U10371 ( .A1(n14086), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8171), 
        .B2(n9408), .ZN(n8006) );
  NAND2_X1 U10372 ( .A1(n8309), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8014) );
  INV_X1 U10373 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8008) );
  OR2_X1 U10374 ( .A1(n8312), .A2(n8008), .ZN(n8013) );
  OR2_X1 U10375 ( .A1(n8009), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U10376 ( .A1(n8031), .A2(n8010), .ZN(n15054) );
  OR2_X1 U10377 ( .A1(n8255), .A2(n15054), .ZN(n8012) );
  INV_X1 U10378 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9403) );
  OR2_X1 U10379 ( .A1(n8267), .A2(n9403), .ZN(n8011) );
  NAND4_X1 U10380 ( .A1(n8014), .A2(n8013), .A3(n8012), .A4(n8011), .ZN(n14328) );
  INV_X1 U10381 ( .A(n14328), .ZN(n8015) );
  OR2_X1 U10382 ( .A1(n15188), .A2(n8015), .ZN(n8017) );
  NAND2_X1 U10383 ( .A1(n15188), .A2(n8015), .ZN(n8016) );
  NAND2_X1 U10384 ( .A1(n8017), .A2(n8016), .ZN(n15056) );
  INV_X1 U10385 ( .A(n8018), .ZN(n8020) );
  NAND2_X1 U10386 ( .A1(n8020), .A2(n8019), .ZN(n8023) );
  NAND2_X1 U10387 ( .A1(n8021), .A2(SI_10_), .ZN(n8022) );
  NAND2_X1 U10388 ( .A1(n8023), .A2(n8022), .ZN(n8027) );
  NAND2_X1 U10389 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  NAND2_X1 U10390 ( .A1(n8100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8044) );
  XNOR2_X1 U10391 ( .A(n8044), .B(P1_IR_REG_11__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U10392 ( .A1(n14086), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8171), 
        .B2(n14406), .ZN(n8029) );
  NAND2_X1 U10393 ( .A1(n14077), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10394 ( .A1(n8031), .A2(n8030), .ZN(n8032) );
  NAND2_X1 U10395 ( .A1(n8049), .A2(n8032), .ZN(n14932) );
  OR2_X1 U10396 ( .A1(n8255), .A2(n14932), .ZN(n8036) );
  INV_X1 U10397 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9404) );
  OR2_X1 U10398 ( .A1(n8267), .A2(n9404), .ZN(n8035) );
  INV_X1 U10399 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8033) );
  OR2_X1 U10400 ( .A1(n14081), .A2(n8033), .ZN(n8034) );
  NAND4_X1 U10401 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), .ZN(n15058) );
  NAND2_X1 U10402 ( .A1(n14927), .A2(n14284), .ZN(n14930) );
  INV_X1 U10403 ( .A(n15058), .ZN(n11268) );
  OR2_X1 U10404 ( .A1(n14934), .A2(n11268), .ZN(n8038) );
  OR2_X1 U10405 ( .A1(n8040), .A2(n8039), .ZN(n8041) );
  NAND2_X1 U10406 ( .A1(n8042), .A2(n8041), .ZN(n10566) );
  NAND2_X1 U10407 ( .A1(n10566), .A2(n14087), .ZN(n8047) );
  INV_X1 U10408 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U10409 ( .A1(n8044), .A2(n8043), .ZN(n8045) );
  NAND2_X1 U10410 ( .A1(n8045), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8060) );
  XNOR2_X1 U10411 ( .A(n8060), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9413) );
  AOI22_X1 U10412 ( .A1(n14086), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9413), 
        .B2(n8171), .ZN(n8046) );
  NAND2_X1 U10413 ( .A1(n14077), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8055) );
  INV_X1 U10414 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10763) );
  OR2_X1 U10415 ( .A1(n8267), .A2(n10763), .ZN(n8054) );
  INV_X1 U10416 ( .A(n8065), .ZN(n8051) );
  NAND2_X1 U10417 ( .A1(n8049), .A2(n8048), .ZN(n8050) );
  NAND2_X1 U10418 ( .A1(n8051), .A2(n8050), .ZN(n11299) );
  OR2_X1 U10419 ( .A1(n8255), .A2(n11299), .ZN(n8053) );
  INV_X1 U10420 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9409) );
  OR2_X1 U10421 ( .A1(n14081), .A2(n9409), .ZN(n8052) );
  NAND4_X1 U10422 ( .A1(n8055), .A2(n8054), .A3(n8053), .A4(n8052), .ZN(n14327) );
  INV_X1 U10423 ( .A(n14327), .ZN(n8056) );
  XNOR2_X1 U10424 ( .A(n14885), .B(n8056), .ZN(n14281) );
  OR2_X1 U10425 ( .A1(n14885), .A2(n8056), .ZN(n8057) );
  XNOR2_X1 U10426 ( .A(n8058), .B(n7692), .ZN(n10818) );
  NAND2_X1 U10427 ( .A1(n10818), .A2(n14087), .ZN(n8064) );
  INV_X1 U10428 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10429 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  NAND2_X1 U10430 ( .A1(n8061), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8075) );
  INV_X1 U10431 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8074) );
  XNOR2_X1 U10432 ( .A(n8075), .B(n8074), .ZN(n15009) );
  OAI22_X1 U10433 ( .A1(n15009), .A2(n8999), .B1(n7896), .B2(n9501), .ZN(n8062) );
  INV_X1 U10434 ( .A(n8062), .ZN(n8063) );
  NOR2_X1 U10435 ( .A1(n8065), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8066) );
  OR2_X1 U10436 ( .A1(n8080), .A2(n8066), .ZN(n11314) );
  OR2_X1 U10437 ( .A1(n11314), .A2(n8255), .ZN(n8071) );
  INV_X1 U10438 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9557) );
  OR2_X1 U10439 ( .A1(n14081), .A2(n9557), .ZN(n8070) );
  INV_X1 U10440 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8067) );
  OR2_X1 U10441 ( .A1(n8312), .A2(n8067), .ZN(n8069) );
  INV_X1 U10442 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9562) );
  OR2_X1 U10443 ( .A1(n8267), .A2(n9562), .ZN(n8068) );
  NAND4_X1 U10444 ( .A1(n8071), .A2(n8070), .A3(n8069), .A4(n8068), .ZN(n14326) );
  XNOR2_X1 U10445 ( .A(n14961), .B(n13926), .ZN(n14283) );
  INV_X1 U10446 ( .A(n14283), .ZN(n11026) );
  OR2_X1 U10447 ( .A1(n14961), .A2(n13926), .ZN(n8072) );
  XNOR2_X1 U10448 ( .A(n8091), .B(SI_14_), .ZN(n8090) );
  XNOR2_X1 U10449 ( .A(n8090), .B(n8073), .ZN(n10899) );
  NAND2_X1 U10450 ( .A1(n10899), .A2(n14087), .ZN(n8079) );
  NAND2_X1 U10451 ( .A1(n8075), .A2(n8074), .ZN(n8076) );
  NAND2_X1 U10452 ( .A1(n8076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8077) );
  XNOR2_X1 U10453 ( .A(n8077), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9563) );
  AOI22_X1 U10454 ( .A1(n9563), .A2(n8171), .B1(n14086), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8078) );
  INV_X1 U10455 ( .A(n8255), .ZN(n8179) );
  OR2_X1 U10456 ( .A1(n8080), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8081) );
  AND2_X1 U10457 ( .A1(n8109), .A2(n8081), .ZN(n13922) );
  NAND2_X1 U10458 ( .A1(n8179), .A2(n13922), .ZN(n8087) );
  INV_X1 U10459 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8082) );
  OR2_X1 U10460 ( .A1(n14081), .A2(n8082), .ZN(n8086) );
  INV_X1 U10461 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8083) );
  OR2_X1 U10462 ( .A1(n8312), .A2(n8083), .ZN(n8085) );
  INV_X1 U10463 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9564) );
  OR2_X1 U10464 ( .A1(n8267), .A2(n9564), .ZN(n8084) );
  OR2_X1 U10465 ( .A1(n14952), .A2(n11683), .ZN(n14165) );
  NAND2_X1 U10466 ( .A1(n14952), .A2(n11683), .ZN(n14166) );
  NAND2_X1 U10467 ( .A1(n8088), .A2(n14166), .ZN(n11211) );
  NAND2_X1 U10468 ( .A1(n8090), .A2(n8089), .ZN(n8094) );
  INV_X1 U10469 ( .A(n8091), .ZN(n8092) );
  NAND2_X1 U10470 ( .A1(n8092), .A2(SI_14_), .ZN(n8093) );
  NAND2_X1 U10471 ( .A1(n8094), .A2(n8093), .ZN(n8099) );
  INV_X1 U10472 ( .A(n8095), .ZN(n8096) );
  NAND2_X1 U10473 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  NAND2_X1 U10474 ( .A1(n11001), .A2(n14087), .ZN(n8107) );
  INV_X1 U10475 ( .A(n8100), .ZN(n8104) );
  NOR2_X1 U10476 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n8101) );
  AND2_X1 U10477 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  NAND2_X1 U10478 ( .A1(n8104), .A2(n8103), .ZN(n8118) );
  NAND2_X1 U10479 ( .A1(n8118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8105) );
  XNOR2_X1 U10480 ( .A(n8105), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U10481 ( .A1(n14086), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10327), 
        .B2(n8171), .ZN(n8106) );
  NAND2_X1 U10482 ( .A1(n8109), .A2(n8108), .ZN(n8110) );
  AND2_X1 U10483 ( .A1(n8128), .A2(n8110), .ZN(n14072) );
  NAND2_X1 U10484 ( .A1(n14072), .A2(n8179), .ZN(n8115) );
  NAND2_X1 U10485 ( .A1(n14077), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8114) );
  INV_X1 U10486 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11207) );
  OR2_X1 U10487 ( .A1(n8267), .A2(n11207), .ZN(n8113) );
  INV_X1 U10488 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8111) );
  OR2_X1 U10489 ( .A1(n14081), .A2(n8111), .ZN(n8112) );
  NAND2_X1 U10490 ( .A1(n14944), .A2(n11690), .ZN(n14174) );
  NAND2_X1 U10491 ( .A1(n14173), .A2(n14174), .ZN(n14288) );
  XNOR2_X1 U10492 ( .A(n8117), .B(n8116), .ZN(n11354) );
  NAND2_X1 U10493 ( .A1(n11354), .A2(n14087), .ZN(n8126) );
  NAND2_X1 U10494 ( .A1(n8120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8119) );
  MUX2_X1 U10495 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8119), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8123) );
  INV_X1 U10496 ( .A(n8120), .ZN(n8122) );
  INV_X1 U10497 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U10498 ( .A1(n8122), .A2(n8121), .ZN(n8137) );
  NAND2_X1 U10499 ( .A1(n8123), .A2(n8137), .ZN(n10488) );
  OAI22_X1 U10500 ( .A1(n10488), .A2(n8999), .B1(n7896), .B2(n13776), .ZN(
        n8124) );
  INV_X1 U10501 ( .A(n8124), .ZN(n8125) );
  AND2_X1 U10502 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  OR2_X1 U10503 ( .A1(n8129), .A2(n8144), .ZN(n13992) );
  AOI22_X1 U10504 ( .A1(n8309), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n14077), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n8131) );
  NAND2_X1 U10505 ( .A1(n14076), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8130) );
  OAI211_X1 U10506 ( .C1(n13992), .C2(n8255), .A(n8131), .B(n8130), .ZN(n14323) );
  XNOR2_X1 U10507 ( .A(n14714), .B(n14323), .ZN(n14285) );
  INV_X1 U10508 ( .A(n14323), .ZN(n14607) );
  NAND2_X1 U10509 ( .A1(n14714), .A2(n14607), .ZN(n8132) );
  XNOR2_X1 U10510 ( .A(n8134), .B(n9512), .ZN(n8135) );
  XNOR2_X1 U10511 ( .A(n8136), .B(n8135), .ZN(n11358) );
  NAND2_X1 U10512 ( .A1(n11358), .A2(n14087), .ZN(n8143) );
  NAND2_X1 U10513 ( .A1(n8137), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8138) );
  MUX2_X1 U10514 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8138), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8141) );
  AND2_X1 U10515 ( .A1(n8141), .A2(n8140), .ZN(n10957) );
  AOI22_X1 U10516 ( .A1(n10957), .A2(n8171), .B1(n14086), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n8142) );
  OR2_X1 U10517 ( .A1(n8144), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10518 ( .A1(n8158), .A2(n8145), .ZN(n14619) );
  AOI22_X1 U10519 ( .A1(n8309), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n14077), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U10520 ( .A1(n14076), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8146) );
  OAI211_X1 U10521 ( .C1(n14619), .C2(n8255), .A(n8147), .B(n8146), .ZN(n14322) );
  NOR2_X1 U10522 ( .A1(n14710), .A2(n14322), .ZN(n14195) );
  INV_X1 U10523 ( .A(n14195), .ZN(n8148) );
  NAND2_X1 U10524 ( .A1(n14710), .A2(n14322), .ZN(n14196) );
  NAND2_X1 U10525 ( .A1(n8148), .A2(n14196), .ZN(n14602) );
  INV_X1 U10526 ( .A(n14602), .ZN(n14604) );
  INV_X1 U10527 ( .A(n14322), .ZN(n13994) );
  OR2_X1 U10528 ( .A1(n14710), .A2(n13994), .ZN(n8149) );
  NAND2_X1 U10529 ( .A1(n8151), .A2(n8150), .ZN(n8152) );
  NAND2_X1 U10530 ( .A1(n8153), .A2(n8152), .ZN(n11369) );
  OR2_X1 U10531 ( .A1(n11369), .A2(n14242), .ZN(n8156) );
  NAND2_X1 U10532 ( .A1(n8140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8154) );
  XNOR2_X1 U10533 ( .A(n8154), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U10534 ( .A1(n14086), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8171), 
        .B2(n15037), .ZN(n8155) );
  NAND2_X1 U10535 ( .A1(n8158), .A2(n8157), .ZN(n8159) );
  NAND2_X1 U10536 ( .A1(n8174), .A2(n8159), .ZN(n14045) );
  OR2_X1 U10537 ( .A1(n14045), .A2(n8255), .ZN(n8166) );
  INV_X1 U10538 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U10539 ( .A1(n14077), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8162) );
  INV_X1 U10540 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8160) );
  OR2_X1 U10541 ( .A1(n8267), .A2(n8160), .ZN(n8161) );
  OAI211_X1 U10542 ( .C1(n14081), .C2(n8163), .A(n8162), .B(n8161), .ZN(n8164)
         );
  INV_X1 U10543 ( .A(n8164), .ZN(n8165) );
  XNOR2_X1 U10544 ( .A(n14705), .B(n14609), .ZN(n14591) );
  INV_X1 U10545 ( .A(n14591), .ZN(n8168) );
  INV_X1 U10546 ( .A(n14609), .ZN(n14321) );
  AND2_X1 U10547 ( .A1(n14198), .A2(n14321), .ZN(n8167) );
  XNOR2_X1 U10548 ( .A(n8170), .B(n8169), .ZN(n11380) );
  NAND2_X1 U10549 ( .A1(n11380), .A2(n14087), .ZN(n8173) );
  AOI22_X1 U10550 ( .A1(n14086), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14598), 
        .B2(n8171), .ZN(n8172) );
  AND2_X1 U10551 ( .A1(n8174), .A2(n13810), .ZN(n8175) );
  OR2_X1 U10552 ( .A1(n8175), .A2(n8186), .ZN(n14578) );
  INV_X1 U10553 ( .A(n14578), .ZN(n13957) );
  INV_X1 U10554 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10954) );
  NAND2_X1 U10555 ( .A1(n14077), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8177) );
  NAND2_X1 U10556 ( .A1(n14076), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8176) );
  OAI211_X1 U10557 ( .C1(n10954), .C2(n14081), .A(n8177), .B(n8176), .ZN(n8178) );
  AOI21_X1 U10558 ( .B1(n13957), .B2(n8179), .A(n8178), .ZN(n11712) );
  OR2_X1 U10559 ( .A1(n14581), .A2(n11712), .ZN(n14202) );
  NAND2_X1 U10560 ( .A1(n14581), .A2(n11712), .ZN(n14203) );
  NAND2_X1 U10561 ( .A1(n14202), .A2(n14203), .ZN(n14291) );
  INV_X1 U10562 ( .A(n14291), .ZN(n14572) );
  NAND2_X1 U10563 ( .A1(n14573), .A2(n14572), .ZN(n14571) );
  NAND2_X1 U10564 ( .A1(n14571), .A2(n14203), .ZN(n14550) );
  INV_X1 U10565 ( .A(n14550), .ZN(n8193) );
  NAND2_X1 U10566 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  NAND2_X1 U10567 ( .A1(n8183), .A2(n8182), .ZN(n11393) );
  OR2_X1 U10568 ( .A1(n11393), .A2(n14242), .ZN(n8185) );
  OR2_X1 U10569 ( .A1(n7896), .A2(n10498), .ZN(n8184) );
  OR2_X1 U10570 ( .A1(n8186), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U10571 ( .A1(n8201), .A2(n8187), .ZN(n14559) );
  OR2_X1 U10572 ( .A1(n14559), .A2(n8255), .ZN(n8192) );
  INV_X1 U10573 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14694) );
  NAND2_X1 U10574 ( .A1(n14077), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10575 ( .A1(n14076), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8188) );
  OAI211_X1 U10576 ( .C1(n14081), .C2(n14694), .A(n8189), .B(n8188), .ZN(n8190) );
  INV_X1 U10577 ( .A(n8190), .ZN(n8191) );
  NAND2_X1 U10578 ( .A1(n8192), .A2(n8191), .ZN(n14577) );
  XNOR2_X1 U10579 ( .A(n14688), .B(n14577), .ZN(n14565) );
  INV_X1 U10580 ( .A(n14565), .ZN(n14549) );
  INV_X1 U10581 ( .A(n14688), .ZN(n8315) );
  NAND2_X1 U10582 ( .A1(n8315), .A2(n14577), .ZN(n8194) );
  OR2_X1 U10583 ( .A1(n8196), .A2(n8195), .ZN(n8197) );
  AND2_X1 U10584 ( .A1(n8198), .A2(n8197), .ZN(n11407) );
  NAND2_X1 U10585 ( .A1(n11407), .A2(n14087), .ZN(n8200) );
  INV_X1 U10586 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10716) );
  OR2_X1 U10587 ( .A1(n7896), .A2(n10716), .ZN(n8199) );
  NAND2_X1 U10588 ( .A1(n8201), .A2(n13973), .ZN(n8203) );
  INV_X1 U10589 ( .A(n8214), .ZN(n8202) );
  NAND2_X1 U10590 ( .A1(n8203), .A2(n8202), .ZN(n14538) );
  OR2_X1 U10591 ( .A1(n14538), .A2(n8255), .ZN(n8208) );
  INV_X1 U10592 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n13783) );
  NAND2_X1 U10593 ( .A1(n8309), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8205) );
  NAND2_X1 U10594 ( .A1(n14076), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8204) );
  OAI211_X1 U10595 ( .C1(n8312), .C2(n13783), .A(n8205), .B(n8204), .ZN(n8206)
         );
  INV_X1 U10596 ( .A(n8206), .ZN(n8207) );
  NAND2_X1 U10597 ( .A1(n8208), .A2(n8207), .ZN(n14553) );
  XNOR2_X1 U10598 ( .A(n14682), .B(n14553), .ZN(n14545) );
  INV_X1 U10599 ( .A(n14553), .ZN(n8209) );
  OR2_X1 U10600 ( .A1(n14682), .A2(n8209), .ZN(n8210) );
  OR2_X1 U10601 ( .A1(n11156), .A2(n13064), .ZN(n8211) );
  NAND2_X1 U10602 ( .A1(n8309), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8219) );
  INV_X1 U10603 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8212) );
  OR2_X1 U10604 ( .A1(n8312), .A2(n8212), .ZN(n8218) );
  OAI21_X1 U10605 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n8214), .A(n8213), .ZN(
        n14036) );
  OR2_X1 U10606 ( .A1(n8255), .A2(n14036), .ZN(n8217) );
  INV_X1 U10607 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8215) );
  OR2_X1 U10608 ( .A1(n8267), .A2(n8215), .ZN(n8216) );
  INV_X1 U10609 ( .A(n14676), .ZN(n14528) );
  NAND2_X1 U10610 ( .A1(n14528), .A2(n14216), .ZN(n8220) );
  XNOR2_X1 U10611 ( .A(n8221), .B(SI_23_), .ZN(n8222) );
  XNOR2_X1 U10612 ( .A(n8223), .B(n8222), .ZN(n11433) );
  NAND2_X1 U10613 ( .A1(n11433), .A2(n14087), .ZN(n8225) );
  INV_X1 U10614 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11178) );
  OR2_X1 U10615 ( .A1(n7896), .A2(n11178), .ZN(n8224) );
  NAND2_X1 U10616 ( .A1(n14077), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8233) );
  INV_X1 U10617 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8226) );
  OR2_X1 U10618 ( .A1(n14081), .A2(n8226), .ZN(n8232) );
  OAI21_X1 U10619 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8228), .A(n8227), .ZN(
        n14516) );
  OR2_X1 U10620 ( .A1(n8255), .A2(n14516), .ZN(n8231) );
  INV_X1 U10621 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n8229) );
  OR2_X1 U10622 ( .A1(n8267), .A2(n8229), .ZN(n8230) );
  NAND4_X1 U10623 ( .A1(n8233), .A2(n8232), .A3(n8231), .A4(n8230), .ZN(n14320) );
  XNOR2_X1 U10624 ( .A(n14668), .B(n14320), .ZN(n14509) );
  INV_X1 U10625 ( .A(n14668), .ZN(n8300) );
  INV_X1 U10626 ( .A(n14512), .ZN(n14476) );
  XNOR2_X1 U10627 ( .A(n14659), .B(n14319), .ZN(n14471) );
  NAND2_X1 U10628 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  NAND2_X1 U10629 ( .A1(n13898), .A2(n14087), .ZN(n8239) );
  INV_X1 U10630 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14750) );
  OR2_X1 U10631 ( .A1(n7896), .A2(n14750), .ZN(n8238) );
  NAND2_X1 U10632 ( .A1(n14076), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8246) );
  INV_X1 U10633 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n13761) );
  OR2_X1 U10634 ( .A1(n8312), .A2(n13761), .ZN(n8245) );
  OAI21_X1 U10635 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n8241), .A(n8240), .ZN(
        n14460) );
  OR2_X1 U10636 ( .A1(n8255), .A2(n14460), .ZN(n8244) );
  INV_X1 U10637 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8242) );
  OR2_X1 U10638 ( .A1(n14081), .A2(n8242), .ZN(n8243) );
  NAND2_X1 U10639 ( .A1(n14652), .A2(n8247), .ZN(n8248) );
  XNOR2_X1 U10640 ( .A(n8249), .B(SI_27_), .ZN(n8250) );
  NAND2_X1 U10641 ( .A1(n13894), .A2(n14087), .ZN(n8252) );
  OR2_X1 U10642 ( .A1(n7896), .A2(n11329), .ZN(n8251) );
  NAND2_X1 U10643 ( .A1(n8309), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8260) );
  INV_X1 U10644 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8253) );
  OR2_X1 U10645 ( .A1(n8312), .A2(n8253), .ZN(n8259) );
  XNOR2_X1 U10646 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n8254), .ZN(n13915) );
  INV_X1 U10647 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8256) );
  OR2_X1 U10648 ( .A1(n8267), .A2(n8256), .ZN(n8257) );
  INV_X1 U10649 ( .A(n14317), .ZN(n8302) );
  INV_X1 U10650 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14745) );
  INV_X1 U10651 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13886) );
  MUX2_X1 U10652 ( .A(n14745), .B(n13886), .S(n13064), .Z(n13056) );
  XNOR2_X1 U10653 ( .A(n13056), .B(SI_29_), .ZN(n13059) );
  NAND2_X1 U10654 ( .A1(n13885), .A2(n14087), .ZN(n8265) );
  OR2_X1 U10655 ( .A1(n7896), .A2(n14745), .ZN(n8264) );
  NAND2_X1 U10656 ( .A1(n8309), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U10657 ( .A1(n14077), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8270) );
  OR2_X1 U10658 ( .A1(n8255), .A2(n14430), .ZN(n8269) );
  INV_X1 U10659 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8266) );
  OR2_X1 U10660 ( .A1(n8267), .A2(n8266), .ZN(n8268) );
  NAND4_X1 U10661 ( .A1(n8271), .A2(n8270), .A3(n8269), .A4(n8268), .ZN(n14315) );
  INV_X1 U10662 ( .A(n14315), .ZN(n8272) );
  XNOR2_X1 U10663 ( .A(n8273), .B(n14299), .ZN(n8275) );
  NAND2_X1 U10664 ( .A1(n14756), .A2(n14598), .ZN(n8274) );
  INV_X1 U10665 ( .A(n14085), .ZN(n8307) );
  NAND2_X1 U10666 ( .A1(n14084), .A2(n8307), .ZN(n14245) );
  INV_X1 U10667 ( .A(n14319), .ZN(n14489) );
  INV_X1 U10668 ( .A(n14320), .ZN(n14490) );
  INV_X1 U10669 ( .A(n15141), .ZN(n14099) );
  NOR2_X1 U10670 ( .A1(n8991), .A2(n14099), .ZN(n9619) );
  INV_X1 U10671 ( .A(n14336), .ZN(n14110) );
  NAND2_X1 U10672 ( .A1(n14110), .A2(n9725), .ZN(n8277) );
  NAND2_X1 U10673 ( .A1(n7206), .A2(n14117), .ZN(n8278) );
  INV_X1 U10674 ( .A(n14275), .ZN(n8279) );
  NAND2_X1 U10675 ( .A1(n9852), .A2(n8279), .ZN(n8281) );
  OR2_X1 U10676 ( .A1(n15160), .A2(n14332), .ZN(n8280) );
  XNOR2_X1 U10677 ( .A(n14135), .B(n14331), .ZN(n14276) );
  INV_X1 U10678 ( .A(n14276), .ZN(n10093) );
  OR2_X1 U10679 ( .A1(n14135), .A2(n14331), .ZN(n8282) );
  NAND2_X1 U10680 ( .A1(n15067), .A2(n14280), .ZN(n8284) );
  OR2_X1 U10681 ( .A1(n15076), .A2(n14329), .ZN(n8283) );
  OR2_X1 U10682 ( .A1(n15188), .A2(n14328), .ZN(n8285) );
  OR2_X1 U10683 ( .A1(n14934), .A2(n15058), .ZN(n8287) );
  OR2_X1 U10684 ( .A1(n14885), .A2(n14327), .ZN(n8288) );
  NAND2_X1 U10685 ( .A1(n8289), .A2(n8288), .ZN(n11024) );
  NAND2_X1 U10686 ( .A1(n11024), .A2(n14283), .ZN(n8291) );
  OR2_X1 U10687 ( .A1(n14961), .A2(n14326), .ZN(n8290) );
  XNOR2_X1 U10688 ( .A(n14952), .B(n11683), .ZN(n14289) );
  INV_X1 U10689 ( .A(n14289), .ZN(n10979) );
  INV_X1 U10690 ( .A(n11683), .ZN(n14325) );
  NAND2_X1 U10691 ( .A1(n14952), .A2(n14325), .ZN(n8292) );
  OR2_X1 U10692 ( .A1(n14944), .A2(n14324), .ZN(n8293) );
  AND2_X1 U10693 ( .A1(n14705), .A2(n14321), .ZN(n14201) );
  OR2_X1 U10694 ( .A1(n14705), .A2(n14321), .ZN(n14200) );
  NAND2_X1 U10695 ( .A1(n14570), .A2(n14291), .ZN(n8295) );
  INV_X1 U10696 ( .A(n11712), .ZN(n14555) );
  OR2_X1 U10697 ( .A1(n14581), .A2(n14555), .ZN(n8294) );
  NAND2_X1 U10698 ( .A1(n8295), .A2(n8294), .ZN(n14566) );
  NAND2_X1 U10699 ( .A1(n14688), .A2(n14577), .ZN(n8296) );
  OR2_X1 U10700 ( .A1(n14682), .A2(n14553), .ZN(n8297) );
  NAND2_X1 U10701 ( .A1(n14676), .A2(n14216), .ZN(n8298) );
  INV_X1 U10702 ( .A(n14471), .ZN(n14468) );
  XNOR2_X1 U10703 ( .A(n14652), .B(n14318), .ZN(n14455) );
  INV_X1 U10704 ( .A(n14455), .ZN(n14453) );
  NAND2_X1 U10705 ( .A1(n14639), .A2(n14316), .ZN(n8304) );
  NAND2_X1 U10706 ( .A1(n8304), .A2(n8303), .ZN(n14295) );
  AND2_X1 U10707 ( .A1(n14092), .A2(n14617), .ZN(n8305) );
  NAND2_X1 U10708 ( .A1(n14756), .A2(n14617), .ZN(n14083) );
  NAND2_X2 U10709 ( .A1(n14083), .A2(n14103), .ZN(n11795) );
  NAND2_X1 U10710 ( .A1(n8305), .A2(n11795), .ZN(n15068) );
  OR2_X1 U10711 ( .A1(n14091), .A2(n14617), .ZN(n15163) );
  INV_X1 U10712 ( .A(n14084), .ZN(n15140) );
  AND2_X1 U10713 ( .A1(n15140), .A2(n8307), .ZN(n14302) );
  NAND2_X1 U10714 ( .A1(n8306), .A2(n14302), .ZN(n15092) );
  NAND3_X1 U10715 ( .A1(n8306), .A2(n14598), .A3(n15140), .ZN(n8308) );
  INV_X1 U10716 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n13606) );
  NAND2_X1 U10717 ( .A1(n14076), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8311) );
  NAND2_X1 U10718 ( .A1(n8309), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8310) );
  OAI211_X1 U10719 ( .C1(n8312), .C2(n13606), .A(n8311), .B(n8310), .ZN(n14314) );
  INV_X1 U10720 ( .A(n11338), .ZN(n9012) );
  OR2_X1 U10721 ( .A1(n14092), .A2(n9012), .ZN(n14608) );
  INV_X1 U10722 ( .A(P1_B_REG_SCAN_IN), .ZN(n8313) );
  NOR2_X1 U10723 ( .A1(n6560), .A2(n8313), .ZN(n8314) );
  NOR2_X1 U10724 ( .A1(n14608), .A2(n8314), .ZN(n14417) );
  NAND2_X1 U10725 ( .A1(n9723), .A2(n14117), .ZN(n9767) );
  INV_X1 U10726 ( .A(n15160), .ZN(n10317) );
  INV_X1 U10727 ( .A(n14135), .ZN(n15171) );
  INV_X1 U10728 ( .A(n14952), .ZN(n10976) );
  NAND2_X1 U10729 ( .A1(n11029), .A2(n10976), .ZN(n11202) );
  NAND2_X1 U10730 ( .A1(n8315), .A2(n14575), .ZN(n14562) );
  INV_X1 U10731 ( .A(n14253), .ZN(n14432) );
  OAI21_X1 U10732 ( .B1(n8316), .B2(n14432), .A(n8988), .ZN(n8317) );
  NAND2_X1 U10733 ( .A1(n14637), .A2(n15197), .ZN(n8318) );
  NAND2_X1 U10734 ( .A1(n8319), .A2(n8318), .ZN(P1_U3525) );
  NAND4_X1 U10735 ( .A1(n8322), .A2(n8321), .A3(n8320), .A4(n13831), .ZN(n8323) );
  INV_X1 U10736 ( .A(n8686), .ZN(n8329) );
  INV_X1 U10737 ( .A(n8408), .ZN(n8339) );
  NAND2_X1 U10738 ( .A1(n8339), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U10739 ( .A1(n8334), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8335) );
  MUX2_X1 U10740 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8335), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8336) );
  NAND2_X1 U10741 ( .A1(n8336), .A2(n6601), .ZN(n9716) );
  NAND2_X1 U10742 ( .A1(n12163), .A2(n9716), .ZN(n8337) );
  NAND2_X1 U10743 ( .A1(n12268), .A2(n8337), .ZN(n8341) );
  NAND2_X1 U10744 ( .A1(n6601), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8338) );
  MUX2_X1 U10745 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8338), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8340) );
  NAND2_X1 U10746 ( .A1(n8341), .A2(n11990), .ZN(n8343) );
  INV_X1 U10747 ( .A(n9716), .ZN(n8933) );
  OAI21_X1 U10748 ( .B1(n8933), .B2(n8876), .A(n8925), .ZN(n8342) );
  NAND2_X1 U10749 ( .A1(n8343), .A2(n8342), .ZN(n9736) );
  NAND2_X1 U10750 ( .A1(n9736), .A2(n15515), .ZN(n9838) );
  INV_X1 U10751 ( .A(n12268), .ZN(n9680) );
  NAND2_X1 U10752 ( .A1(n9680), .A2(n9716), .ZN(n12152) );
  OR2_X1 U10753 ( .A1(n9838), .A2(n12152), .ZN(n8344) );
  OR3_X1 U10754 ( .A1(n12268), .A2(n8925), .A3(n9716), .ZN(n8924) );
  OR2_X1 U10755 ( .A1(n12151), .A2(n12163), .ZN(n15497) );
  AND2_X1 U10756 ( .A1(n11601), .A2(n15497), .ZN(n12500) );
  XNOR2_X1 U10757 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8460) );
  NAND2_X1 U10758 ( .A1(n9301), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8459) );
  INV_X1 U10759 ( .A(n8459), .ZN(n8345) );
  NAND2_X1 U10760 ( .A1(n8460), .A2(n8345), .ZN(n8347) );
  NAND2_X1 U10761 ( .A1(n9048), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U10762 ( .A1(n8347), .A2(n8346), .ZN(n8477) );
  NAND2_X1 U10763 ( .A1(n9054), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10764 ( .A1(n8477), .A2(n8348), .ZN(n8350) );
  NAND2_X1 U10765 ( .A1(n9453), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U10766 ( .A1(n8350), .A2(n8349), .ZN(n8492) );
  NAND2_X1 U10767 ( .A1(n9056), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8352) );
  INV_X1 U10768 ( .A(n8504), .ZN(n8353) );
  INV_X1 U10769 ( .A(n8519), .ZN(n8354) );
  NAND2_X1 U10770 ( .A1(n8520), .A2(n8354), .ZN(n8356) );
  NAND2_X1 U10771 ( .A1(n9074), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U10772 ( .A1(n13630), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8357) );
  INV_X1 U10773 ( .A(n8537), .ZN(n8358) );
  NAND2_X1 U10774 ( .A1(n9087), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10775 ( .A1(n9094), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8361) );
  XNOR2_X1 U10776 ( .A(n13821), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n8564) );
  INV_X1 U10777 ( .A(n8564), .ZN(n8363) );
  NAND2_X1 U10778 ( .A1(n13821), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U10779 ( .A1(n9131), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U10780 ( .A1(n8366), .A2(n8365), .ZN(n8578) );
  NAND2_X1 U10781 ( .A1(n9450), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U10782 ( .A1(n9448), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10783 ( .A1(n9446), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U10784 ( .A1(n9444), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U10785 ( .A1(n8372), .A2(n8371), .ZN(n8622) );
  NAND2_X1 U10786 ( .A1(n9617), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U10787 ( .A1(n9615), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8376) );
  INV_X1 U10788 ( .A(n8653), .ZN(n8380) );
  NAND2_X1 U10789 ( .A1(n9653), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8381) );
  INV_X1 U10790 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U10791 ( .A1(n9651), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U10792 ( .A1(n8381), .A2(n8378), .ZN(n8652) );
  INV_X1 U10793 ( .A(n8652), .ZN(n8379) );
  NAND2_X1 U10794 ( .A1(n13776), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U10795 ( .A1(n9600), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U10796 ( .A1(n9655), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U10797 ( .A1(n13792), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U10798 ( .A1(n9835), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10799 ( .A1(n9837), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8386) );
  INV_X1 U10800 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10153) );
  NAND2_X1 U10801 ( .A1(n10153), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8389) );
  INV_X1 U10802 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10151) );
  NAND2_X1 U10803 ( .A1(n10151), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10804 ( .A1(n10498), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10805 ( .A1(n11394), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8390) );
  AND2_X1 U10806 ( .A1(n8391), .A2(n8390), .ZN(n8724) );
  NAND2_X1 U10807 ( .A1(n10716), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8393) );
  INV_X1 U10808 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11408) );
  NAND2_X1 U10809 ( .A1(n11408), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8392) );
  AND2_X1 U10810 ( .A1(n8393), .A2(n8392), .ZN(n8737) );
  NAND2_X1 U10811 ( .A1(n8394), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10812 ( .A1(n13738), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10813 ( .A1(n8397), .A2(n8395), .ZN(n8749) );
  INV_X1 U10814 ( .A(n8749), .ZN(n8396) );
  XNOR2_X1 U10815 ( .A(n11434), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U10816 ( .A1(n11434), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8398) );
  INV_X1 U10817 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13906) );
  NAND2_X1 U10818 ( .A1(n8400), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10819 ( .A1(n14754), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8774) );
  INV_X1 U10820 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13903) );
  NAND2_X1 U10821 ( .A1(n13903), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10822 ( .A1(n8774), .A2(n8403), .ZN(n8404) );
  NAND2_X1 U10823 ( .A1(n8405), .A2(n8404), .ZN(n8406) );
  NAND2_X1 U10824 ( .A1(n8775), .A2(n8406), .ZN(n10681) );
  NAND2_X2 U10825 ( .A1(n6563), .A2(n9293), .ZN(n8503) );
  INV_X1 U10826 ( .A(SI_25_), .ZN(n10680) );
  INV_X2 U10827 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U10828 ( .A1(n8485), .A2(n8418), .ZN(n8512) );
  INV_X1 U10829 ( .A(n8512), .ZN(n8420) );
  NAND2_X1 U10830 ( .A1(n8420), .A2(n8419), .ZN(n8527) );
  OR2_X2 U10831 ( .A1(n8557), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8568) );
  OR2_X2 U10832 ( .A1(n8597), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8611) );
  INV_X1 U10833 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8427) );
  OR2_X2 U10834 ( .A1(n8646), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8662) );
  INV_X1 U10835 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8429) );
  OR2_X2 U10836 ( .A1(n8676), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8690) );
  INV_X1 U10837 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8431) );
  OR2_X2 U10838 ( .A1(n8704), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8718) );
  INV_X1 U10839 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8433) );
  OR2_X2 U10840 ( .A1(n8730), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8743) );
  INV_X1 U10841 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8435) );
  OR2_X2 U10842 ( .A1(n8753), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8761) );
  OR2_X2 U10843 ( .A1(n8761), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8768) );
  INV_X1 U10844 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8437) );
  INV_X1 U10845 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10846 ( .A1(n8770), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10847 ( .A1(n8782), .A2(n8441), .ZN(n12309) );
  NAND2_X1 U10848 ( .A1(n12309), .A2(n8484), .ZN(n8449) );
  AND2_X4 U10849 ( .A1(n8443), .A2(n12628), .ZN(n8827) );
  INV_X1 U10850 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n13801) );
  NAND2_X1 U10851 ( .A1(n8877), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10852 ( .A1(n6568), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8445) );
  OAI211_X1 U10853 ( .C1(n10337), .C2(n13801), .A(n8446), .B(n8445), .ZN(n8447) );
  INV_X1 U10854 ( .A(n8447), .ZN(n8448) );
  INV_X1 U10855 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9904) );
  OR2_X1 U10856 ( .A1(n8458), .A2(n9904), .ZN(n8453) );
  NAND2_X1 U10857 ( .A1(n6568), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10858 ( .A1(n8484), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U10859 ( .A1(n8827), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8450) );
  INV_X1 U10860 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9648) );
  MUX2_X1 U10861 ( .A(n9648), .B(n9302), .S(n6563), .Z(n8457) );
  NAND2_X1 U10862 ( .A1(n8454), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8455) );
  AND2_X1 U10863 ( .A1(n8459), .A2(n8455), .ZN(n9030) );
  OR2_X1 U10864 ( .A1(n8503), .A2(n9030), .ZN(n8456) );
  INV_X1 U10865 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15468) );
  OR2_X1 U10866 ( .A1(n8458), .A2(n15468), .ZN(n8469) );
  NAND2_X1 U10867 ( .A1(n8827), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10868 ( .A1(n8486), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10869 ( .A1(n6566), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8467) );
  NAND4_X1 U10870 ( .A1(n8469), .A2(n8470), .A3(n8468), .A4(n8467), .ZN(n9514)
         );
  INV_X1 U10871 ( .A(n8518), .ZN(n8659) );
  XNOR2_X1 U10872 ( .A(n8460), .B(n8459), .ZN(n9068) );
  INV_X1 U10873 ( .A(n8461), .ZN(n8462) );
  OR2_X1 U10874 ( .A1(n6563), .A2(n9546), .ZN(n8464) );
  NAND2_X1 U10875 ( .A1(n9514), .A2(n10290), .ZN(n11995) );
  NAND2_X1 U10876 ( .A1(n11991), .A2(n11995), .ZN(n9864) );
  INV_X1 U10877 ( .A(n10290), .ZN(n8471) );
  NAND2_X2 U10878 ( .A1(n8471), .A2(n10076), .ZN(n11996) );
  NAND2_X1 U10879 ( .A1(n9864), .A2(n11996), .ZN(n11543) );
  NAND2_X1 U10880 ( .A1(n6567), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10881 ( .A1(n8543), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U10882 ( .A1(n8827), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10883 ( .A1(n8484), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8472) );
  OR2_X1 U10884 ( .A1(n8518), .A2(SI_2_), .ZN(n8482) );
  XNOR2_X1 U10885 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8476) );
  XNOR2_X1 U10886 ( .A(n8477), .B(n8476), .ZN(n9036) );
  OR2_X1 U10887 ( .A1(n8503), .A2(n9036), .ZN(n8481) );
  NOR2_X1 U10888 ( .A1(n8461), .A2(n12619), .ZN(n8478) );
  OR2_X1 U10889 ( .A1(n6563), .A2(n9664), .ZN(n8480) );
  NAND3_X1 U10890 ( .A1(n8482), .A2(n8481), .A3(n8480), .ZN(n10083) );
  NAND2_X1 U10891 ( .A1(n11543), .A2(n11971), .ZN(n8483) );
  INV_X1 U10892 ( .A(n12180), .ZN(n11998) );
  NAND2_X1 U10893 ( .A1(n11998), .A2(n11997), .ZN(n12003) );
  NAND2_X1 U10894 ( .A1(n8484), .A2(n8485), .ZN(n8490) );
  NAND2_X1 U10895 ( .A1(n6567), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10896 ( .A1(n8543), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10897 ( .A1(n8827), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8487) );
  OR2_X1 U10898 ( .A1(n8518), .A2(SI_3_), .ZN(n8496) );
  XNOR2_X1 U10899 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8491) );
  XNOR2_X1 U10900 ( .A(n8492), .B(n8491), .ZN(n9033) );
  NAND2_X1 U10901 ( .A1(n8479), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8493) );
  XNOR2_X1 U10902 ( .A(n8493), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9697) );
  OR2_X1 U10903 ( .A1(n6563), .A2(n9697), .ZN(n8494) );
  INV_X1 U10904 ( .A(n8837), .ZN(n9508) );
  AND2_X1 U10905 ( .A1(n12002), .A2(n12010), .ZN(n10224) );
  NAND2_X1 U10906 ( .A1(n8497), .A2(n12002), .ZN(n10459) );
  NAND2_X1 U10907 ( .A1(n6567), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U10908 ( .A1(n8827), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U10909 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8498) );
  NAND2_X1 U10910 ( .A1(n8512), .A2(n8498), .ZN(n10508) );
  NAND2_X1 U10911 ( .A1(n6566), .A2(n10508), .ZN(n8500) );
  NAND2_X1 U10912 ( .A1(n8543), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8499) );
  NAND4_X1 U10913 ( .A1(n8502), .A2(n8501), .A3(n8500), .A4(n8499), .ZN(n12179) );
  OR2_X1 U10914 ( .A1(n11951), .A2(SI_4_), .ZN(n8509) );
  XNOR2_X1 U10915 ( .A(n8505), .B(n8504), .ZN(n9064) );
  OR2_X1 U10916 ( .A1(n8813), .A2(n9064), .ZN(n8508) );
  NAND2_X1 U10917 ( .A1(n8521), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8506) );
  OR2_X1 U10918 ( .A1(n9535), .A2(n9816), .ZN(n8507) );
  AND3_X2 U10919 ( .A1(n8509), .A2(n8508), .A3(n8507), .ZN(n12015) );
  NAND2_X1 U10920 ( .A1(n10459), .A2(n12008), .ZN(n8511) );
  INV_X1 U10921 ( .A(n12179), .ZN(n10559) );
  NAND2_X1 U10922 ( .A1(n10559), .A2(n12015), .ZN(n8510) );
  NAND2_X1 U10923 ( .A1(n8511), .A2(n8510), .ZN(n10520) );
  NAND2_X1 U10924 ( .A1(n6568), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U10925 ( .A1(n8827), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U10926 ( .A1(n8512), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U10927 ( .A1(n8527), .A2(n8513), .ZN(n10548) );
  NAND2_X1 U10928 ( .A1(n6566), .A2(n10548), .ZN(n8515) );
  NAND2_X1 U10929 ( .A1(n8877), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8514) );
  OR2_X1 U10930 ( .A1(n11951), .A2(SI_5_), .ZN(n8525) );
  XNOR2_X1 U10931 ( .A(n8520), .B(n8519), .ZN(n9041) );
  OR2_X1 U10932 ( .A1(n8813), .A2(n9041), .ZN(n8524) );
  NOR2_X1 U10933 ( .A1(n8521), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8533) );
  OR2_X1 U10934 ( .A1(n8533), .A2(n12619), .ZN(n8522) );
  XNOR2_X1 U10935 ( .A(n8522), .B(P3_IR_REG_5__SCAN_IN), .ZN(n9882) );
  OR2_X1 U10936 ( .A1(n9535), .A2(n9882), .ZN(n8523) );
  NAND2_X1 U10937 ( .A1(n10734), .A2(n10562), .ZN(n12018) );
  INV_X1 U10938 ( .A(n10734), .ZN(n10748) );
  INV_X1 U10939 ( .A(n10562), .ZN(n15486) );
  NAND2_X1 U10940 ( .A1(n10748), .A2(n15486), .ZN(n12011) );
  NAND2_X1 U10941 ( .A1(n10520), .A2(n12012), .ZN(n8526) );
  NAND2_X1 U10942 ( .A1(n8526), .A2(n12018), .ZN(n10741) );
  NAND2_X1 U10943 ( .A1(n6567), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U10944 ( .A1(n8827), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8531) );
  NAND2_X1 U10945 ( .A1(n8527), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10946 ( .A1(n8541), .A2(n8528), .ZN(n10753) );
  NAND2_X1 U10947 ( .A1(n8484), .A2(n10753), .ZN(n8530) );
  NAND2_X1 U10948 ( .A1(n8543), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U10949 ( .A1(n8533), .A2(n13831), .ZN(n8535) );
  NAND2_X1 U10950 ( .A1(n8535), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8534) );
  MUX2_X1 U10951 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8534), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n8536) );
  NAND2_X1 U10952 ( .A1(n8536), .A2(n8550), .ZN(n10172) );
  INV_X1 U10953 ( .A(SI_6_), .ZN(n9031) );
  OR2_X1 U10954 ( .A1(n11951), .A2(n9031), .ZN(n8540) );
  XNOR2_X1 U10955 ( .A(n8538), .B(n8537), .ZN(n9032) );
  OR2_X1 U10956 ( .A1(n8813), .A2(n9032), .ZN(n8539) );
  NAND2_X1 U10957 ( .A1(n10844), .A2(n10754), .ZN(n12024) );
  INV_X1 U10958 ( .A(n10844), .ZN(n12178) );
  NAND2_X1 U10959 ( .A1(n12178), .A2(n15491), .ZN(n12025) );
  AND2_X1 U10960 ( .A1(n12024), .A2(n12025), .ZN(n10743) );
  NAND2_X1 U10961 ( .A1(n6568), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10962 ( .A1(n8827), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U10963 ( .A1(n8541), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U10964 ( .A1(n8557), .A2(n8542), .ZN(n10797) );
  NAND2_X1 U10965 ( .A1(n8484), .A2(n10797), .ZN(n8545) );
  NAND2_X1 U10966 ( .A1(n8543), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8544) );
  NAND4_X1 U10967 ( .A1(n8547), .A2(n8546), .A3(n8545), .A4(n8544), .ZN(n12177) );
  OR2_X1 U10968 ( .A1(n11951), .A2(SI_7_), .ZN(n8556) );
  XNOR2_X1 U10969 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8548) );
  XNOR2_X1 U10970 ( .A(n8549), .B(n8548), .ZN(n9069) );
  OR2_X1 U10971 ( .A1(n8813), .A2(n9069), .ZN(n8555) );
  NAND2_X1 U10972 ( .A1(n8550), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8551) );
  MUX2_X1 U10973 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8551), .S(
        P3_IR_REG_7__SCAN_IN), .Z(n8553) );
  NAND2_X1 U10974 ( .A1(n8553), .A2(n8552), .ZN(n10259) );
  OR2_X1 U10975 ( .A1(n6563), .A2(n10254), .ZN(n8554) );
  INV_X1 U10976 ( .A(n12177), .ZN(n11074) );
  NAND2_X1 U10977 ( .A1(n11074), .A2(n10796), .ZN(n12030) );
  NAND2_X1 U10978 ( .A1(n6568), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U10979 ( .A1(n8827), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10980 ( .A1(n8557), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10981 ( .A1(n8568), .A2(n8558), .ZN(n11077) );
  NAND2_X1 U10982 ( .A1(n8484), .A2(n11077), .ZN(n8560) );
  NAND2_X1 U10983 ( .A1(n8877), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8559) );
  NAND4_X1 U10984 ( .A1(n8562), .A2(n8561), .A3(n8560), .A4(n8559), .ZN(n12176) );
  NAND2_X1 U10985 ( .A1(n8552), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8563) );
  XNOR2_X1 U10986 ( .A(n8563), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10612) );
  INV_X1 U10987 ( .A(SI_8_), .ZN(n9039) );
  OR2_X1 U10988 ( .A1(n11951), .A2(n9039), .ZN(n8567) );
  XNOR2_X1 U10989 ( .A(n8565), .B(n8564), .ZN(n9040) );
  OR2_X1 U10990 ( .A1(n8503), .A2(n9040), .ZN(n8566) );
  OAI211_X1 U10991 ( .C1(n9535), .C2(n10631), .A(n8567), .B(n8566), .ZN(n12034) );
  XNOR2_X1 U10992 ( .A(n12176), .B(n12034), .ZN(n12032) );
  INV_X1 U10993 ( .A(n12176), .ZN(n10890) );
  NAND2_X1 U10994 ( .A1(n10890), .A2(n12034), .ZN(n12035) );
  NAND2_X1 U10995 ( .A1(n8827), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U10996 ( .A1(n6567), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U10997 ( .A1(n8568), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10998 ( .A1(n8584), .A2(n8569), .ZN(n10892) );
  NAND2_X1 U10999 ( .A1(n8484), .A2(n10892), .ZN(n8570) );
  NOR2_X1 U11000 ( .A1(n8573), .A2(n12619), .ZN(n8574) );
  MUX2_X1 U11001 ( .A(n12619), .B(n8574), .S(P3_IR_REG_9__SCAN_IN), .Z(n8575)
         );
  INV_X1 U11002 ( .A(n8575), .ZN(n8577) );
  INV_X1 U11003 ( .A(n8325), .ZN(n8576) );
  NAND2_X1 U11004 ( .A1(n8577), .A2(n8576), .ZN(n15453) );
  INV_X1 U11005 ( .A(n15453), .ZN(n10632) );
  NAND2_X1 U11006 ( .A1(n8579), .A2(n8578), .ZN(n8580) );
  AND2_X1 U11007 ( .A1(n8581), .A2(n8580), .ZN(n9051) );
  OR2_X1 U11008 ( .A1(n8813), .A2(n9051), .ZN(n8583) );
  OR2_X1 U11009 ( .A1(n11951), .A2(SI_9_), .ZN(n8582) );
  OAI211_X1 U11010 ( .C1(n10632), .C2(n9535), .A(n8583), .B(n8582), .ZN(n10860) );
  NAND2_X1 U11011 ( .A1(n12175), .A2(n10860), .ZN(n12040) );
  NAND2_X1 U11012 ( .A1(n8827), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U11013 ( .A1(n6567), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U11014 ( .A1(n8584), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U11015 ( .A1(n8597), .A2(n8585), .ZN(n10842) );
  NAND2_X1 U11016 ( .A1(n8484), .A2(n10842), .ZN(n8587) );
  NAND2_X1 U11017 ( .A1(n8877), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8586) );
  XNOR2_X1 U11018 ( .A(n9450), .B(P2_DATAO_REG_10__SCAN_IN), .ZN(n8590) );
  XNOR2_X1 U11019 ( .A(n8591), .B(n8590), .ZN(n9072) );
  OR2_X1 U11020 ( .A1(n8813), .A2(n9072), .ZN(n8595) );
  OR2_X1 U11021 ( .A1(n11951), .A2(SI_10_), .ZN(n8594) );
  OR2_X1 U11022 ( .A1(n8325), .A2(n12619), .ZN(n8592) );
  INV_X1 U11023 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8605) );
  XNOR2_X1 U11024 ( .A(n8592), .B(n8605), .ZN(n10802) );
  INV_X1 U11025 ( .A(n10802), .ZN(n10805) );
  OR2_X1 U11026 ( .A1(n9535), .A2(n10805), .ZN(n8593) );
  NAND2_X1 U11027 ( .A1(n11086), .A2(n10869), .ZN(n12044) );
  NAND2_X1 U11028 ( .A1(n12174), .A2(n15514), .ZN(n12049) );
  INV_X1 U11029 ( .A(n12049), .ZN(n8596) );
  NAND2_X1 U11030 ( .A1(n8827), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U11031 ( .A1(n6568), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U11032 ( .A1(n8597), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U11033 ( .A1(n8611), .A2(n8598), .ZN(n11131) );
  NAND2_X1 U11034 ( .A1(n8484), .A2(n11131), .ZN(n8600) );
  NAND2_X1 U11035 ( .A1(n8877), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8599) );
  XNOR2_X1 U11036 ( .A(n7317), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8603) );
  XNOR2_X1 U11037 ( .A(n8604), .B(n8603), .ZN(n9078) );
  OR2_X1 U11038 ( .A1(n8813), .A2(n9078), .ZN(n8610) );
  OR2_X1 U11039 ( .A1(n11951), .A2(SI_11_), .ZN(n8609) );
  NAND2_X1 U11040 ( .A1(n8325), .A2(n8605), .ZN(n8617) );
  NAND2_X1 U11041 ( .A1(n8617), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8607) );
  INV_X1 U11042 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8606) );
  XNOR2_X1 U11043 ( .A(n8607), .B(n8606), .ZN(n10929) );
  INV_X1 U11044 ( .A(n10929), .ZN(n10936) );
  OR2_X1 U11045 ( .A1(n9535), .A2(n10936), .ZN(n8608) );
  XNOR2_X1 U11046 ( .A(n12173), .B(n11133), .ZN(n12050) );
  NAND2_X1 U11047 ( .A1(n11113), .A2(n12050), .ZN(n11112) );
  NAND2_X1 U11048 ( .A1(n11149), .A2(n11133), .ZN(n12057) );
  NAND2_X1 U11049 ( .A1(n8827), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U11050 ( .A1(n6567), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U11051 ( .A1(n8611), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U11052 ( .A1(n8634), .A2(n8612), .ZN(n11170) );
  NAND2_X1 U11053 ( .A1(n6566), .A2(n11170), .ZN(n8614) );
  NAND2_X1 U11054 ( .A1(n8877), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8613) );
  NOR2_X1 U11055 ( .A1(n8617), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8620) );
  OR2_X1 U11056 ( .A1(n8620), .A2(n12619), .ZN(n8618) );
  MUX2_X1 U11057 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8618), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8621) );
  INV_X1 U11058 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U11059 ( .A1(n8620), .A2(n8619), .ZN(n8631) );
  NAND2_X1 U11060 ( .A1(n8621), .A2(n8631), .ZN(n11230) );
  NAND2_X1 U11061 ( .A1(n8623), .A2(n8622), .ZN(n8624) );
  NAND2_X1 U11062 ( .A1(n8625), .A2(n8624), .ZN(n9086) );
  OR2_X1 U11063 ( .A1(n8813), .A2(n9086), .ZN(n8627) );
  OR2_X1 U11064 ( .A1(n11951), .A2(n13820), .ZN(n8626) );
  OAI211_X1 U11065 ( .C1(n9535), .C2(n11230), .A(n8627), .B(n8626), .ZN(n11171) );
  NOR2_X1 U11066 ( .A1(n11144), .A2(n11171), .ZN(n12054) );
  INV_X1 U11067 ( .A(n11171), .ZN(n12614) );
  NOR2_X1 U11068 ( .A1(n12481), .A2(n12614), .ZN(n12055) );
  NOR2_X1 U11069 ( .A1(n12054), .A2(n12055), .ZN(n11164) );
  INV_X1 U11070 ( .A(n12055), .ZN(n12058) );
  NAND2_X1 U11071 ( .A1(n6667), .A2(n9505), .ZN(n8628) );
  NAND2_X1 U11072 ( .A1(n8629), .A2(n8628), .ZN(n9127) );
  NAND2_X1 U11073 ( .A1(n8631), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8630) );
  MUX2_X1 U11074 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8630), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8632) );
  NAND2_X1 U11075 ( .A1(n8632), .A2(n8656), .ZN(n11257) );
  INV_X1 U11076 ( .A(n11257), .ZN(n11235) );
  OAI22_X1 U11077 ( .A1(n11951), .A2(SI_13_), .B1(n11235), .B2(n9535), .ZN(
        n8633) );
  AOI21_X1 U11078 ( .B1(n9127), .B2(n11948), .A(n8633), .ZN(n11105) );
  NAND2_X1 U11079 ( .A1(n6568), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8639) );
  NAND2_X1 U11080 ( .A1(n8827), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U11081 ( .A1(n8634), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U11082 ( .A1(n8646), .A2(n8635), .ZN(n12484) );
  NAND2_X1 U11083 ( .A1(n8484), .A2(n12484), .ZN(n8637) );
  NAND2_X1 U11084 ( .A1(n8877), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8636) );
  AND2_X1 U11085 ( .A1(n11105), .A2(n11099), .ZN(n12059) );
  INV_X1 U11086 ( .A(n11105), .ZN(n12609) );
  NAND2_X1 U11087 ( .A1(n12609), .A2(n12464), .ZN(n12063) );
  XNOR2_X1 U11088 ( .A(n8641), .B(n8640), .ZN(n9184) );
  NAND2_X1 U11089 ( .A1(n9184), .A2(n11948), .ZN(n8645) );
  INV_X1 U11090 ( .A(n9535), .ZN(n8715) );
  NAND2_X1 U11091 ( .A1(n8656), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8643) );
  INV_X1 U11092 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8642) );
  XNOR2_X1 U11093 ( .A(n8643), .B(n8642), .ZN(n11225) );
  AOI22_X1 U11094 ( .A1(n8659), .A2(n9183), .B1(n8715), .B2(n11225), .ZN(n8644) );
  NAND2_X1 U11095 ( .A1(n8827), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U11096 ( .A1(n6568), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U11097 ( .A1(n8646), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U11098 ( .A1(n8662), .A2(n8647), .ZN(n12467) );
  NAND2_X1 U11099 ( .A1(n8484), .A2(n12467), .ZN(n8649) );
  NAND2_X1 U11100 ( .A1(n8877), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8648) );
  NAND4_X1 U11101 ( .A1(n8651), .A2(n8650), .A3(n8649), .A4(n8648), .ZN(n12478) );
  OR2_X1 U11102 ( .A1(n12605), .A2(n12478), .ZN(n12068) );
  NAND2_X1 U11103 ( .A1(n8653), .A2(n8652), .ZN(n8655) );
  NAND2_X1 U11104 ( .A1(n8655), .A2(n8654), .ZN(n9451) );
  NAND2_X1 U11105 ( .A1(n9451), .A2(n11948), .ZN(n8661) );
  INV_X1 U11106 ( .A(SI_15_), .ZN(n13727) );
  OAI21_X1 U11107 ( .B1(n8656), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8658) );
  INV_X1 U11108 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8657) );
  XNOR2_X1 U11109 ( .A(n8658), .B(n8657), .ZN(n12222) );
  AOI22_X1 U11110 ( .A1(n8659), .A2(n13727), .B1(n8715), .B2(n12222), .ZN(
        n8660) );
  NAND2_X1 U11111 ( .A1(n8661), .A2(n8660), .ZN(n12543) );
  NAND2_X1 U11112 ( .A1(n8827), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11113 ( .A1(n6568), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U11114 ( .A1(n8662), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U11115 ( .A1(n8676), .A2(n8663), .ZN(n12447) );
  NAND2_X1 U11116 ( .A1(n8484), .A2(n12447), .ZN(n8665) );
  NAND2_X1 U11117 ( .A1(n8877), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8664) );
  NAND4_X1 U11118 ( .A1(n8667), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n12463) );
  NAND2_X1 U11119 ( .A1(n12543), .A2(n12463), .ZN(n12071) );
  OR2_X1 U11120 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  AND2_X1 U11121 ( .A1(n8671), .A2(n8670), .ZN(n9506) );
  NAND2_X1 U11122 ( .A1(n9506), .A2(n11948), .ZN(n8675) );
  MUX2_X1 U11123 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8672), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8673) );
  AND2_X1 U11124 ( .A1(n8673), .A2(n8686), .ZN(n12220) );
  AOI22_X1 U11125 ( .A1(n8659), .A2(SI_16_), .B1(n8715), .B2(n12220), .ZN(
        n8674) );
  NAND2_X1 U11126 ( .A1(n8827), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11127 ( .A1(n6567), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11128 ( .A1(n8676), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U11129 ( .A1(n8690), .A2(n8677), .ZN(n12437) );
  NAND2_X1 U11130 ( .A1(n8484), .A2(n12437), .ZN(n8679) );
  NAND2_X1 U11131 ( .A1(n8877), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8678) );
  NAND4_X1 U11132 ( .A1(n8681), .A2(n8680), .A3(n8679), .A4(n8678), .ZN(n12452) );
  NAND2_X1 U11133 ( .A1(n12539), .A2(n12452), .ZN(n12078) );
  INV_X1 U11134 ( .A(n12539), .ZN(n12439) );
  INV_X1 U11135 ( .A(n12452), .ZN(n11934) );
  NAND2_X1 U11136 ( .A1(n12439), .A2(n11934), .ZN(n12074) );
  NAND2_X1 U11137 ( .A1(n12428), .A2(n12074), .ZN(n12416) );
  OR2_X1 U11138 ( .A1(n8683), .A2(n8682), .ZN(n8684) );
  NAND2_X1 U11139 ( .A1(n8685), .A2(n8684), .ZN(n9511) );
  NAND2_X1 U11140 ( .A1(n9511), .A2(n11948), .ZN(n8689) );
  NAND2_X1 U11141 ( .A1(n8686), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8687) );
  XNOR2_X1 U11142 ( .A(n8687), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14906) );
  INV_X1 U11143 ( .A(n14906), .ZN(n12252) );
  AOI22_X1 U11144 ( .A1(n8659), .A2(n9512), .B1(n8715), .B2(n12252), .ZN(n8688) );
  NAND2_X1 U11145 ( .A1(n8827), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U11146 ( .A1(n6567), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U11147 ( .A1(n8690), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11148 ( .A1(n8704), .A2(n8691), .ZN(n12417) );
  NAND2_X1 U11149 ( .A1(n6566), .A2(n12417), .ZN(n8693) );
  NAND2_X1 U11150 ( .A1(n8877), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8692) );
  NAND4_X1 U11151 ( .A1(n8695), .A2(n8694), .A3(n8693), .A4(n8692), .ZN(n12434) );
  NAND2_X1 U11152 ( .A1(n12535), .A2(n12434), .ZN(n12093) );
  OR2_X1 U11153 ( .A1(n8697), .A2(n8696), .ZN(n8698) );
  NAND2_X1 U11154 ( .A1(n8699), .A2(n8698), .ZN(n9618) );
  NAND2_X1 U11155 ( .A1(n8700), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8701) );
  XNOR2_X1 U11156 ( .A(n8701), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U11157 ( .A1(n8659), .A2(SI_18_), .B1(n8715), .B2(n12267), .ZN(
        n8702) );
  NAND2_X1 U11158 ( .A1(n8827), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U11159 ( .A1(n6567), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11160 ( .A1(n8704), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U11161 ( .A1(n8718), .A2(n8705), .ZN(n12409) );
  NAND2_X1 U11162 ( .A1(n8484), .A2(n12409), .ZN(n8707) );
  NAND2_X1 U11163 ( .A1(n8877), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8706) );
  NAND4_X1 U11164 ( .A1(n8709), .A2(n8708), .A3(n8707), .A4(n8706), .ZN(n12422) );
  NAND2_X1 U11165 ( .A1(n12598), .A2(n12422), .ZN(n8710) );
  INV_X1 U11166 ( .A(n12598), .ZN(n8855) );
  INV_X1 U11167 ( .A(n12422), .ZN(n12382) );
  NAND2_X1 U11168 ( .A1(n8855), .A2(n12382), .ZN(n12096) );
  NAND2_X1 U11169 ( .A1(n8710), .A2(n12096), .ZN(n12398) );
  INV_X1 U11170 ( .A(n8710), .ZN(n12083) );
  OR2_X1 U11171 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  NAND2_X1 U11172 ( .A1(n8714), .A2(n8713), .ZN(n9679) );
  AOI22_X1 U11173 ( .A1(n8659), .A2(SI_19_), .B1(n12268), .B2(n8715), .ZN(
        n8716) );
  NAND2_X1 U11174 ( .A1(n8827), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U11175 ( .A1(n6568), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U11176 ( .A1(n8718), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11177 ( .A1(n8730), .A2(n8719), .ZN(n12386) );
  NAND2_X1 U11178 ( .A1(n6566), .A2(n12386), .ZN(n8721) );
  NAND2_X1 U11179 ( .A1(n8877), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8720) );
  OR2_X1 U11180 ( .A1(n12390), .A2(n12407), .ZN(n12082) );
  NAND2_X1 U11181 ( .A1(n12390), .A2(n12407), .ZN(n12101) );
  OR2_X1 U11182 ( .A1(n8725), .A2(n8724), .ZN(n8726) );
  NAND2_X1 U11183 ( .A1(n8727), .A2(n8726), .ZN(n9718) );
  NAND2_X1 U11184 ( .A1(n8827), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U11185 ( .A1(n6568), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U11186 ( .A1(n8730), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11187 ( .A1(n8743), .A2(n8731), .ZN(n12375) );
  NAND2_X1 U11188 ( .A1(n6566), .A2(n12375), .ZN(n8733) );
  NAND2_X1 U11189 ( .A1(n8877), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8732) );
  XNOR2_X1 U11190 ( .A(n12104), .B(n12381), .ZN(n12370) );
  OR2_X1 U11191 ( .A1(n8738), .A2(n8737), .ZN(n8739) );
  NAND2_X1 U11192 ( .A1(n8740), .A2(n8739), .ZN(n9834) );
  INV_X1 U11193 ( .A(SI_21_), .ZN(n9833) );
  NAND2_X1 U11194 ( .A1(n6568), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11195 ( .A1(n8877), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U11196 ( .A1(n8743), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11197 ( .A1(n8753), .A2(n8744), .ZN(n12361) );
  NAND2_X1 U11198 ( .A1(n6566), .A2(n12361), .ZN(n8746) );
  NAND2_X1 U11199 ( .A1(n8827), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8745) );
  AND2_X1 U11200 ( .A1(n8856), .A2(n12348), .ZN(n12109) );
  XNOR2_X1 U11201 ( .A(n8750), .B(n8749), .ZN(n9876) );
  NAND2_X1 U11202 ( .A1(n9876), .A2(n11948), .ZN(n8752) );
  NAND2_X1 U11203 ( .A1(n8753), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U11204 ( .A1(n8761), .A2(n8754), .ZN(n12350) );
  AOI22_X1 U11205 ( .A1(n12350), .A2(n8484), .B1(n8877), .B2(
        P3_REG0_REG_22__SCAN_IN), .ZN(n8756) );
  AOI22_X1 U11206 ( .A1(n8827), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n6567), .B2(
        P3_REG1_REG_22__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11207 ( .A1(n11905), .A2(n12360), .ZN(n12117) );
  XNOR2_X1 U11208 ( .A(n8758), .B(n8757), .ZN(n10154) );
  NAND2_X1 U11209 ( .A1(n10154), .A2(n11948), .ZN(n8760) );
  INV_X1 U11210 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12579) );
  NAND2_X1 U11211 ( .A1(n8761), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U11212 ( .A1(n8768), .A2(n8762), .ZN(n12339) );
  NAND2_X1 U11213 ( .A1(n12339), .A2(n8484), .ZN(n8764) );
  AOI22_X1 U11214 ( .A1(n8827), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n6568), .B2(
        P3_REG1_REG_23__SCAN_IN), .ZN(n8763) );
  INV_X1 U11215 ( .A(n12320), .ZN(n12349) );
  NOR2_X1 U11216 ( .A1(n12338), .A2(n12349), .ZN(n12121) );
  XNOR2_X1 U11217 ( .A(n8765), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n10544) );
  NAND2_X1 U11218 ( .A1(n10544), .A2(n11948), .ZN(n8767) );
  INV_X1 U11219 ( .A(SI_24_), .ZN(n10545) );
  NAND2_X1 U11220 ( .A1(n8768), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U11221 ( .A1(n8770), .A2(n8769), .ZN(n12324) );
  NAND2_X1 U11222 ( .A1(n12324), .A2(n6566), .ZN(n8773) );
  AOI22_X1 U11223 ( .A1(n8827), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n6567), .B2(
        P3_REG1_REG_24__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U11224 ( .A1(n8877), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U11225 ( .A1(n11878), .A2(n12335), .ZN(n12120) );
  NAND2_X1 U11226 ( .A1(n12316), .A2(n12315), .ZN(n12314) );
  NAND2_X1 U11227 ( .A1(n14750), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8789) );
  INV_X1 U11228 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13899) );
  NAND2_X1 U11229 ( .A1(n13899), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8776) );
  AND2_X1 U11230 ( .A1(n8789), .A2(n8776), .ZN(n8777) );
  OR2_X1 U11231 ( .A1(n8778), .A2(n8777), .ZN(n8779) );
  NAND2_X1 U11232 ( .A1(n8790), .A2(n8779), .ZN(n10873) );
  INV_X1 U11233 ( .A(SI_26_), .ZN(n10874) );
  OR2_X2 U11234 ( .A1(n8782), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U11235 ( .A1(n8782), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8783) );
  NAND2_X1 U11236 ( .A1(n8796), .A2(n8783), .ZN(n12291) );
  NAND2_X1 U11237 ( .A1(n12291), .A2(n6566), .ZN(n8788) );
  INV_X1 U11238 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U11239 ( .A1(n8877), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U11240 ( .A1(n6568), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8784) );
  OAI211_X1 U11241 ( .C1(n10337), .C2(n12292), .A(n8785), .B(n8784), .ZN(n8786) );
  INV_X1 U11242 ( .A(n8786), .ZN(n8787) );
  NAND2_X1 U11243 ( .A1(n12295), .A2(n11860), .ZN(n12137) );
  NAND2_X1 U11244 ( .A1(n12135), .A2(n12137), .ZN(n11340) );
  NAND2_X1 U11245 ( .A1(n11329), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U11246 ( .A1(n13897), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U11247 ( .A1(n8807), .A2(n8791), .ZN(n8804) );
  XNOR2_X1 U11248 ( .A(n8806), .B(n8804), .ZN(n11160) );
  NAND2_X1 U11249 ( .A1(n11160), .A2(n11948), .ZN(n8793) );
  INV_X1 U11250 ( .A(n8796), .ZN(n8795) );
  INV_X1 U11251 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11252 ( .A1(n8795), .A2(n8794), .ZN(n8815) );
  NAND2_X1 U11253 ( .A1(n8796), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U11254 ( .A1(n8815), .A2(n8797), .ZN(n11668) );
  NAND2_X1 U11255 ( .A1(n11668), .A2(n6566), .ZN(n8802) );
  INV_X1 U11256 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n11608) );
  NAND2_X1 U11257 ( .A1(n8877), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U11258 ( .A1(n6568), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8798) );
  OAI211_X1 U11259 ( .C1(n10337), .C2(n11608), .A(n8799), .B(n8798), .ZN(n8800) );
  INV_X1 U11260 ( .A(n8800), .ZN(n8801) );
  AND2_X2 U11261 ( .A1(n8802), .A2(n8801), .ZN(n11923) );
  NAND2_X1 U11262 ( .A1(n11622), .A2(n11923), .ZN(n8945) );
  OR2_X2 U11263 ( .A1(n11622), .A2(n11923), .ZN(n8803) );
  NAND2_X2 U11264 ( .A1(n8945), .A2(n8803), .ZN(n11983) );
  INV_X1 U11265 ( .A(n8804), .ZN(n8805) );
  NAND2_X1 U11266 ( .A1(n8808), .A2(n8807), .ZN(n8811) );
  NAND2_X1 U11267 ( .A1(n13588), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U11268 ( .A1(n11484), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8809) );
  AND2_X1 U11269 ( .A1(n8821), .A2(n8809), .ZN(n8810) );
  NAND2_X1 U11270 ( .A1(n8811), .A2(n8810), .ZN(n8822) );
  OR2_X1 U11271 ( .A1(n8811), .A2(n8810), .ZN(n8812) );
  NAND2_X1 U11272 ( .A1(n8822), .A2(n8812), .ZN(n11083) );
  OR2_X1 U11273 ( .A1(n11951), .A2(n11082), .ZN(n8814) );
  NAND2_X1 U11274 ( .A1(n8815), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11275 ( .A1(n8826), .A2(n8816), .ZN(n11811) );
  INV_X1 U11276 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n11575) );
  NAND2_X1 U11277 ( .A1(n6567), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U11278 ( .A1(n8877), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8817) );
  OAI211_X1 U11279 ( .C1(n11575), .C2(n10337), .A(n8818), .B(n8817), .ZN(n8819) );
  INV_X1 U11280 ( .A(n8945), .ZN(n8820) );
  NOR2_X1 U11281 ( .A1(n8862), .A2(n8820), .ZN(n11982) );
  NOR2_X1 U11282 ( .A1(n11819), .A2(n11666), .ZN(n8861) );
  NAND2_X1 U11283 ( .A1(n8822), .A2(n8821), .ZN(n11332) );
  XNOR2_X1 U11284 ( .A(n13886), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n8823) );
  XNOR2_X1 U11285 ( .A(n11332), .B(n8823), .ZN(n12625) );
  NAND2_X1 U11286 ( .A1(n12625), .A2(n11948), .ZN(n8825) );
  INV_X1 U11287 ( .A(SI_29_), .ZN(n12630) );
  OR2_X1 U11288 ( .A1(n11951), .A2(n12630), .ZN(n8824) );
  NAND2_X1 U11289 ( .A1(n8825), .A2(n8824), .ZN(n8931) );
  NAND2_X1 U11290 ( .A1(n11615), .A2(n8484), .ZN(n10340) );
  INV_X1 U11291 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U11292 ( .A1(n8877), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8829) );
  NAND2_X1 U11293 ( .A1(n8827), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8828) );
  OAI211_X1 U11294 ( .C1(n8831), .C2(n8830), .A(n8829), .B(n8828), .ZN(n8832)
         );
  INV_X1 U11295 ( .A(n8832), .ZN(n8833) );
  INV_X1 U11296 ( .A(n8872), .ZN(n8834) );
  INV_X1 U11297 ( .A(n12390), .ZN(n12527) );
  INV_X1 U11298 ( .A(n10860), .ZN(n15507) );
  INV_X1 U11299 ( .A(n11559), .ZN(n9843) );
  NAND2_X1 U11300 ( .A1(n10076), .A2(n10290), .ZN(n8836) );
  NOR2_X1 U11301 ( .A1(n12180), .A2(n11997), .ZN(n10225) );
  OR2_X1 U11302 ( .A1(n8837), .A2(n15475), .ZN(n8838) );
  NAND2_X1 U11303 ( .A1(n10227), .A2(n8838), .ZN(n10461) );
  INV_X1 U11304 ( .A(n12008), .ZN(n10460) );
  NAND2_X1 U11305 ( .A1(n10461), .A2(n10460), .ZN(n8840) );
  NAND2_X1 U11306 ( .A1(n12179), .A2(n12015), .ZN(n8839) );
  OR2_X1 U11307 ( .A1(n10844), .A2(n15491), .ZN(n8841) );
  INV_X1 U11308 ( .A(n8841), .ZN(n10783) );
  OR2_X1 U11309 ( .A1(n12012), .A2(n10783), .ZN(n8843) );
  AND2_X1 U11310 ( .A1(n10734), .A2(n15486), .ZN(n10744) );
  AOI21_X1 U11311 ( .B1(n10742), .B2(n8841), .A(n12027), .ZN(n8842) );
  NAND2_X1 U11312 ( .A1(n12177), .A2(n10796), .ZN(n8844) );
  NAND2_X1 U11313 ( .A1(n8845), .A2(n8844), .ZN(n10987) );
  INV_X1 U11314 ( .A(n10987), .ZN(n8846) );
  INV_X1 U11315 ( .A(n8847), .ZN(n12041) );
  NOR2_X1 U11316 ( .A1(n12176), .A2(n12034), .ZN(n10770) );
  NOR2_X1 U11317 ( .A1(n12038), .A2(n10770), .ZN(n8848) );
  INV_X1 U11318 ( .A(n11108), .ZN(n8849) );
  NAND2_X1 U11319 ( .A1(n12481), .A2(n11171), .ZN(n8850) );
  NAND2_X1 U11320 ( .A1(n7610), .A2(n12063), .ZN(n12476) );
  INV_X1 U11321 ( .A(n12478), .ZN(n11625) );
  INV_X1 U11322 ( .A(n12463), .ZN(n11829) );
  INV_X1 U11323 ( .A(n12429), .ZN(n12432) );
  INV_X1 U11324 ( .A(n12398), .ZN(n12402) );
  NAND2_X1 U11325 ( .A1(n12358), .A2(n11965), .ZN(n8857) );
  NAND2_X1 U11326 ( .A1(n8856), .A2(n12372), .ZN(n11964) );
  INV_X1 U11327 ( .A(n11905), .ZN(n12585) );
  NOR2_X1 U11328 ( .A1(n12585), .A2(n12360), .ZN(n8858) );
  NAND2_X1 U11329 ( .A1(n12338), .A2(n12320), .ZN(n8859) );
  INV_X1 U11330 ( .A(n12335), .ZN(n12170) );
  NAND2_X1 U11331 ( .A1(n11878), .A2(n12170), .ZN(n8860) );
  INV_X1 U11332 ( .A(n8861), .ZN(n11986) );
  NAND2_X1 U11333 ( .A1(n11671), .A2(n11923), .ZN(n8865) );
  INV_X1 U11334 ( .A(n11983), .ZN(n8864) );
  NAND2_X1 U11335 ( .A1(n11927), .A2(n11860), .ZN(n11586) );
  AND2_X2 U11336 ( .A1(n8865), .A2(n11592), .ZN(n8947) );
  AND2_X2 U11337 ( .A1(n11984), .A2(n8947), .ZN(n8867) );
  AND2_X1 U11338 ( .A1(n12304), .A2(n8867), .ZN(n8866) );
  NAND2_X1 U11339 ( .A1(n12305), .A2(n8866), .ZN(n8952) );
  INV_X1 U11340 ( .A(n8867), .ZN(n8869) );
  NAND2_X1 U11341 ( .A1(n11650), .A2(n12321), .ZN(n12127) );
  NAND2_X1 U11342 ( .A1(n12295), .A2(n12306), .ZN(n8868) );
  AND2_X1 U11343 ( .A1(n12127), .A2(n8868), .ZN(n11587) );
  AND2_X1 U11344 ( .A1(n11587), .A2(n11983), .ZN(n11593) );
  INV_X1 U11345 ( .A(n11666), .ZN(n12168) );
  NAND2_X1 U11346 ( .A1(n11819), .A2(n12168), .ZN(n8870) );
  AND2_X1 U11347 ( .A1(n8951), .A2(n8870), .ZN(n8871) );
  NAND2_X1 U11348 ( .A1(n8952), .A2(n8871), .ZN(n8873) );
  XNOR2_X1 U11349 ( .A(n8873), .B(n8872), .ZN(n8887) );
  NAND2_X1 U11350 ( .A1(n12268), .A2(n12163), .ZN(n8934) );
  NOR2_X1 U11351 ( .A1(n11990), .A2(n9716), .ZN(n12157) );
  INV_X1 U11352 ( .A(n12157), .ZN(n8874) );
  INV_X1 U11353 ( .A(n11081), .ZN(n12160) );
  INV_X1 U11354 ( .A(n8875), .ZN(n9531) );
  NAND2_X1 U11355 ( .A1(n12160), .A2(n9531), .ZN(n9541) );
  AND2_X1 U11356 ( .A1(n9535), .A2(n9541), .ZN(n8883) );
  INV_X1 U11357 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11358 ( .A1(n8877), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U11359 ( .A1(n6568), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8878) );
  OAI211_X1 U11360 ( .C1(n10337), .C2(n8880), .A(n8879), .B(n8878), .ZN(n8881)
         );
  INV_X1 U11361 ( .A(n8881), .ZN(n8882) );
  AND2_X1 U11362 ( .A1(n10340), .A2(n8882), .ZN(n11958) );
  INV_X1 U11363 ( .A(P3_B_REG_SCAN_IN), .ZN(n8884) );
  NOR2_X1 U11364 ( .A1(n11081), .A2(n8884), .ZN(n8885) );
  OR2_X1 U11365 ( .A1(n12408), .A2(n8885), .ZN(n12283) );
  OAI22_X1 U11366 ( .A1(n11666), .A2(n12406), .B1(n11958), .B2(n12283), .ZN(
        n8886) );
  AOI21_X2 U11367 ( .B1(n8887), .B2(n12474), .A(n8886), .ZN(n11614) );
  OAI21_X1 U11368 ( .B1(n12500), .B2(n11621), .A(n11614), .ZN(n8942) );
  INV_X1 U11369 ( .A(n8888), .ZN(n8897) );
  NAND2_X1 U11370 ( .A1(n8897), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8889) );
  MUX2_X1 U11371 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8889), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8891) );
  NAND2_X1 U11372 ( .A1(n8892), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8893) );
  MUX2_X1 U11373 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8893), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8895) );
  NAND2_X1 U11374 ( .A1(n8895), .A2(n6742), .ZN(n10547) );
  XNOR2_X1 U11375 ( .A(n10547), .B(P3_B_REG_SCAN_IN), .ZN(n8899) );
  NAND2_X1 U11376 ( .A1(n6742), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8896) );
  MUX2_X1 U11377 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8896), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8898) );
  NAND2_X1 U11378 ( .A1(n8898), .A2(n8897), .ZN(n10682) );
  NAND2_X1 U11379 ( .A1(n8899), .A2(n10682), .ZN(n8900) );
  NAND2_X1 U11380 ( .A1(n10875), .A2(n10547), .ZN(n8901) );
  INV_X1 U11381 ( .A(n8915), .ZN(n9336) );
  INV_X1 U11382 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U11383 ( .A1(n9336), .A2(n9111), .ZN(n8904) );
  NAND2_X1 U11384 ( .A1(n10875), .A2(n10682), .ZN(n8903) );
  XNOR2_X1 U11385 ( .A(n12616), .B(n10235), .ZN(n8923) );
  NOR3_X1 U11386 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .ZN(n13799) );
  NOR3_X1 U11387 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .A3(
        P3_D_REG_8__SCAN_IN), .ZN(n8907) );
  NOR4_X1 U11388 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n8906) );
  NOR4_X1 U11389 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8905) );
  NAND4_X1 U11390 ( .A1(n13799), .A2(n8907), .A3(n8906), .A4(n8905), .ZN(n8913) );
  NOR4_X1 U11391 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8911) );
  NOR4_X1 U11392 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n8910) );
  NOR4_X1 U11393 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8909) );
  NOR4_X1 U11394 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8908) );
  NAND4_X1 U11395 ( .A1(n8911), .A2(n8910), .A3(n8909), .A4(n8908), .ZN(n8912)
         );
  NOR2_X1 U11396 ( .A1(n8913), .A2(n8912), .ZN(n8914) );
  NOR2_X1 U11397 ( .A1(n10682), .A2(n10547), .ZN(n8916) );
  INV_X1 U11398 ( .A(n8918), .ZN(n8919) );
  NAND2_X1 U11399 ( .A1(n8919), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8920) );
  MUX2_X1 U11400 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8920), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8921) );
  NAND2_X1 U11401 ( .A1(n8921), .A2(n8892), .ZN(n9536) );
  INV_X1 U11402 ( .A(n12615), .ZN(n9110) );
  AND2_X1 U11403 ( .A1(n8936), .A2(n12159), .ZN(n8922) );
  NAND2_X1 U11404 ( .A1(n12152), .A2(n12103), .ZN(n10231) );
  NAND2_X1 U11405 ( .A1(n8924), .A2(n12129), .ZN(n10233) );
  AND2_X1 U11406 ( .A1(n10231), .A2(n10233), .ZN(n8928) );
  OAI22_X1 U11407 ( .A1(n15515), .A2(n8933), .B1(n12268), .B2(n8925), .ZN(
        n8926) );
  AOI21_X1 U11408 ( .B1(n8926), .B2(n12152), .A(n12103), .ZN(n8927) );
  MUX2_X1 U11409 ( .A(n8928), .B(n8927), .S(n10235), .Z(n8929) );
  MUX2_X1 U11410 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n8942), .S(n15540), .Z(
        n8930) );
  INV_X1 U11411 ( .A(n8930), .ZN(n8932) );
  INV_X1 U11412 ( .A(n8931), .ZN(n11617) );
  NAND2_X1 U11413 ( .A1(n8932), .A2(n7696), .ZN(P3_U3488) );
  INV_X1 U11414 ( .A(n10235), .ZN(n9108) );
  NAND2_X1 U11415 ( .A1(n11990), .A2(n8933), .ZN(n12155) );
  OR2_X1 U11416 ( .A1(n8934), .A2(n12155), .ZN(n9744) );
  OAI21_X1 U11417 ( .B1(n12129), .B2(n12152), .A(n9744), .ZN(n8935) );
  NAND2_X1 U11418 ( .A1(n9752), .A2(n8935), .ZN(n8940) );
  INV_X1 U11419 ( .A(n8936), .ZN(n8937) );
  NOR2_X1 U11420 ( .A1(n12616), .A2(n8937), .ZN(n8938) );
  AND2_X1 U11421 ( .A1(n8938), .A2(n10235), .ZN(n9750) );
  NAND2_X1 U11422 ( .A1(n9750), .A2(n9736), .ZN(n8939) );
  NAND2_X1 U11423 ( .A1(n8940), .A2(n8939), .ZN(n8941) );
  MUX2_X1 U11424 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n8942), .S(n15519), .Z(
        n8943) );
  INV_X1 U11425 ( .A(n8943), .ZN(n8944) );
  NAND2_X1 U11426 ( .A1(n15519), .A2(n15508), .ZN(n12613) );
  NAND2_X1 U11427 ( .A1(n8944), .A2(n7695), .ZN(P3_U3456) );
  INV_X1 U11428 ( .A(n11819), .ZN(n8956) );
  NAND2_X1 U11429 ( .A1(n11584), .A2(n8945), .ZN(n8946) );
  NAND2_X1 U11430 ( .A1(n12303), .A2(n11593), .ZN(n8948) );
  NAND2_X1 U11431 ( .A1(n8948), .A2(n8947), .ZN(n8950) );
  INV_X1 U11432 ( .A(n11984), .ZN(n8949) );
  AOI21_X1 U11433 ( .B1(n8950), .B2(n8949), .A(n12404), .ZN(n8955) );
  AND2_X1 U11434 ( .A1(n8952), .A2(n8951), .ZN(n8954) );
  OAI22_X1 U11435 ( .A1(n11814), .A2(n12408), .B1(n11923), .B2(n12406), .ZN(
        n8953) );
  OAI21_X1 U11436 ( .B1(n11581), .B2(n12500), .A(n11577), .ZN(n8957) );
  NAND2_X1 U11437 ( .A1(n8966), .A2(n8965), .ZN(n9205) );
  INV_X1 U11438 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8970) );
  NOR2_X1 U11439 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8972) );
  NOR3_X1 U11440 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .A3(P2_IR_REG_21__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U11441 ( .A1(n8979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8978) );
  MUX2_X1 U11442 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8978), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8980) );
  NAND2_X1 U11443 ( .A1(n8980), .A2(n9211), .ZN(n13900) );
  NAND2_X1 U11444 ( .A1(n8981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8982) );
  MUX2_X1 U11445 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8982), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8983) );
  NAND2_X1 U11446 ( .A1(n8983), .A2(n8979), .ZN(n13902) );
  NOR2_X1 U11447 ( .A1(n13900), .A2(n13902), .ZN(n8984) );
  NAND2_X1 U11448 ( .A1(n13904), .A2(n8984), .ZN(n9263) );
  XNOR2_X1 U11449 ( .A(n8986), .B(n8985), .ZN(n9262) );
  INV_X1 U11450 ( .A(n9262), .ZN(n11179) );
  NOR2_X1 U11451 ( .A1(n9263), .A2(n11179), .ZN(n9214) );
  INV_X1 U11452 ( .A(n9102), .ZN(n8987) );
  OR2_X2 U11453 ( .A1(n10044), .A2(n8987), .ZN(n14337) );
  AND2_X1 U11454 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14340) );
  INV_X1 U11455 ( .A(n14340), .ZN(n8994) );
  INV_X1 U11456 ( .A(n14103), .ZN(n9765) );
  NAND2_X2 U11457 ( .A1(n10044), .A2(n9765), .ZN(n11798) );
  INV_X1 U11458 ( .A(n10044), .ZN(n8992) );
  OR2_X1 U11459 ( .A1(n8991), .A2(n11798), .ZN(n8993) );
  OAI21_X1 U11460 ( .B1(n6717), .B2(n9605), .A(n9604), .ZN(n9394) );
  MUX2_X1 U11461 ( .A(n8994), .B(n9394), .S(n6560), .Z(n8997) );
  NOR2_X1 U11462 ( .A1(n6560), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8995) );
  OR2_X1 U11463 ( .A1(n11338), .A2(n8995), .ZN(n14999) );
  AOI21_X1 U11464 ( .B1(n7503), .B2(n14999), .A(n14337), .ZN(n8996) );
  OAI21_X1 U11465 ( .B1(n8997), .B2(n11338), .A(n8996), .ZN(n14363) );
  INV_X1 U11466 ( .A(n14363), .ZN(n9028) );
  NAND2_X1 U11467 ( .A1(n8998), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14311) );
  NAND2_X1 U11468 ( .A1(n9395), .A2(n14311), .ZN(n9003) );
  OR2_X1 U11469 ( .A1(n14092), .A2(n8998), .ZN(n9000) );
  AND2_X1 U11470 ( .A1(n9000), .A2(n8999), .ZN(n9002) );
  INV_X1 U11471 ( .A(n9002), .ZN(n9001) );
  NAND2_X1 U11472 ( .A1(n9003), .A2(n9002), .ZN(n15004) );
  OR2_X1 U11473 ( .A1(n11338), .A2(n6560), .ZN(n9004) );
  OR2_X1 U11474 ( .A1(n15004), .A2(n9004), .ZN(n15025) );
  MUX2_X1 U11475 ( .A(n9006), .B(P1_REG2_REG_2__SCAN_IN), .S(n14351), .Z(
        n14359) );
  XNOR2_X1 U11476 ( .A(n14342), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n14341) );
  NAND2_X1 U11477 ( .A1(n14341), .A2(n14340), .ZN(n14339) );
  INV_X1 U11478 ( .A(n14342), .ZN(n14346) );
  NAND2_X1 U11479 ( .A1(n14346), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U11480 ( .A1(n14339), .A2(n9005), .ZN(n14358) );
  AND2_X1 U11481 ( .A1(n14359), .A2(n14358), .ZN(n14376) );
  NOR2_X1 U11482 ( .A1(n14351), .A2(n9006), .ZN(n14375) );
  MUX2_X1 U11483 ( .A(n10100), .B(P1_REG2_REG_3__SCAN_IN), .S(n14368), .Z(
        n14374) );
  OAI21_X1 U11484 ( .B1(n14376), .B2(n14375), .A(n14374), .ZN(n14378) );
  INV_X1 U11485 ( .A(n14368), .ZN(n14367) );
  NAND2_X1 U11486 ( .A1(n14367), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9008) );
  MUX2_X1 U11487 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9763), .S(n9116), .Z(n9007)
         );
  AOI21_X1 U11488 ( .B1(n14378), .B2(n9008), .A(n9007), .ZN(n9119) );
  INV_X1 U11489 ( .A(n9119), .ZN(n9010) );
  NAND3_X1 U11490 ( .A1(n14378), .A2(n9008), .A3(n9007), .ZN(n9009) );
  NAND3_X1 U11491 ( .A1(n15040), .A2(n9010), .A3(n9009), .ZN(n9011) );
  NAND2_X1 U11492 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10050) );
  OAI211_X1 U11493 ( .C1(n6823), .C2(n15047), .A(n9011), .B(n10050), .ZN(n9027) );
  OR2_X1 U11494 ( .A1(n15004), .A2(n9012), .ZN(n15029) );
  MUX2_X1 U11496 ( .A(n9017), .B(P1_REG1_REG_2__SCAN_IN), .S(n14351), .Z(
        n14356) );
  MUX2_X1 U11497 ( .A(n9013), .B(P1_REG1_REG_1__SCAN_IN), .S(n14342), .Z(n9015) );
  AND2_X1 U11498 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9014) );
  NAND2_X1 U11499 ( .A1(n9015), .A2(n9014), .ZN(n14345) );
  NAND2_X1 U11500 ( .A1(n14346), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9016) );
  NAND2_X1 U11501 ( .A1(n14345), .A2(n9016), .ZN(n14355) );
  NAND2_X1 U11502 ( .A1(n14356), .A2(n14355), .ZN(n14371) );
  OR2_X1 U11503 ( .A1(n14351), .A2(n9017), .ZN(n14370) );
  NAND2_X1 U11504 ( .A1(n14371), .A2(n14370), .ZN(n9019) );
  MUX2_X1 U11505 ( .A(n9020), .B(P1_REG1_REG_3__SCAN_IN), .S(n14368), .Z(n9018) );
  NAND2_X1 U11506 ( .A1(n9019), .A2(n9018), .ZN(n14373) );
  OR2_X1 U11507 ( .A1(n14368), .A2(n9020), .ZN(n9021) );
  MUX2_X1 U11508 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7917), .S(n9116), .Z(n9022)
         );
  AOI21_X1 U11509 ( .B1(n14373), .B2(n9021), .A(n9022), .ZN(n9112) );
  INV_X1 U11510 ( .A(n9112), .ZN(n9024) );
  NAND3_X1 U11511 ( .A1(n14373), .A2(n9022), .A3(n9021), .ZN(n9023) );
  NAND2_X1 U11512 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  OAI22_X1 U11513 ( .A1(n9116), .A2(n15029), .B1(n15027), .B2(n9025), .ZN(
        n9026) );
  OR3_X1 U11514 ( .A1(n9028), .A2(n9027), .A3(n9026), .ZN(P1_U3247) );
  NOR2_X1 U11515 ( .A1(n13064), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12617) );
  MUX2_X1 U11516 ( .A(n9302), .B(n9648), .S(P3_STATE_REG_SCAN_IN), .Z(n9029)
         );
  OAI21_X1 U11517 ( .B1(n9030), .B2(n12627), .A(n9029), .ZN(P3_U3295) );
  OAI222_X1 U11518 ( .A1(P3_U3151), .A2(n10172), .B1(n12627), .B2(n9032), .C1(
        n9031), .C2(n12623), .ZN(P3_U3289) );
  INV_X1 U11519 ( .A(n9033), .ZN(n9035) );
  INV_X1 U11520 ( .A(SI_3_), .ZN(n9034) );
  OAI222_X1 U11521 ( .A1(n7338), .A2(P3_U3151), .B1(n12627), .B2(n9035), .C1(
        n9034), .C2(n12623), .ZN(P3_U3292) );
  INV_X1 U11522 ( .A(n9664), .ZN(n9670) );
  INV_X1 U11523 ( .A(n9036), .ZN(n9037) );
  INV_X1 U11524 ( .A(SI_2_), .ZN(n13830) );
  OAI222_X1 U11525 ( .A1(n9670), .A2(P3_U3151), .B1(n12627), .B2(n9037), .C1(
        n13830), .C2(n12623), .ZN(P3_U3293) );
  NAND2_X1 U11526 ( .A1(n13064), .A2(P1_U3086), .ZN(n14755) );
  AND2_X1 U11527 ( .A1(n9293), .A2(P1_U3086), .ZN(n11176) );
  INV_X2 U11528 ( .A(n11176), .ZN(n14753) );
  OAI222_X1 U11529 ( .A1(n14755), .A2(n9038), .B1(n14753), .B2(n9292), .C1(
        P1_U3086), .C2(n14342), .ZN(P1_U3354) );
  OAI222_X1 U11530 ( .A1(P3_U3151), .A2(n10631), .B1(n12627), .B2(n9040), .C1(
        n9039), .C2(n12623), .ZN(P3_U3287) );
  INV_X1 U11531 ( .A(SI_5_), .ZN(n9043) );
  INV_X1 U11532 ( .A(n9041), .ZN(n9042) );
  OAI222_X1 U11533 ( .A1(P3_U3151), .A2(n9895), .B1(n12623), .B2(n9043), .C1(
        n12627), .C2(n9042), .ZN(P3_U3290) );
  NOR2_X1 U11534 ( .A1(n13064), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13890) );
  INV_X2 U11535 ( .A(n13890), .ZN(n13905) );
  AND2_X1 U11536 ( .A1(n13064), .A2(P2_U3088), .ZN(n13893) );
  INV_X2 U11537 ( .A(n13893), .ZN(n13908) );
  OR2_X1 U11538 ( .A1(n9044), .A2(n13881), .ZN(n9046) );
  XNOR2_X1 U11539 ( .A(n9046), .B(n9045), .ZN(n9456) );
  OAI222_X1 U11540 ( .A1(n13905), .A2(n9453), .B1(n13908), .B2(n9452), .C1(
        P2_U3088), .C2(n9456), .ZN(P2_U3325) );
  NAND2_X1 U11541 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9047) );
  INV_X1 U11542 ( .A(n9781), .ZN(n9055) );
  OR2_X1 U11543 ( .A1(n9049), .A2(n13881), .ZN(n9050) );
  XNOR2_X1 U11544 ( .A(n9050), .B(n9057), .ZN(n15224) );
  OAI222_X1 U11545 ( .A1(n13905), .A2(n9782), .B1(n13908), .B2(n9055), .C1(
        P2_U3088), .C2(n15224), .ZN(P2_U3324) );
  INV_X1 U11546 ( .A(SI_9_), .ZN(n9053) );
  INV_X1 U11547 ( .A(n9051), .ZN(n9052) );
  OAI222_X1 U11548 ( .A1(P3_U3151), .A2(n15453), .B1(n12623), .B2(n9053), .C1(
        n12627), .C2(n9052), .ZN(P3_U3286) );
  INV_X1 U11549 ( .A(n14755), .ZN(n14739) );
  INV_X1 U11550 ( .A(n14739), .ZN(n11330) );
  OAI222_X1 U11551 ( .A1(n11330), .A2(n9054), .B1(n14753), .B2(n9452), .C1(
        P1_U3086), .C2(n14351), .ZN(P1_U3353) );
  OAI222_X1 U11552 ( .A1(n11330), .A2(n9056), .B1(n14753), .B2(n9055), .C1(
        P1_U3086), .C2(n14368), .ZN(P1_U3352) );
  INV_X1 U11553 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9061) );
  INV_X1 U11554 ( .A(n9950), .ZN(n9062) );
  NAND2_X1 U11555 ( .A1(n9049), .A2(n9057), .ZN(n9059) );
  NAND2_X1 U11556 ( .A1(n9059), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9058) );
  MUX2_X1 U11557 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9058), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9060) );
  AND2_X1 U11558 ( .A1(n9060), .A2(n9374), .ZN(n9951) );
  INV_X1 U11559 ( .A(n9951), .ZN(n15236) );
  OAI222_X1 U11560 ( .A1(n13905), .A2(n9061), .B1(n13908), .B2(n9062), .C1(
        P2_U3088), .C2(n15236), .ZN(P2_U3323) );
  OAI222_X1 U11561 ( .A1(n11330), .A2(n9063), .B1(n14753), .B2(n9062), .C1(
        P1_U3086), .C2(n9116), .ZN(P1_U3351) );
  INV_X1 U11562 ( .A(n9816), .ZN(n9821) );
  INV_X1 U11563 ( .A(SI_4_), .ZN(n9066) );
  INV_X1 U11564 ( .A(n9064), .ZN(n9065) );
  OAI222_X1 U11565 ( .A1(P3_U3151), .A2(n9821), .B1(n12623), .B2(n9066), .C1(
        n12627), .C2(n9065), .ZN(P3_U3291) );
  OAI222_X1 U11566 ( .A1(n12627), .A2(n9068), .B1(n12623), .B2(n9067), .C1(
        P3_U3151), .C2(n9546), .ZN(P3_U3294) );
  INV_X1 U11567 ( .A(n9069), .ZN(n9071) );
  INV_X1 U11568 ( .A(SI_7_), .ZN(n9070) );
  OAI222_X1 U11569 ( .A1(n10259), .A2(P3_U3151), .B1(n12627), .B2(n9071), .C1(
        n9070), .C2(n12623), .ZN(P3_U3288) );
  INV_X1 U11570 ( .A(n9072), .ZN(n9073) );
  OAI222_X1 U11571 ( .A1(P3_U3151), .A2(n10802), .B1(n12623), .B2(n13829), 
        .C1(n12627), .C2(n9073), .ZN(P3_U3285) );
  INV_X1 U11572 ( .A(n9957), .ZN(n9076) );
  INV_X1 U11573 ( .A(n9138), .ZN(n9126) );
  OAI222_X1 U11574 ( .A1(n11330), .A2(n9074), .B1(n14753), .B2(n9076), .C1(
        P1_U3086), .C2(n9126), .ZN(P1_U3350) );
  INV_X1 U11575 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U11576 ( .A1(n9374), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9075) );
  XNOR2_X1 U11577 ( .A(n9075), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9958) );
  INV_X1 U11578 ( .A(n9958), .ZN(n9441) );
  OAI222_X1 U11579 ( .A1(n13905), .A2(n9077), .B1(n13908), .B2(n9076), .C1(
        P2_U3088), .C2(n9441), .ZN(P2_U3322) );
  INV_X1 U11580 ( .A(n9078), .ZN(n9079) );
  OAI222_X1 U11581 ( .A1(P3_U3151), .A2(n10929), .B1(n12623), .B2(n9080), .C1(
        n12627), .C2(n9079), .ZN(P3_U3284) );
  INV_X1 U11582 ( .A(n9971), .ZN(n9085) );
  INV_X1 U11583 ( .A(n9374), .ZN(n9082) );
  INV_X1 U11584 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U11585 ( .A1(n9082), .A2(n9081), .ZN(n9088) );
  NAND2_X1 U11586 ( .A1(n9088), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9083) );
  XNOR2_X1 U11587 ( .A(n9083), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9972) );
  INV_X1 U11588 ( .A(n9972), .ZN(n9428) );
  OAI222_X1 U11589 ( .A1(n13905), .A2(n9084), .B1(n13908), .B2(n9085), .C1(
        P2_U3088), .C2(n9428), .ZN(P2_U3321) );
  INV_X1 U11590 ( .A(n9139), .ZN(n9156) );
  OAI222_X1 U11591 ( .A1(n11330), .A2(n13630), .B1(n14753), .B2(n9085), .C1(
        P1_U3086), .C2(n9156), .ZN(P1_U3349) );
  OAI222_X1 U11592 ( .A1(P3_U3151), .A2(n11230), .B1(n12623), .B2(n13820), 
        .C1(n12627), .C2(n9086), .ZN(P3_U3283) );
  NOR2_X1 U11593 ( .A1(n15006), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11594 ( .A(n9984), .ZN(n9093) );
  INV_X1 U11595 ( .A(n14391), .ZN(n9151) );
  OAI222_X1 U11596 ( .A1(n11330), .A2(n9087), .B1(n14753), .B2(n9093), .C1(
        P1_U3086), .C2(n9151), .ZN(P1_U3348) );
  INV_X1 U11597 ( .A(n9088), .ZN(n9090) );
  NAND2_X1 U11598 ( .A1(n9090), .A2(n9089), .ZN(n9095) );
  NAND2_X1 U11599 ( .A1(n9095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9091) );
  XNOR2_X1 U11600 ( .A(n9091), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13220) );
  INV_X1 U11601 ( .A(n13220), .ZN(n9092) );
  OAI222_X1 U11602 ( .A1(n13905), .A2(n9094), .B1(n13908), .B2(n9093), .C1(
        P2_U3088), .C2(n9092), .ZN(P2_U3320) );
  INV_X1 U11603 ( .A(n9997), .ZN(n9098) );
  NAND2_X1 U11604 ( .A1(n9129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9096) );
  XNOR2_X1 U11605 ( .A(n9096), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9998) );
  INV_X1 U11606 ( .A(n9998), .ZN(n9097) );
  OAI222_X1 U11607 ( .A1(n13905), .A2(n13821), .B1(n13908), .B2(n9098), .C1(
        P2_U3088), .C2(n9097), .ZN(P2_U3319) );
  INV_X1 U11608 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9099) );
  INV_X1 U11609 ( .A(n9175), .ZN(n9166) );
  OAI222_X1 U11610 ( .A1(n11330), .A2(n9099), .B1(n14753), .B2(n9098), .C1(
        P1_U3086), .C2(n9166), .ZN(P1_U3347) );
  INV_X1 U11611 ( .A(n9395), .ZN(n9101) );
  AND2_X2 U11612 ( .A1(n9101), .A2(n9100), .ZN(n15137) );
  INV_X1 U11613 ( .A(n14751), .ZN(n9103) );
  NAND2_X1 U11614 ( .A1(n9102), .A2(n14748), .ZN(n9105) );
  OAI22_X1 U11615 ( .A1(n15137), .A2(P1_D_REG_1__SCAN_IN), .B1(n9103), .B2(
        n9105), .ZN(n9104) );
  INV_X1 U11616 ( .A(n9104), .ZN(P1_U3446) );
  INV_X1 U11617 ( .A(n7730), .ZN(n9106) );
  OAI22_X1 U11618 ( .A1(n15137), .A2(P1_D_REG_0__SCAN_IN), .B1(n9106), .B2(
        n9105), .ZN(n9107) );
  INV_X1 U11619 ( .A(n9107), .ZN(P1_U3445) );
  NAND2_X1 U11620 ( .A1(n9108), .A2(n9110), .ZN(n9109) );
  OAI21_X1 U11621 ( .B1(n9111), .B2(n9110), .A(n9109), .ZN(P3_U3377) );
  MUX2_X1 U11622 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7933), .S(n9138), .Z(n9115)
         );
  AOI21_X1 U11623 ( .B1(n9113), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9112), .ZN(
        n9114) );
  NAND2_X1 U11624 ( .A1(n9114), .A2(n9115), .ZN(n9135) );
  OAI21_X1 U11625 ( .B1(n9115), .B2(n9114), .A(n9135), .ZN(n9123) );
  NOR2_X1 U11626 ( .A1(n9116), .A2(n9763), .ZN(n9118) );
  MUX2_X1 U11627 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9935), .S(n9138), .Z(n9117)
         );
  OAI21_X1 U11628 ( .B1(n9119), .B2(n9118), .A(n9117), .ZN(n9142) );
  INV_X1 U11629 ( .A(n9142), .ZN(n9121) );
  NOR3_X1 U11630 ( .A1(n9119), .A2(n9118), .A3(n9117), .ZN(n9120) );
  NOR3_X1 U11631 ( .A1(n15025), .A2(n9121), .A3(n9120), .ZN(n9122) );
  AOI21_X1 U11632 ( .B1(n15035), .B2(n9123), .A(n9122), .ZN(n9125) );
  AND2_X1 U11633 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10194) );
  AOI21_X1 U11634 ( .B1(n15006), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10194), .ZN(
        n9124) );
  OAI211_X1 U11635 ( .C1(n9126), .C2(n15029), .A(n9125), .B(n9124), .ZN(
        P1_U3248) );
  OAI222_X1 U11636 ( .A1(P3_U3151), .A2(n11257), .B1(n12623), .B2(n9128), .C1(
        n12627), .C2(n9127), .ZN(P3_U3282) );
  INV_X1 U11637 ( .A(n10128), .ZN(n9133) );
  OAI21_X1 U11638 ( .B1(n9129), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9130) );
  XNOR2_X1 U11639 ( .A(n9130), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10129) );
  INV_X1 U11640 ( .A(n10129), .ZN(n9383) );
  OAI222_X1 U11641 ( .A1(n13905), .A2(n9131), .B1(n13908), .B2(n9133), .C1(
        P2_U3088), .C2(n9383), .ZN(P2_U3318) );
  INV_X1 U11642 ( .A(n9188), .ZN(n9132) );
  OAI222_X1 U11643 ( .A1(n11330), .A2(n9134), .B1(n14753), .B2(n9133), .C1(
        P1_U3086), .C2(n9132), .ZN(P1_U3346) );
  OAI21_X1 U11644 ( .B1(n9138), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9135), .ZN(
        n9137) );
  MUX2_X1 U11645 ( .A(n9149), .B(P1_REG1_REG_6__SCAN_IN), .S(n9139), .Z(n9136)
         );
  NOR2_X1 U11646 ( .A1(n9137), .A2(n9136), .ZN(n14396) );
  AOI211_X1 U11647 ( .C1(n9137), .C2(n9136), .A(n15027), .B(n14396), .ZN(n9145) );
  NAND2_X1 U11648 ( .A1(n9138), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9141) );
  MUX2_X1 U11649 ( .A(n9858), .B(P1_REG2_REG_6__SCAN_IN), .S(n9139), .Z(n9140)
         );
  AOI21_X1 U11650 ( .B1(n9142), .B2(n9141), .A(n9140), .ZN(n14389) );
  AND3_X1 U11651 ( .A1(n9142), .A2(n9141), .A3(n9140), .ZN(n9143) );
  NOR3_X1 U11652 ( .A1(n15025), .A2(n14389), .A3(n9143), .ZN(n9144) );
  NOR2_X1 U11653 ( .A1(n9145), .A2(n9144), .ZN(n9147) );
  AND2_X1 U11654 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10313) );
  AOI21_X1 U11655 ( .B1(n15006), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10313), .ZN(
        n9146) );
  OAI211_X1 U11656 ( .C1(n9156), .C2(n15029), .A(n9147), .B(n9146), .ZN(
        P1_U3249) );
  MUX2_X1 U11657 ( .A(n9148), .B(P1_REG1_REG_8__SCAN_IN), .S(n9175), .Z(n9153)
         );
  INV_X1 U11658 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15202) );
  NOR2_X1 U11659 ( .A1(n9156), .A2(n9149), .ZN(n14390) );
  MUX2_X1 U11660 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n15202), .S(n14391), .Z(
        n9150) );
  OAI21_X1 U11661 ( .B1(n14396), .B2(n14390), .A(n9150), .ZN(n14394) );
  OAI21_X1 U11662 ( .B1(n15202), .B2(n9151), .A(n14394), .ZN(n9152) );
  NOR2_X1 U11663 ( .A1(n9152), .A2(n9153), .ZN(n9178) );
  AOI21_X1 U11664 ( .B1(n9153), .B2(n9152), .A(n9178), .ZN(n9165) );
  NOR2_X1 U11665 ( .A1(n9154), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10701) );
  NOR2_X1 U11666 ( .A1(n15029), .A2(n9166), .ZN(n9155) );
  AOI211_X1 U11667 ( .C1(n15006), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10701), .B(
        n9155), .ZN(n9164) );
  NOR2_X1 U11668 ( .A1(n9156), .A2(n9858), .ZN(n14384) );
  MUX2_X1 U11669 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9157), .S(n14391), .Z(n9158) );
  OAI21_X1 U11670 ( .B1(n14389), .B2(n14384), .A(n9158), .ZN(n14387) );
  NAND2_X1 U11671 ( .A1(n14391), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9160) );
  MUX2_X1 U11672 ( .A(n7979), .B(P1_REG2_REG_8__SCAN_IN), .S(n9175), .Z(n9159)
         );
  AOI21_X1 U11673 ( .B1(n14387), .B2(n9160), .A(n9159), .ZN(n9170) );
  INV_X1 U11674 ( .A(n9170), .ZN(n9162) );
  NAND3_X1 U11675 ( .A1(n14387), .A2(n9160), .A3(n9159), .ZN(n9161) );
  NAND3_X1 U11676 ( .A1(n9162), .A2(n15040), .A3(n9161), .ZN(n9163) );
  OAI211_X1 U11677 ( .C1(n9165), .C2(n15027), .A(n9164), .B(n9163), .ZN(
        P1_U3251) );
  INV_X1 U11678 ( .A(n15029), .ZN(n15038) );
  INV_X1 U11679 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14780) );
  NAND2_X1 U11680 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10884) );
  OAI21_X1 U11681 ( .B1(n15047), .B2(n14780), .A(n10884), .ZN(n9174) );
  NOR2_X1 U11682 ( .A1(n9166), .A2(n7979), .ZN(n9169) );
  MUX2_X1 U11683 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9167), .S(n9188), .Z(n9168)
         );
  OAI21_X1 U11684 ( .B1(n9170), .B2(n9169), .A(n9168), .ZN(n9191) );
  INV_X1 U11685 ( .A(n9191), .ZN(n9172) );
  NOR3_X1 U11686 ( .A1(n9170), .A2(n9169), .A3(n9168), .ZN(n9171) );
  NOR3_X1 U11687 ( .A1(n9172), .A2(n9171), .A3(n15025), .ZN(n9173) );
  AOI211_X1 U11688 ( .C1(n15038), .C2(n9188), .A(n9174), .B(n9173), .ZN(n9182)
         );
  NOR2_X1 U11689 ( .A1(n9175), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9176) );
  MUX2_X1 U11690 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7993), .S(n9188), .Z(n9177)
         );
  OAI21_X1 U11691 ( .B1(n9178), .B2(n9176), .A(n9177), .ZN(n9185) );
  INV_X1 U11692 ( .A(n9185), .ZN(n9180) );
  NOR3_X1 U11693 ( .A1(n9178), .A2(n9177), .A3(n9176), .ZN(n9179) );
  OAI21_X1 U11694 ( .B1(n9180), .B2(n9179), .A(n15035), .ZN(n9181) );
  NAND2_X1 U11695 ( .A1(n9182), .A2(n9181), .ZN(P1_U3252) );
  OAI222_X1 U11696 ( .A1(n11225), .A2(P3_U3151), .B1(n12627), .B2(n9184), .C1(
        n9183), .C2(n12623), .ZN(P3_U3281) );
  OAI21_X1 U11697 ( .B1(n9188), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9185), .ZN(
        n9187) );
  INV_X1 U11698 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15207) );
  MUX2_X1 U11699 ( .A(n15207), .B(P1_REG1_REG_10__SCAN_IN), .S(n9408), .Z(
        n9186) );
  NOR2_X1 U11700 ( .A1(n9187), .A2(n9186), .ZN(n9407) );
  AOI211_X1 U11701 ( .C1(n9187), .C2(n9186), .A(n15027), .B(n9407), .ZN(n9197)
         );
  INV_X1 U11702 ( .A(n9408), .ZN(n9447) );
  NAND2_X1 U11703 ( .A1(n9188), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9190) );
  MUX2_X1 U11704 ( .A(n9403), .B(P1_REG2_REG_10__SCAN_IN), .S(n9408), .Z(n9189) );
  AOI21_X1 U11705 ( .B1(n9191), .B2(n9190), .A(n9189), .ZN(n14409) );
  INV_X1 U11706 ( .A(n14409), .ZN(n9193) );
  NAND3_X1 U11707 ( .A1(n9191), .A2(n9190), .A3(n9189), .ZN(n9192) );
  NAND3_X1 U11708 ( .A1(n9193), .A2(n15040), .A3(n9192), .ZN(n9195) );
  AND2_X1 U11709 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11125) );
  AOI21_X1 U11710 ( .B1(n15006), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11125), 
        .ZN(n9194) );
  OAI211_X1 U11711 ( .C1(n15029), .C2(n9447), .A(n9195), .B(n9194), .ZN(n9196)
         );
  OR2_X1 U11712 ( .A1(n9197), .A2(n9196), .ZN(P1_U3253) );
  INV_X1 U11713 ( .A(n15224), .ZN(n9229) );
  INV_X1 U11714 ( .A(n9456), .ZN(n9226) );
  INV_X1 U11715 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13474) );
  NAND3_X1 U11716 ( .A1(n15213), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n15212) );
  NAND2_X1 U11717 ( .A1(n9224), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9246) );
  INV_X1 U11718 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10500) );
  MUX2_X1 U11719 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10500), .S(n9456), .Z(n9247) );
  INV_X1 U11720 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9198) );
  MUX2_X1 U11721 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9198), .S(n15224), .Z(
        n15230) );
  INV_X1 U11722 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9199) );
  MUX2_X1 U11723 ( .A(n9199), .B(P2_REG2_REG_4__SCAN_IN), .S(n9951), .Z(n15244) );
  NOR2_X1 U11724 ( .A1(n15245), .A2(n15244), .ZN(n15243) );
  AND2_X1 U11725 ( .A1(n9951), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9435) );
  INV_X1 U11726 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10424) );
  MUX2_X1 U11727 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10424), .S(n9958), .Z(n9434) );
  OAI21_X1 U11728 ( .B1(n15243), .B2(n9435), .A(n9434), .ZN(n9433) );
  NAND2_X1 U11729 ( .A1(n9958), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9423) );
  INV_X1 U11730 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9200) );
  MUX2_X1 U11731 ( .A(n9200), .B(P2_REG2_REG_6__SCAN_IN), .S(n9972), .Z(n9422)
         );
  AOI21_X1 U11732 ( .B1(n9433), .B2(n9423), .A(n9422), .ZN(n13216) );
  NOR2_X1 U11733 ( .A1(n9428), .A2(n9200), .ZN(n13215) );
  INV_X1 U11734 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9201) );
  MUX2_X1 U11735 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9201), .S(n13220), .Z(
        n13214) );
  NAND2_X1 U11736 ( .A1(n13220), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9204) );
  INV_X1 U11737 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9202) );
  MUX2_X1 U11738 ( .A(n9202), .B(P2_REG2_REG_8__SCAN_IN), .S(n9998), .Z(n9203)
         );
  NAND3_X1 U11739 ( .A1(n13213), .A2(n9204), .A3(n9203), .ZN(n9217) );
  NAND2_X1 U11740 ( .A1(n9205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9207) );
  INV_X1 U11741 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9206) );
  XNOR2_X1 U11742 ( .A(n9207), .B(n9206), .ZN(n12867) );
  NAND2_X1 U11743 ( .A1(n9208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9209) );
  XNOR2_X2 U11744 ( .A(n9210), .B(n9279), .ZN(n9215) );
  AOI21_X1 U11745 ( .B1(n9805), .B2(n9262), .A(n11381), .ZN(n9213) );
  OR2_X1 U11746 ( .A1(n9214), .A2(n9213), .ZN(n9222) );
  INV_X1 U11747 ( .A(n9220), .ZN(n13169) );
  NAND2_X1 U11748 ( .A1(n13169), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13895) );
  NOR2_X1 U11749 ( .A1(n13895), .A2(n9215), .ZN(n9216) );
  NAND2_X1 U11750 ( .A1(n9217), .A2(n15296), .ZN(n9245) );
  NAND2_X1 U11751 ( .A1(n9222), .A2(n9215), .ZN(n15237) );
  INV_X1 U11752 ( .A(n15273), .ZN(n15299) );
  OR2_X1 U11753 ( .A1(n9222), .A2(P2_U3088), .ZN(n13249) );
  INV_X1 U11754 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9218) );
  NAND2_X1 U11755 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10282) );
  OAI21_X1 U11756 ( .B1(n13249), .B2(n9218), .A(n10282), .ZN(n9219) );
  AOI21_X1 U11757 ( .B1(n9998), .B2(n15299), .A(n9219), .ZN(n9244) );
  NOR2_X1 U11758 ( .A1(n9215), .A2(P2_U3088), .ZN(n13889) );
  AND2_X1 U11759 ( .A1(n13889), .A2(n9220), .ZN(n9221) );
  NAND2_X1 U11760 ( .A1(n9222), .A2(n9221), .ZN(n13239) );
  INV_X1 U11761 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9223) );
  MUX2_X1 U11762 ( .A(n9223), .B(P2_REG1_REG_3__SCAN_IN), .S(n15224), .Z(
        n15227) );
  AND2_X1 U11763 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15216) );
  NAND2_X1 U11764 ( .A1(n15217), .A2(n15216), .ZN(n15215) );
  NAND2_X1 U11765 ( .A1(n9224), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U11766 ( .A1(n15215), .A2(n9225), .ZN(n9251) );
  XNOR2_X1 U11767 ( .A(n9456), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11768 ( .A1(n9251), .A2(n9252), .ZN(n9228) );
  NAND2_X1 U11769 ( .A1(n9226), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9227) );
  NAND2_X1 U11770 ( .A1(n9228), .A2(n9227), .ZN(n15228) );
  NAND2_X1 U11771 ( .A1(n15227), .A2(n15228), .ZN(n15226) );
  NAND2_X1 U11772 ( .A1(n9229), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U11773 ( .A1(n15226), .A2(n9230), .ZN(n15241) );
  INV_X1 U11774 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9231) );
  MUX2_X1 U11775 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9231), .S(n9951), .Z(n15240) );
  NAND2_X1 U11776 ( .A1(n15241), .A2(n15240), .ZN(n15239) );
  NAND2_X1 U11777 ( .A1(n9951), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11778 ( .A1(n15239), .A2(n9232), .ZN(n9431) );
  INV_X1 U11779 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9233) );
  MUX2_X1 U11780 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9233), .S(n9958), .Z(n9430)
         );
  NAND2_X1 U11781 ( .A1(n9431), .A2(n9430), .ZN(n9429) );
  NAND2_X1 U11782 ( .A1(n9958), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U11783 ( .A1(n9429), .A2(n9234), .ZN(n9420) );
  INV_X1 U11784 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9235) );
  MUX2_X1 U11785 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9235), .S(n9972), .Z(n9419)
         );
  NAND2_X1 U11786 ( .A1(n9420), .A2(n9419), .ZN(n13223) );
  NAND2_X1 U11787 ( .A1(n9972), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13222) );
  NAND2_X1 U11788 ( .A1(n13223), .A2(n13222), .ZN(n9238) );
  INV_X1 U11789 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9236) );
  MUX2_X1 U11790 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9236), .S(n13220), .Z(n9237) );
  NAND2_X1 U11791 ( .A1(n9238), .A2(n9237), .ZN(n13225) );
  NAND2_X1 U11792 ( .A1(n13220), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9240) );
  INV_X1 U11793 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10033) );
  MUX2_X1 U11794 ( .A(n10033), .B(P2_REG1_REG_8__SCAN_IN), .S(n9998), .Z(n9239) );
  AOI21_X1 U11795 ( .B1(n13225), .B2(n9240), .A(n9239), .ZN(n9330) );
  INV_X1 U11796 ( .A(n9330), .ZN(n9242) );
  NAND3_X1 U11797 ( .A1(n13225), .A2(n9240), .A3(n9239), .ZN(n9241) );
  NAND3_X1 U11798 ( .A1(n15302), .A2(n9242), .A3(n9241), .ZN(n9243) );
  OAI211_X1 U11799 ( .C1(n9322), .C2(n9245), .A(n9244), .B(n9243), .ZN(
        P2_U3222) );
  AND3_X1 U11800 ( .A1(n9247), .A2(n15212), .A3(n9246), .ZN(n9248) );
  NOR3_X1 U11801 ( .A1(n15242), .A2(n9249), .A3(n9248), .ZN(n9250) );
  AOI21_X1 U11802 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .A(n9250), 
        .ZN(n9255) );
  INV_X1 U11803 ( .A(n13249), .ZN(n15294) );
  XOR2_X1 U11804 ( .A(n9252), .B(n9251), .Z(n9253) );
  AOI22_X1 U11805 ( .A1(n15294), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n15302), 
        .B2(n9253), .ZN(n9254) );
  OAI211_X1 U11806 ( .C1(n9456), .C2(n15273), .A(n9255), .B(n9254), .ZN(
        P2_U3216) );
  INV_X1 U11807 ( .A(P2_B_REG_SCAN_IN), .ZN(n9256) );
  XNOR2_X1 U11808 ( .A(n13904), .B(n9256), .ZN(n9257) );
  NAND2_X1 U11809 ( .A1(n9257), .A2(n13902), .ZN(n9258) );
  INV_X1 U11810 ( .A(n13900), .ZN(n9277) );
  INV_X1 U11811 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15356) );
  NAND2_X1 U11812 ( .A1(n15321), .A2(n15356), .ZN(n9260) );
  NAND2_X1 U11813 ( .A1(n13900), .A2(n13902), .ZN(n9259) );
  NAND2_X1 U11814 ( .A1(n15357), .A2(n9784), .ZN(n9275) );
  NAND2_X1 U11815 ( .A1(n6561), .A2(n13244), .ZN(n13163) );
  NAND2_X1 U11816 ( .A1(n9805), .A2(n13163), .ZN(n9786) );
  AND2_X1 U11817 ( .A1(n15358), .A2(n9786), .ZN(n9274) );
  NOR4_X1 U11818 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9272) );
  INV_X1 U11819 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15342) );
  INV_X1 U11820 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15341) );
  INV_X1 U11821 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15348) );
  INV_X1 U11822 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15345) );
  NAND4_X1 U11823 ( .A1(n15342), .A2(n15341), .A3(n15348), .A4(n15345), .ZN(
        n13841) );
  NOR4_X1 U11824 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n9268) );
  NOR4_X1 U11825 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9267) );
  NOR4_X1 U11826 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n9266) );
  NOR4_X1 U11827 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9265) );
  NAND4_X1 U11828 ( .A1(n9268), .A2(n9267), .A3(n9266), .A4(n9265), .ZN(n9269)
         );
  NOR4_X1 U11829 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        n13841), .A4(n9269), .ZN(n9271) );
  NOR4_X1 U11830 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9270) );
  NAND3_X1 U11831 ( .A1(n9272), .A2(n9271), .A3(n9270), .ZN(n9273) );
  NAND2_X1 U11832 ( .A1(n15321), .A2(n9273), .ZN(n9773) );
  NAND2_X1 U11833 ( .A1(n9274), .A2(n9773), .ZN(n10343) );
  OR2_X1 U11834 ( .A1(n9275), .A2(n10343), .ZN(n9943) );
  INV_X1 U11835 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11836 ( .A1(n15321), .A2(n9276), .ZN(n9278) );
  OR2_X1 U11837 ( .A1(n13904), .A2(n9277), .ZN(n15354) );
  NAND2_X1 U11838 ( .A1(n9281), .A2(n9280), .ZN(n13880) );
  INV_X1 U11839 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U11840 ( .A1(n9464), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9291) );
  NAND2_X1 U11841 ( .A1(n9306), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11842 ( .A1(n9305), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9288) );
  NOR2_X1 U11843 ( .A1(n9285), .A2(n9286), .ZN(n9307) );
  NAND2_X1 U11844 ( .A1(n9307), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9287) );
  AND2_X1 U11845 ( .A1(n9288), .A2(n9287), .ZN(n9289) );
  NAND3_X2 U11846 ( .A1(n9291), .A2(n9290), .A3(n9289), .ZN(n13212) );
  OR2_X1 U11847 ( .A1(n6565), .A2(n9048), .ZN(n9294) );
  INV_X1 U11848 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15364) );
  NAND2_X1 U11849 ( .A1(n9305), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U11850 ( .A1(n9307), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9297) );
  NAND4_X1 U11851 ( .A1(n9300), .A2(n9299), .A3(n9298), .A4(n9297), .ZN(n9847)
         );
  INV_X1 U11852 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n15211) );
  XNOR2_X1 U11853 ( .A(n9302), .B(n9301), .ZN(n13910) );
  OR2_X1 U11854 ( .A1(n9847), .A2(n12876), .ZN(n9848) );
  INV_X1 U11855 ( .A(n9848), .ZN(n9458) );
  XNOR2_X1 U11856 ( .A(n6954), .B(n9458), .ZN(n9315) );
  OR2_X1 U11857 ( .A1(n12867), .A2(n13244), .ZN(n9304) );
  INV_X1 U11858 ( .A(n6561), .ZN(n13157) );
  NAND2_X1 U11859 ( .A1(n10346), .A2(n13157), .ZN(n9303) );
  NAND2_X1 U11860 ( .A1(n9805), .A2(n9215), .ZN(n12808) );
  NAND2_X1 U11861 ( .A1(n9305), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11862 ( .A1(n9306), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U11863 ( .A1(n9307), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11864 ( .A1(n9464), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9308) );
  NAND4_X1 U11865 ( .A1(n9311), .A2(n9310), .A3(n9309), .A4(n9308), .ZN(n13211) );
  NAND2_X1 U11866 ( .A1(n12848), .A2(n13211), .ZN(n9314) );
  INV_X1 U11867 ( .A(n9215), .ZN(n9312) );
  AND2_X2 U11868 ( .A1(n9805), .A2(n9312), .ZN(n13167) );
  NAND2_X1 U11869 ( .A1(n13167), .A2(n9847), .ZN(n9313) );
  NAND2_X1 U11870 ( .A1(n9314), .A2(n9313), .ZN(n9914) );
  AOI21_X1 U11871 ( .B1(n9315), .B2(n15409), .A(n9914), .ZN(n13473) );
  INV_X1 U11872 ( .A(n12876), .ZN(n15312) );
  NAND2_X1 U11873 ( .A1(n15312), .A2(n13470), .ZN(n9316) );
  AND3_X1 U11874 ( .A1(n13431), .A2(n9471), .A3(n9316), .ZN(n13466) );
  INV_X1 U11875 ( .A(n9778), .ZN(n15313) );
  AND2_X1 U11876 ( .A1(n15421), .A2(n13470), .ZN(n9317) );
  NOR2_X1 U11877 ( .A1(n13466), .A2(n9317), .ZN(n9320) );
  XNOR2_X1 U11878 ( .A(n12867), .B(n12872), .ZN(n9318) );
  NAND2_X1 U11879 ( .A1(n9318), .A2(n13244), .ZN(n10347) );
  INV_X1 U11880 ( .A(n10347), .ZN(n15428) );
  INV_X1 U11881 ( .A(n15423), .ZN(n15363) );
  AND2_X1 U11882 ( .A1(n9847), .A2(n15312), .ZN(n9911) );
  XNOR2_X1 U11883 ( .A(n6954), .B(n9911), .ZN(n13468) );
  OAI21_X1 U11884 ( .B1(n15428), .B2(n15363), .A(n13468), .ZN(n9319) );
  AND3_X1 U11885 ( .A1(n13473), .A2(n9320), .A3(n9319), .ZN(n15366) );
  NAND2_X1 U11886 ( .A1(n15441), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9321) );
  OAI21_X1 U11887 ( .B1(n15441), .B2(n15366), .A(n9321), .ZN(P2_U3500) );
  INV_X1 U11888 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9323) );
  MUX2_X1 U11889 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9323), .S(n10129), .Z(n9324) );
  OAI21_X1 U11890 ( .B1(n9325), .B2(n9324), .A(n9376), .ZN(n9329) );
  INV_X1 U11891 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10142) );
  NOR2_X1 U11892 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10142), .ZN(n9326) );
  AOI21_X1 U11893 ( .B1(n15294), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n9326), .ZN(
        n9327) );
  OAI21_X1 U11894 ( .B1(n9383), .B2(n15273), .A(n9327), .ZN(n9328) );
  AOI21_X1 U11895 ( .B1(n9329), .B2(n15296), .A(n9328), .ZN(n9335) );
  AOI21_X1 U11896 ( .B1(n9998), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9330), .ZN(
        n9332) );
  INV_X1 U11897 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n15439) );
  MUX2_X1 U11898 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n15439), .S(n10129), .Z(
        n9331) );
  AND2_X1 U11899 ( .A1(n9332), .A2(n9331), .ZN(n9382) );
  NOR2_X1 U11900 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  OAI21_X1 U11901 ( .B1(n9382), .B2(n9333), .A(n15302), .ZN(n9334) );
  NAND2_X1 U11902 ( .A1(n9335), .A2(n9334), .ZN(P2_U3223) );
  NOR2_X1 U11903 ( .A1(n9336), .A2(n12615), .ZN(n9339) );
  CLKBUF_X1 U11904 ( .A(n9339), .Z(n9363) );
  INV_X1 U11905 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9337) );
  NOR2_X1 U11906 ( .A1(n9363), .A2(n9337), .ZN(P3_U3257) );
  INV_X1 U11907 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9338) );
  NOR2_X1 U11908 ( .A1(n9363), .A2(n9338), .ZN(P3_U3261) );
  INV_X1 U11909 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9340) );
  NOR2_X1 U11910 ( .A1(n9363), .A2(n9340), .ZN(P3_U3239) );
  INV_X1 U11911 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9341) );
  NOR2_X1 U11912 ( .A1(n9339), .A2(n9341), .ZN(P3_U3244) );
  INV_X1 U11913 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n13642) );
  NOR2_X1 U11914 ( .A1(n9339), .A2(n13642), .ZN(P3_U3258) );
  INV_X1 U11915 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9342) );
  NOR2_X1 U11916 ( .A1(n9339), .A2(n9342), .ZN(P3_U3245) );
  INV_X1 U11917 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9343) );
  NOR2_X1 U11918 ( .A1(n9339), .A2(n9343), .ZN(P3_U3237) );
  INV_X1 U11919 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9344) );
  NOR2_X1 U11920 ( .A1(n9339), .A2(n9344), .ZN(P3_U3238) );
  INV_X1 U11921 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9345) );
  NOR2_X1 U11922 ( .A1(n9339), .A2(n9345), .ZN(P3_U3241) );
  INV_X1 U11923 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n13617) );
  NOR2_X1 U11924 ( .A1(n9339), .A2(n13617), .ZN(P3_U3260) );
  INV_X1 U11925 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9346) );
  NOR2_X1 U11926 ( .A1(n9363), .A2(n9346), .ZN(P3_U3259) );
  INV_X1 U11927 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n13645) );
  NOR2_X1 U11928 ( .A1(n9363), .A2(n13645), .ZN(P3_U3249) );
  INV_X1 U11929 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9347) );
  NOR2_X1 U11930 ( .A1(n9363), .A2(n9347), .ZN(P3_U3254) );
  INV_X1 U11931 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9348) );
  NOR2_X1 U11932 ( .A1(n9363), .A2(n9348), .ZN(P3_U3256) );
  INV_X1 U11933 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n13763) );
  NOR2_X1 U11934 ( .A1(n9363), .A2(n13763), .ZN(P3_U3255) );
  INV_X1 U11935 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9349) );
  NOR2_X1 U11936 ( .A1(n9363), .A2(n9349), .ZN(P3_U3263) );
  INV_X1 U11937 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9350) );
  NOR2_X1 U11938 ( .A1(n9339), .A2(n9350), .ZN(P3_U3262) );
  INV_X1 U11939 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9351) );
  NOR2_X1 U11940 ( .A1(n9339), .A2(n9351), .ZN(P3_U3234) );
  INV_X1 U11941 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9352) );
  NOR2_X1 U11942 ( .A1(n9339), .A2(n9352), .ZN(P3_U3235) );
  INV_X1 U11943 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9353) );
  NOR2_X1 U11944 ( .A1(n9339), .A2(n9353), .ZN(P3_U3236) );
  INV_X1 U11945 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9354) );
  NOR2_X1 U11946 ( .A1(n9363), .A2(n9354), .ZN(P3_U3253) );
  INV_X1 U11947 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9355) );
  NOR2_X1 U11948 ( .A1(n9363), .A2(n9355), .ZN(P3_U3252) );
  INV_X1 U11949 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9356) );
  NOR2_X1 U11950 ( .A1(n9363), .A2(n9356), .ZN(P3_U3246) );
  INV_X1 U11951 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9357) );
  NOR2_X1 U11952 ( .A1(n9363), .A2(n9357), .ZN(P3_U3240) );
  INV_X1 U11953 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9358) );
  NOR2_X1 U11954 ( .A1(n9363), .A2(n9358), .ZN(P3_U3248) );
  INV_X1 U11955 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9359) );
  NOR2_X1 U11956 ( .A1(n9363), .A2(n9359), .ZN(P3_U3242) );
  INV_X1 U11957 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9360) );
  NOR2_X1 U11958 ( .A1(n9363), .A2(n9360), .ZN(P3_U3243) );
  INV_X1 U11959 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9361) );
  NOR2_X1 U11960 ( .A1(n9363), .A2(n9361), .ZN(P3_U3251) );
  INV_X1 U11961 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n13644) );
  NOR2_X1 U11962 ( .A1(n9363), .A2(n13644), .ZN(P3_U3247) );
  INV_X1 U11963 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9362) );
  NOR2_X1 U11964 ( .A1(n9363), .A2(n9362), .ZN(P3_U3250) );
  INV_X1 U11965 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9371) );
  INV_X1 U11966 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11967 ( .A1(n15296), .A2(n9364), .ZN(n9365) );
  OAI211_X1 U11968 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n13239), .A(n15273), .B(
        n9365), .ZN(n9366) );
  INV_X1 U11969 ( .A(n9366), .ZN(n9368) );
  AOI22_X1 U11970 ( .A1(n15302), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15296), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9367) );
  MUX2_X1 U11971 ( .A(n9368), .B(n9367), .S(n15211), .Z(n9370) );
  NAND2_X1 U11972 ( .A1(P2_U3088), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9369) );
  OAI211_X1 U11973 ( .C1(n13249), .C2(n9371), .A(n9370), .B(n9369), .ZN(
        P2_U3214) );
  INV_X1 U11974 ( .A(n9372), .ZN(n9373) );
  OAI21_X1 U11975 ( .B1(n9374), .B2(n9373), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9375) );
  XNOR2_X1 U11976 ( .A(n9375), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10377) );
  NAND2_X1 U11977 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10707)
         );
  OAI21_X1 U11978 ( .B1(n13249), .B2(n7450), .A(n10707), .ZN(n9381) );
  OAI21_X1 U11979 ( .B1(n10129), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9376), .ZN(
        n9379) );
  INV_X1 U11980 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9377) );
  MUX2_X1 U11981 ( .A(n9377), .B(P2_REG2_REG_10__SCAN_IN), .S(n10377), .Z(
        n9378) );
  AOI211_X1 U11982 ( .C1(n9379), .C2(n9378), .A(n15242), .B(n9487), .ZN(n9380)
         );
  AOI211_X1 U11983 ( .C1(n15299), .C2(n10377), .A(n9381), .B(n9380), .ZN(n9388) );
  AOI21_X1 U11984 ( .B1(n15439), .B2(n9383), .A(n9382), .ZN(n9386) );
  INV_X1 U11985 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9384) );
  MUX2_X1 U11986 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9384), .S(n10377), .Z(
        n9385) );
  NAND2_X1 U11987 ( .A1(n9386), .A2(n9385), .ZN(n9481) );
  OAI211_X1 U11988 ( .C1(n9386), .C2(n9385), .A(n9481), .B(n15302), .ZN(n9387)
         );
  NAND2_X1 U11989 ( .A1(n9388), .A2(n9387), .ZN(P2_U3224) );
  INV_X1 U11990 ( .A(n9389), .ZN(n9762) );
  NAND3_X1 U11991 ( .A1(n9390), .A2(n9762), .A3(n9760), .ZN(n9400) );
  OR2_X1 U11992 ( .A1(n9400), .A2(n9395), .ZN(n9397) );
  INV_X1 U11993 ( .A(n9397), .ZN(n9393) );
  NOR2_X1 U11994 ( .A1(n15159), .A2(n9391), .ZN(n9392) );
  NAND2_X1 U11995 ( .A1(n9400), .A2(n9396), .ZN(n10047) );
  NAND2_X1 U11996 ( .A1(n10047), .A2(n14309), .ZN(n13964) );
  AOI22_X1 U11997 ( .A1(n9394), .A2(n14052), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n13964), .ZN(n9402) );
  INV_X1 U11998 ( .A(n14309), .ZN(n9399) );
  NOR2_X2 U11999 ( .A1(n14055), .A2(n14608), .ZN(n14023) );
  AOI22_X1 U12000 ( .A1(n15141), .A2(n9398), .B1(n14023), .B2(n14624), .ZN(
        n9401) );
  NAND2_X1 U12001 ( .A1(n9402), .A2(n9401), .ZN(P1_U3232) );
  MUX2_X1 U12002 ( .A(n10763), .B(P1_REG2_REG_12__SCAN_IN), .S(n9413), .Z(
        n9406) );
  INV_X1 U12003 ( .A(n14406), .ZN(n9497) );
  NOR2_X1 U12004 ( .A1(n9447), .A2(n9403), .ZN(n14408) );
  MUX2_X1 U12005 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n9404), .S(n14406), .Z(
        n14407) );
  OAI21_X1 U12006 ( .B1(n14409), .B2(n14408), .A(n14407), .ZN(n14411) );
  OAI21_X1 U12007 ( .B1(n9404), .B2(n9497), .A(n14411), .ZN(n9405) );
  NOR2_X1 U12008 ( .A1(n9405), .A2(n9406), .ZN(n9560) );
  AOI21_X1 U12009 ( .B1(n9406), .B2(n9405), .A(n9560), .ZN(n9418) );
  AOI21_X1 U12010 ( .B1(n9408), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9407), .ZN(
        n14401) );
  MUX2_X1 U12011 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n8033), .S(n14406), .Z(
        n14402) );
  NAND2_X1 U12012 ( .A1(n14401), .A2(n14402), .ZN(n14400) );
  NAND2_X1 U12013 ( .A1(n9497), .A2(n8033), .ZN(n9410) );
  MUX2_X1 U12014 ( .A(n9409), .B(P1_REG1_REG_12__SCAN_IN), .S(n9413), .Z(n9411) );
  AOI21_X1 U12015 ( .B1(n14400), .B2(n9410), .A(n9411), .ZN(n9556) );
  AND3_X1 U12016 ( .A1(n14400), .A2(n9411), .A3(n9410), .ZN(n9412) );
  OAI21_X1 U12017 ( .B1(n9556), .B2(n9412), .A(n15035), .ZN(n9417) );
  NOR2_X1 U12018 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8048), .ZN(n9415) );
  INV_X1 U12019 ( .A(n9413), .ZN(n9561) );
  NOR2_X1 U12020 ( .A1(n15029), .A2(n9561), .ZN(n9414) );
  AOI211_X1 U12021 ( .C1(n15006), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9415), .B(
        n9414), .ZN(n9416) );
  OAI211_X1 U12022 ( .C1(n9418), .C2(n15025), .A(n9417), .B(n9416), .ZN(
        P1_U3255) );
  NAND2_X1 U12023 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n12841) );
  OAI211_X1 U12024 ( .C1(n9420), .C2(n9419), .A(n15302), .B(n13223), .ZN(n9421) );
  NAND2_X1 U12025 ( .A1(n12841), .A2(n9421), .ZN(n9426) );
  AND3_X1 U12026 ( .A1(n9433), .A2(n9423), .A3(n9422), .ZN(n9424) );
  NOR3_X1 U12027 ( .A1(n15242), .A2(n13216), .A3(n9424), .ZN(n9425) );
  AOI211_X1 U12028 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n15294), .A(n9426), .B(
        n9425), .ZN(n9427) );
  OAI21_X1 U12029 ( .B1(n9428), .B2(n15273), .A(n9427), .ZN(P2_U3220) );
  NAND2_X1 U12030 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10073) );
  OAI211_X1 U12031 ( .C1(n9431), .C2(n9430), .A(n15302), .B(n9429), .ZN(n9432)
         );
  NAND2_X1 U12032 ( .A1(n10073), .A2(n9432), .ZN(n9439) );
  INV_X1 U12033 ( .A(n9433), .ZN(n9437) );
  NOR3_X1 U12034 ( .A1(n15243), .A2(n9435), .A3(n9434), .ZN(n9436) );
  NOR3_X1 U12035 ( .A1(n15242), .A2(n9437), .A3(n9436), .ZN(n9438) );
  AOI211_X1 U12036 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n15294), .A(n9439), .B(
        n9438), .ZN(n9440) );
  OAI21_X1 U12037 ( .B1(n9441), .B2(n15273), .A(n9440), .ZN(P2_U3219) );
  INV_X1 U12038 ( .A(n10566), .ZN(n9445) );
  NAND2_X1 U12039 ( .A1(n9442), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9443) );
  XNOR2_X1 U12040 ( .A(n9443), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10567) );
  INV_X1 U12041 ( .A(n10567), .ZN(n11046) );
  OAI222_X1 U12042 ( .A1(n13905), .A2(n9444), .B1(n13908), .B2(n9445), .C1(
        P2_U3088), .C2(n11046), .ZN(P2_U3315) );
  OAI222_X1 U12043 ( .A1(n11330), .A2(n9446), .B1(n14753), .B2(n9445), .C1(
        P1_U3086), .C2(n9561), .ZN(P1_U3343) );
  INV_X1 U12044 ( .A(n10376), .ZN(n9449) );
  OAI222_X1 U12045 ( .A1(n11330), .A2(n9448), .B1(n14753), .B2(n9449), .C1(
        P1_U3086), .C2(n9447), .ZN(P1_U3345) );
  INV_X1 U12046 ( .A(n10377), .ZN(n9482) );
  OAI222_X1 U12047 ( .A1(n13905), .A2(n9450), .B1(n13908), .B2(n9449), .C1(
        P2_U3088), .C2(n9482), .ZN(P2_U3317) );
  OAI222_X1 U12048 ( .A1(P3_U3151), .A2(n12222), .B1(n12623), .B2(n13727), 
        .C1(n12627), .C2(n9451), .ZN(P3_U3280) );
  OR2_X1 U12049 ( .A1(n13082), .A2(n9452), .ZN(n9455) );
  OR2_X1 U12050 ( .A1(n13083), .A2(n9453), .ZN(n9454) );
  NAND2_X1 U12051 ( .A1(n13211), .A2(n9473), .ZN(n9457) );
  INV_X1 U12052 ( .A(n9944), .ZN(n13121) );
  NAND2_X1 U12053 ( .A1(n6954), .A2(n9458), .ZN(n9461) );
  OR2_X1 U12054 ( .A1(n13212), .A2(n9459), .ZN(n9460) );
  NAND2_X1 U12055 ( .A1(n9461), .A2(n9460), .ZN(n9462) );
  NAND2_X1 U12056 ( .A1(n9462), .A2(n13121), .ZN(n10476) );
  OAI21_X1 U12057 ( .B1(n13121), .B2(n9462), .A(n10476), .ZN(n9463) );
  NAND2_X1 U12058 ( .A1(n9463), .A2(n15409), .ZN(n9470) );
  NAND2_X1 U12059 ( .A1(n13072), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9467) );
  INV_X1 U12060 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U12061 ( .A1(n11502), .A2(n9465), .ZN(n9466) );
  NAND2_X1 U12062 ( .A1(n12848), .A2(n13210), .ZN(n9469) );
  NAND2_X1 U12063 ( .A1(n13167), .A2(n13212), .ZN(n9468) );
  AND2_X1 U12064 ( .A1(n9469), .A2(n9468), .ZN(n10202) );
  NAND2_X1 U12065 ( .A1(n9470), .A2(n10202), .ZN(n10504) );
  NAND2_X1 U12066 ( .A1(n9471), .A2(n12888), .ZN(n9472) );
  NAND3_X1 U12067 ( .A1(n10471), .A2(n13431), .A3(n9472), .ZN(n10507) );
  OAI21_X1 U12068 ( .B1(n15379), .B2(n9473), .A(n10507), .ZN(n9474) );
  NOR2_X1 U12069 ( .A1(n10504), .A2(n9474), .ZN(n9479) );
  OR2_X1 U12070 ( .A1(n13212), .A2(n13470), .ZN(n9475) );
  NAND2_X1 U12071 ( .A1(n9476), .A2(n9475), .ZN(n9945) );
  XNOR2_X1 U12072 ( .A(n9945), .B(n13121), .ZN(n10501) );
  INV_X1 U12073 ( .A(n10501), .ZN(n9477) );
  NAND2_X1 U12074 ( .A1(n9477), .A2(n13571), .ZN(n9478) );
  AND2_X1 U12075 ( .A1(n9479), .A2(n9478), .ZN(n15368) );
  NAND2_X1 U12076 ( .A1(n15441), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9480) );
  OAI21_X1 U12077 ( .B1(n15368), .B2(n15441), .A(n9480), .ZN(P2_U3501) );
  OAI21_X1 U12078 ( .B1(n9384), .B2(n9482), .A(n9481), .ZN(n9517) );
  NAND2_X1 U12079 ( .A1(n9483), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9484) );
  XNOR2_X1 U12080 ( .A(n9484), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10580) );
  INV_X1 U12081 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9485) );
  XNOR2_X1 U12082 ( .A(n10580), .B(n9485), .ZN(n9516) );
  XNOR2_X1 U12083 ( .A(n9517), .B(n9516), .ZN(n9496) );
  INV_X1 U12084 ( .A(n10580), .ZN(n9499) );
  INV_X1 U12085 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9486) );
  OR2_X1 U12086 ( .A1(n9499), .A2(n9486), .ZN(n9488) );
  NAND2_X1 U12087 ( .A1(n9499), .A2(n9486), .ZN(n9522) );
  AOI21_X1 U12088 ( .B1(n9488), .B2(n9522), .A(n9489), .ZN(n9491) );
  INV_X1 U12089 ( .A(n9524), .ZN(n9490) );
  OAI21_X1 U12090 ( .B1(n9491), .B2(n9490), .A(n15296), .ZN(n9495) );
  INV_X1 U12091 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9492) );
  NAND2_X1 U12092 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10668)
         );
  OAI21_X1 U12093 ( .B1(n13249), .B2(n9492), .A(n10668), .ZN(n9493) );
  AOI21_X1 U12094 ( .B1(n10580), .B2(n15299), .A(n9493), .ZN(n9494) );
  OAI211_X1 U12095 ( .C1(n9496), .C2(n13239), .A(n9495), .B(n9494), .ZN(
        P2_U3225) );
  INV_X1 U12096 ( .A(n10579), .ZN(n9500) );
  OAI222_X1 U12097 ( .A1(n11330), .A2(n9498), .B1(n14753), .B2(n9500), .C1(
        P1_U3086), .C2(n9497), .ZN(P1_U3344) );
  OAI222_X1 U12098 ( .A1(n13905), .A2(n7317), .B1(n13908), .B2(n9500), .C1(
        P2_U3088), .C2(n9499), .ZN(P2_U3316) );
  INV_X1 U12099 ( .A(n10818), .ZN(n9504) );
  OAI222_X1 U12100 ( .A1(n14755), .A2(n9501), .B1(n14753), .B2(n9504), .C1(
        n15009), .C2(P1_U3086), .ZN(P1_U3342) );
  OR2_X1 U12101 ( .A1(n9502), .A2(n13881), .ZN(n9503) );
  XNOR2_X1 U12102 ( .A(n9503), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15257) );
  INV_X1 U12103 ( .A(n15257), .ZN(n11050) );
  OAI222_X1 U12104 ( .A1(n13905), .A2(n9505), .B1(n13908), .B2(n9504), .C1(
        n11050), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12105 ( .A(n12220), .ZN(n12249) );
  INV_X1 U12106 ( .A(n9506), .ZN(n9507) );
  OAI222_X1 U12107 ( .A1(P3_U3151), .A2(n12249), .B1(n12623), .B2(n13778), 
        .C1(n12627), .C2(n9507), .ZN(P3_U3279) );
  INV_X1 U12108 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n9510) );
  NAND2_X1 U12109 ( .A1(n9508), .A2(P3_U3897), .ZN(n9509) );
  OAI21_X1 U12110 ( .B1(P3_U3897), .B2(n9510), .A(n9509), .ZN(P3_U3494) );
  OAI222_X1 U12111 ( .A1(P3_U3151), .A2(n12252), .B1(n12623), .B2(n9512), .C1(
        n12627), .C2(n9511), .ZN(P3_U3278) );
  NAND2_X1 U12112 ( .A1(n12181), .A2(P3_DATAO_REG_19__SCAN_IN), .ZN(n9513) );
  OAI21_X1 U12113 ( .B1(n12407), .B2(n12181), .A(n9513), .ZN(P3_U3510) );
  INV_X1 U12114 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n13608) );
  INV_X1 U12115 ( .A(n9514), .ZN(n11547) );
  NAND2_X1 U12116 ( .A1(n9514), .A2(P3_U3897), .ZN(n9515) );
  OAI21_X1 U12117 ( .B1(P3_U3897), .B2(n13608), .A(n9515), .ZN(P3_U3492) );
  INV_X1 U12118 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11045) );
  XNOR2_X1 U12119 ( .A(n10567), .B(n11045), .ZN(n11047) );
  AOI22_X1 U12120 ( .A1(n9517), .A2(n9516), .B1(P2_REG1_REG_11__SCAN_IN), .B2(
        n10580), .ZN(n11048) );
  XOR2_X1 U12121 ( .A(n11047), .B(n11048), .Z(n9530) );
  INV_X1 U12122 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U12123 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n9518) );
  OAI21_X1 U12124 ( .B1(n13249), .B2(n9519), .A(n9518), .ZN(n9528) );
  INV_X1 U12125 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11037) );
  NAND2_X1 U12126 ( .A1(n10567), .A2(n11037), .ZN(n9520) );
  OAI21_X1 U12127 ( .B1(n10567), .B2(n11037), .A(n9520), .ZN(n9521) );
  INV_X1 U12128 ( .A(n9521), .ZN(n9523) );
  INV_X1 U12129 ( .A(n11036), .ZN(n9526) );
  NAND3_X1 U12130 ( .A1(n9524), .A2(n9523), .A3(n9522), .ZN(n9525) );
  AOI21_X1 U12131 ( .B1(n9526), .B2(n9525), .A(n15242), .ZN(n9527) );
  AOI211_X1 U12132 ( .C1(n15299), .C2(n10567), .A(n9528), .B(n9527), .ZN(n9529) );
  OAI21_X1 U12133 ( .B1(n9530), .B2(n13239), .A(n9529), .ZN(P2_U3226) );
  AND2_X1 U12134 ( .A1(P3_U3897), .A2(n11081), .ZN(n12280) );
  INV_X1 U12135 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11557) );
  INV_X1 U12136 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9532) );
  MUX2_X1 U12137 ( .A(n11557), .B(n9532), .S(n12275), .Z(n9533) );
  AND2_X1 U12138 ( .A1(n9533), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9646) );
  MUX2_X1 U12139 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12275), .Z(n9573) );
  INV_X1 U12140 ( .A(n9546), .ZN(n9574) );
  XNOR2_X1 U12141 ( .A(n9573), .B(n9574), .ZN(n9572) );
  XOR2_X1 U12142 ( .A(n9646), .B(n9572), .Z(n9555) );
  NAND2_X1 U12143 ( .A1(n12103), .A2(n9536), .ZN(n9534) );
  AND2_X1 U12144 ( .A1(n9535), .A2(n9534), .ZN(n9543) );
  INV_X1 U12145 ( .A(n9536), .ZN(n9537) );
  NAND2_X1 U12146 ( .A1(n9537), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12165) );
  INV_X1 U12147 ( .A(n12165), .ZN(n10211) );
  OR2_X1 U12148 ( .A1(n12159), .A2(n10211), .ZN(n9544) );
  MUX2_X1 U12149 ( .A(n9548), .B(P3_U3897), .S(n12160), .Z(n14907) );
  INV_X1 U12150 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9540) );
  NOR2_X1 U12151 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11557), .ZN(n9637) );
  NAND2_X1 U12152 ( .A1(n8461), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9538) );
  OAI21_X1 U12153 ( .B1(n9546), .B2(n9637), .A(n9538), .ZN(n9539) );
  NOR2_X1 U12154 ( .A1(n9539), .A2(n9540), .ZN(n9578) );
  AOI21_X1 U12155 ( .B1(n9540), .B2(n9539), .A(n9578), .ZN(n9552) );
  INV_X1 U12156 ( .A(n9541), .ZN(n9542) );
  INV_X1 U12157 ( .A(n9543), .ZN(n9545) );
  AOI22_X1 U12158 ( .A1(n15458), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9551) );
  NAND2_X1 U12159 ( .A1(n9648), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9582) );
  NOR2_X1 U12160 ( .A1(n9547), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9549) );
  OAI21_X1 U12161 ( .B1(n9583), .B2(n9549), .A(n15461), .ZN(n9550) );
  OAI211_X1 U12162 ( .C1(n9552), .C2(n15465), .A(n9551), .B(n9550), .ZN(n9553)
         );
  AOI21_X1 U12163 ( .B1(n9574), .B2(n14907), .A(n9553), .ZN(n9554) );
  OAI21_X1 U12164 ( .B1(n15454), .B2(n9555), .A(n9554), .ZN(P3_U3183) );
  INV_X1 U12165 ( .A(n9563), .ZN(n10325) );
  AOI22_X1 U12166 ( .A1(n9563), .A2(n8082), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n10325), .ZN(n9559) );
  AOI21_X1 U12167 ( .B1(n9409), .B2(n9561), .A(n9556), .ZN(n15013) );
  MUX2_X1 U12168 ( .A(n9557), .B(P1_REG1_REG_13__SCAN_IN), .S(n15009), .Z(
        n15012) );
  NAND2_X1 U12169 ( .A1(n15013), .A2(n15012), .ZN(n15011) );
  OAI21_X1 U12170 ( .B1(n15009), .B2(n9557), .A(n15011), .ZN(n9558) );
  NOR2_X1 U12171 ( .A1(n9559), .A2(n9558), .ZN(n10324) );
  AOI21_X1 U12172 ( .B1(n9559), .B2(n9558), .A(n10324), .ZN(n9571) );
  AOI21_X1 U12173 ( .B1(n10763), .B2(n9561), .A(n9560), .ZN(n15016) );
  MUX2_X1 U12174 ( .A(n9562), .B(P1_REG2_REG_13__SCAN_IN), .S(n15009), .Z(
        n15015) );
  NAND2_X1 U12175 ( .A1(n15016), .A2(n15015), .ZN(n15014) );
  OAI21_X1 U12176 ( .B1(n9562), .B2(n15009), .A(n15014), .ZN(n9566) );
  MUX2_X1 U12177 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n9564), .S(n9563), .Z(n9565) );
  NAND2_X1 U12178 ( .A1(n9565), .A2(n9566), .ZN(n10318) );
  OAI211_X1 U12179 ( .C1(n9566), .C2(n9565), .A(n15040), .B(n10318), .ZN(n9568) );
  AND2_X1 U12180 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13923) );
  AOI21_X1 U12181 ( .B1(n15006), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n13923), 
        .ZN(n9567) );
  OAI211_X1 U12182 ( .C1(n15029), .C2(n10325), .A(n9568), .B(n9567), .ZN(n9569) );
  INV_X1 U12183 ( .A(n9569), .ZN(n9570) );
  OAI21_X1 U12184 ( .B1(n9571), .B2(n15027), .A(n9570), .ZN(P1_U3257) );
  MUX2_X1 U12185 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12275), .Z(n9663) );
  XNOR2_X1 U12186 ( .A(n9663), .B(n9664), .ZN(n9661) );
  NAND2_X1 U12187 ( .A1(n9572), .A2(n9646), .ZN(n9577) );
  INV_X1 U12188 ( .A(n9573), .ZN(n9575) );
  NAND2_X1 U12189 ( .A1(n9575), .A2(n9574), .ZN(n9576) );
  NAND2_X1 U12190 ( .A1(n9577), .A2(n9576), .ZN(n9662) );
  XOR2_X1 U12191 ( .A(n9661), .B(n9662), .Z(n9592) );
  INV_X1 U12192 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11553) );
  XNOR2_X1 U12193 ( .A(n9664), .B(n11553), .ZN(n9580) );
  AOI21_X1 U12194 ( .B1(n8461), .B2(P3_REG2_REG_0__SCAN_IN), .A(n9578), .ZN(
        n9579) );
  AOI21_X1 U12195 ( .B1(n9580), .B2(n9579), .A(n9669), .ZN(n9581) );
  NOR2_X1 U12196 ( .A1(n15465), .A2(n9581), .ZN(n9590) );
  INV_X1 U12197 ( .A(n15461), .ZN(n12258) );
  INV_X1 U12198 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15522) );
  AOI21_X1 U12199 ( .B1(n9586), .B2(n9585), .A(n9668), .ZN(n9588) );
  AOI22_X1 U12200 ( .A1(n15458), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n9587) );
  OAI21_X1 U12201 ( .B1(n12258), .B2(n9588), .A(n9587), .ZN(n9589) );
  AOI211_X1 U12202 ( .C1(n14907), .C2(n9664), .A(n9590), .B(n9589), .ZN(n9591)
         );
  OAI21_X1 U12203 ( .B1(n9592), .B2(n15454), .A(n9591), .ZN(P3_U3184) );
  INV_X1 U12204 ( .A(n11354), .ZN(n9599) );
  OAI222_X1 U12205 ( .A1(n14755), .A2(n13776), .B1(n14753), .B2(n9599), .C1(
        n10488), .C2(P1_U3086), .ZN(P1_U3339) );
  NAND2_X1 U12206 ( .A1(n9502), .A2(n9593), .ZN(n9613) );
  OR2_X1 U12207 ( .A1(n9613), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n9649) );
  NOR2_X1 U12208 ( .A1(n9649), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n9597) );
  INV_X1 U12209 ( .A(n9597), .ZN(n9594) );
  NAND2_X1 U12210 ( .A1(n9594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9595) );
  MUX2_X1 U12211 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9595), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9598) );
  INV_X1 U12212 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U12213 ( .A1(n9597), .A2(n9596), .ZN(n9657) );
  AND2_X1 U12214 ( .A1(n9598), .A2(n9657), .ZN(n15283) );
  INV_X1 U12215 ( .A(n15283), .ZN(n11058) );
  OAI222_X1 U12216 ( .A1(n13905), .A2(n9600), .B1(n13908), .B2(n9599), .C1(
        n11058), .C2(P2_U3088), .ZN(P2_U3311) );
  XNOR2_X1 U12217 ( .A(n9601), .B(n11795), .ZN(n9603) );
  NOR2_X1 U12218 ( .A1(n9603), .A2(n9602), .ZN(n9606) );
  AOI21_X1 U12219 ( .B1(n9603), .B2(n9602), .A(n9606), .ZN(n13961) );
  OAI21_X1 U12220 ( .B1(n11765), .B2(n9605), .A(n9604), .ZN(n13960) );
  AND2_X1 U12221 ( .A1(n13961), .A2(n13960), .ZN(n13962) );
  AOI22_X1 U12222 ( .A1(n11787), .A2(n14336), .B1(n10307), .B2(n14111), .ZN(
        n10036) );
  OAI22_X1 U12223 ( .A1(n14110), .A2(n11798), .B1(n9725), .B2(n11794), .ZN(
        n9607) );
  XNOR2_X1 U12224 ( .A(n9607), .B(n11795), .ZN(n10035) );
  XOR2_X1 U12225 ( .A(n10036), .B(n10035), .Z(n9608) );
  AOI21_X1 U12226 ( .B1(n9609), .B2(n9608), .A(n10038), .ZN(n9612) );
  AOI22_X1 U12227 ( .A1(n14023), .A2(n14335), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n13964), .ZN(n9611) );
  NOR2_X2 U12228 ( .A1(n14055), .A2(n14606), .ZN(n14064) );
  AOI22_X1 U12229 ( .A1(n14111), .A2(n9398), .B1(n14064), .B2(n14624), .ZN(
        n9610) );
  OAI211_X1 U12230 ( .C1(n9612), .C2(n14074), .A(n9611), .B(n9610), .ZN(
        P1_U3237) );
  INV_X1 U12231 ( .A(n10899), .ZN(n9616) );
  NAND2_X1 U12232 ( .A1(n9613), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9614) );
  XNOR2_X1 U12233 ( .A(n9614), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11053) );
  INV_X1 U12234 ( .A(n11053), .ZN(n15272) );
  OAI222_X1 U12235 ( .A1(n13905), .A2(n9615), .B1(n13908), .B2(n9616), .C1(
        n15272), .C2(P2_U3088), .ZN(P2_U3313) );
  OAI222_X1 U12236 ( .A1(n14755), .A2(n9617), .B1(n14753), .B2(n9616), .C1(
        n10325), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U12237 ( .A(n12267), .ZN(n12273) );
  OAI222_X1 U12238 ( .A1(P3_U3151), .A2(n12273), .B1(n12623), .B2(n13597), 
        .C1(n12627), .C2(n9618), .ZN(P3_U3277) );
  INV_X1 U12239 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12240 ( .A1(n14271), .A2(n9619), .ZN(n9620) );
  NAND2_X1 U12241 ( .A1(n9621), .A2(n9620), .ZN(n9925) );
  INV_X1 U12242 ( .A(n9925), .ZN(n9630) );
  AND2_X1 U12243 ( .A1(n13965), .A2(n15141), .ZN(n9622) );
  OR2_X1 U12244 ( .A1(n9622), .A2(n9722), .ZN(n9628) );
  MUX2_X1 U12245 ( .A(n9623), .B(n14271), .S(n14338), .Z(n9626) );
  AOI22_X1 U12246 ( .A1(n14338), .A2(n14554), .B1(n15059), .B2(n14336), .ZN(
        n9625) );
  INV_X1 U12247 ( .A(n15068), .ZN(n15167) );
  NAND2_X1 U12248 ( .A1(n9925), .A2(n15167), .ZN(n9624) );
  OAI211_X1 U12249 ( .C1(n9626), .C2(n15084), .A(n9625), .B(n9624), .ZN(n9627)
         );
  INV_X1 U12250 ( .A(n9627), .ZN(n9927) );
  INV_X1 U12251 ( .A(n9628), .ZN(n9920) );
  AOI22_X1 U12252 ( .A1(n9920), .A2(n8988), .B1(n13965), .B2(n15159), .ZN(
        n9629) );
  OAI211_X1 U12253 ( .C1(n9630), .C2(n15163), .A(n9927), .B(n9629), .ZN(n9634)
         );
  NAND2_X1 U12254 ( .A1(n9634), .A2(n15197), .ZN(n9631) );
  OAI21_X1 U12255 ( .B1(n15197), .B2(n9632), .A(n9631), .ZN(P1_U3462) );
  INV_X2 U12256 ( .A(n15206), .ZN(n15209) );
  NAND2_X1 U12257 ( .A1(n9634), .A2(n15209), .ZN(n9635) );
  OAI21_X1 U12258 ( .B1(n15209), .B2(n9013), .A(n9635), .ZN(P1_U3529) );
  INV_X1 U12259 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n13742) );
  NAND2_X1 U12260 ( .A1(n10748), .A2(P3_U3897), .ZN(n9636) );
  OAI21_X1 U12261 ( .B1(P3_U3897), .B2(n13742), .A(n9636), .ZN(P3_U3496) );
  INV_X1 U12262 ( .A(n14907), .ZN(n15452) );
  NAND3_X1 U12263 ( .A1(n12258), .A2(n15465), .A3(n15454), .ZN(n9645) );
  INV_X1 U12264 ( .A(n9637), .ZN(n9643) );
  INV_X1 U12265 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9757) );
  MUX2_X1 U12266 ( .A(n9637), .B(n6949), .S(n12275), .Z(n9638) );
  NAND2_X1 U12267 ( .A1(n12280), .A2(n9638), .ZN(n9639) );
  OAI21_X1 U12268 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n9757), .A(n9639), .ZN(
        n9640) );
  AOI21_X1 U12269 ( .B1(n15458), .B2(P3_ADDR_REG_0__SCAN_IN), .A(n9640), .ZN(
        n9642) );
  NAND2_X1 U12270 ( .A1(n15461), .A2(n6949), .ZN(n9641) );
  OAI211_X1 U12271 ( .C1(n9643), .C2(n15465), .A(n9642), .B(n9641), .ZN(n9644)
         );
  AOI21_X1 U12272 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9647) );
  OAI21_X1 U12273 ( .B1(n9648), .B2(n15452), .A(n9647), .ZN(P3_U3182) );
  INV_X1 U12274 ( .A(n11001), .ZN(n9652) );
  NAND2_X1 U12275 ( .A1(n9649), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9650) );
  XNOR2_X1 U12276 ( .A(n9650), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15274) );
  INV_X1 U12277 ( .A(n15274), .ZN(n11054) );
  OAI222_X1 U12278 ( .A1(n13905), .A2(n9651), .B1(n13908), .B2(n9652), .C1(
        P2_U3088), .C2(n11054), .ZN(P2_U3312) );
  INV_X1 U12279 ( .A(n10327), .ZN(n15028) );
  OAI222_X1 U12280 ( .A1(n14755), .A2(n9653), .B1(n14753), .B2(n9652), .C1(
        P1_U3086), .C2(n15028), .ZN(P1_U3340) );
  INV_X1 U12281 ( .A(n11358), .ZN(n9660) );
  INV_X1 U12282 ( .A(n10957), .ZN(n9654) );
  OAI222_X1 U12283 ( .A1(n14755), .A2(n9655), .B1(n14753), .B2(n9660), .C1(
        n9654), .C2(P1_U3086), .ZN(P1_U3338) );
  NAND2_X1 U12284 ( .A1(n9657), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9658) );
  MUX2_X1 U12285 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9658), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n9659) );
  AND2_X1 U12286 ( .A1(n9656), .A2(n9659), .ZN(n15300) );
  INV_X1 U12287 ( .A(n15300), .ZN(n11060) );
  OAI222_X1 U12288 ( .A1(n13905), .A2(n13792), .B1(n13908), .B2(n9660), .C1(
        n11060), .C2(P2_U3088), .ZN(P2_U3310) );
  MUX2_X1 U12289 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12275), .Z(n9696) );
  XNOR2_X1 U12290 ( .A(n9696), .B(n9697), .ZN(n9694) );
  NAND2_X1 U12291 ( .A1(n9662), .A2(n9661), .ZN(n9667) );
  INV_X1 U12292 ( .A(n9663), .ZN(n9665) );
  NAND2_X1 U12293 ( .A1(n9665), .A2(n9664), .ZN(n9666) );
  NAND2_X1 U12294 ( .A1(n9667), .A2(n9666), .ZN(n9695) );
  XOR2_X1 U12295 ( .A(n9694), .B(n9695), .Z(n9678) );
  XOR2_X1 U12296 ( .A(P3_REG1_REG_3__SCAN_IN), .B(n9703), .Z(n9675) );
  NOR2_X1 U12297 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8485), .ZN(n10220) );
  AOI21_X1 U12298 ( .B1(n15458), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10220), .ZN(
        n9674) );
  OAI21_X1 U12299 ( .B1(n9671), .B2(P3_REG2_REG_3__SCAN_IN), .A(n9706), .ZN(
        n9672) );
  NAND2_X1 U12300 ( .A1(n7334), .A2(n9672), .ZN(n9673) );
  OAI211_X1 U12301 ( .C1(n12258), .C2(n9675), .A(n9674), .B(n9673), .ZN(n9676)
         );
  AOI21_X1 U12302 ( .B1(n9697), .B2(n14907), .A(n9676), .ZN(n9677) );
  OAI21_X1 U12303 ( .B1(n9678), .B2(n15454), .A(n9677), .ZN(P3_U3185) );
  OAI222_X1 U12304 ( .A1(n12623), .A2(n9681), .B1(P3_U3151), .B2(n9680), .C1(
        n12627), .C2(n9679), .ZN(P3_U3276) );
  INV_X1 U12305 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9691) );
  XNOR2_X1 U12306 ( .A(n9682), .B(n9684), .ZN(n10108) );
  OAI21_X1 U12307 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n10106) );
  OAI211_X1 U12308 ( .C1(n9723), .C2(n14117), .A(n8988), .B(n9767), .ZN(n10104) );
  OR2_X1 U12309 ( .A1(n14122), .A2(n14608), .ZN(n9687) );
  NAND2_X1 U12310 ( .A1(n14336), .A2(n14554), .ZN(n9686) );
  AND2_X1 U12311 ( .A1(n9687), .A2(n9686), .ZN(n10101) );
  OAI211_X1 U12312 ( .C1(n14117), .C2(n15191), .A(n10104), .B(n10101), .ZN(
        n9688) );
  AOI21_X1 U12313 ( .B1(n10106), .B2(n15195), .A(n9688), .ZN(n9689) );
  OAI21_X1 U12314 ( .B1(n15084), .B2(n10108), .A(n9689), .ZN(n9692) );
  NAND2_X1 U12315 ( .A1(n9692), .A2(n15197), .ZN(n9690) );
  OAI21_X1 U12316 ( .B1(n15197), .B2(n9691), .A(n9690), .ZN(P1_U3468) );
  NAND2_X1 U12317 ( .A1(n9692), .A2(n15209), .ZN(n9693) );
  OAI21_X1 U12318 ( .B1(n15209), .B2(n9020), .A(n9693), .ZN(P1_U3531) );
  MUX2_X1 U12319 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12275), .Z(n9815) );
  XNOR2_X1 U12320 ( .A(n9815), .B(n9816), .ZN(n9813) );
  NAND2_X1 U12321 ( .A1(n9695), .A2(n9694), .ZN(n9700) );
  INV_X1 U12322 ( .A(n9696), .ZN(n9698) );
  NAND2_X1 U12323 ( .A1(n9698), .A2(n9697), .ZN(n9699) );
  NAND2_X1 U12324 ( .A1(n9700), .A2(n9699), .ZN(n9814) );
  XOR2_X1 U12325 ( .A(n9813), .B(n9814), .Z(n9715) );
  INV_X1 U12326 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15526) );
  MUX2_X1 U12327 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n15526), .S(n9816), .Z(n9705) );
  INV_X1 U12328 ( .A(n9701), .ZN(n9702) );
  AOI21_X1 U12329 ( .B1(n9705), .B2(n9704), .A(n9820), .ZN(n9712) );
  AND2_X1 U12330 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10515) );
  AOI21_X1 U12331 ( .B1(n15458), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10515), .ZN(
        n9711) );
  INV_X1 U12332 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10466) );
  NOR2_X1 U12333 ( .A1(n9816), .A2(n10466), .ZN(n9822) );
  AOI21_X1 U12334 ( .B1(n9816), .B2(n10466), .A(n9822), .ZN(n9708) );
  NAND2_X1 U12335 ( .A1(n9706), .A2(n6726), .ZN(n9707) );
  OAI21_X1 U12336 ( .B1(n9708), .B2(n9707), .A(n9824), .ZN(n9709) );
  NAND2_X1 U12337 ( .A1(n7334), .A2(n9709), .ZN(n9710) );
  OAI211_X1 U12338 ( .C1(n12258), .C2(n9712), .A(n9711), .B(n9710), .ZN(n9713)
         );
  AOI21_X1 U12339 ( .B1(n9816), .B2(n14907), .A(n9713), .ZN(n9714) );
  OAI21_X1 U12340 ( .B1(n9715), .B2(n15454), .A(n9714), .ZN(P3_U3186) );
  OAI222_X1 U12341 ( .A1(n12627), .A2(n9718), .B1(n12623), .B2(n9717), .C1(
        P3_U3151), .C2(n9716), .ZN(P3_U3275) );
  INV_X1 U12342 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9732) );
  INV_X1 U12343 ( .A(n15163), .ZN(n15186) );
  OAI21_X1 U12344 ( .B1(n9721), .B2(n9720), .A(n9719), .ZN(n10162) );
  OAI21_X1 U12345 ( .B1(n9722), .B2(n9725), .A(n8988), .ZN(n9724) );
  OR2_X1 U12346 ( .A1(n9724), .A2(n9723), .ZN(n10158) );
  OAI21_X1 U12347 ( .B1(n9725), .B2(n15191), .A(n10158), .ZN(n9730) );
  XNOR2_X1 U12348 ( .A(n9726), .B(n14268), .ZN(n9729) );
  NAND2_X1 U12349 ( .A1(n10162), .A2(n15167), .ZN(n9728) );
  AOI22_X1 U12350 ( .A1(n14624), .A2(n14554), .B1(n15059), .B2(n14335), .ZN(
        n9727) );
  OAI211_X1 U12351 ( .C1(n15084), .C2(n9729), .A(n9728), .B(n9727), .ZN(n10159) );
  AOI211_X1 U12352 ( .C1(n15186), .C2(n10162), .A(n9730), .B(n10159), .ZN(
        n9733) );
  OR2_X1 U12353 ( .A1(n9733), .A2(n15196), .ZN(n9731) );
  OAI21_X1 U12354 ( .B1(n15197), .B2(n9732), .A(n9731), .ZN(P1_U3465) );
  OR2_X1 U12355 ( .A1(n9733), .A2(n15206), .ZN(n9734) );
  OAI21_X1 U12356 ( .B1(n15209), .B2(n9017), .A(n9734), .ZN(P1_U3530) );
  OAI211_X1 U12357 ( .C1(n9750), .C2(n9744), .A(n9735), .B(n10231), .ZN(n9739)
         );
  INV_X1 U12358 ( .A(n9736), .ZN(n9737) );
  NOR2_X1 U12359 ( .A1(n9752), .A2(n9737), .ZN(n9738) );
  OAI21_X1 U12360 ( .B1(n9739), .B2(n9738), .A(P3_STATE_REG_SCAN_IN), .ZN(
        n9742) );
  INV_X1 U12361 ( .A(n9750), .ZN(n9740) );
  NAND3_X1 U12362 ( .A1(n9740), .A2(n12159), .A3(n12103), .ZN(n9741) );
  NAND2_X1 U12363 ( .A1(n9742), .A2(n9741), .ZN(n10212) );
  NOR2_X1 U12364 ( .A1(n10212), .A2(n12615), .ZN(n10088) );
  INV_X1 U12365 ( .A(n9838), .ZN(n9743) );
  NAND2_X1 U12366 ( .A1(n9752), .A2(n9743), .ZN(n9747) );
  INV_X1 U12367 ( .A(n9744), .ZN(n9745) );
  NAND2_X1 U12368 ( .A1(n9750), .A2(n9745), .ZN(n9746) );
  NAND2_X1 U12369 ( .A1(n9747), .A2(n9746), .ZN(n9748) );
  INV_X1 U12370 ( .A(n11991), .ZN(n9867) );
  NAND2_X1 U12371 ( .A1(n12182), .A2(n11559), .ZN(n11988) );
  NAND2_X1 U12372 ( .A1(n9867), .A2(n11988), .ZN(n11966) );
  INV_X1 U12373 ( .A(n12152), .ZN(n12161) );
  AND2_X1 U12374 ( .A1(n12159), .A2(n12161), .ZN(n9749) );
  AND2_X1 U12375 ( .A1(n9750), .A2(n9749), .ZN(n9871) );
  AND2_X1 U12376 ( .A1(n12159), .A2(n15508), .ZN(n9751) );
  NAND2_X1 U12377 ( .A1(n9752), .A2(n9751), .ZN(n9754) );
  NOR2_X1 U12378 ( .A1(n12151), .A2(n15515), .ZN(n9753) );
  OAI22_X1 U12379 ( .A1(n11547), .A2(n11933), .B1(n11935), .B2(n11559), .ZN(
        n9755) );
  AOI21_X1 U12380 ( .B1(n11920), .B2(n11966), .A(n9755), .ZN(n9756) );
  OAI21_X1 U12381 ( .B1(n10088), .B2(n9757), .A(n9756), .ZN(P3_U3172) );
  INV_X1 U12382 ( .A(n14122), .ZN(n14334) );
  XNOR2_X1 U12383 ( .A(n15147), .B(n14334), .ZN(n14273) );
  XOR2_X1 U12384 ( .A(n9758), .B(n14273), .Z(n9759) );
  AOI222_X1 U12385 ( .A1(n15139), .A2(n9759), .B1(n14335), .B2(n14554), .C1(
        n14333), .C2(n15059), .ZN(n15146) );
  NAND4_X1 U12386 ( .A1(n9762), .A2(n14309), .A3(n9761), .A4(n9760), .ZN(
        n14431) );
  MUX2_X1 U12387 ( .A(n9763), .B(n15146), .S(n15104), .Z(n9772) );
  XNOR2_X1 U12388 ( .A(n9764), .B(n14273), .ZN(n15149) );
  NAND2_X1 U12389 ( .A1(n9765), .A2(n14598), .ZN(n14094) );
  NAND2_X1 U12390 ( .A1(n15068), .A2(n14094), .ZN(n9766) );
  INV_X1 U12391 ( .A(n14623), .ZN(n15102) );
  OAI211_X1 U12392 ( .C1(n6818), .C2(n15147), .A(n8988), .B(n9937), .ZN(n15145) );
  NOR2_X1 U12393 ( .A1(n15145), .A2(n14583), .ZN(n9770) );
  INV_X1 U12394 ( .A(n15092), .ZN(n9768) );
  OAI22_X1 U12395 ( .A1(n14541), .A2(n15147), .B1(n10054), .B2(n15091), .ZN(
        n9769) );
  AOI211_X1 U12396 ( .C1(n15149), .C2(n15102), .A(n9770), .B(n9769), .ZN(n9771) );
  NAND2_X1 U12397 ( .A1(n9772), .A2(n9771), .ZN(P1_U3289) );
  INV_X1 U12398 ( .A(n9773), .ZN(n9774) );
  INV_X1 U12399 ( .A(n13163), .ZN(n13168) );
  INV_X1 U12400 ( .A(n13167), .ZN(n12806) );
  NAND2_X1 U12401 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9962) );
  OAI21_X1 U12402 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9962), .ZN(n12788) );
  NAND2_X1 U12403 ( .A1(n9306), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U12404 ( .A1(n13072), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U12405 ( .A1(n6551), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9775) );
  OAI22_X1 U12406 ( .A1(n7410), .A2(n12806), .B1(n10065), .B2(n12808), .ZN(
        n10479) );
  NOR2_X1 U12407 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9465), .ZN(n15222) );
  NOR2_X1 U12408 ( .A1(n9778), .A2(n6561), .ZN(n13459) );
  NAND2_X1 U12409 ( .A1(n9807), .A2(n13459), .ZN(n9780) );
  INV_X1 U12410 ( .A(n9784), .ZN(n9779) );
  NAND2_X1 U12411 ( .A1(n9785), .A2(n9784), .ZN(n9789) );
  AND2_X1 U12412 ( .A1(n9787), .A2(n9786), .ZN(n9788) );
  NAND2_X1 U12413 ( .A1(n9789), .A2(n9788), .ZN(n9846) );
  NAND2_X1 U12414 ( .A1(n9846), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12825) );
  OAI22_X1 U12415 ( .A1(n12866), .A2(n10472), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n12825), .ZN(n9790) );
  AOI211_X1 U12416 ( .C1(n12838), .C2(n10479), .A(n15222), .B(n9790), .ZN(
        n9812) );
  NAND2_X1 U12417 ( .A1(n10347), .A2(n13164), .ZN(n9796) );
  XNOR2_X1 U12418 ( .A(n9796), .B(n13470), .ZN(n10203) );
  OR2_X2 U12419 ( .A1(n6550), .A2(n6984), .ZN(n9845) );
  NAND2_X1 U12420 ( .A1(n9845), .A2(n13212), .ZN(n9793) );
  XNOR2_X1 U12421 ( .A(n10203), .B(n9793), .ZN(n9912) );
  OR2_X1 U12422 ( .A1(n9796), .A2(n15312), .ZN(n9907) );
  NAND2_X1 U12423 ( .A1(n9911), .A2(n9845), .ZN(n9791) );
  AND2_X1 U12424 ( .A1(n9907), .A2(n9791), .ZN(n9792) );
  NAND2_X1 U12425 ( .A1(n9912), .A2(n9792), .ZN(n9908) );
  INV_X1 U12426 ( .A(n10203), .ZN(n9794) );
  NAND2_X1 U12427 ( .A1(n9794), .A2(n9793), .ZN(n9795) );
  XNOR2_X1 U12428 ( .A(n9796), .B(n12888), .ZN(n9797) );
  NAND2_X1 U12429 ( .A1(n9845), .A2(n13211), .ZN(n9798) );
  XNOR2_X1 U12430 ( .A(n9797), .B(n9798), .ZN(n10204) );
  INV_X1 U12431 ( .A(n9797), .ZN(n9799) );
  NAND2_X1 U12432 ( .A1(n9799), .A2(n9798), .ZN(n9800) );
  XNOR2_X1 U12433 ( .A(n9796), .B(n15370), .ZN(n12791) );
  NAND2_X1 U12434 ( .A1(n9845), .A2(n13210), .ZN(n9802) );
  INV_X1 U12435 ( .A(n9802), .ZN(n9801) );
  NAND2_X1 U12436 ( .A1(n12791), .A2(n9801), .ZN(n10058) );
  INV_X1 U12437 ( .A(n12791), .ZN(n9803) );
  NAND2_X1 U12438 ( .A1(n9803), .A2(n9802), .ZN(n9804) );
  NAND2_X1 U12439 ( .A1(n10058), .A2(n9804), .ZN(n9808) );
  NOR2_X1 U12440 ( .A1(n15421), .A2(n9805), .ZN(n9806) );
  AOI21_X1 U12441 ( .B1(n9809), .B2(n9808), .A(n12854), .ZN(n9810) );
  NAND2_X1 U12442 ( .A1(n9810), .A2(n12785), .ZN(n9811) );
  NAND2_X1 U12443 ( .A1(n9812), .A2(n9811), .ZN(P2_U3190) );
  MUX2_X1 U12444 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12275), .Z(n9881) );
  XNOR2_X1 U12445 ( .A(n9881), .B(n9882), .ZN(n9879) );
  NAND2_X1 U12446 ( .A1(n9814), .A2(n9813), .ZN(n9819) );
  INV_X1 U12447 ( .A(n9815), .ZN(n9817) );
  NAND2_X1 U12448 ( .A1(n9817), .A2(n9816), .ZN(n9818) );
  NAND2_X1 U12449 ( .A1(n9819), .A2(n9818), .ZN(n9880) );
  XOR2_X1 U12450 ( .A(n9879), .B(n9880), .Z(n9832) );
  XNOR2_X1 U12451 ( .A(n9896), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U12452 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8419), .ZN(n10561) );
  INV_X1 U12453 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10525) );
  INV_X1 U12454 ( .A(n9822), .ZN(n9823) );
  AOI21_X1 U12455 ( .B1(n10525), .B2(n9825), .A(n9888), .ZN(n9826) );
  NOR2_X1 U12456 ( .A1(n9826), .A2(n15465), .ZN(n9827) );
  AOI211_X1 U12457 ( .C1(n15458), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n10561), .B(
        n9827), .ZN(n9828) );
  OAI21_X1 U12458 ( .B1(n9895), .B2(n15452), .A(n9828), .ZN(n9829) );
  AOI21_X1 U12459 ( .B1(n15461), .B2(n9830), .A(n9829), .ZN(n9831) );
  OAI21_X1 U12460 ( .B1(n9832), .B2(n15454), .A(n9831), .ZN(P3_U3187) );
  OAI222_X1 U12461 ( .A1(n12627), .A2(n9834), .B1(n12623), .B2(n9833), .C1(
        P3_U3151), .C2(n11990), .ZN(P3_U3274) );
  INV_X1 U12462 ( .A(n15037), .ZN(n10960) );
  OAI222_X1 U12463 ( .A1(n14755), .A2(n9835), .B1(n14753), .B2(n11369), .C1(
        n10960), .C2(P1_U3086), .ZN(P1_U3337) );
  NAND2_X1 U12464 ( .A1(n9656), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9836) );
  XNOR2_X1 U12465 ( .A(n9836), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13234) );
  INV_X1 U12466 ( .A(n13234), .ZN(n11061) );
  OAI222_X1 U12467 ( .A1(n13905), .A2(n9837), .B1(n13908), .B2(n11369), .C1(
        n11061), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U12468 ( .A(n12556), .ZN(n12494) );
  NAND2_X1 U12469 ( .A1(n9838), .A2(n12404), .ZN(n9839) );
  NAND2_X1 U12470 ( .A1(n11966), .A2(n9839), .ZN(n9841) );
  NAND2_X1 U12471 ( .A1(n9514), .A2(n12479), .ZN(n9840) );
  NAND2_X1 U12472 ( .A1(n9841), .A2(n9840), .ZN(n11555) );
  MUX2_X1 U12473 ( .A(P3_REG1_REG_0__SCAN_IN), .B(n11555), .S(n15540), .Z(
        n9842) );
  AOI21_X1 U12474 ( .B1(n12494), .B2(n9843), .A(n9842), .ZN(n9844) );
  INV_X1 U12475 ( .A(n9844), .ZN(P3_U3459) );
  INV_X1 U12476 ( .A(n9845), .ZN(n12677) );
  AOI21_X1 U12477 ( .B1(n12677), .B2(n12846), .A(n12831), .ZN(n9851) );
  NOR2_X1 U12478 ( .A1(n9846), .A2(P2_U3088), .ZN(n10201) );
  INV_X1 U12479 ( .A(n10201), .ZN(n9915) );
  AND2_X1 U12480 ( .A1(n12848), .A2(n13212), .ZN(n15309) );
  AOI22_X1 U12481 ( .A1(n9915), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n12838), .B2(
        n15309), .ZN(n9850) );
  INV_X1 U12482 ( .A(n12852), .ZN(n12818) );
  NAND2_X1 U12483 ( .A1(n9847), .A2(n12876), .ZN(n12871) );
  NAND2_X1 U12484 ( .A1(n9848), .A2(n12871), .ZN(n15362) );
  NAND2_X1 U12485 ( .A1(n12818), .A2(n15362), .ZN(n9849) );
  OAI211_X1 U12486 ( .C1(n9851), .C2(n12876), .A(n9850), .B(n9849), .ZN(
        P2_U3204) );
  XNOR2_X1 U12487 ( .A(n9852), .B(n14275), .ZN(n15164) );
  OAI21_X1 U12488 ( .B1(n9853), .B2(n14275), .A(n9854), .ZN(n9857) );
  NAND2_X1 U12489 ( .A1(n14333), .A2(n14554), .ZN(n9856) );
  NAND2_X1 U12490 ( .A1(n14331), .A2(n15059), .ZN(n9855) );
  NAND2_X1 U12491 ( .A1(n9856), .A2(n9855), .ZN(n10314) );
  AOI21_X1 U12492 ( .B1(n9857), .B2(n15139), .A(n10314), .ZN(n15162) );
  MUX2_X1 U12493 ( .A(n9858), .B(n15162), .S(n15104), .Z(n9862) );
  INV_X1 U12494 ( .A(n9936), .ZN(n9859) );
  AOI211_X1 U12495 ( .C1(n15160), .C2(n9859), .A(n14589), .B(n10095), .ZN(
        n15158) );
  OAI22_X1 U12496 ( .A1(n14541), .A2(n10317), .B1(n10311), .B2(n15091), .ZN(
        n9860) );
  AOI21_X1 U12497 ( .B1(n15158), .B2(n15101), .A(n9860), .ZN(n9861) );
  OAI211_X1 U12498 ( .C1(n14623), .C2(n15164), .A(n9862), .B(n9861), .ZN(
        P1_U3287) );
  INV_X1 U12499 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n9875) );
  AOI21_X1 U12500 ( .B1(n11544), .B2(n11990), .A(n12157), .ZN(n9863) );
  OAI21_X1 U12501 ( .B1(n10291), .B2(n11807), .A(n9864), .ZN(n9865) );
  NAND3_X1 U12502 ( .A1(n11967), .A2(n11807), .A3(n9867), .ZN(n9868) );
  OAI211_X1 U12503 ( .C1(n9869), .C2(n8835), .A(n10079), .B(n9868), .ZN(n9870)
         );
  NAND2_X1 U12504 ( .A1(n9870), .A2(n11920), .ZN(n9874) );
  OAI22_X1 U12505 ( .A1(n11998), .A2(n11933), .B1(n11935), .B2(n10290), .ZN(
        n9872) );
  AOI21_X1 U12506 ( .B1(n11931), .B2(n12182), .A(n9872), .ZN(n9873) );
  OAI211_X1 U12507 ( .C1(n10088), .C2(n9875), .A(n9874), .B(n9873), .ZN(
        P3_U3162) );
  INV_X1 U12508 ( .A(n9876), .ZN(n9878) );
  OAI22_X1 U12509 ( .A1(n12163), .A2(P3_U3151), .B1(SI_22_), .B2(n12623), .ZN(
        n9877) );
  AOI21_X1 U12510 ( .B1(n9878), .B2(n12617), .A(n9877), .ZN(P3_U3273) );
  MUX2_X1 U12511 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12275), .Z(n10166) );
  INV_X1 U12512 ( .A(n10172), .ZN(n10167) );
  XNOR2_X1 U12513 ( .A(n10166), .B(n10167), .ZN(n10164) );
  NAND2_X1 U12514 ( .A1(n9880), .A2(n9879), .ZN(n9885) );
  INV_X1 U12515 ( .A(n9881), .ZN(n9883) );
  NAND2_X1 U12516 ( .A1(n9883), .A2(n9882), .ZN(n9884) );
  NAND2_X1 U12517 ( .A1(n9885), .A2(n9884), .ZN(n10165) );
  XOR2_X1 U12518 ( .A(n10164), .B(n10165), .Z(n9903) );
  NAND2_X1 U12519 ( .A1(n10172), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10175) );
  OAI21_X1 U12520 ( .B1(n10172), .B2(P3_REG2_REG_6__SCAN_IN), .A(n10175), .ZN(
        n9889) );
  AOI21_X1 U12521 ( .B1(n6715), .B2(n9889), .A(n10177), .ZN(n9892) );
  INV_X1 U12522 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n9890) );
  NOR2_X1 U12523 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9890), .ZN(n10736) );
  AOI21_X1 U12524 ( .B1(n15458), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10736), .ZN(
        n9891) );
  OAI21_X1 U12525 ( .B1(n9892), .B2(n15465), .A(n9891), .ZN(n9901) );
  INV_X1 U12526 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15530) );
  MUX2_X1 U12527 ( .A(n15530), .B(P3_REG1_REG_6__SCAN_IN), .S(n10172), .Z(
        n9898) );
  INV_X1 U12528 ( .A(n9893), .ZN(n9894) );
  AOI21_X1 U12529 ( .B1(n9898), .B2(n9897), .A(n10171), .ZN(n9899) );
  NOR2_X1 U12530 ( .A1(n9899), .A2(n12258), .ZN(n9900) );
  AOI211_X1 U12531 ( .C1(n14907), .C2(n10167), .A(n9901), .B(n9900), .ZN(n9902) );
  OAI21_X1 U12532 ( .B1(n9903), .B2(n15454), .A(n9902), .ZN(P3_U3188) );
  OAI22_X1 U12533 ( .A1(n12613), .A2(n11559), .B1(n15519), .B2(n9904), .ZN(
        n9905) );
  AOI21_X1 U12534 ( .B1(n11555), .B2(n15519), .A(n9905), .ZN(n9906) );
  INV_X1 U12535 ( .A(n9906), .ZN(P3_U3390) );
  INV_X1 U12536 ( .A(n9907), .ZN(n9910) );
  INV_X1 U12537 ( .A(n9912), .ZN(n9909) );
  INV_X1 U12538 ( .A(n9908), .ZN(n10205) );
  AOI21_X1 U12539 ( .B1(n9910), .B2(n9909), .A(n10205), .ZN(n9918) );
  NOR3_X1 U12540 ( .A1(n12852), .A2(n9912), .A3(n6938), .ZN(n9913) );
  AOI21_X1 U12541 ( .B1(n13470), .B2(n12831), .A(n9913), .ZN(n9917) );
  AOI22_X1 U12542 ( .A1(n9915), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n12838), .B2(
        n9914), .ZN(n9916) );
  OAI211_X1 U12543 ( .C1(n9918), .C2(n12854), .A(n9917), .B(n9916), .ZN(
        P2_U3194) );
  INV_X1 U12544 ( .A(n14094), .ZN(n9919) );
  NAND2_X1 U12545 ( .A1(n15104), .A2(n9919), .ZN(n9941) );
  INV_X1 U12546 ( .A(n9941), .ZN(n15081) );
  INV_X1 U12547 ( .A(n15091), .ZN(n15073) );
  AOI22_X1 U12548 ( .A1(n15106), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n15073), .ZN(n9922) );
  NOR2_X1 U12549 ( .A1(n14583), .A2(n14589), .ZN(n14628) );
  NAND2_X1 U12550 ( .A1(n14628), .A2(n9920), .ZN(n9921) );
  OAI211_X1 U12551 ( .C1(n9923), .C2(n14541), .A(n9922), .B(n9921), .ZN(n9924)
         );
  AOI21_X1 U12552 ( .B1(n15081), .B2(n9925), .A(n9924), .ZN(n9926) );
  OAI21_X1 U12553 ( .B1(n15106), .B2(n9927), .A(n9926), .ZN(P1_U3292) );
  XNOR2_X1 U12554 ( .A(n9928), .B(n14272), .ZN(n9934) );
  INV_X1 U12555 ( .A(n9934), .ZN(n15155) );
  NAND2_X1 U12556 ( .A1(n9929), .A2(n14272), .ZN(n9930) );
  AOI21_X1 U12557 ( .B1(n9931), .B2(n9930), .A(n15084), .ZN(n9933) );
  OAI22_X1 U12558 ( .A1(n10305), .A2(n14608), .B1(n14122), .B2(n14606), .ZN(
        n9932) );
  AOI211_X1 U12559 ( .C1(n9934), .C2(n15167), .A(n9933), .B(n9932), .ZN(n15154) );
  MUX2_X1 U12560 ( .A(n9935), .B(n15154), .S(n15104), .Z(n9940) );
  AOI211_X1 U12561 ( .C1(n15152), .C2(n9937), .A(n14589), .B(n9936), .ZN(
        n15151) );
  INV_X1 U12562 ( .A(n15152), .ZN(n10190) );
  OAI22_X1 U12563 ( .A1(n14541), .A2(n10190), .B1(n15091), .B2(n10197), .ZN(
        n9938) );
  AOI21_X1 U12564 ( .B1(n15151), .B2(n15101), .A(n9938), .ZN(n9939) );
  OAI211_X1 U12565 ( .C1(n15155), .C2(n9941), .A(n9940), .B(n9939), .ZN(
        P1_U3288) );
  INV_X1 U12566 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10030) );
  NAND2_X1 U12567 ( .A1(n9945), .A2(n9944), .ZN(n9947) );
  OR2_X1 U12568 ( .A1(n13211), .A2(n12888), .ZN(n9946) );
  NAND2_X1 U12569 ( .A1(n9947), .A2(n9946), .ZN(n10469) );
  NAND2_X1 U12570 ( .A1(n10469), .A2(n10475), .ZN(n9949) );
  OR2_X1 U12571 ( .A1(n13210), .A2(n15370), .ZN(n9948) );
  NAND2_X1 U12572 ( .A1(n9949), .A2(n9948), .ZN(n10367) );
  NAND2_X1 U12573 ( .A1(n9950), .A2(n13068), .ZN(n9953) );
  AOI22_X1 U12574 ( .A1(n11382), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n11381), 
        .B2(n9951), .ZN(n9952) );
  NAND2_X1 U12575 ( .A1(n9953), .A2(n9952), .ZN(n12900) );
  NAND2_X1 U12576 ( .A1(n13209), .A2(n15380), .ZN(n9954) );
  NAND2_X1 U12577 ( .A1(n10418), .A2(n9954), .ZN(n13124) );
  NAND2_X1 U12578 ( .A1(n10367), .A2(n13124), .ZN(n9956) );
  NAND2_X1 U12579 ( .A1(n10065), .A2(n15380), .ZN(n9955) );
  NAND2_X1 U12580 ( .A1(n9957), .A2(n13068), .ZN(n9960) );
  AOI22_X1 U12581 ( .A1(n11382), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n11381), 
        .B2(n9958), .ZN(n9959) );
  NAND2_X1 U12582 ( .A1(n9960), .A2(n9959), .ZN(n15385) );
  INV_X1 U12583 ( .A(n15385), .ZN(n10429) );
  INV_X1 U12584 ( .A(n9962), .ZN(n9961) );
  NAND2_X1 U12585 ( .A1(n9961), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9976) );
  INV_X1 U12586 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n13814) );
  NAND2_X1 U12587 ( .A1(n9962), .A2(n13814), .ZN(n9963) );
  NAND2_X1 U12588 ( .A1(n9976), .A2(n9963), .ZN(n10428) );
  OR2_X1 U12589 ( .A1(n11492), .A2(n10428), .ZN(n9967) );
  NAND2_X1 U12590 ( .A1(n7659), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U12591 ( .A1(n13072), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U12592 ( .A1(n6551), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9964) );
  NAND4_X1 U12593 ( .A1(n9967), .A2(n9966), .A3(n9965), .A4(n9964), .ZN(n13208) );
  NAND2_X1 U12594 ( .A1(n10429), .A2(n13208), .ZN(n9968) );
  INV_X1 U12595 ( .A(n13208), .ZN(n10372) );
  NAND2_X1 U12596 ( .A1(n10372), .A2(n15385), .ZN(n10022) );
  NAND2_X1 U12597 ( .A1(n9968), .A2(n10022), .ZN(n13125) );
  NAND2_X1 U12598 ( .A1(n10417), .A2(n13125), .ZN(n9970) );
  NAND2_X1 U12599 ( .A1(n10429), .A2(n10372), .ZN(n9969) );
  AOI22_X1 U12600 ( .A1(n11382), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n11381), 
        .B2(n9972), .ZN(n9973) );
  NAND2_X1 U12601 ( .A1(n9306), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U12602 ( .A1(n6551), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9980) );
  INV_X1 U12603 ( .A(n9976), .ZN(n9974) );
  NAND2_X1 U12604 ( .A1(n9974), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9989) );
  INV_X1 U12605 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U12606 ( .A1(n9976), .A2(n9975), .ZN(n9977) );
  AND2_X1 U12607 ( .A1(n9989), .A2(n9977), .ZN(n12836) );
  NAND2_X1 U12608 ( .A1(n11502), .A2(n12836), .ZN(n9979) );
  NAND2_X1 U12609 ( .A1(n13072), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9978) );
  NAND4_X1 U12610 ( .A1(n9981), .A2(n9980), .A3(n9979), .A4(n9978), .ZN(n13207) );
  XNOR2_X1 U12611 ( .A(n15393), .B(n13207), .ZN(n13127) );
  INV_X1 U12612 ( .A(n13127), .ZN(n9982) );
  OR2_X1 U12613 ( .A1(n15393), .A2(n13207), .ZN(n9983) );
  NAND2_X1 U12614 ( .A1(n9984), .A2(n13068), .ZN(n9986) );
  AOI22_X1 U12615 ( .A1(n11382), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11381), 
        .B2(n13220), .ZN(n9985) );
  NAND2_X1 U12616 ( .A1(n9986), .A2(n9985), .ZN(n15402) );
  NAND2_X1 U12617 ( .A1(n6551), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U12618 ( .A1(n7659), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9993) );
  INV_X1 U12619 ( .A(n9989), .ZN(n9987) );
  NAND2_X1 U12620 ( .A1(n9987), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10002) );
  INV_X1 U12621 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U12622 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  AND2_X1 U12623 ( .A1(n10002), .A2(n9990), .ZN(n12638) );
  NAND2_X1 U12624 ( .A1(n11502), .A2(n12638), .ZN(n9992) );
  NAND2_X1 U12625 ( .A1(n13072), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9991) );
  NAND4_X1 U12626 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n13206) );
  XNOR2_X1 U12627 ( .A(n15402), .B(n13206), .ZN(n13128) );
  INV_X1 U12628 ( .A(n13128), .ZN(n9995) );
  OR2_X1 U12629 ( .A1(n15402), .A2(n13206), .ZN(n9996) );
  NAND2_X1 U12630 ( .A1(n9997), .A2(n13068), .ZN(n10000) );
  AOI22_X1 U12631 ( .A1(n11382), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11381), 
        .B2(n9998), .ZN(n9999) );
  NAND2_X1 U12632 ( .A1(n10000), .A2(n9999), .ZN(n12924) );
  NAND2_X1 U12633 ( .A1(n9306), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U12634 ( .A1(n13072), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10006) );
  INV_X1 U12635 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U12636 ( .A1(n10002), .A2(n10001), .ZN(n10003) );
  AND2_X1 U12637 ( .A1(n10009), .A2(n10003), .ZN(n10281) );
  NAND2_X1 U12638 ( .A1(n11502), .A2(n10281), .ZN(n10005) );
  NAND2_X1 U12639 ( .A1(n6551), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10004) );
  NAND4_X1 U12640 ( .A1(n10007), .A2(n10006), .A3(n10005), .A4(n10004), .ZN(
        n13205) );
  XNOR2_X1 U12641 ( .A(n12924), .B(n13205), .ZN(n13130) );
  XNOR2_X1 U12642 ( .A(n10349), .B(n13130), .ZN(n10445) );
  NAND2_X1 U12643 ( .A1(n9306), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U12644 ( .A1(n6551), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10013) );
  INV_X1 U12645 ( .A(n10009), .ZN(n10008) );
  NAND2_X1 U12646 ( .A1(n10008), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U12647 ( .A1(n10009), .A2(n10142), .ZN(n10010) );
  AND2_X1 U12648 ( .A1(n10134), .A2(n10010), .ZN(n10360) );
  NAND2_X1 U12649 ( .A1(n11502), .A2(n10360), .ZN(n10012) );
  NAND2_X1 U12650 ( .A1(n13072), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10011) );
  NAND4_X1 U12651 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n13203) );
  NAND2_X1 U12652 ( .A1(n12848), .A2(n13203), .ZN(n10016) );
  NAND2_X1 U12653 ( .A1(n13167), .A2(n13206), .ZN(n10015) );
  NAND2_X1 U12654 ( .A1(n10016), .A2(n10015), .ZN(n10435) );
  NAND2_X1 U12655 ( .A1(n10470), .A2(n15380), .ZN(n10425) );
  OR2_X1 U12656 ( .A1(n10425), .A2(n15385), .ZN(n10426) );
  INV_X1 U12657 ( .A(n15402), .ZN(n10453) );
  INV_X1 U12658 ( .A(n10017), .ZN(n10448) );
  INV_X1 U12659 ( .A(n12924), .ZN(n10438) );
  INV_X1 U12660 ( .A(n10358), .ZN(n10018) );
  AOI211_X1 U12661 ( .C1(n12924), .C2(n10448), .A(n13562), .B(n10018), .ZN(
        n10440) );
  AOI211_X1 U12662 ( .C1(n15421), .C2(n12924), .A(n10435), .B(n10440), .ZN(
        n10028) );
  NAND2_X1 U12663 ( .A1(n10476), .A2(n10474), .ZN(n10019) );
  INV_X1 U12664 ( .A(n10475), .ZN(n13122) );
  NAND2_X1 U12665 ( .A1(n10019), .A2(n13122), .ZN(n10478) );
  NAND2_X1 U12666 ( .A1(n10478), .A2(n10370), .ZN(n10020) );
  INV_X1 U12667 ( .A(n13124), .ZN(n10366) );
  NAND2_X1 U12668 ( .A1(n10020), .A2(n10366), .ZN(n10419) );
  NAND2_X1 U12669 ( .A1(n10419), .A2(n10418), .ZN(n10021) );
  INV_X1 U12670 ( .A(n13125), .ZN(n10416) );
  NAND2_X1 U12671 ( .A1(n10021), .A2(n10416), .ZN(n10421) );
  NAND2_X1 U12672 ( .A1(n10421), .A2(n10022), .ZN(n10405) );
  NAND2_X1 U12673 ( .A1(n10405), .A2(n13127), .ZN(n10404) );
  INV_X1 U12674 ( .A(n13207), .ZN(n12633) );
  NAND2_X1 U12675 ( .A1(n15393), .A2(n12633), .ZN(n10023) );
  INV_X1 U12676 ( .A(n13206), .ZN(n12918) );
  OR2_X1 U12677 ( .A1(n15402), .A2(n12918), .ZN(n10024) );
  INV_X1 U12678 ( .A(n13130), .ZN(n10025) );
  NAND2_X1 U12679 ( .A1(n10026), .A2(n10025), .ZN(n10441) );
  NAND3_X1 U12680 ( .A1(n10442), .A2(n10441), .A3(n15409), .ZN(n10027) );
  OAI211_X1 U12681 ( .C1(n15405), .C2(n10445), .A(n10028), .B(n10027), .ZN(
        n10031) );
  NAND2_X1 U12682 ( .A1(n10031), .A2(n15431), .ZN(n10029) );
  OAI21_X1 U12683 ( .B1(n15431), .B2(n10030), .A(n10029), .ZN(P2_U3454) );
  NAND2_X1 U12684 ( .A1(n10031), .A2(n15443), .ZN(n10032) );
  OAI21_X1 U12685 ( .B1(n15443), .B2(n10033), .A(n10032), .ZN(P2_U3507) );
  OAI22_X1 U12686 ( .A1(n7206), .A2(n11797), .B1(n14117), .B2(n11798), .ZN(
        n10040) );
  NAND2_X1 U12687 ( .A1(n11783), .A2(n14116), .ZN(n10034) );
  INV_X1 U12688 ( .A(n10035), .ZN(n10037) );
  OAI22_X1 U12689 ( .A1(n14122), .A2(n11797), .B1(n15147), .B2(n11798), .ZN(
        n10185) );
  INV_X1 U12690 ( .A(n10185), .ZN(n10041) );
  OAI22_X1 U12691 ( .A1(n14122), .A2(n11798), .B1(n15147), .B2(n11794), .ZN(
        n10042) );
  XNOR2_X1 U12692 ( .A(n10042), .B(n11795), .ZN(n10186) );
  XNOR2_X1 U12693 ( .A(n10187), .B(n10186), .ZN(n10057) );
  INV_X1 U12694 ( .A(n10043), .ZN(n10045) );
  AND2_X1 U12695 ( .A1(n10045), .A2(n10044), .ZN(n10046) );
  NAND2_X1 U12696 ( .A1(n10047), .A2(n10046), .ZN(n10049) );
  INV_X1 U12697 ( .A(n14311), .ZN(n10048) );
  AOI21_X2 U12698 ( .B1(n10049), .B2(P1_STATE_REG_SCAN_IN), .A(n10048), .ZN(
        n14026) );
  INV_X1 U12699 ( .A(n10050), .ZN(n10051) );
  AOI21_X1 U12700 ( .B1(n14023), .B2(n14333), .A(n10051), .ZN(n10053) );
  NAND2_X1 U12701 ( .A1(n14064), .A2(n14335), .ZN(n10052) );
  OAI211_X1 U12702 ( .C1(n14026), .C2(n10054), .A(n10053), .B(n10052), .ZN(
        n10055) );
  AOI21_X1 U12703 ( .B1(n14124), .B2(n9398), .A(n10055), .ZN(n10056) );
  OAI21_X1 U12704 ( .B1(n10057), .B2(n14074), .A(n10056), .ZN(P1_U3230) );
  XNOR2_X1 U12705 ( .A(n12732), .B(n12900), .ZN(n10060) );
  NAND2_X1 U12706 ( .A1(n9845), .A2(n13209), .ZN(n10061) );
  XNOR2_X1 U12707 ( .A(n10060), .B(n10061), .ZN(n12790) );
  AND2_X1 U12708 ( .A1(n12790), .A2(n10058), .ZN(n10059) );
  NAND2_X1 U12709 ( .A1(n12785), .A2(n10059), .ZN(n12784) );
  INV_X1 U12710 ( .A(n10060), .ZN(n10064) );
  NAND2_X1 U12711 ( .A1(n10064), .A2(n10061), .ZN(n10062) );
  NAND2_X1 U12712 ( .A1(n12784), .A2(n10062), .ZN(n10063) );
  INV_X2 U12713 ( .A(n12667), .ZN(n12684) );
  XNOR2_X1 U12714 ( .A(n12684), .B(n15385), .ZN(n10109) );
  NAND2_X1 U12715 ( .A1(n9845), .A2(n13208), .ZN(n10110) );
  XNOR2_X1 U12716 ( .A(n10109), .B(n10110), .ZN(n10066) );
  OAI22_X1 U12717 ( .A1(n12852), .A2(n10065), .B1(n10064), .B2(n12854), .ZN(
        n10067) );
  NAND3_X1 U12718 ( .A1(n10067), .A2(n7484), .A3(n12784), .ZN(n10074) );
  INV_X1 U12719 ( .A(n12825), .ZN(n12862) );
  INV_X1 U12720 ( .A(n10428), .ZN(n10068) );
  AOI22_X1 U12721 ( .A1(n15385), .A2(n12831), .B1(n12862), .B2(n10068), .ZN(
        n10072) );
  NAND2_X1 U12722 ( .A1(n12848), .A2(n13207), .ZN(n10070) );
  NAND2_X1 U12723 ( .A1(n13167), .A2(n13209), .ZN(n10069) );
  NAND2_X1 U12724 ( .A1(n10070), .A2(n10069), .ZN(n10422) );
  NAND2_X1 U12725 ( .A1(n12838), .A2(n10422), .ZN(n10071) );
  AND4_X1 U12726 ( .A1(n10074), .A2(n10073), .A3(n10072), .A4(n10071), .ZN(
        n10075) );
  OAI21_X1 U12727 ( .B1(n10113), .B2(n12854), .A(n10075), .ZN(P2_U3199) );
  INV_X1 U12728 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10087) );
  XNOR2_X1 U12729 ( .A(n10290), .B(n11655), .ZN(n10077) );
  NAND2_X1 U12730 ( .A1(n10077), .A2(n10076), .ZN(n10078) );
  NAND2_X1 U12731 ( .A1(n10079), .A2(n10078), .ZN(n10080) );
  OAI21_X1 U12732 ( .B1(n10081), .B2(n10080), .A(n10215), .ZN(n10082) );
  NAND2_X1 U12733 ( .A1(n10082), .A2(n11920), .ZN(n10086) );
  OAI22_X1 U12734 ( .A1(n8837), .A2(n11933), .B1(n11935), .B2(n10083), .ZN(
        n10084) );
  AOI21_X1 U12735 ( .B1(n11931), .B2(n9514), .A(n10084), .ZN(n10085) );
  OAI211_X1 U12736 ( .C1(n10088), .C2(n10087), .A(n10086), .B(n10085), .ZN(
        P3_U3177) );
  XNOR2_X1 U12737 ( .A(n10089), .B(n14276), .ZN(n10092) );
  NAND2_X1 U12738 ( .A1(n14332), .A2(n14554), .ZN(n10091) );
  NAND2_X1 U12739 ( .A1(n14330), .A2(n15059), .ZN(n10090) );
  NAND2_X1 U12740 ( .A1(n10091), .A2(n10090), .ZN(n10541) );
  AOI21_X1 U12741 ( .B1(n10092), .B2(n15139), .A(n10541), .ZN(n15170) );
  XNOR2_X1 U12742 ( .A(n10094), .B(n10093), .ZN(n15173) );
  NAND2_X1 U12743 ( .A1(n15173), .A2(n15102), .ZN(n10099) );
  OAI22_X1 U12744 ( .A1(n15104), .A2(n9157), .B1(n10539), .B2(n15091), .ZN(
        n10097) );
  OAI211_X1 U12745 ( .C1(n10095), .C2(n15171), .A(n8988), .B(n15097), .ZN(
        n15169) );
  NOR2_X1 U12746 ( .A1(n15169), .A2(n14583), .ZN(n10096) );
  AOI211_X1 U12747 ( .C1(n15075), .C2(n14135), .A(n10097), .B(n10096), .ZN(
        n10098) );
  OAI211_X1 U12748 ( .C1(n15170), .C2(n15106), .A(n10099), .B(n10098), .ZN(
        P1_U3286) );
  INV_X1 U12749 ( .A(n14627), .ZN(n14532) );
  INV_X1 U12750 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13943) );
  AOI22_X1 U12751 ( .A1(n15075), .A2(n14116), .B1(n13943), .B2(n15073), .ZN(
        n10103) );
  MUX2_X1 U12752 ( .A(n10101), .B(n10100), .S(n15106), .Z(n10102) );
  OAI211_X1 U12753 ( .C1(n10104), .C2(n14583), .A(n10103), .B(n10102), .ZN(
        n10105) );
  AOI21_X1 U12754 ( .B1(n10106), .B2(n15102), .A(n10105), .ZN(n10107) );
  OAI21_X1 U12755 ( .B1(n10108), .B2(n14532), .A(n10107), .ZN(P1_U3290) );
  INV_X1 U12756 ( .A(n10109), .ZN(n10111) );
  NAND2_X1 U12757 ( .A1(n10111), .A2(n10110), .ZN(n10112) );
  NAND2_X1 U12758 ( .A1(n9845), .A2(n13207), .ZN(n10116) );
  INV_X1 U12759 ( .A(n10116), .ZN(n10114) );
  NAND2_X1 U12760 ( .A1(n10115), .A2(n10114), .ZN(n10118) );
  NAND2_X1 U12761 ( .A1(n12634), .A2(n10116), .ZN(n10117) );
  XNOR2_X1 U12762 ( .A(n15402), .B(n12684), .ZN(n10120) );
  NAND2_X1 U12763 ( .A1(n9845), .A2(n13206), .ZN(n10121) );
  INV_X1 U12764 ( .A(n10121), .ZN(n10119) );
  NAND2_X1 U12765 ( .A1(n10120), .A2(n10119), .ZN(n10123) );
  INV_X1 U12766 ( .A(n10120), .ZN(n10278) );
  NAND2_X1 U12767 ( .A1(n10278), .A2(n10121), .ZN(n10122) );
  AND2_X1 U12768 ( .A1(n10123), .A2(n10122), .ZN(n12631) );
  XNOR2_X1 U12769 ( .A(n12924), .B(n12684), .ZN(n10125) );
  NAND2_X1 U12770 ( .A1(n9845), .A2(n13205), .ZN(n10126) );
  XNOR2_X1 U12771 ( .A(n10125), .B(n10126), .ZN(n10288) );
  AND2_X1 U12772 ( .A1(n10288), .A2(n10123), .ZN(n10124) );
  INV_X1 U12773 ( .A(n10125), .ZN(n10146) );
  NAND2_X1 U12774 ( .A1(n10146), .A2(n10126), .ZN(n10127) );
  NAND2_X1 U12775 ( .A1(n10128), .A2(n13068), .ZN(n10131) );
  AOI22_X1 U12776 ( .A1(n11382), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n11381), 
        .B2(n10129), .ZN(n10130) );
  XNOR2_X1 U12777 ( .A(n15412), .B(n12684), .ZN(n10657) );
  NAND2_X1 U12778 ( .A1(n9845), .A2(n13203), .ZN(n10658) );
  XNOR2_X1 U12779 ( .A(n10657), .B(n10658), .ZN(n10145) );
  NAND2_X1 U12780 ( .A1(n10132), .A2(n10145), .ZN(n10661) );
  NAND2_X1 U12781 ( .A1(n7659), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U12782 ( .A1(n6551), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10138) );
  INV_X1 U12783 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U12784 ( .A1(n10134), .A2(n10133), .ZN(n10135) );
  AND2_X1 U12785 ( .A1(n10392), .A2(n10135), .ZN(n10706) );
  NAND2_X1 U12786 ( .A1(n11502), .A2(n10706), .ZN(n10137) );
  NAND2_X1 U12787 ( .A1(n13072), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10136) );
  NAND4_X1 U12788 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n13202) );
  NAND2_X1 U12789 ( .A1(n12848), .A2(n13202), .ZN(n10141) );
  NAND2_X1 U12790 ( .A1(n13167), .A2(n13205), .ZN(n10140) );
  AND2_X1 U12791 ( .A1(n10141), .A2(n10140), .ZN(n10355) );
  OAI22_X1 U12792 ( .A1(n12860), .A2(n10355), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10142), .ZN(n10144) );
  INV_X1 U12793 ( .A(n15412), .ZN(n10359) );
  NOR2_X1 U12794 ( .A1(n12866), .A2(n10359), .ZN(n10143) );
  AOI211_X1 U12795 ( .C1(n12862), .C2(n10360), .A(n10144), .B(n10143), .ZN(
        n10150) );
  INV_X1 U12796 ( .A(n10145), .ZN(n10148) );
  INV_X1 U12797 ( .A(n13205), .ZN(n10352) );
  OAI22_X1 U12798 ( .A1(n12852), .A2(n10352), .B1(n10146), .B2(n12854), .ZN(
        n10147) );
  NAND3_X1 U12799 ( .A1(n10284), .A2(n10148), .A3(n10147), .ZN(n10149) );
  OAI211_X1 U12800 ( .C1(n10661), .C2(n12854), .A(n10150), .B(n10149), .ZN(
        P2_U3203) );
  INV_X1 U12801 ( .A(n11380), .ZN(n10152) );
  OAI222_X1 U12802 ( .A1(n13905), .A2(n10151), .B1(n13908), .B2(n10152), .C1(
        n13244), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U12803 ( .A1(n14755), .A2(n10153), .B1(n14753), .B2(n10152), .C1(
        P1_U3086), .C2(n14617), .ZN(P1_U3336) );
  NAND2_X1 U12804 ( .A1(n10154), .A2(n12617), .ZN(n10155) );
  OAI211_X1 U12805 ( .C1(n10156), .C2(n12623), .A(n10155), .B(n12165), .ZN(
        P3_U3272) );
  AOI22_X1 U12806 ( .A1(n15075), .A2(n14111), .B1(n15073), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10157) );
  OAI21_X1 U12807 ( .B1(n14583), .B2(n10158), .A(n10157), .ZN(n10161) );
  MUX2_X1 U12808 ( .A(n10159), .B(P1_REG2_REG_2__SCAN_IN), .S(n15106), .Z(
        n10160) );
  AOI211_X1 U12809 ( .C1(n15081), .C2(n10162), .A(n10161), .B(n10160), .ZN(
        n10163) );
  INV_X1 U12810 ( .A(n10163), .ZN(P1_U3291) );
  MUX2_X1 U12811 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12275), .Z(n10253) );
  XNOR2_X1 U12812 ( .A(n10253), .B(n10254), .ZN(n10251) );
  NAND2_X1 U12813 ( .A1(n10165), .A2(n10164), .ZN(n10170) );
  INV_X1 U12814 ( .A(n10166), .ZN(n10168) );
  NAND2_X1 U12815 ( .A1(n10168), .A2(n10167), .ZN(n10169) );
  NAND2_X1 U12816 ( .A1(n10170), .A2(n10169), .ZN(n10252) );
  XOR2_X1 U12817 ( .A(n10251), .B(n10252), .Z(n10184) );
  NAND2_X1 U12818 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10173), .ZN(n10260) );
  OAI21_X1 U12819 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10173), .A(n10260), .ZN(
        n10182) );
  AND2_X1 U12820 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10795) );
  AOI21_X1 U12821 ( .B1(n15458), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10795), .ZN(
        n10174) );
  OAI21_X1 U12822 ( .B1(n15452), .B2(n10259), .A(n10174), .ZN(n10181) );
  INV_X1 U12823 ( .A(n10175), .ZN(n10176) );
  NOR2_X1 U12824 ( .A1(n10177), .A2(n10176), .ZN(n10178) );
  NOR2_X1 U12825 ( .A1(n10178), .A2(n10254), .ZN(n10268) );
  INV_X1 U12826 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10267) );
  XNOR2_X1 U12827 ( .A(n10266), .B(n10267), .ZN(n10179) );
  NOR2_X1 U12828 ( .A1(n10179), .A2(n15465), .ZN(n10180) );
  AOI211_X1 U12829 ( .C1(n15461), .C2(n10182), .A(n10181), .B(n10180), .ZN(
        n10183) );
  OAI21_X1 U12830 ( .B1(n10184), .B2(n15454), .A(n10183), .ZN(P3_U3189) );
  AOI22_X1 U12831 ( .A1(n15152), .A2(n11783), .B1(n10307), .B2(n14333), .ZN(
        n10188) );
  XOR2_X1 U12832 ( .A(n11795), .B(n10188), .Z(n10192) );
  OAI22_X1 U12833 ( .A1(n10190), .A2(n11798), .B1(n10189), .B2(n11797), .ZN(
        n10191) );
  NAND2_X1 U12834 ( .A1(n10192), .A2(n10191), .ZN(n10304) );
  NAND2_X1 U12835 ( .A1(n6712), .A2(n10304), .ZN(n10193) );
  XNOR2_X1 U12836 ( .A(n6598), .B(n10193), .ZN(n10200) );
  AOI21_X1 U12837 ( .B1(n14023), .B2(n14332), .A(n10194), .ZN(n10196) );
  NAND2_X1 U12838 ( .A1(n14064), .A2(n14334), .ZN(n10195) );
  OAI211_X1 U12839 ( .C1(n14026), .C2(n10197), .A(n10196), .B(n10195), .ZN(
        n10198) );
  AOI21_X1 U12840 ( .B1(n15152), .B2(n9398), .A(n10198), .ZN(n10199) );
  OAI21_X1 U12841 ( .B1(n10200), .B2(n14074), .A(n10199), .ZN(P1_U3227) );
  INV_X1 U12842 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10499) );
  OAI22_X1 U12843 ( .A1(n12860), .A2(n10202), .B1(n10201), .B2(n10499), .ZN(
        n10208) );
  AOI22_X1 U12844 ( .A1(n12818), .A2(n13212), .B1(n12846), .B2(n10203), .ZN(
        n10206) );
  NOR3_X1 U12845 ( .A1(n10206), .A2(n10205), .A3(n10204), .ZN(n10207) );
  AOI211_X1 U12846 ( .C1(n12888), .C2(n12831), .A(n10208), .B(n10207), .ZN(
        n10209) );
  OAI21_X1 U12847 ( .B1(n10210), .B2(n12854), .A(n10209), .ZN(P2_U3209) );
  NAND2_X1 U12848 ( .A1(n10213), .A2(n11998), .ZN(n10214) );
  XNOR2_X1 U12849 ( .A(n10244), .B(n11807), .ZN(n10509) );
  XNOR2_X1 U12850 ( .A(n10509), .B(n8837), .ZN(n10216) );
  INV_X1 U12851 ( .A(n11920), .ZN(n11940) );
  AOI21_X1 U12852 ( .B1(n10217), .B2(n10216), .A(n11940), .ZN(n10218) );
  NAND2_X1 U12853 ( .A1(n10218), .A2(n6704), .ZN(n10222) );
  INV_X1 U12854 ( .A(n11931), .ZN(n11895) );
  OAI22_X1 U12855 ( .A1(n11895), .A2(n11998), .B1(n10559), .B2(n11933), .ZN(
        n10219) );
  AOI211_X1 U12856 ( .C1(n10244), .C2(n11904), .A(n10220), .B(n10219), .ZN(
        n10221) );
  OAI211_X1 U12857 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n10872), .A(n10222), .B(
        n10221), .ZN(P3_U3158) );
  NAND2_X1 U12858 ( .A1(n12181), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10223) );
  OAI21_X1 U12859 ( .B1(n11814), .B2(n12181), .A(n10223), .ZN(P3_U3520) );
  INV_X1 U12860 ( .A(n11545), .ZN(n10226) );
  OAI21_X1 U12861 ( .B1(n10226), .B2(n10225), .A(n10224), .ZN(n10228) );
  NAND3_X1 U12862 ( .A1(n10228), .A2(n12474), .A3(n10227), .ZN(n10230) );
  AOI22_X1 U12863 ( .A1(n12480), .A2(n12180), .B1(n12179), .B2(n12479), .ZN(
        n10229) );
  OAI211_X1 U12864 ( .C1(n11601), .C2(n15476), .A(n10230), .B(n10229), .ZN(
        n15478) );
  INV_X1 U12865 ( .A(n15478), .ZN(n10250) );
  NAND2_X1 U12866 ( .A1(n10235), .A2(n10231), .ZN(n10232) );
  NAND2_X1 U12867 ( .A1(n10232), .A2(n10233), .ZN(n10237) );
  INV_X1 U12868 ( .A(n10233), .ZN(n10234) );
  NAND2_X1 U12869 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  NAND2_X1 U12870 ( .A1(n10239), .A2(n10238), .ZN(n10241) );
  INV_X2 U12871 ( .A(n12490), .ZN(n12486) );
  INV_X1 U12872 ( .A(n15476), .ZN(n10248) );
  OR2_X1 U12873 ( .A1(n12151), .A2(n11990), .ZN(n10300) );
  INV_X1 U12874 ( .A(n10300), .ZN(n10240) );
  NAND2_X1 U12875 ( .A1(n12490), .A2(n10240), .ZN(n12299) );
  INV_X1 U12876 ( .A(n12299), .ZN(n10780) );
  INV_X1 U12877 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10246) );
  INV_X1 U12878 ( .A(n10241), .ZN(n10243) );
  AND2_X1 U12879 ( .A1(n15508), .A2(n12151), .ZN(n10242) );
  AOI22_X1 U12880 ( .A1(n12438), .A2(n10244), .B1(n12485), .B2(n8485), .ZN(
        n10245) );
  OAI21_X1 U12881 ( .B1(n10246), .B2(n12490), .A(n10245), .ZN(n10247) );
  AOI21_X1 U12882 ( .B1(n10248), .B2(n10780), .A(n10247), .ZN(n10249) );
  OAI21_X1 U12883 ( .B1(n10250), .B2(n12486), .A(n10249), .ZN(P3_U3230) );
  MUX2_X1 U12884 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12275), .Z(n10611) );
  XNOR2_X1 U12885 ( .A(n10611), .B(n10612), .ZN(n10609) );
  NAND2_X1 U12886 ( .A1(n10252), .A2(n10251), .ZN(n10257) );
  INV_X1 U12887 ( .A(n10253), .ZN(n10255) );
  NAND2_X1 U12888 ( .A1(n10255), .A2(n10254), .ZN(n10256) );
  NAND2_X1 U12889 ( .A1(n10257), .A2(n10256), .ZN(n10610) );
  XOR2_X1 U12890 ( .A(n10609), .B(n10610), .Z(n10277) );
  INV_X1 U12891 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15534) );
  AOI22_X1 U12892 ( .A1(n10612), .A2(n15534), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n10631), .ZN(n10263) );
  NAND2_X1 U12893 ( .A1(n10259), .A2(n10258), .ZN(n10261) );
  NAND2_X1 U12894 ( .A1(n10261), .A2(n10260), .ZN(n10262) );
  OAI21_X1 U12895 ( .B1(n10263), .B2(n10262), .A(n10622), .ZN(n10275) );
  INV_X1 U12896 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10264) );
  NOR2_X1 U12897 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10264), .ZN(n11076) );
  AOI21_X1 U12898 ( .B1(n15458), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11076), .ZN(
        n10265) );
  OAI21_X1 U12899 ( .B1(n15452), .B2(n10631), .A(n10265), .ZN(n10274) );
  NAND2_X1 U12900 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10631), .ZN(n10269) );
  OAI21_X1 U12901 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10631), .A(n10269), .ZN(
        n10270) );
  NOR2_X1 U12902 ( .A1(n10271), .A2(n10270), .ZN(n10630) );
  AOI21_X1 U12903 ( .B1(n10271), .B2(n10270), .A(n10630), .ZN(n10272) );
  NOR2_X1 U12904 ( .A1(n10272), .A2(n15465), .ZN(n10273) );
  AOI211_X1 U12905 ( .C1(n15461), .C2(n10275), .A(n10274), .B(n10273), .ZN(
        n10276) );
  OAI21_X1 U12906 ( .B1(n10277), .B2(n15454), .A(n10276), .ZN(P3_U3190) );
  INV_X1 U12907 ( .A(n12635), .ZN(n10280) );
  NOR3_X1 U12908 ( .A1(n12852), .A2(n10278), .A3(n12918), .ZN(n10279) );
  AOI21_X1 U12909 ( .B1(n10280), .B2(n12846), .A(n10279), .ZN(n10289) );
  INV_X1 U12910 ( .A(n10281), .ZN(n10433) );
  NAND2_X1 U12911 ( .A1(n12838), .A2(n10435), .ZN(n10283) );
  OAI211_X1 U12912 ( .C1(n12825), .C2(n10433), .A(n10283), .B(n10282), .ZN(
        n10286) );
  NOR2_X1 U12913 ( .A1(n10284), .A2(n12854), .ZN(n10285) );
  AOI211_X1 U12914 ( .C1(n12924), .C2(n12831), .A(n10286), .B(n10285), .ZN(
        n10287) );
  OAI21_X1 U12915 ( .B1(n10289), .B2(n10288), .A(n10287), .ZN(P2_U3193) );
  OR2_X1 U12916 ( .A1(n10290), .A2(n15515), .ZN(n12558) );
  NAND2_X1 U12917 ( .A1(n11987), .A2(n10291), .ZN(n10292) );
  NAND2_X1 U12918 ( .A1(n10293), .A2(n10292), .ZN(n10297) );
  NAND2_X1 U12919 ( .A1(n12180), .A2(n12479), .ZN(n10295) );
  NAND2_X1 U12920 ( .A1(n12182), .A2(n12480), .ZN(n10294) );
  NAND2_X1 U12921 ( .A1(n10295), .A2(n10294), .ZN(n10296) );
  AOI21_X1 U12922 ( .B1(n10297), .B2(n12474), .A(n10296), .ZN(n12560) );
  OAI21_X1 U12923 ( .B1(n11544), .B2(n12558), .A(n12560), .ZN(n10298) );
  MUX2_X1 U12924 ( .A(n10298), .B(P3_REG2_REG_1__SCAN_IN), .S(n12486), .Z(
        n10299) );
  INV_X1 U12925 ( .A(n10299), .ZN(n10303) );
  XNOR2_X1 U12926 ( .A(n11987), .B(n11991), .ZN(n12557) );
  NAND2_X1 U12927 ( .A1(n11601), .A2(n10300), .ZN(n10301) );
  INV_X1 U12928 ( .A(n12493), .ZN(n12457) );
  AOI22_X1 U12929 ( .A1(n12557), .A2(n12457), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n12485), .ZN(n10302) );
  NAND2_X1 U12930 ( .A1(n10303), .A2(n10302), .ZN(P3_U3232) );
  INV_X1 U12931 ( .A(n9398), .ZN(n14067) );
  OAI22_X1 U12932 ( .A1(n10317), .A2(n11794), .B1(n10305), .B2(n11798), .ZN(
        n10306) );
  XNOR2_X1 U12933 ( .A(n10306), .B(n11795), .ZN(n10529) );
  AND2_X1 U12934 ( .A1(n11787), .A2(n14332), .ZN(n10308) );
  AOI21_X1 U12935 ( .B1(n15160), .B2(n10307), .A(n10308), .ZN(n10532) );
  XNOR2_X1 U12936 ( .A(n10529), .B(n10532), .ZN(n10309) );
  NAND2_X1 U12937 ( .A1(n10310), .A2(n10309), .ZN(n10530) );
  OAI211_X1 U12938 ( .C1(n10310), .C2(n10309), .A(n10530), .B(n14052), .ZN(
        n10316) );
  INV_X1 U12939 ( .A(n14055), .ZN(n11282) );
  NOR2_X1 U12940 ( .A1(n14026), .A2(n10311), .ZN(n10312) );
  AOI211_X1 U12941 ( .C1(n11282), .C2(n10314), .A(n10313), .B(n10312), .ZN(
        n10315) );
  OAI211_X1 U12942 ( .C1(n10317), .C2(n14067), .A(n10316), .B(n10315), .ZN(
        P1_U3239) );
  OAI21_X1 U12943 ( .B1(n9564), .B2(n10325), .A(n10318), .ZN(n10319) );
  NOR2_X1 U12944 ( .A1(n10327), .A2(n10319), .ZN(n10320) );
  XNOR2_X1 U12945 ( .A(n10327), .B(n10319), .ZN(n15023) );
  NOR2_X1 U12946 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15023), .ZN(n15022) );
  NOR2_X1 U12947 ( .A1(n10320), .A2(n15022), .ZN(n10323) );
  INV_X1 U12948 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10321) );
  MUX2_X1 U12949 ( .A(n10321), .B(P1_REG2_REG_16__SCAN_IN), .S(n10488), .Z(
        n10322) );
  NAND2_X1 U12950 ( .A1(n10323), .A2(n10322), .ZN(n10483) );
  OAI211_X1 U12951 ( .C1(n10323), .C2(n10322), .A(n10483), .B(n15040), .ZN(
        n10333) );
  NAND2_X1 U12952 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13993)
         );
  XNOR2_X1 U12953 ( .A(n10488), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10486) );
  AOI21_X1 U12954 ( .B1(n10325), .B2(n8082), .A(n10324), .ZN(n10326) );
  NOR2_X1 U12955 ( .A1(n10327), .A2(n10326), .ZN(n10328) );
  XNOR2_X1 U12956 ( .A(n10327), .B(n10326), .ZN(n15021) );
  NOR2_X1 U12957 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n15021), .ZN(n15020) );
  NOR2_X1 U12958 ( .A1(n10328), .A2(n15020), .ZN(n10487) );
  XOR2_X1 U12959 ( .A(n10486), .B(n10487), .Z(n10329) );
  NAND2_X1 U12960 ( .A1(n15035), .A2(n10329), .ZN(n10330) );
  NAND2_X1 U12961 ( .A1(n13993), .A2(n10330), .ZN(n10331) );
  AOI21_X1 U12962 ( .B1(n15006), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10331), 
        .ZN(n10332) );
  OAI211_X1 U12963 ( .C1(n15029), .C2(n10488), .A(n10333), .B(n10332), .ZN(
        P1_U3259) );
  INV_X1 U12964 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n10342) );
  INV_X1 U12965 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n10336) );
  NAND2_X1 U12966 ( .A1(n8877), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U12967 ( .A1(n6567), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10334) );
  OAI211_X1 U12968 ( .C1(n10337), .C2(n10336), .A(n10335), .B(n10334), .ZN(
        n10338) );
  INV_X1 U12969 ( .A(n10338), .ZN(n10339) );
  INV_X1 U12970 ( .A(n12284), .ZN(n11961) );
  NAND2_X1 U12971 ( .A1(n11961), .A2(P3_U3897), .ZN(n10341) );
  OAI21_X1 U12972 ( .B1(P3_U3897), .B2(n10342), .A(n10341), .ZN(P3_U3522) );
  OR3_X1 U12973 ( .A1(n10344), .A2(n10343), .A3(n15357), .ZN(n10345) );
  INV_X1 U12974 ( .A(n12868), .ZN(n15315) );
  NAND2_X1 U12975 ( .A1(n10347), .A2(n15315), .ZN(n10348) );
  NAND2_X1 U12976 ( .A1(n12924), .A2(n13205), .ZN(n10350) );
  INV_X1 U12977 ( .A(n13203), .ZN(n12930) );
  XNOR2_X1 U12978 ( .A(n15412), .B(n12930), .ZN(n13132) );
  OAI21_X1 U12979 ( .B1(n10351), .B2(n13132), .A(n10381), .ZN(n15414) );
  INV_X1 U12980 ( .A(n13132), .ZN(n10353) );
  OAI211_X1 U12981 ( .C1(n10354), .C2(n10353), .A(n10388), .B(n15409), .ZN(
        n10356) );
  NAND2_X1 U12982 ( .A1(n10356), .A2(n10355), .ZN(n15416) );
  NAND2_X1 U12983 ( .A1(n15416), .A2(n13472), .ZN(n10365) );
  INV_X1 U12984 ( .A(n10384), .ZN(n10357) );
  AOI211_X1 U12985 ( .C1(n15412), .C2(n10358), .A(n13562), .B(n10357), .ZN(
        n15411) );
  NOR2_X1 U12986 ( .A1(n13420), .A2(n10359), .ZN(n10363) );
  INV_X1 U12987 ( .A(n10360), .ZN(n10361) );
  OAI22_X1 U12988 ( .A1(n13472), .A2(n9323), .B1(n10361), .B2(n13397), .ZN(
        n10362) );
  AOI211_X1 U12989 ( .C1(n15411), .C2(n13467), .A(n10363), .B(n10362), .ZN(
        n10364) );
  OAI211_X1 U12990 ( .C1(n13465), .C2(n15414), .A(n10365), .B(n10364), .ZN(
        P2_U3256) );
  XNOR2_X1 U12991 ( .A(n10367), .B(n10366), .ZN(n15376) );
  OAI211_X1 U12992 ( .C1(n10470), .C2(n15380), .A(n10425), .B(n13431), .ZN(
        n15377) );
  INV_X1 U12993 ( .A(n15377), .ZN(n10369) );
  OAI22_X1 U12994 ( .A1(n13420), .A2(n15380), .B1(n12788), .B2(n13397), .ZN(
        n10368) );
  AOI21_X1 U12995 ( .B1(n13467), .B2(n10369), .A(n10368), .ZN(n10375) );
  NAND3_X1 U12996 ( .A1(n10478), .A2(n13124), .A3(n10370), .ZN(n10371) );
  AOI21_X1 U12997 ( .B1(n10419), .B2(n10371), .A(n13575), .ZN(n10373) );
  OAI22_X1 U12998 ( .A1(n7155), .A2(n12806), .B1(n10372), .B2(n12808), .ZN(
        n12787) );
  NOR2_X1 U12999 ( .A1(n10373), .A2(n12787), .ZN(n15378) );
  MUX2_X1 U13000 ( .A(n9199), .B(n15378), .S(n13472), .Z(n10374) );
  OAI211_X1 U13001 ( .C1(n15376), .C2(n13465), .A(n10375), .B(n10374), .ZN(
        P2_U3261) );
  NAND2_X1 U13002 ( .A1(n10376), .A2(n13068), .ZN(n10379) );
  AOI22_X1 U13003 ( .A1(n11382), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n11381), 
        .B2(n10377), .ZN(n10378) );
  XNOR2_X1 U13004 ( .A(n15420), .B(n13202), .ZN(n13134) );
  NAND2_X1 U13005 ( .A1(n15412), .A2(n13203), .ZN(n10380) );
  NAND2_X1 U13006 ( .A1(n10381), .A2(n10380), .ZN(n10383) );
  INV_X1 U13007 ( .A(n10578), .ZN(n10382) );
  AOI21_X1 U13008 ( .B1(n13134), .B2(n10383), .A(n10382), .ZN(n15424) );
  AOI211_X1 U13009 ( .C1(n15420), .C2(n10384), .A(n13562), .B(n10651), .ZN(
        n15419) );
  INV_X2 U13010 ( .A(n13472), .ZN(n15320) );
  INV_X1 U13011 ( .A(n13397), .ZN(n15318) );
  AOI22_X1 U13012 ( .A1(n15320), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10706), 
        .B2(n15318), .ZN(n10385) );
  OAI21_X1 U13013 ( .B1(n7229), .B2(n13420), .A(n10385), .ZN(n10386) );
  AOI21_X1 U13014 ( .B1(n15419), .B2(n13467), .A(n10386), .ZN(n10402) );
  OR2_X1 U13015 ( .A1(n15412), .A2(n12930), .ZN(n10387) );
  NAND2_X1 U13016 ( .A1(n10388), .A2(n10387), .ZN(n10389) );
  NAND2_X1 U13017 ( .A1(n10389), .A2(n13134), .ZN(n10599) );
  OAI211_X1 U13018 ( .C1(n10389), .C2(n13134), .A(n10599), .B(n15409), .ZN(
        n10400) );
  NAND2_X1 U13019 ( .A1(n6551), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U13020 ( .A1(n9306), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10396) );
  INV_X1 U13021 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U13022 ( .A1(n10392), .A2(n10391), .ZN(n10393) );
  AND2_X1 U13023 ( .A1(n10571), .A2(n10393), .ZN(n10667) );
  NAND2_X1 U13024 ( .A1(n11502), .A2(n10667), .ZN(n10395) );
  NAND2_X1 U13025 ( .A1(n13072), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10394) );
  NAND4_X1 U13026 ( .A1(n10397), .A2(n10396), .A3(n10395), .A4(n10394), .ZN(
        n13201) );
  NAND2_X1 U13027 ( .A1(n12848), .A2(n13201), .ZN(n10399) );
  NAND2_X1 U13028 ( .A1(n13167), .A2(n13203), .ZN(n10398) );
  AND2_X1 U13029 ( .A1(n10399), .A2(n10398), .ZN(n10709) );
  NAND2_X1 U13030 ( .A1(n10400), .A2(n10709), .ZN(n15426) );
  NAND2_X1 U13031 ( .A1(n15426), .A2(n13472), .ZN(n10401) );
  OAI211_X1 U13032 ( .C1(n15424), .C2(n13465), .A(n10402), .B(n10401), .ZN(
        P2_U3255) );
  XNOR2_X1 U13033 ( .A(n10403), .B(n13127), .ZN(n15396) );
  OAI21_X1 U13034 ( .B1(n10405), .B2(n13127), .A(n10404), .ZN(n10408) );
  NAND2_X1 U13035 ( .A1(n12848), .A2(n13206), .ZN(n10407) );
  NAND2_X1 U13036 ( .A1(n13167), .A2(n13208), .ZN(n10406) );
  NAND2_X1 U13037 ( .A1(n10407), .A2(n10406), .ZN(n12837) );
  AOI21_X1 U13038 ( .B1(n10408), .B2(n15409), .A(n12837), .ZN(n15399) );
  MUX2_X1 U13039 ( .A(n9200), .B(n15399), .S(n13472), .Z(n10415) );
  NAND2_X1 U13040 ( .A1(n10426), .A2(n15393), .ZN(n10409) );
  NAND2_X1 U13041 ( .A1(n10409), .A2(n13431), .ZN(n10410) );
  NOR2_X1 U13042 ( .A1(n10449), .A2(n10410), .ZN(n15395) );
  INV_X1 U13043 ( .A(n15393), .ZN(n10412) );
  INV_X1 U13044 ( .A(n12836), .ZN(n10411) );
  OAI22_X1 U13045 ( .A1(n13420), .A2(n10412), .B1(n13397), .B2(n10411), .ZN(
        n10413) );
  AOI21_X1 U13046 ( .B1(n13467), .B2(n15395), .A(n10413), .ZN(n10414) );
  OAI211_X1 U13047 ( .C1(n13465), .C2(n15396), .A(n10415), .B(n10414), .ZN(
        P2_U3259) );
  XNOR2_X1 U13048 ( .A(n10417), .B(n10416), .ZN(n15388) );
  NAND3_X1 U13049 ( .A1(n10419), .A2(n13125), .A3(n10418), .ZN(n10420) );
  NAND2_X1 U13050 ( .A1(n10421), .A2(n10420), .ZN(n10423) );
  AOI21_X1 U13051 ( .B1(n10423), .B2(n15409), .A(n10422), .ZN(n15391) );
  MUX2_X1 U13052 ( .A(n10424), .B(n15391), .S(n13472), .Z(n10432) );
  AOI21_X1 U13053 ( .B1(n10425), .B2(n15385), .A(n13562), .ZN(n10427) );
  AND2_X1 U13054 ( .A1(n10427), .A2(n10426), .ZN(n15387) );
  OAI22_X1 U13055 ( .A1(n13420), .A2(n10429), .B1(n13397), .B2(n10428), .ZN(
        n10430) );
  AOI21_X1 U13056 ( .B1(n13467), .B2(n15387), .A(n10430), .ZN(n10431) );
  OAI211_X1 U13057 ( .C1(n15388), .C2(n13465), .A(n10432), .B(n10431), .ZN(
        P2_U3260) );
  NAND2_X1 U13058 ( .A1(n15320), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10437) );
  NOR2_X1 U13059 ( .A1(n13397), .A2(n10433), .ZN(n10434) );
  AOI21_X1 U13060 ( .B1(n13472), .B2(n10435), .A(n10434), .ZN(n10436) );
  OAI211_X1 U13061 ( .C1(n13420), .C2(n10438), .A(n10437), .B(n10436), .ZN(
        n10439) );
  AOI21_X1 U13062 ( .B1(n10440), .B2(n13467), .A(n10439), .ZN(n10444) );
  NAND3_X1 U13063 ( .A1(n10442), .A2(n10441), .A3(n13406), .ZN(n10443) );
  OAI211_X1 U13064 ( .C1(n10445), .C2(n13465), .A(n10444), .B(n10443), .ZN(
        P2_U3257) );
  XNOR2_X1 U13065 ( .A(n10446), .B(n13128), .ZN(n15406) );
  XNOR2_X1 U13066 ( .A(n10447), .B(n13128), .ZN(n15408) );
  NAND2_X1 U13067 ( .A1(n15408), .A2(n13406), .ZN(n10458) );
  OAI211_X1 U13068 ( .C1(n10453), .C2(n10449), .A(n10448), .B(n13431), .ZN(
        n15403) );
  INV_X1 U13069 ( .A(n15403), .ZN(n10456) );
  NAND2_X1 U13070 ( .A1(n12848), .A2(n13205), .ZN(n10451) );
  NAND2_X1 U13071 ( .A1(n13167), .A2(n13207), .ZN(n10450) );
  NAND2_X1 U13072 ( .A1(n10451), .A2(n10450), .ZN(n15401) );
  MUX2_X1 U13073 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n15401), .S(n13472), .Z(
        n10455) );
  INV_X1 U13074 ( .A(n12638), .ZN(n10452) );
  OAI22_X1 U13075 ( .A1(n13420), .A2(n10453), .B1(n13397), .B2(n10452), .ZN(
        n10454) );
  AOI211_X1 U13076 ( .C1(n10456), .C2(n13467), .A(n10455), .B(n10454), .ZN(
        n10457) );
  OAI211_X1 U13077 ( .C1(n15406), .C2(n13465), .A(n10458), .B(n10457), .ZN(
        P2_U3258) );
  XNOR2_X1 U13078 ( .A(n10459), .B(n10460), .ZN(n15481) );
  XNOR2_X1 U13079 ( .A(n10461), .B(n12008), .ZN(n10463) );
  OAI22_X1 U13080 ( .A1(n8837), .A2(n12406), .B1(n10734), .B2(n12408), .ZN(
        n10462) );
  AOI21_X1 U13081 ( .B1(n10463), .B2(n12474), .A(n10462), .ZN(n10464) );
  OAI21_X1 U13082 ( .B1(n11601), .B2(n15481), .A(n10464), .ZN(n15483) );
  INV_X1 U13083 ( .A(n15483), .ZN(n10465) );
  MUX2_X1 U13084 ( .A(n10466), .B(n10465), .S(n12490), .Z(n10468) );
  AOI22_X1 U13085 ( .A1(n12438), .A2(n12015), .B1(n12485), .B2(n10508), .ZN(
        n10467) );
  OAI211_X1 U13086 ( .C1(n15481), .C2(n12299), .A(n10468), .B(n10467), .ZN(
        P3_U3229) );
  XNOR2_X1 U13087 ( .A(n10469), .B(n13122), .ZN(n15373) );
  AOI211_X1 U13088 ( .C1(n15370), .C2(n10471), .A(n13562), .B(n10470), .ZN(
        n15369) );
  OAI22_X1 U13089 ( .A1(n13420), .A2(n10472), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13397), .ZN(n10473) );
  AOI21_X1 U13090 ( .B1(n13467), .B2(n15369), .A(n10473), .ZN(n10482) );
  NAND3_X1 U13091 ( .A1(n10476), .A2(n10475), .A3(n10474), .ZN(n10477) );
  AOI21_X1 U13092 ( .B1(n10478), .B2(n10477), .A(n13575), .ZN(n10480) );
  NOR2_X1 U13093 ( .A1(n10480), .A2(n10479), .ZN(n15372) );
  MUX2_X1 U13094 ( .A(n9198), .B(n15372), .S(n13472), .Z(n10481) );
  OAI211_X1 U13095 ( .C1(n15373), .C2(n13465), .A(n10482), .B(n10481), .ZN(
        P2_U3262) );
  OAI21_X1 U13096 ( .B1(n10321), .B2(n10488), .A(n10483), .ZN(n10956) );
  INV_X1 U13097 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10484) );
  XNOR2_X1 U13098 ( .A(n10957), .B(n10484), .ZN(n10955) );
  XNOR2_X1 U13099 ( .A(n10956), .B(n10955), .ZN(n10497) );
  NAND2_X1 U13100 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14005)
         );
  INV_X1 U13101 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10485) );
  XNOR2_X1 U13102 ( .A(n10957), .B(n10485), .ZN(n10947) );
  NAND2_X1 U13103 ( .A1(n10487), .A2(n10486), .ZN(n10491) );
  INV_X1 U13104 ( .A(n10488), .ZN(n10489) );
  NAND2_X1 U13105 ( .A1(n10489), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U13106 ( .A1(n10491), .A2(n10490), .ZN(n10948) );
  XOR2_X1 U13107 ( .A(n10947), .B(n10948), .Z(n10492) );
  NAND2_X1 U13108 ( .A1(n15035), .A2(n10492), .ZN(n10493) );
  NAND2_X1 U13109 ( .A1(n14005), .A2(n10493), .ZN(n10494) );
  AOI21_X1 U13110 ( .B1(n15006), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n10494), 
        .ZN(n10496) );
  NAND2_X1 U13111 ( .A1(n15038), .A2(n10957), .ZN(n10495) );
  OAI211_X1 U13112 ( .C1(n10497), .C2(n15025), .A(n10496), .B(n10495), .ZN(
        P1_U3260) );
  OAI222_X1 U13113 ( .A1(n14755), .A2(n10498), .B1(n14753), .B2(n11393), .C1(
        n14085), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI22_X1 U13114 ( .A1(n13472), .A2(n10500), .B1(n10499), .B2(n13397), .ZN(
        n10503) );
  NOR2_X1 U13115 ( .A1(n13465), .A2(n10501), .ZN(n10502) );
  AOI211_X1 U13116 ( .C1(n13472), .C2(n10504), .A(n10503), .B(n10502), .ZN(
        n10506) );
  NAND2_X1 U13117 ( .A1(n13471), .A2(n12888), .ZN(n10505) );
  OAI211_X1 U13118 ( .C1(n10507), .C2(n13440), .A(n10506), .B(n10505), .ZN(
        P2_U3263) );
  OAI222_X1 U13119 ( .A1(n13905), .A2(n11394), .B1(P2_U3088), .B2(n6561), .C1(
        n13908), .C2(n11393), .ZN(P2_U3307) );
  INV_X1 U13120 ( .A(n10508), .ZN(n10518) );
  XNOR2_X1 U13121 ( .A(n12015), .B(n11807), .ZN(n10510) );
  NAND2_X1 U13122 ( .A1(n10510), .A2(n10559), .ZN(n10555) );
  INV_X1 U13123 ( .A(n10510), .ZN(n10511) );
  NAND2_X1 U13124 ( .A1(n10511), .A2(n12179), .ZN(n10512) );
  AND2_X1 U13125 ( .A1(n10555), .A2(n10512), .ZN(n10552) );
  NAND2_X1 U13126 ( .A1(n6596), .A2(n10552), .ZN(n10549) );
  OAI21_X1 U13127 ( .B1(n6596), .B2(n10552), .A(n10549), .ZN(n10513) );
  NAND2_X1 U13128 ( .A1(n10513), .A2(n11920), .ZN(n10517) );
  OAI22_X1 U13129 ( .A1(n11895), .A2(n8837), .B1(n10734), .B2(n11933), .ZN(
        n10514) );
  AOI211_X1 U13130 ( .C1(n12015), .C2(n11904), .A(n10515), .B(n10514), .ZN(
        n10516) );
  OAI211_X1 U13131 ( .C1(n10518), .C2(n10872), .A(n10517), .B(n10516), .ZN(
        P3_U3170) );
  NOR2_X1 U13132 ( .A1(n10519), .A2(n12012), .ZN(n10745) );
  AOI21_X1 U13133 ( .B1(n12012), .B2(n10519), .A(n10745), .ZN(n10523) );
  AOI22_X1 U13134 ( .A1(n12178), .A2(n12479), .B1(n12480), .B2(n12179), .ZN(
        n10522) );
  XNOR2_X1 U13135 ( .A(n10520), .B(n12012), .ZN(n15485) );
  INV_X1 U13136 ( .A(n11601), .ZN(n10988) );
  NAND2_X1 U13137 ( .A1(n15485), .A2(n10988), .ZN(n10521) );
  OAI211_X1 U13138 ( .C1(n10523), .C2(n12404), .A(n10522), .B(n10521), .ZN(
        n15489) );
  INV_X1 U13139 ( .A(n15489), .ZN(n10528) );
  AOI22_X1 U13140 ( .A1(n12438), .A2(n10562), .B1(n12485), .B2(n10548), .ZN(
        n10524) );
  OAI21_X1 U13141 ( .B1(n10525), .B2(n12490), .A(n10524), .ZN(n10526) );
  AOI21_X1 U13142 ( .B1(n15485), .B2(n10780), .A(n10526), .ZN(n10527) );
  OAI21_X1 U13143 ( .B1(n10528), .B2(n12486), .A(n10527), .ZN(P3_U3228) );
  INV_X1 U13144 ( .A(n10529), .ZN(n10531) );
  OAI22_X1 U13145 ( .A1(n15171), .A2(n11794), .B1(n10533), .B2(n11798), .ZN(
        n10534) );
  XNOR2_X1 U13146 ( .A(n10534), .B(n11795), .ZN(n10692) );
  AND2_X1 U13147 ( .A1(n11787), .A2(n14331), .ZN(n10535) );
  AOI21_X1 U13148 ( .B1(n14135), .B2(n10307), .A(n10535), .ZN(n10693) );
  XNOR2_X1 U13149 ( .A(n10692), .B(n10693), .ZN(n10536) );
  OAI211_X1 U13150 ( .C1(n10537), .C2(n10536), .A(n10696), .B(n14052), .ZN(
        n10543) );
  NOR2_X1 U13151 ( .A1(n10538), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14383) );
  NOR2_X1 U13152 ( .A1(n14026), .A2(n10539), .ZN(n10540) );
  AOI211_X1 U13153 ( .C1(n11282), .C2(n10541), .A(n14383), .B(n10540), .ZN(
        n10542) );
  OAI211_X1 U13154 ( .C1(n15171), .C2(n14067), .A(n10543), .B(n10542), .ZN(
        P1_U3213) );
  INV_X1 U13155 ( .A(n10544), .ZN(n10546) );
  OAI222_X1 U13156 ( .A1(n10547), .A2(P3_U3151), .B1(n12627), .B2(n10546), 
        .C1(n10545), .C2(n12623), .ZN(P3_U3271) );
  INV_X1 U13157 ( .A(n10548), .ZN(n10565) );
  INV_X1 U13158 ( .A(n10549), .ZN(n10551) );
  INV_X1 U13159 ( .A(n10555), .ZN(n10550) );
  XNOR2_X1 U13160 ( .A(n10562), .B(n11655), .ZN(n10730) );
  XNOR2_X1 U13161 ( .A(n10730), .B(n10734), .ZN(n10554) );
  NOR3_X1 U13162 ( .A1(n10551), .A2(n10550), .A3(n10554), .ZN(n10558) );
  AND2_X1 U13163 ( .A1(n10552), .A2(n10554), .ZN(n10553) );
  INV_X1 U13164 ( .A(n10554), .ZN(n10556) );
  OR2_X1 U13165 ( .A1(n10556), .A2(n10555), .ZN(n10557) );
  OAI21_X1 U13166 ( .B1(n10558), .B2(n7077), .A(n11920), .ZN(n10564) );
  OAI22_X1 U13167 ( .A1(n11895), .A2(n10559), .B1(n10844), .B2(n11933), .ZN(
        n10560) );
  AOI211_X1 U13168 ( .C1(n10562), .C2(n11904), .A(n10561), .B(n10560), .ZN(
        n10563) );
  OAI211_X1 U13169 ( .C1(n10565), .C2(n10872), .A(n10564), .B(n10563), .ZN(
        P3_U3167) );
  NAND2_X1 U13170 ( .A1(n10566), .A2(n13068), .ZN(n10569) );
  AOI22_X1 U13171 ( .A1(n11382), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11381), 
        .B2(n10567), .ZN(n10568) );
  INV_X1 U13172 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10570) );
  NAND2_X1 U13173 ( .A1(n10571), .A2(n10570), .ZN(n10572) );
  NAND2_X1 U13174 ( .A1(n10586), .A2(n10572), .ZN(n10721) );
  OR2_X1 U13175 ( .A1(n11492), .A2(n10721), .ZN(n10576) );
  NAND2_X1 U13176 ( .A1(n9306), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10575) );
  NAND2_X1 U13177 ( .A1(n6551), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10574) );
  NAND2_X1 U13178 ( .A1(n13072), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10573) );
  NAND4_X1 U13179 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n13200) );
  XNOR2_X1 U13180 ( .A(n13855), .B(n13200), .ZN(n13133) );
  OR2_X1 U13181 ( .A1(n15420), .A2(n13202), .ZN(n10577) );
  NAND2_X1 U13182 ( .A1(n10579), .A2(n13068), .ZN(n10582) );
  AOI22_X1 U13183 ( .A1(n11382), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11381), 
        .B2(n10580), .ZN(n10581) );
  NOR2_X1 U13184 ( .A1(n12941), .A2(n13201), .ZN(n10583) );
  NAND2_X1 U13185 ( .A1(n12941), .A2(n13201), .ZN(n10584) );
  XOR2_X1 U13186 ( .A(n13133), .B(n10838), .Z(n13859) );
  INV_X1 U13187 ( .A(n12941), .ZN(n10684) );
  OR2_X2 U13188 ( .A1(n10650), .A2(n13855), .ZN(n10834) );
  INV_X1 U13189 ( .A(n10834), .ZN(n10585) );
  AOI211_X1 U13190 ( .C1(n13855), .C2(n10650), .A(n13562), .B(n10585), .ZN(
        n13853) );
  NAND2_X1 U13191 ( .A1(n13471), .A2(n13855), .ZN(n10596) );
  NAND2_X1 U13192 ( .A1(n7659), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10591) );
  NAND2_X1 U13193 ( .A1(n13072), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10590) );
  INV_X1 U13194 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n13591) );
  NAND2_X1 U13195 ( .A1(n10586), .A2(n13591), .ZN(n10587) );
  AND2_X1 U13196 ( .A1(n10825), .A2(n10587), .ZN(n11181) );
  NAND2_X1 U13197 ( .A1(n11502), .A2(n11181), .ZN(n10589) );
  NAND2_X1 U13198 ( .A1(n6551), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10588) );
  NAND4_X1 U13199 ( .A1(n10591), .A2(n10590), .A3(n10589), .A4(n10588), .ZN(
        n13199) );
  NAND2_X1 U13200 ( .A1(n12848), .A2(n13199), .ZN(n10593) );
  NAND2_X1 U13201 ( .A1(n13167), .A2(n13201), .ZN(n10592) );
  NAND2_X1 U13202 ( .A1(n10593), .A2(n10592), .ZN(n13854) );
  NOR2_X1 U13203 ( .A1(n13397), .A2(n10721), .ZN(n10594) );
  AOI21_X1 U13204 ( .B1(n13472), .B2(n13854), .A(n10594), .ZN(n10595) );
  OAI211_X1 U13205 ( .C1(n13472), .C2(n11037), .A(n10596), .B(n10595), .ZN(
        n10597) );
  AOI21_X1 U13206 ( .B1(n13853), .B2(n13467), .A(n10597), .ZN(n10603) );
  INV_X1 U13207 ( .A(n13202), .ZN(n10672) );
  OR2_X1 U13208 ( .A1(n15420), .A2(n10672), .ZN(n10598) );
  INV_X1 U13209 ( .A(n13201), .ZN(n10600) );
  XNOR2_X1 U13210 ( .A(n12941), .B(n10600), .ZN(n13138) );
  NAND2_X1 U13211 ( .A1(n12941), .A2(n10600), .ZN(n10601) );
  XNOR2_X1 U13212 ( .A(n10821), .B(n13133), .ZN(n13856) );
  NAND2_X1 U13213 ( .A1(n13856), .A2(n13406), .ZN(n10602) );
  OAI211_X1 U13214 ( .C1(n13859), .C2(n13465), .A(n10603), .B(n10602), .ZN(
        P2_U3253) );
  INV_X1 U13215 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10605) );
  INV_X1 U13216 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10604) );
  MUX2_X1 U13217 ( .A(n10605), .B(n10604), .S(n12275), .Z(n10606) );
  NAND2_X1 U13218 ( .A1(n10606), .A2(n10805), .ZN(n10810) );
  INV_X1 U13219 ( .A(n10606), .ZN(n10607) );
  NAND2_X1 U13220 ( .A1(n10607), .A2(n10802), .ZN(n10608) );
  NAND2_X1 U13221 ( .A1(n10810), .A2(n10608), .ZN(n10621) );
  NAND2_X1 U13222 ( .A1(n10610), .A2(n10609), .ZN(n10615) );
  INV_X1 U13223 ( .A(n10611), .ZN(n10613) );
  NAND2_X1 U13224 ( .A1(n10613), .A2(n10612), .ZN(n10614) );
  NAND2_X1 U13225 ( .A1(n10615), .A2(n10614), .ZN(n15451) );
  INV_X1 U13226 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15446) );
  INV_X1 U13227 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15536) );
  MUX2_X1 U13228 ( .A(n15446), .B(n15536), .S(n12275), .Z(n10616) );
  AND2_X1 U13229 ( .A1(n10616), .A2(n10632), .ZN(n15447) );
  INV_X1 U13230 ( .A(n10616), .ZN(n10617) );
  NAND2_X1 U13231 ( .A1(n10617), .A2(n15453), .ZN(n15448) );
  NAND2_X1 U13232 ( .A1(n10618), .A2(n15448), .ZN(n10620) );
  INV_X1 U13233 ( .A(n10811), .ZN(n10619) );
  AOI21_X1 U13234 ( .B1(n10621), .B2(n10620), .A(n10619), .ZN(n10642) );
  AOI22_X1 U13235 ( .A1(n10805), .A2(n10604), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n10802), .ZN(n10627) );
  NAND2_X1 U13236 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10631), .ZN(n10623) );
  NAND2_X1 U13237 ( .A1(n15453), .A2(n10624), .ZN(n10625) );
  XNOR2_X1 U13238 ( .A(n10624), .B(n10632), .ZN(n15460) );
  OAI21_X1 U13239 ( .B1(n10627), .B2(n10626), .A(n10804), .ZN(n10640) );
  INV_X1 U13240 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n10628) );
  NOR2_X1 U13241 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10628), .ZN(n10868) );
  AOI21_X1 U13242 ( .B1(n15458), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n10868), 
        .ZN(n10629) );
  OAI21_X1 U13243 ( .B1(n15452), .B2(n10802), .A(n10629), .ZN(n10639) );
  NOR2_X1 U13244 ( .A1(n10632), .A2(n10633), .ZN(n10634) );
  XOR2_X1 U13245 ( .A(n10633), .B(n15453), .Z(n15445) );
  AOI22_X1 U13246 ( .A1(n10805), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n10605), 
        .B2(n10802), .ZN(n10635) );
  AOI21_X1 U13247 ( .B1(n10636), .B2(n10635), .A(n10801), .ZN(n10637) );
  NOR2_X1 U13248 ( .A1(n10637), .A2(n15465), .ZN(n10638) );
  AOI211_X1 U13249 ( .C1(n15461), .C2(n10640), .A(n10639), .B(n10638), .ZN(
        n10641) );
  OAI21_X1 U13250 ( .B1(n10642), .B2(n15454), .A(n10641), .ZN(P3_U3192) );
  XNOR2_X1 U13251 ( .A(n10643), .B(n13138), .ZN(n10687) );
  INV_X1 U13252 ( .A(n10687), .ZN(n10656) );
  INV_X1 U13253 ( .A(n10644), .ZN(n10645) );
  AOI21_X1 U13254 ( .B1(n13138), .B2(n10646), .A(n10645), .ZN(n10649) );
  NAND2_X1 U13255 ( .A1(n12848), .A2(n13200), .ZN(n10648) );
  NAND2_X1 U13256 ( .A1(n13167), .A2(n13202), .ZN(n10647) );
  AND2_X1 U13257 ( .A1(n10648), .A2(n10647), .ZN(n10670) );
  OAI21_X1 U13258 ( .B1(n10649), .B2(n13575), .A(n10670), .ZN(n10685) );
  OAI211_X1 U13259 ( .C1(n10684), .C2(n10651), .A(n13431), .B(n10650), .ZN(
        n10683) );
  AOI22_X1 U13260 ( .A1(n15320), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10667), 
        .B2(n15318), .ZN(n10653) );
  NAND2_X1 U13261 ( .A1(n12941), .A2(n13471), .ZN(n10652) );
  OAI211_X1 U13262 ( .C1(n10683), .C2(n13440), .A(n10653), .B(n10652), .ZN(
        n10654) );
  AOI21_X1 U13263 ( .B1(n10685), .B2(n13472), .A(n10654), .ZN(n10655) );
  OAI21_X1 U13264 ( .B1(n13465), .B2(n10656), .A(n10655), .ZN(P2_U3254) );
  INV_X1 U13265 ( .A(n10657), .ZN(n10659) );
  NAND2_X1 U13266 ( .A1(n10659), .A2(n10658), .ZN(n10660) );
  NAND2_X1 U13267 ( .A1(n10661), .A2(n10660), .ZN(n10711) );
  XNOR2_X1 U13268 ( .A(n15420), .B(n12684), .ZN(n10663) );
  NAND2_X1 U13269 ( .A1(n9845), .A2(n13202), .ZN(n10664) );
  INV_X1 U13270 ( .A(n10664), .ZN(n10662) );
  NAND2_X1 U13271 ( .A1(n10663), .A2(n10662), .ZN(n10666) );
  INV_X1 U13272 ( .A(n10663), .ZN(n10673) );
  NAND2_X1 U13273 ( .A1(n10673), .A2(n10664), .ZN(n10665) );
  NAND2_X1 U13274 ( .A1(n10666), .A2(n10665), .ZN(n10712) );
  XNOR2_X1 U13275 ( .A(n12941), .B(n12684), .ZN(n10723) );
  NAND2_X1 U13276 ( .A1(n9845), .A2(n13201), .ZN(n10717) );
  XNOR2_X1 U13277 ( .A(n10723), .B(n10717), .ZN(n10675) );
  NAND2_X1 U13278 ( .A1(n12862), .A2(n10667), .ZN(n10669) );
  OAI211_X1 U13279 ( .C1(n12860), .C2(n10670), .A(n10669), .B(n10668), .ZN(
        n10678) );
  INV_X1 U13280 ( .A(n10671), .ZN(n10710) );
  NOR3_X1 U13281 ( .A1(n10673), .A2(n10672), .A3(n12852), .ZN(n10674) );
  AOI21_X1 U13282 ( .B1(n10710), .B2(n12846), .A(n10674), .ZN(n10676) );
  NOR2_X1 U13283 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  AOI211_X1 U13284 ( .C1(n12941), .C2(n12831), .A(n10678), .B(n10677), .ZN(
        n10679) );
  OAI21_X1 U13285 ( .B1(n10722), .B2(n12854), .A(n10679), .ZN(P2_U3208) );
  OAI222_X1 U13286 ( .A1(P3_U3151), .A2(n10682), .B1(n12627), .B2(n10681), 
        .C1(n10680), .C2(n12623), .ZN(P3_U3270) );
  OAI21_X1 U13287 ( .B1(n10684), .B2(n15379), .A(n10683), .ZN(n10686) );
  AOI211_X1 U13288 ( .C1(n10687), .C2(n13571), .A(n10686), .B(n10685), .ZN(
        n10690) );
  NAND2_X1 U13289 ( .A1(n15441), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10688) );
  OAI21_X1 U13290 ( .B1(n10690), .B2(n15441), .A(n10688), .ZN(P2_U3510) );
  NAND2_X1 U13291 ( .A1(n15429), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10689) );
  OAI21_X1 U13292 ( .B1(n10690), .B2(n15429), .A(n10689), .ZN(P2_U3463) );
  AOI22_X1 U13293 ( .A1(n15089), .A2(n11783), .B1(n10307), .B2(n14330), .ZN(
        n10691) );
  XNOR2_X1 U13294 ( .A(n10691), .B(n11795), .ZN(n10876) );
  AOI22_X1 U13295 ( .A1(n15089), .A2(n10307), .B1(n11787), .B2(n14330), .ZN(
        n10877) );
  XNOR2_X1 U13296 ( .A(n10876), .B(n10877), .ZN(n10698) );
  INV_X1 U13297 ( .A(n10693), .ZN(n10694) );
  AOI21_X1 U13298 ( .B1(n10698), .B2(n10697), .A(n6705), .ZN(n10705) );
  NAND2_X1 U13299 ( .A1(n14331), .A2(n14554), .ZN(n10700) );
  NAND2_X1 U13300 ( .A1(n14329), .A2(n15059), .ZN(n10699) );
  NAND2_X1 U13301 ( .A1(n10700), .A2(n10699), .ZN(n15086) );
  AOI21_X1 U13302 ( .B1(n11282), .B2(n15086), .A(n10701), .ZN(n10702) );
  OAI21_X1 U13303 ( .B1(n14026), .B2(n15090), .A(n10702), .ZN(n10703) );
  AOI21_X1 U13304 ( .B1(n15089), .B2(n9398), .A(n10703), .ZN(n10704) );
  OAI21_X1 U13305 ( .B1(n10705), .B2(n14074), .A(n10704), .ZN(P1_U3221) );
  NAND2_X1 U13306 ( .A1(n12862), .A2(n10706), .ZN(n10708) );
  OAI211_X1 U13307 ( .C1(n12860), .C2(n10709), .A(n10708), .B(n10707), .ZN(
        n10714) );
  AOI211_X1 U13308 ( .C1(n10712), .C2(n10711), .A(n12854), .B(n10710), .ZN(
        n10713) );
  AOI211_X1 U13309 ( .C1(n15420), .C2(n12831), .A(n10714), .B(n10713), .ZN(
        n10715) );
  INV_X1 U13310 ( .A(n10715), .ZN(P2_U3189) );
  INV_X1 U13311 ( .A(n11407), .ZN(n10740) );
  OAI222_X1 U13312 ( .A1(n14755), .A2(n10716), .B1(n14753), .B2(n10740), .C1(
        n15140), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U13313 ( .A(n10723), .ZN(n10718) );
  NAND2_X1 U13314 ( .A1(n10718), .A2(n10717), .ZN(n10719) );
  XNOR2_X1 U13315 ( .A(n13855), .B(n12684), .ZN(n11189) );
  NAND2_X1 U13316 ( .A1(n9845), .A2(n13200), .ZN(n11190) );
  XNOR2_X1 U13317 ( .A(n11189), .B(n11190), .ZN(n10724) );
  AOI22_X1 U13318 ( .A1(n12838), .A2(n13854), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10720) );
  OAI21_X1 U13319 ( .B1(n10721), .B2(n12825), .A(n10720), .ZN(n10728) );
  INV_X1 U13320 ( .A(n10722), .ZN(n10726) );
  AOI22_X1 U13321 ( .A1(n10723), .A2(n12846), .B1(n12818), .B2(n13201), .ZN(
        n10725) );
  NOR3_X1 U13322 ( .A1(n10726), .A2(n10725), .A3(n10724), .ZN(n10727) );
  AOI211_X1 U13323 ( .C1(n13855), .C2(n12831), .A(n10728), .B(n10727), .ZN(
        n10729) );
  OAI21_X1 U13324 ( .B1(n11193), .B2(n12854), .A(n10729), .ZN(P2_U3196) );
  INV_X1 U13325 ( .A(n10753), .ZN(n10739) );
  XNOR2_X1 U13326 ( .A(n10754), .B(n11807), .ZN(n10843) );
  XNOR2_X1 U13327 ( .A(n12178), .B(n10843), .ZN(n10732) );
  INV_X1 U13328 ( .A(n10730), .ZN(n10731) );
  NAND2_X1 U13329 ( .A1(n10731), .A2(n10734), .ZN(n10846) );
  AOI21_X1 U13330 ( .B1(n10849), .B2(n10846), .A(n10732), .ZN(n10733) );
  OR3_X1 U13331 ( .A1(n10793), .A2(n10733), .A3(n11940), .ZN(n10738) );
  OAI22_X1 U13332 ( .A1(n11895), .A2(n10734), .B1(n11074), .B2(n11933), .ZN(
        n10735) );
  OAI211_X1 U13333 ( .C1(n10739), .C2(n10872), .A(n10738), .B(n10737), .ZN(
        P3_U3179) );
  OAI222_X1 U13334 ( .A1(n13905), .A2(n11408), .B1(P2_U3088), .B2(n13155), 
        .C1(n13908), .C2(n10740), .ZN(P2_U3306) );
  INV_X1 U13335 ( .A(n10743), .ZN(n11968) );
  XNOR2_X1 U13336 ( .A(n10741), .B(n11968), .ZN(n15492) );
  INV_X1 U13337 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10752) );
  NOR2_X1 U13338 ( .A1(n10745), .A2(n10742), .ZN(n10784) );
  INV_X1 U13339 ( .A(n10784), .ZN(n10747) );
  OAI21_X1 U13340 ( .B1(n10745), .B2(n10744), .A(n10743), .ZN(n10746) );
  NAND3_X1 U13341 ( .A1(n10747), .A2(n12474), .A3(n10746), .ZN(n10750) );
  AOI22_X1 U13342 ( .A1(n10748), .A2(n12480), .B1(n12479), .B2(n12177), .ZN(
        n10749) );
  OAI211_X1 U13343 ( .C1(n11601), .C2(n15492), .A(n10750), .B(n10749), .ZN(
        n15494) );
  INV_X1 U13344 ( .A(n15494), .ZN(n10751) );
  MUX2_X1 U13345 ( .A(n10752), .B(n10751), .S(n12490), .Z(n10756) );
  AOI22_X1 U13346 ( .A1(n12438), .A2(n10754), .B1(n12485), .B2(n10753), .ZN(
        n10755) );
  OAI211_X1 U13347 ( .C1(n15492), .C2(n12299), .A(n10756), .B(n10755), .ZN(
        P3_U3227) );
  XNOR2_X1 U13348 ( .A(n10757), .B(n6869), .ZN(n14887) );
  OAI211_X1 U13349 ( .C1(n10759), .C2(n6869), .A(n10758), .B(n15139), .ZN(
        n10761) );
  AOI22_X1 U13350 ( .A1(n15059), .A2(n14326), .B1(n15058), .B2(n14554), .ZN(
        n10760) );
  NAND2_X1 U13351 ( .A1(n10761), .A2(n10760), .ZN(n14883) );
  AOI21_X1 U13352 ( .B1(n14937), .B2(n14885), .A(n14589), .ZN(n10762) );
  AND2_X1 U13353 ( .A1(n10762), .A2(n11030), .ZN(n14884) );
  NAND2_X1 U13354 ( .A1(n14884), .A2(n15101), .ZN(n10766) );
  OAI22_X1 U13355 ( .A1(n15104), .A2(n10763), .B1(n11299), .B2(n15091), .ZN(
        n10764) );
  AOI21_X1 U13356 ( .B1(n14885), .B2(n15075), .A(n10764), .ZN(n10765) );
  NAND2_X1 U13357 ( .A1(n10766), .A2(n10765), .ZN(n10767) );
  AOI21_X1 U13358 ( .B1(n14883), .B2(n15104), .A(n10767), .ZN(n10768) );
  OAI21_X1 U13359 ( .B1(n14623), .B2(n14887), .A(n10768), .ZN(P1_U3281) );
  XNOR2_X1 U13360 ( .A(n10769), .B(n12038), .ZN(n15510) );
  INV_X1 U13361 ( .A(n10770), .ZN(n10772) );
  INV_X1 U13362 ( .A(n12038), .ZN(n10771) );
  AOI21_X1 U13363 ( .B1(n10985), .B2(n10772), .A(n10771), .ZN(n10773) );
  OR3_X1 U13364 ( .A1(n10774), .A2(n12404), .A3(n10773), .ZN(n10776) );
  AOI22_X1 U13365 ( .A1(n12174), .A2(n12479), .B1(n12480), .B2(n12176), .ZN(
        n10775) );
  NAND2_X1 U13366 ( .A1(n10776), .A2(n10775), .ZN(n10777) );
  AOI21_X1 U13367 ( .B1(n15510), .B2(n10988), .A(n10777), .ZN(n15512) );
  AOI22_X1 U13368 ( .A1(n12438), .A2(n15507), .B1(n12485), .B2(n10892), .ZN(
        n10778) );
  OAI21_X1 U13369 ( .B1(n15446), .B2(n12490), .A(n10778), .ZN(n10779) );
  AOI21_X1 U13370 ( .B1(n15510), .B2(n10780), .A(n10779), .ZN(n10781) );
  OAI21_X1 U13371 ( .B1(n15512), .B2(n12486), .A(n10781), .ZN(P3_U3224) );
  XOR2_X1 U13372 ( .A(n10782), .B(n12027), .Z(n15498) );
  NOR2_X1 U13373 ( .A1(n10784), .A2(n10783), .ZN(n10785) );
  XOR2_X1 U13374 ( .A(n12027), .B(n10785), .Z(n10787) );
  OAI22_X1 U13375 ( .A1(n10890), .A2(n12408), .B1(n10844), .B2(n12406), .ZN(
        n10786) );
  AOI21_X1 U13376 ( .B1(n10787), .B2(n12474), .A(n10786), .ZN(n10788) );
  OAI21_X1 U13377 ( .B1(n11601), .B2(n15498), .A(n10788), .ZN(n15500) );
  NAND2_X1 U13378 ( .A1(n15500), .A2(n12490), .ZN(n10792) );
  INV_X1 U13379 ( .A(n10796), .ZN(n15496) );
  INV_X1 U13380 ( .A(n10797), .ZN(n10789) );
  OAI22_X1 U13381 ( .A1(n12488), .A2(n15496), .B1(n10789), .B2(n12387), .ZN(
        n10790) );
  AOI21_X1 U13382 ( .B1(n12486), .B2(P3_REG2_REG_7__SCAN_IN), .A(n10790), .ZN(
        n10791) );
  OAI211_X1 U13383 ( .C1(n15498), .C2(n12299), .A(n10792), .B(n10791), .ZN(
        P3_U3226) );
  NOR2_X1 U13384 ( .A1(n10844), .A2(n10843), .ZN(n10851) );
  NOR2_X1 U13385 ( .A1(n10793), .A2(n10851), .ZN(n11070) );
  XNOR2_X1 U13386 ( .A(n12027), .B(n11655), .ZN(n10850) );
  XNOR2_X1 U13387 ( .A(n11070), .B(n10850), .ZN(n10800) );
  OAI22_X1 U13388 ( .A1(n11895), .A2(n10844), .B1(n10890), .B2(n11933), .ZN(
        n10794) );
  AOI211_X1 U13389 ( .C1(n10796), .C2(n11904), .A(n10795), .B(n10794), .ZN(
        n10799) );
  NAND2_X1 U13390 ( .A1(n11938), .A2(n10797), .ZN(n10798) );
  OAI211_X1 U13391 ( .C1(n10800), .C2(n11940), .A(n10799), .B(n10798), .ZN(
        P3_U3153) );
  INV_X1 U13392 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n13794) );
  AOI21_X1 U13393 ( .B1(n13794), .B2(n10803), .A(n10923), .ZN(n10817) );
  OAI21_X1 U13394 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n10806), .A(n10930), 
        .ZN(n10809) );
  AND2_X1 U13395 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11132) );
  AOI21_X1 U13396 ( .B1(n15458), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11132), 
        .ZN(n10807) );
  OAI21_X1 U13397 ( .B1(n15452), .B2(n10929), .A(n10807), .ZN(n10808) );
  AOI21_X1 U13398 ( .B1(n10809), .B2(n15461), .A(n10808), .ZN(n10816) );
  NAND2_X1 U13399 ( .A1(n10811), .A2(n10810), .ZN(n10813) );
  MUX2_X1 U13400 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12275), .Z(n10935) );
  XNOR2_X1 U13401 ( .A(n10935), .B(n10936), .ZN(n10812) );
  NAND2_X1 U13402 ( .A1(n10813), .A2(n10812), .ZN(n10941) );
  OAI21_X1 U13403 ( .B1(n10813), .B2(n10812), .A(n10941), .ZN(n10814) );
  NAND2_X1 U13404 ( .A1(n10814), .A2(n12280), .ZN(n10815) );
  OAI211_X1 U13405 ( .C1(n10817), .C2(n15465), .A(n10816), .B(n10815), .ZN(
        P3_U3193) );
  NAND2_X1 U13406 ( .A1(n10818), .A2(n13068), .ZN(n10820) );
  AOI22_X1 U13407 ( .A1(n11382), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11381), 
        .B2(n15257), .ZN(n10819) );
  XNOR2_X1 U13408 ( .A(n13582), .B(n13199), .ZN(n13136) );
  INV_X1 U13409 ( .A(n13200), .ZN(n12949) );
  OR2_X1 U13410 ( .A1(n13855), .A2(n12949), .ZN(n10822) );
  XOR2_X1 U13411 ( .A(n13136), .B(n10904), .Z(n10833) );
  NAND2_X1 U13412 ( .A1(n6551), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10830) );
  NAND2_X1 U13413 ( .A1(n7659), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10829) );
  INV_X1 U13414 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10824) );
  NAND2_X1 U13415 ( .A1(n10825), .A2(n10824), .ZN(n10826) );
  AND2_X1 U13416 ( .A1(n10906), .A2(n10826), .ZN(n10902) );
  NAND2_X1 U13417 ( .A1(n11502), .A2(n10902), .ZN(n10828) );
  NAND2_X1 U13418 ( .A1(n13072), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10827) );
  NAND4_X1 U13419 ( .A1(n10830), .A2(n10829), .A3(n10828), .A4(n10827), .ZN(
        n13198) );
  NAND2_X1 U13420 ( .A1(n12848), .A2(n13198), .ZN(n10832) );
  NAND2_X1 U13421 ( .A1(n13167), .A2(n13200), .ZN(n10831) );
  NAND2_X1 U13422 ( .A1(n10832), .A2(n10831), .ZN(n11182) );
  AOI21_X1 U13423 ( .B1(n10833), .B2(n15409), .A(n11182), .ZN(n13584) );
  AOI211_X1 U13424 ( .C1(n13582), .C2(n10834), .A(n13562), .B(n7228), .ZN(
        n13581) );
  INV_X1 U13425 ( .A(n13582), .ZN(n10836) );
  AOI22_X1 U13426 ( .A1(n15320), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11181), 
        .B2(n15318), .ZN(n10835) );
  OAI21_X1 U13427 ( .B1(n10836), .B2(n13420), .A(n10835), .ZN(n10840) );
  AND2_X1 U13428 ( .A1(n13855), .A2(n13200), .ZN(n10837) );
  XNOR2_X1 U13429 ( .A(n10896), .B(n13136), .ZN(n13585) );
  NOR2_X1 U13430 ( .A1(n13585), .A2(n13465), .ZN(n10839) );
  AOI211_X1 U13431 ( .C1(n13581), .C2(n13467), .A(n10840), .B(n10839), .ZN(
        n10841) );
  OAI21_X1 U13432 ( .B1(n15320), .B2(n13584), .A(n10841), .ZN(P2_U3252) );
  INV_X1 U13433 ( .A(n10842), .ZN(n11019) );
  XNOR2_X1 U13434 ( .A(n12034), .B(n11807), .ZN(n10854) );
  XNOR2_X1 U13435 ( .A(n10854), .B(n12176), .ZN(n10852) );
  NAND2_X1 U13436 ( .A1(n10844), .A2(n10843), .ZN(n10845) );
  NAND3_X1 U13437 ( .A1(n10852), .A2(n10846), .A3(n10845), .ZN(n10847) );
  NOR2_X1 U13438 ( .A1(n10850), .A2(n10847), .ZN(n10848) );
  INV_X1 U13439 ( .A(n10852), .ZN(n11071) );
  OAI21_X1 U13440 ( .B1(n11074), .B2(n11071), .A(n10850), .ZN(n10857) );
  INV_X1 U13441 ( .A(n10850), .ZN(n11069) );
  NAND2_X1 U13442 ( .A1(n10852), .A2(n10851), .ZN(n10853) );
  NAND2_X1 U13443 ( .A1(n11069), .A2(n10853), .ZN(n10856) );
  INV_X1 U13444 ( .A(n10854), .ZN(n10855) );
  AOI22_X1 U13445 ( .A1(n10857), .A2(n10856), .B1(n12176), .B2(n10855), .ZN(
        n10858) );
  XNOR2_X1 U13446 ( .A(n10860), .B(n11807), .ZN(n10861) );
  XNOR2_X1 U13447 ( .A(n10861), .B(n12175), .ZN(n11087) );
  OR2_X1 U13448 ( .A1(n11088), .A2(n11087), .ZN(n10888) );
  INV_X1 U13449 ( .A(n12175), .ZN(n11073) );
  INV_X1 U13450 ( .A(n10861), .ZN(n10862) );
  NAND2_X1 U13451 ( .A1(n11073), .A2(n10862), .ZN(n10863) );
  AND2_X1 U13452 ( .A1(n10888), .A2(n10863), .ZN(n10866) );
  XNOR2_X1 U13453 ( .A(n10869), .B(n11655), .ZN(n11084) );
  XNOR2_X1 U13454 ( .A(n11084), .B(n11086), .ZN(n10865) );
  AND2_X1 U13455 ( .A1(n10863), .A2(n10865), .ZN(n11089) );
  NAND2_X1 U13456 ( .A1(n10888), .A2(n11089), .ZN(n10864) );
  OAI211_X1 U13457 ( .C1(n10866), .C2(n10865), .A(n10864), .B(n11920), .ZN(
        n10871) );
  OAI22_X1 U13458 ( .A1(n11895), .A2(n11073), .B1(n11149), .B2(n11933), .ZN(
        n10867) );
  AOI211_X1 U13459 ( .C1(n10869), .C2(n11904), .A(n10868), .B(n10867), .ZN(
        n10870) );
  OAI211_X1 U13460 ( .C1(n11019), .C2(n10872), .A(n10871), .B(n10870), .ZN(
        P3_U3157) );
  OAI222_X1 U13461 ( .A1(P3_U3151), .A2(n10875), .B1(n12623), .B2(n10874), 
        .C1(n12627), .C2(n10873), .ZN(P3_U3269) );
  AOI22_X1 U13462 ( .A1(n15076), .A2(n11783), .B1(n10307), .B2(n14329), .ZN(
        n10878) );
  XOR2_X1 U13463 ( .A(n11795), .B(n10878), .Z(n11116) );
  INV_X1 U13464 ( .A(n15076), .ZN(n15181) );
  OAI22_X1 U13465 ( .A1(n15181), .A2(n11798), .B1(n10879), .B2(n11797), .ZN(
        n11117) );
  INV_X1 U13466 ( .A(n11117), .ZN(n11119) );
  XNOR2_X1 U13467 ( .A(n11116), .B(n11119), .ZN(n10880) );
  XNOR2_X1 U13468 ( .A(n11118), .B(n10880), .ZN(n10887) );
  NAND2_X1 U13469 ( .A1(n14330), .A2(n14554), .ZN(n10882) );
  NAND2_X1 U13470 ( .A1(n14328), .A2(n15059), .ZN(n10881) );
  NAND2_X1 U13471 ( .A1(n10882), .A2(n10881), .ZN(n15070) );
  NAND2_X1 U13472 ( .A1(n11282), .A2(n15070), .ZN(n10883) );
  OAI211_X1 U13473 ( .C1(n14026), .C2(n15072), .A(n10884), .B(n10883), .ZN(
        n10885) );
  AOI21_X1 U13474 ( .B1(n15076), .B2(n9398), .A(n10885), .ZN(n10886) );
  OAI21_X1 U13475 ( .B1(n10887), .B2(n14074), .A(n10886), .ZN(P1_U3231) );
  INV_X1 U13476 ( .A(n10888), .ZN(n10889) );
  AOI21_X1 U13477 ( .B1(n11087), .B2(n11088), .A(n10889), .ZN(n10895) );
  NOR2_X1 U13478 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8423), .ZN(n15457) );
  OAI22_X1 U13479 ( .A1(n11895), .A2(n10890), .B1(n11086), .B2(n11933), .ZN(
        n10891) );
  AOI211_X1 U13480 ( .C1(n15507), .C2(n11904), .A(n15457), .B(n10891), .ZN(
        n10894) );
  NAND2_X1 U13481 ( .A1(n11938), .A2(n10892), .ZN(n10893) );
  OAI211_X1 U13482 ( .C1(n10895), .C2(n11940), .A(n10894), .B(n10893), .ZN(
        P3_U3171) );
  NAND2_X1 U13483 ( .A1(n13582), .A2(n13199), .ZN(n10897) );
  NAND2_X1 U13484 ( .A1(n10899), .A2(n13068), .ZN(n10901) );
  AOI22_X1 U13485 ( .A1(n11382), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n11381), 
        .B2(n11053), .ZN(n10900) );
  INV_X1 U13486 ( .A(n13198), .ZN(n12962) );
  XNOR2_X1 U13487 ( .A(n13577), .B(n12962), .ZN(n13140) );
  XNOR2_X1 U13488 ( .A(n11005), .B(n13140), .ZN(n13580) );
  INV_X1 U13489 ( .A(n10902), .ZN(n12699) );
  INV_X1 U13490 ( .A(n13199), .ZN(n12694) );
  NOR2_X1 U13491 ( .A1(n13582), .A2(n12694), .ZN(n10903) );
  INV_X1 U13492 ( .A(n13140), .ZN(n11004) );
  XNOR2_X1 U13493 ( .A(n10998), .B(n11004), .ZN(n10914) );
  INV_X1 U13494 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12859) );
  NAND2_X1 U13495 ( .A1(n10906), .A2(n12859), .ZN(n10907) );
  NAND2_X1 U13496 ( .A1(n11363), .A2(n10907), .ZN(n12858) );
  OR2_X1 U13497 ( .A1(n11492), .A2(n12858), .ZN(n10911) );
  NAND2_X1 U13498 ( .A1(n9306), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n10910) );
  NAND2_X1 U13499 ( .A1(n13072), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n10909) );
  NAND2_X1 U13500 ( .A1(n6551), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n10908) );
  NAND4_X1 U13501 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n13197) );
  NAND2_X1 U13502 ( .A1(n12848), .A2(n13197), .ZN(n10913) );
  NAND2_X1 U13503 ( .A1(n13167), .A2(n13199), .ZN(n10912) );
  NAND2_X1 U13504 ( .A1(n10913), .A2(n10912), .ZN(n12697) );
  AOI21_X1 U13505 ( .B1(n10914), .B2(n15409), .A(n12697), .ZN(n13579) );
  OAI21_X1 U13506 ( .B1(n12699), .B2(n13397), .A(n13579), .ZN(n10915) );
  NAND2_X1 U13507 ( .A1(n10915), .A2(n13472), .ZN(n10921) );
  INV_X1 U13508 ( .A(n11007), .ZN(n10916) );
  AOI211_X1 U13509 ( .C1(n13577), .C2(n10917), .A(n13562), .B(n10916), .ZN(
        n13576) );
  INV_X1 U13510 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10918) );
  OAI22_X1 U13511 ( .A1(n7227), .A2(n13420), .B1(n13472), .B2(n10918), .ZN(
        n10919) );
  AOI21_X1 U13512 ( .B1(n13576), .B2(n13467), .A(n10919), .ZN(n10920) );
  OAI211_X1 U13513 ( .C1(n13580), .C2(n13465), .A(n10921), .B(n10920), .ZN(
        P2_U3251) );
  NOR2_X1 U13514 ( .A1(n10936), .A2(n10922), .ZN(n10924) );
  INV_X1 U13515 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n10925) );
  MUX2_X1 U13516 ( .A(n10925), .B(P3_REG2_REG_12__SCAN_IN), .S(n11230), .Z(
        n10926) );
  AOI21_X1 U13517 ( .B1(n10927), .B2(n10926), .A(n6694), .ZN(n10946) );
  NAND2_X1 U13518 ( .A1(n10929), .A2(n10928), .ZN(n10931) );
  NAND2_X1 U13519 ( .A1(n10931), .A2(n10930), .ZN(n11219) );
  INV_X1 U13520 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12554) );
  XNOR2_X1 U13521 ( .A(n11230), .B(n12554), .ZN(n11218) );
  XNOR2_X1 U13522 ( .A(n11219), .B(n11218), .ZN(n10934) );
  INV_X1 U13523 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14834) );
  INV_X1 U13524 ( .A(n15458), .ZN(n14910) );
  INV_X1 U13525 ( .A(n11230), .ZN(n10938) );
  NAND2_X1 U13526 ( .A1(n14907), .A2(n10938), .ZN(n10932) );
  NAND2_X1 U13527 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11148)
         );
  OAI211_X1 U13528 ( .C1(n14834), .C2(n14910), .A(n10932), .B(n11148), .ZN(
        n10933) );
  AOI21_X1 U13529 ( .B1(n10934), .B2(n15461), .A(n10933), .ZN(n10945) );
  INV_X1 U13530 ( .A(n10935), .ZN(n10937) );
  NAND2_X1 U13531 ( .A1(n10937), .A2(n10936), .ZN(n10939) );
  AND2_X1 U13532 ( .A1(n10941), .A2(n10939), .ZN(n10943) );
  MUX2_X1 U13533 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12275), .Z(n11231) );
  XNOR2_X1 U13534 ( .A(n11231), .B(n10938), .ZN(n10942) );
  AND2_X1 U13535 ( .A1(n10942), .A2(n10939), .ZN(n10940) );
  NAND2_X1 U13536 ( .A1(n10941), .A2(n10940), .ZN(n11233) );
  OAI211_X1 U13537 ( .C1(n10943), .C2(n10942), .A(n12280), .B(n11233), .ZN(
        n10944) );
  OAI211_X1 U13538 ( .C1(n10946), .C2(n15465), .A(n10945), .B(n10944), .ZN(
        P3_U3194) );
  NAND2_X1 U13539 ( .A1(n10948), .A2(n10947), .ZN(n10950) );
  NAND2_X1 U13540 ( .A1(n10957), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n10949) );
  NAND2_X1 U13541 ( .A1(n10950), .A2(n10949), .ZN(n10951) );
  NAND2_X1 U13542 ( .A1(n10951), .A2(n15037), .ZN(n10952) );
  XNOR2_X1 U13543 ( .A(n10951), .B(n10960), .ZN(n15036) );
  NAND2_X1 U13544 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n15036), .ZN(n15034) );
  NAND2_X1 U13545 ( .A1(n10952), .A2(n15034), .ZN(n10953) );
  XNOR2_X1 U13546 ( .A(n10954), .B(n10953), .ZN(n10967) );
  INV_X1 U13547 ( .A(n10967), .ZN(n10965) );
  NAND2_X1 U13548 ( .A1(n10956), .A2(n10955), .ZN(n10959) );
  NAND2_X1 U13549 ( .A1(n10957), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10958) );
  NAND2_X1 U13550 ( .A1(n10959), .A2(n10958), .ZN(n10961) );
  XNOR2_X1 U13551 ( .A(n10961), .B(n10960), .ZN(n15041) );
  NAND2_X1 U13552 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15041), .ZN(n15039) );
  NAND2_X1 U13553 ( .A1(n10961), .A2(n15037), .ZN(n10962) );
  NAND2_X1 U13554 ( .A1(n15039), .A2(n10962), .ZN(n10963) );
  XOR2_X1 U13555 ( .A(n10963), .B(P1_REG2_REG_19__SCAN_IN), .Z(n10966) );
  OAI21_X1 U13556 ( .B1(n10966), .B2(n15025), .A(n15029), .ZN(n10964) );
  AOI21_X1 U13557 ( .B1(n10965), .B2(n15035), .A(n10964), .ZN(n10969) );
  AOI22_X1 U13558 ( .A1(n10967), .A2(n15035), .B1(n15040), .B2(n10966), .ZN(
        n10968) );
  MUX2_X1 U13559 ( .A(n10969), .B(n10968), .S(n14617), .Z(n10970) );
  NAND2_X1 U13560 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13953)
         );
  OAI211_X1 U13561 ( .C1(n10971), .C2(n15047), .A(n10970), .B(n13953), .ZN(
        P1_U3262) );
  XNOR2_X1 U13562 ( .A(n10972), .B(n14289), .ZN(n14957) );
  INV_X1 U13563 ( .A(n14957), .ZN(n10983) );
  OR2_X1 U13564 ( .A1(n11690), .A2(n14608), .ZN(n10974) );
  NAND2_X1 U13565 ( .A1(n14326), .A2(n14554), .ZN(n10973) );
  NAND2_X1 U13566 ( .A1(n10974), .A2(n10973), .ZN(n14951) );
  AOI22_X1 U13567 ( .A1(n15104), .A2(n14951), .B1(n13922), .B2(n15073), .ZN(
        n10975) );
  OAI21_X1 U13568 ( .B1(n9564), .B2(n15104), .A(n10975), .ZN(n10978) );
  OAI211_X1 U13569 ( .C1(n11029), .C2(n10976), .A(n8988), .B(n11202), .ZN(
        n14953) );
  NOR2_X1 U13570 ( .A1(n14953), .A2(n14583), .ZN(n10977) );
  AOI211_X1 U13571 ( .C1(n15075), .C2(n14952), .A(n10978), .B(n10977), .ZN(
        n10982) );
  NAND2_X1 U13572 ( .A1(n10980), .A2(n10979), .ZN(n14949) );
  NAND3_X1 U13573 ( .A1(n14950), .A2(n14949), .A3(n15102), .ZN(n10981) );
  OAI211_X1 U13574 ( .C1(n10983), .C2(n14532), .A(n10982), .B(n10981), .ZN(
        P1_U3279) );
  XNOR2_X1 U13575 ( .A(n10984), .B(n12032), .ZN(n15505) );
  INV_X1 U13576 ( .A(n15505), .ZN(n10996) );
  INV_X1 U13577 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10993) );
  INV_X1 U13578 ( .A(n10985), .ZN(n10986) );
  AOI21_X1 U13579 ( .B1(n12032), .B2(n10987), .A(n10986), .ZN(n10991) );
  AOI22_X1 U13580 ( .A1(n12480), .A2(n12177), .B1(n12175), .B2(n12479), .ZN(
        n10990) );
  NAND2_X1 U13581 ( .A1(n15505), .A2(n10988), .ZN(n10989) );
  OAI211_X1 U13582 ( .C1(n10991), .C2(n12404), .A(n10990), .B(n10989), .ZN(
        n15503) );
  INV_X1 U13583 ( .A(n15503), .ZN(n10992) );
  MUX2_X1 U13584 ( .A(n10993), .B(n10992), .S(n12490), .Z(n10995) );
  AOI22_X1 U13585 ( .A1(n12438), .A2(n12034), .B1(n12485), .B2(n11077), .ZN(
        n10994) );
  OAI211_X1 U13586 ( .C1(n10996), .C2(n12299), .A(n10995), .B(n10994), .ZN(
        P3_U3225) );
  OR2_X1 U13587 ( .A1(n13577), .A2(n12962), .ZN(n10997) );
  NAND2_X1 U13588 ( .A1(n13577), .A2(n12962), .ZN(n10999) );
  NAND2_X1 U13589 ( .A1(n11000), .A2(n10999), .ZN(n11353) );
  NAND2_X1 U13590 ( .A1(n11001), .A2(n13068), .ZN(n11003) );
  AOI22_X1 U13591 ( .A1(n11382), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n11381), 
        .B2(n15274), .ZN(n11002) );
  INV_X1 U13592 ( .A(n13197), .ZN(n12853) );
  XNOR2_X1 U13593 ( .A(n12973), .B(n12853), .ZN(n13141) );
  XNOR2_X1 U13594 ( .A(n11353), .B(n13141), .ZN(n13574) );
  INV_X1 U13595 ( .A(n13406), .ZN(n13443) );
  OAI21_X1 U13596 ( .B1(n11006), .B2(n13141), .A(n11522), .ZN(n13572) );
  INV_X1 U13597 ( .A(n13465), .ZN(n13469) );
  INV_X1 U13598 ( .A(n12973), .ZN(n13568) );
  AOI211_X1 U13599 ( .C1(n12973), .C2(n11007), .A(n13562), .B(n13455), .ZN(
        n13570) );
  NAND2_X1 U13600 ( .A1(n13570), .A2(n13467), .ZN(n11014) );
  INV_X1 U13601 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11035) );
  NAND2_X1 U13602 ( .A1(n6551), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U13603 ( .A1(n9306), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n11008) );
  AND2_X1 U13604 ( .A1(n11009), .A2(n11008), .ZN(n11011) );
  XNOR2_X1 U13605 ( .A(n11363), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n13458) );
  NAND2_X1 U13606 ( .A1(n13458), .A2(n11502), .ZN(n11010) );
  OAI211_X1 U13607 ( .C1(n11513), .C2(n11035), .A(n11011), .B(n11010), .ZN(
        n13196) );
  AOI22_X1 U13608 ( .A1(n13196), .A2(n12848), .B1(n13167), .B2(n13198), .ZN(
        n13567) );
  OAI22_X1 U13609 ( .A1(n15320), .A2(n13567), .B1(n12858), .B2(n13397), .ZN(
        n11012) );
  AOI21_X1 U13610 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n15320), .A(n11012), 
        .ZN(n11013) );
  OAI211_X1 U13611 ( .C1(n13568), .C2(n13420), .A(n11014), .B(n11013), .ZN(
        n11015) );
  AOI21_X1 U13612 ( .B1(n13572), .B2(n13469), .A(n11015), .ZN(n11016) );
  OAI21_X1 U13613 ( .B1(n13574), .B2(n13443), .A(n11016), .ZN(P2_U3250) );
  XNOR2_X1 U13614 ( .A(n11017), .B(n7346), .ZN(n11018) );
  AOI222_X1 U13615 ( .A1(n12474), .A2(n11018), .B1(n12173), .B2(n12479), .C1(
        n12175), .C2(n12480), .ZN(n15513) );
  OAI22_X1 U13616 ( .A1(n12488), .A2(n15514), .B1(n11019), .B2(n12387), .ZN(
        n11020) );
  AOI21_X1 U13617 ( .B1(n12486), .B2(P3_REG2_REG_10__SCAN_IN), .A(n11020), 
        .ZN(n11023) );
  XNOR2_X1 U13618 ( .A(n11021), .B(n7346), .ZN(n15517) );
  NAND2_X1 U13619 ( .A1(n15517), .A2(n12457), .ZN(n11022) );
  OAI211_X1 U13620 ( .C1(n15513), .C2(n12486), .A(n11023), .B(n11022), .ZN(
        P3_U3223) );
  XNOR2_X1 U13621 ( .A(n11024), .B(n11026), .ZN(n14965) );
  OAI211_X1 U13622 ( .C1(n11027), .C2(n11026), .A(n15139), .B(n11025), .ZN(
        n14962) );
  AOI22_X1 U13623 ( .A1(n14325), .A2(n15059), .B1(n14554), .B2(n14327), .ZN(
        n14958) );
  OAI211_X1 U13624 ( .C1(n15091), .C2(n11314), .A(n14962), .B(n14958), .ZN(
        n11028) );
  NAND2_X1 U13625 ( .A1(n11028), .A2(n15104), .ZN(n11034) );
  AOI211_X1 U13626 ( .C1(n14961), .C2(n11030), .A(n14589), .B(n11029), .ZN(
        n14959) );
  INV_X1 U13627 ( .A(n14961), .ZN(n11031) );
  OAI22_X1 U13628 ( .A1(n11031), .A2(n14541), .B1(n9562), .B2(n15104), .ZN(
        n11032) );
  AOI21_X1 U13629 ( .B1(n14959), .B2(n15101), .A(n11032), .ZN(n11033) );
  OAI211_X1 U13630 ( .C1(n14965), .C2(n14623), .A(n11034), .B(n11033), .ZN(
        P1_U3280) );
  INV_X1 U13631 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11043) );
  MUX2_X1 U13632 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n11043), .S(n15300), .Z(
        n15297) );
  MUX2_X1 U13633 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n11035), .S(n15283), .Z(
        n15285) );
  INV_X1 U13634 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13732) );
  AOI21_X1 U13635 ( .B1(n11046), .B2(n11037), .A(n11036), .ZN(n15253) );
  NOR2_X1 U13636 ( .A1(n15257), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11038) );
  AOI21_X1 U13637 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n15257), .A(n11038), 
        .ZN(n15252) );
  NAND2_X1 U13638 ( .A1(n15253), .A2(n15252), .ZN(n15251) );
  OAI21_X1 U13639 ( .B1(n13732), .B2(n11050), .A(n15251), .ZN(n11039) );
  NAND2_X1 U13640 ( .A1(n11053), .A2(n11039), .ZN(n11040) );
  AOI22_X1 U13641 ( .A1(n15275), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n15274), 
        .B2(n11041), .ZN(n11042) );
  OAI21_X1 U13642 ( .B1(n11060), .B2(n11043), .A(n15295), .ZN(n13230) );
  AOI21_X1 U13643 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11044), .A(n13232), 
        .ZN(n11068) );
  INV_X1 U13644 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n11373) );
  NOR2_X1 U13645 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11373), .ZN(n11065) );
  INV_X1 U13646 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11059) );
  XNOR2_X1 U13647 ( .A(n11060), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15304) );
  INV_X1 U13648 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11057) );
  XNOR2_X1 U13649 ( .A(n11058), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15289) );
  XNOR2_X1 U13650 ( .A(n15272), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15268) );
  INV_X1 U13651 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11051) );
  AOI22_X1 U13652 ( .A1(n11048), .A2(n11047), .B1(n11046), .B2(n11045), .ZN(
        n15256) );
  NOR2_X1 U13653 ( .A1(n11050), .A2(n11051), .ZN(n11049) );
  AOI21_X1 U13654 ( .B1(n11051), .B2(n11050), .A(n11049), .ZN(n15255) );
  NAND2_X1 U13655 ( .A1(n15256), .A2(n15255), .ZN(n15254) );
  OAI21_X1 U13656 ( .B1(n11051), .B2(n11050), .A(n15254), .ZN(n15269) );
  NAND2_X1 U13657 ( .A1(n15268), .A2(n15269), .ZN(n15267) );
  INV_X1 U13658 ( .A(n15267), .ZN(n11052) );
  AOI21_X1 U13659 ( .B1(n11053), .B2(P2_REG1_REG_14__SCAN_IN), .A(n11052), 
        .ZN(n11055) );
  XNOR2_X1 U13660 ( .A(n11055), .B(n11054), .ZN(n15277) );
  INV_X1 U13661 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11056) );
  OAI22_X1 U13662 ( .A1(n15277), .A2(n11056), .B1(n11055), .B2(n11054), .ZN(
        n15288) );
  NAND2_X1 U13663 ( .A1(n15289), .A2(n15288), .ZN(n15287) );
  OAI21_X1 U13664 ( .B1(n11058), .B2(n11057), .A(n15287), .ZN(n15303) );
  NAND2_X1 U13665 ( .A1(n15304), .A2(n15303), .ZN(n15301) );
  OAI21_X1 U13666 ( .B1(n11060), .B2(n11059), .A(n15301), .ZN(n13233) );
  XNOR2_X1 U13667 ( .A(n11061), .B(n13233), .ZN(n11062) );
  NAND2_X1 U13668 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11062), .ZN(n13235) );
  OAI211_X1 U13669 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n11062), .A(n15302), 
        .B(n13235), .ZN(n11063) );
  INV_X1 U13670 ( .A(n11063), .ZN(n11064) );
  AOI211_X1 U13671 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n15294), .A(n11065), 
        .B(n11064), .ZN(n11067) );
  NAND2_X1 U13672 ( .A1(n15299), .A2(n13234), .ZN(n11066) );
  OAI211_X1 U13673 ( .C1(n11068), .C2(n15242), .A(n11067), .B(n11066), .ZN(
        P2_U3232) );
  MUX2_X1 U13674 ( .A(n11074), .B(n11070), .S(n11069), .Z(n11072) );
  XNOR2_X1 U13675 ( .A(n11072), .B(n11071), .ZN(n11080) );
  OAI22_X1 U13676 ( .A1(n11895), .A2(n11074), .B1(n11073), .B2(n11933), .ZN(
        n11075) );
  AOI211_X1 U13677 ( .C1(n12034), .C2(n11904), .A(n11076), .B(n11075), .ZN(
        n11079) );
  NAND2_X1 U13678 ( .A1(n11938), .A2(n11077), .ZN(n11078) );
  OAI211_X1 U13679 ( .C1(n11080), .C2(n11940), .A(n11079), .B(n11078), .ZN(
        P3_U3161) );
  OAI222_X1 U13680 ( .A1(n12627), .A2(n11083), .B1(n12623), .B2(n11082), .C1(
        P3_U3151), .C2(n11081), .ZN(P3_U3267) );
  INV_X1 U13681 ( .A(n11084), .ZN(n11085) );
  NOR2_X1 U13682 ( .A1(n11086), .A2(n11085), .ZN(n11090) );
  OR2_X1 U13683 ( .A1(n11090), .A2(n11089), .ZN(n11091) );
  XNOR2_X1 U13684 ( .A(n11133), .B(n11807), .ZN(n11130) );
  XNOR2_X1 U13685 ( .A(n11171), .B(n11655), .ZN(n11093) );
  INV_X1 U13686 ( .A(n11130), .ZN(n11142) );
  AOI21_X1 U13687 ( .B1(n11142), .B2(n12173), .A(n12481), .ZN(n11094) );
  INV_X1 U13688 ( .A(n11093), .ZN(n11145) );
  NAND3_X1 U13689 ( .A1(n12481), .A2(n11142), .A3(n12173), .ZN(n11095) );
  XNOR2_X1 U13690 ( .A(n11105), .B(n11807), .ZN(n11100) );
  NOR2_X1 U13691 ( .A1(n11100), .A2(n11099), .ZN(n11623) );
  NOR2_X1 U13692 ( .A1(n11623), .A2(n6713), .ZN(n11101) );
  XNOR2_X1 U13693 ( .A(n11624), .B(n11101), .ZN(n11107) );
  NAND2_X1 U13694 ( .A1(n11938), .A2(n12484), .ZN(n11103) );
  AND2_X1 U13695 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n11255) );
  AOI21_X1 U13696 ( .B1(n12481), .B2(n11931), .A(n11255), .ZN(n11102) );
  OAI211_X1 U13697 ( .C1(n11625), .C2(n11933), .A(n11103), .B(n11102), .ZN(
        n11104) );
  AOI21_X1 U13698 ( .B1(n11105), .B2(n11904), .A(n11104), .ZN(n11106) );
  OAI21_X1 U13699 ( .B1(n11107), .B2(n11940), .A(n11106), .ZN(P3_U3174) );
  XNOR2_X1 U13700 ( .A(n11108), .B(n12050), .ZN(n11109) );
  AOI222_X1 U13701 ( .A1(n12474), .A2(n11109), .B1(n12481), .B2(n12479), .C1(
        n12174), .C2(n12480), .ZN(n14921) );
  INV_X1 U13702 ( .A(n11131), .ZN(n11110) );
  OAI22_X1 U13703 ( .A1(n12488), .A2(n6739), .B1(n11110), .B2(n12387), .ZN(
        n11111) );
  AOI21_X1 U13704 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n12486), .A(n11111), 
        .ZN(n11115) );
  OAI21_X1 U13705 ( .B1(n11113), .B2(n12050), .A(n11112), .ZN(n14923) );
  NAND2_X1 U13706 ( .A1(n14923), .A2(n12457), .ZN(n11114) );
  OAI211_X1 U13707 ( .C1(n14921), .C2(n12486), .A(n11115), .B(n11114), .ZN(
        P3_U3222) );
  AND2_X1 U13708 ( .A1(n11787), .A2(n14328), .ZN(n11122) );
  AOI21_X1 U13709 ( .B1(n15188), .B2(n10307), .A(n11122), .ZN(n11272) );
  AOI22_X1 U13710 ( .A1(n15188), .A2(n11783), .B1(n10307), .B2(n14328), .ZN(
        n11123) );
  XNOR2_X1 U13711 ( .A(n11123), .B(n11795), .ZN(n11271) );
  XOR2_X1 U13712 ( .A(n11272), .B(n11271), .Z(n11269) );
  XNOR2_X1 U13713 ( .A(n11270), .B(n11269), .ZN(n11129) );
  NAND2_X1 U13714 ( .A1(n14329), .A2(n14554), .ZN(n15050) );
  NOR2_X1 U13715 ( .A1(n14055), .A2(n15050), .ZN(n11124) );
  AOI211_X1 U13716 ( .C1(n14023), .C2(n15058), .A(n11125), .B(n11124), .ZN(
        n11126) );
  OAI21_X1 U13717 ( .B1(n14026), .B2(n15054), .A(n11126), .ZN(n11127) );
  AOI21_X1 U13718 ( .B1(n15188), .B2(n9398), .A(n11127), .ZN(n11128) );
  OAI21_X1 U13719 ( .B1(n11129), .B2(n14074), .A(n11128), .ZN(P1_U3217) );
  XNOR2_X1 U13720 ( .A(n11141), .B(n11130), .ZN(n11143) );
  XNOR2_X1 U13721 ( .A(n11143), .B(n11149), .ZN(n11139) );
  NAND2_X1 U13722 ( .A1(n11938), .A2(n11131), .ZN(n11137) );
  INV_X1 U13723 ( .A(n11933), .ZN(n11893) );
  AOI21_X1 U13724 ( .B1(n12481), .B2(n11893), .A(n11132), .ZN(n11136) );
  NAND2_X1 U13725 ( .A1(n11904), .A2(n11133), .ZN(n11135) );
  NAND2_X1 U13726 ( .A1(n12174), .A2(n11931), .ZN(n11134) );
  NAND4_X1 U13727 ( .A1(n11137), .A2(n11136), .A3(n11135), .A4(n11134), .ZN(
        n11138) );
  AOI21_X1 U13728 ( .B1(n11139), .B2(n11920), .A(n11138), .ZN(n11140) );
  INV_X1 U13729 ( .A(n11140), .ZN(P3_U3176) );
  AOI22_X1 U13730 ( .A1(n11143), .A2(n12173), .B1(n11142), .B2(n11141), .ZN(
        n11147) );
  XNOR2_X1 U13731 ( .A(n11145), .B(n11144), .ZN(n11146) );
  XNOR2_X1 U13732 ( .A(n11147), .B(n11146), .ZN(n11154) );
  OAI21_X1 U13733 ( .B1(n11895), .B2(n11149), .A(n11148), .ZN(n11150) );
  AOI21_X1 U13734 ( .B1(n11893), .B2(n12464), .A(n11150), .ZN(n11151) );
  OAI21_X1 U13735 ( .B1(n12614), .B2(n11935), .A(n11151), .ZN(n11152) );
  AOI21_X1 U13736 ( .B1(n11170), .B2(n11938), .A(n11152), .ZN(n11153) );
  OAI21_X1 U13737 ( .B1(n11154), .B2(n11940), .A(n11153), .ZN(P3_U3164) );
  NAND2_X1 U13738 ( .A1(n11156), .A2(n11155), .ZN(n11157) );
  AND2_X1 U13739 ( .A1(n11158), .A2(n11157), .ZN(n11418) );
  INV_X1 U13740 ( .A(n11418), .ZN(n11159) );
  OAI222_X1 U13741 ( .A1(n13905), .A2(n13738), .B1(P2_U3088), .B2(n12867), 
        .C1(n13908), .C2(n11159), .ZN(P2_U3305) );
  INV_X1 U13742 ( .A(n11160), .ZN(n11162) );
  OAI222_X1 U13743 ( .A1(P3_U3151), .A2(n12275), .B1(n12627), .B2(n11162), 
        .C1(n11161), .C2(n12623), .ZN(P3_U3268) );
  OAI21_X1 U13744 ( .B1(n11165), .B2(n11164), .A(n11163), .ZN(n12553) );
  INV_X1 U13745 ( .A(n12553), .ZN(n11175) );
  OAI211_X1 U13746 ( .C1(n11167), .C2(n7607), .A(n11166), .B(n12474), .ZN(
        n11169) );
  AOI22_X1 U13747 ( .A1(n12464), .A2(n12479), .B1(n12480), .B2(n12173), .ZN(
        n11168) );
  NAND2_X1 U13748 ( .A1(n11169), .A2(n11168), .ZN(n12552) );
  AOI22_X1 U13749 ( .A1(n12438), .A2(n11171), .B1(n12485), .B2(n11170), .ZN(
        n11172) );
  OAI21_X1 U13750 ( .B1(n10925), .B2(n12490), .A(n11172), .ZN(n11173) );
  AOI21_X1 U13751 ( .B1(n12552), .B2(n12490), .A(n11173), .ZN(n11174) );
  OAI21_X1 U13752 ( .B1(n11175), .B2(n12493), .A(n11174), .ZN(P3_U3221) );
  NAND2_X1 U13753 ( .A1(n11433), .A2(n11176), .ZN(n11177) );
  OAI211_X1 U13754 ( .C1(n11178), .C2(n11330), .A(n11177), .B(n14311), .ZN(
        P1_U3332) );
  NAND2_X1 U13755 ( .A1(n11433), .A2(n13893), .ZN(n11180) );
  AND2_X1 U13756 ( .A1(n11179), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13177) );
  INV_X1 U13757 ( .A(n13177), .ZN(n13171) );
  OAI211_X1 U13758 ( .C1(n11434), .C2(n13905), .A(n11180), .B(n13171), .ZN(
        P2_U3304) );
  INV_X1 U13759 ( .A(n11181), .ZN(n11184) );
  AOI22_X1 U13760 ( .A1(n12838), .A2(n11182), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11183) );
  OAI21_X1 U13761 ( .B1(n11184), .B2(n12825), .A(n11183), .ZN(n11197) );
  XNOR2_X1 U13762 ( .A(n13582), .B(n12684), .ZN(n11186) );
  NAND2_X1 U13763 ( .A1(n9845), .A2(n13199), .ZN(n11187) );
  INV_X1 U13764 ( .A(n11187), .ZN(n11185) );
  NAND2_X1 U13765 ( .A1(n11186), .A2(n11185), .ZN(n12642) );
  INV_X1 U13766 ( .A(n11186), .ZN(n12695) );
  NAND2_X1 U13767 ( .A1(n12695), .A2(n11187), .ZN(n11188) );
  NAND2_X1 U13768 ( .A1(n12642), .A2(n11188), .ZN(n11195) );
  INV_X1 U13769 ( .A(n11189), .ZN(n11191) );
  NAND2_X1 U13770 ( .A1(n11191), .A2(n11190), .ZN(n11192) );
  AOI211_X1 U13771 ( .C1(n11195), .C2(n11194), .A(n12854), .B(n6691), .ZN(
        n11196) );
  AOI211_X1 U13772 ( .C1(n13582), .C2(n12831), .A(n11197), .B(n11196), .ZN(
        n11198) );
  INV_X1 U13773 ( .A(n11198), .ZN(P2_U3206) );
  INV_X1 U13774 ( .A(n11199), .ZN(n11200) );
  AOI21_X1 U13775 ( .B1(n11210), .B2(n11201), .A(n11200), .ZN(n14946) );
  AOI211_X1 U13776 ( .C1(n14944), .C2(n11202), .A(n14589), .B(n7634), .ZN(
        n14942) );
  INV_X1 U13777 ( .A(n14942), .ZN(n11206) );
  NAND2_X1 U13778 ( .A1(n14323), .A2(n15059), .ZN(n11204) );
  OR2_X1 U13779 ( .A1(n11683), .A2(n14606), .ZN(n11203) );
  NAND2_X1 U13780 ( .A1(n11204), .A2(n11203), .ZN(n14943) );
  AOI21_X1 U13781 ( .B1(n14072), .B2(n15073), .A(n14943), .ZN(n11205) );
  OAI21_X1 U13782 ( .B1(n11206), .B2(n14598), .A(n11205), .ZN(n11209) );
  INV_X1 U13783 ( .A(n14944), .ZN(n14068) );
  OAI22_X1 U13784 ( .A1(n14068), .A2(n14541), .B1(n15104), .B2(n11207), .ZN(
        n11208) );
  AOI21_X1 U13785 ( .B1(n11209), .B2(n15104), .A(n11208), .ZN(n11213) );
  XNOR2_X1 U13786 ( .A(n11211), .B(n11210), .ZN(n14948) );
  NAND2_X1 U13787 ( .A1(n14948), .A2(n14627), .ZN(n11212) );
  OAI211_X1 U13788 ( .C1(n14946), .C2(n14623), .A(n11213), .B(n11212), .ZN(
        P1_U3278) );
  NAND2_X1 U13789 ( .A1(n11230), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n11214) );
  INV_X1 U13790 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11252) );
  NAND2_X1 U13791 ( .A1(n11225), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12193) );
  OR2_X1 U13792 ( .A1(n11225), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n11216) );
  NAND2_X1 U13793 ( .A1(n12193), .A2(n11216), .ZN(n11240) );
  AOI21_X1 U13794 ( .B1(n11217), .B2(n11240), .A(n12183), .ZN(n11249) );
  AOI22_X1 U13795 ( .A1(n11219), .A2(n11218), .B1(P3_REG1_REG_12__SCAN_IN), 
        .B2(n11230), .ZN(n11220) );
  NAND2_X1 U13796 ( .A1(n11257), .A2(n11221), .ZN(n11222) );
  NAND2_X1 U13797 ( .A1(n11225), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12192) );
  OR2_X1 U13798 ( .A1(n11225), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n11223) );
  AND2_X1 U13799 ( .A1(n12192), .A2(n11223), .ZN(n11241) );
  OAI21_X1 U13800 ( .B1(n11224), .B2(n11241), .A(n12186), .ZN(n11229) );
  INV_X1 U13801 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14848) );
  INV_X1 U13802 ( .A(n11225), .ZN(n11226) );
  NAND2_X1 U13803 ( .A1(n14907), .A2(n11226), .ZN(n11227) );
  NAND2_X1 U13804 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n11827)
         );
  OAI211_X1 U13805 ( .C1(n14848), .C2(n14910), .A(n11227), .B(n11827), .ZN(
        n11228) );
  AOI21_X1 U13806 ( .B1(n11229), .B2(n15461), .A(n11228), .ZN(n11248) );
  NAND2_X1 U13807 ( .A1(n11231), .A2(n11230), .ZN(n11232) );
  NAND2_X1 U13808 ( .A1(n11233), .A2(n11232), .ZN(n11259) );
  MUX2_X1 U13809 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12275), .Z(n11234) );
  XNOR2_X1 U13810 ( .A(n11234), .B(n11257), .ZN(n11258) );
  INV_X1 U13811 ( .A(n11234), .ZN(n11236) );
  NAND2_X1 U13812 ( .A1(n11236), .A2(n11235), .ZN(n11244) );
  NAND2_X1 U13813 ( .A1(n11261), .A2(n11244), .ZN(n11239) );
  INV_X1 U13814 ( .A(n11241), .ZN(n11237) );
  MUX2_X1 U13815 ( .A(n11240), .B(n11237), .S(n12275), .Z(n11238) );
  NAND2_X1 U13816 ( .A1(n11239), .A2(n11238), .ZN(n11246) );
  INV_X1 U13817 ( .A(n11240), .ZN(n11242) );
  MUX2_X1 U13818 ( .A(n11242), .B(n11241), .S(n12275), .Z(n11243) );
  AND2_X1 U13819 ( .A1(n11244), .A2(n11243), .ZN(n11245) );
  NAND2_X1 U13820 ( .A1(n11261), .A2(n11245), .ZN(n12195) );
  NAND3_X1 U13821 ( .A1(n11246), .A2(n12280), .A3(n12195), .ZN(n11247) );
  OAI211_X1 U13822 ( .C1(n11249), .C2(n15465), .A(n11248), .B(n11247), .ZN(
        P3_U3196) );
  AOI21_X1 U13823 ( .B1(n11252), .B2(n11251), .A(n11250), .ZN(n11266) );
  OAI21_X1 U13824 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11254), .A(n11253), 
        .ZN(n11264) );
  AOI21_X1 U13825 ( .B1(n15458), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n11255), 
        .ZN(n11256) );
  OAI21_X1 U13826 ( .B1(n15452), .B2(n11257), .A(n11256), .ZN(n11263) );
  NAND2_X1 U13827 ( .A1(n11259), .A2(n11258), .ZN(n11260) );
  AOI21_X1 U13828 ( .B1(n11261), .B2(n11260), .A(n15454), .ZN(n11262) );
  AOI211_X1 U13829 ( .C1(n15461), .C2(n11264), .A(n11263), .B(n11262), .ZN(
        n11265) );
  OAI21_X1 U13830 ( .B1(n11266), .B2(n15465), .A(n11265), .ZN(P3_U3195) );
  OAI22_X1 U13831 ( .A1(n14969), .A2(n11794), .B1(n11268), .B2(n11798), .ZN(
        n11267) );
  XNOR2_X1 U13832 ( .A(n11267), .B(n11795), .ZN(n11288) );
  OAI22_X1 U13833 ( .A1(n14969), .A2(n11798), .B1(n11268), .B2(n11797), .ZN(
        n11287) );
  XNOR2_X1 U13834 ( .A(n11288), .B(n11287), .ZN(n11279) );
  INV_X1 U13835 ( .A(n11271), .ZN(n11274) );
  INV_X1 U13836 ( .A(n11272), .ZN(n11273) );
  NAND2_X1 U13837 ( .A1(n11274), .A2(n11273), .ZN(n11275) );
  INV_X1 U13838 ( .A(n11279), .ZN(n11277) );
  INV_X1 U13839 ( .A(n11297), .ZN(n11293) );
  AOI21_X1 U13840 ( .B1(n11279), .B2(n11278), .A(n11293), .ZN(n11286) );
  NAND2_X1 U13841 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14404)
         );
  NAND2_X1 U13842 ( .A1(n14327), .A2(n15059), .ZN(n11281) );
  NAND2_X1 U13843 ( .A1(n14328), .A2(n14554), .ZN(n11280) );
  NAND2_X1 U13844 ( .A1(n11281), .A2(n11280), .ZN(n14929) );
  NAND2_X1 U13845 ( .A1(n11282), .A2(n14929), .ZN(n11283) );
  OAI211_X1 U13846 ( .C1(n14026), .C2(n14932), .A(n14404), .B(n11283), .ZN(
        n11284) );
  AOI21_X1 U13847 ( .B1(n14934), .B2(n9398), .A(n11284), .ZN(n11285) );
  OAI21_X1 U13848 ( .B1(n11286), .B2(n14074), .A(n11285), .ZN(P1_U3236) );
  NOR2_X1 U13849 ( .A1(n11288), .A2(n11287), .ZN(n11295) );
  NAND2_X1 U13850 ( .A1(n14885), .A2(n11783), .ZN(n11290) );
  NAND2_X1 U13851 ( .A1(n14327), .A2(n10307), .ZN(n11289) );
  NAND2_X1 U13852 ( .A1(n11290), .A2(n11289), .ZN(n11291) );
  XNOR2_X1 U13853 ( .A(n11291), .B(n11765), .ZN(n11304) );
  AND2_X1 U13854 ( .A1(n11787), .A2(n14327), .ZN(n11292) );
  AOI21_X1 U13855 ( .B1(n14885), .B2(n10307), .A(n11292), .ZN(n11305) );
  XNOR2_X1 U13856 ( .A(n11304), .B(n11305), .ZN(n11294) );
  OAI21_X1 U13857 ( .B1(n11293), .B2(n11295), .A(n11294), .ZN(n11298) );
  NOR2_X1 U13858 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  NAND3_X1 U13859 ( .A1(n11298), .A2(n14052), .A3(n11309), .ZN(n11303) );
  NOR2_X1 U13860 ( .A1(n14026), .A2(n11299), .ZN(n11301) );
  INV_X1 U13861 ( .A(n14023), .ZN(n14066) );
  OAI22_X1 U13862 ( .A1(n14066), .A2(n13926), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8048), .ZN(n11300) );
  AOI211_X1 U13863 ( .C1(n14064), .C2(n15058), .A(n11301), .B(n11300), .ZN(
        n11302) );
  OAI211_X1 U13864 ( .C1(n7632), .C2(n14067), .A(n11303), .B(n11302), .ZN(
        P1_U3224) );
  INV_X1 U13865 ( .A(n11304), .ZN(n11307) );
  INV_X1 U13866 ( .A(n11305), .ZN(n11306) );
  NAND2_X1 U13867 ( .A1(n11307), .A2(n11306), .ZN(n11308) );
  AND2_X1 U13868 ( .A1(n11787), .A2(n14326), .ZN(n11310) );
  AOI21_X1 U13869 ( .B1(n14961), .B2(n10307), .A(n11310), .ZN(n11675) );
  AOI22_X1 U13870 ( .A1(n14961), .A2(n11783), .B1(n10307), .B2(n14326), .ZN(
        n11311) );
  XNOR2_X1 U13871 ( .A(n11311), .B(n11795), .ZN(n11674) );
  XOR2_X1 U13872 ( .A(n11675), .B(n11674), .Z(n11672) );
  XNOR2_X1 U13873 ( .A(n11673), .B(n11672), .ZN(n11317) );
  NAND2_X1 U13874 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n15008)
         );
  OAI21_X1 U13875 ( .B1(n14066), .B2(n11683), .A(n15008), .ZN(n11312) );
  AOI21_X1 U13876 ( .B1(n14064), .B2(n14327), .A(n11312), .ZN(n11313) );
  OAI21_X1 U13877 ( .B1(n14026), .B2(n11314), .A(n11313), .ZN(n11315) );
  AOI21_X1 U13878 ( .B1(n14961), .B2(n9398), .A(n11315), .ZN(n11316) );
  OAI21_X1 U13879 ( .B1(n11317), .B2(n14074), .A(n11316), .ZN(P1_U3234) );
  XNOR2_X1 U13880 ( .A(n11319), .B(n11318), .ZN(n11320) );
  AOI222_X1 U13881 ( .A1(n15139), .A2(n11320), .B1(n14322), .B2(n15059), .C1(
        n14324), .C2(n14554), .ZN(n14717) );
  XNOR2_X1 U13882 ( .A(n11321), .B(n7633), .ZN(n14715) );
  INV_X1 U13883 ( .A(n13992), .ZN(n11322) );
  AOI22_X1 U13884 ( .A1(n15106), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11322), 
        .B2(n15073), .ZN(n11323) );
  OAI21_X1 U13885 ( .B1(n7633), .B2(n14541), .A(n11323), .ZN(n11326) );
  XNOR2_X1 U13886 ( .A(n11324), .B(n14285), .ZN(n14718) );
  NOR2_X1 U13887 ( .A1(n14718), .A2(n14623), .ZN(n11325) );
  AOI211_X1 U13888 ( .C1(n14715), .C2(n14628), .A(n11326), .B(n11325), .ZN(
        n11327) );
  OAI21_X1 U13889 ( .B1(n14717), .B2(n15106), .A(n11327), .ZN(P1_U3277) );
  INV_X1 U13890 ( .A(n13894), .ZN(n11328) );
  OAI222_X1 U13891 ( .A1(n11330), .A2(n11329), .B1(n14753), .B2(n11328), .C1(
        P1_U3086), .C2(n6560), .ZN(P1_U3328) );
  INV_X1 U13892 ( .A(SI_30_), .ZN(n11950) );
  NAND2_X1 U13893 ( .A1(n13886), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U13894 ( .A1(n11332), .A2(n11331), .ZN(n11334) );
  NAND2_X1 U13895 ( .A1(n14745), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11333) );
  NAND2_X1 U13896 ( .A1(n11334), .A2(n11333), .ZN(n11943) );
  INV_X1 U13897 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13884) );
  XNOR2_X1 U13898 ( .A(n13884), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11335) );
  XNOR2_X1 U13899 ( .A(n11943), .B(n11335), .ZN(n11949) );
  INV_X1 U13900 ( .A(n11949), .ZN(n11336) );
  INV_X1 U13901 ( .A(n11444), .ZN(n13907) );
  OAI222_X1 U13902 ( .A1(n14755), .A2(n7291), .B1(n14753), .B2(n13907), .C1(
        n7730), .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U13903 ( .A(n11483), .ZN(n13892) );
  OAI222_X1 U13904 ( .A1(n14755), .A2(n13588), .B1(n14753), .B2(n13892), .C1(
        P1_U3086), .C2(n11338), .ZN(P1_U3327) );
  INV_X1 U13905 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n11346) );
  INV_X1 U13906 ( .A(n15497), .ZN(n15509) );
  INV_X1 U13907 ( .A(n11339), .ZN(n11342) );
  XNOR2_X1 U13908 ( .A(n11343), .B(n12132), .ZN(n11345) );
  OAI22_X1 U13909 ( .A1(n11923), .A2(n12408), .B1(n6554), .B2(n12406), .ZN(
        n11344) );
  OAI21_X1 U13910 ( .B1(n11927), .B2(n12556), .A(n11347), .ZN(P3_U3485) );
  INV_X1 U13911 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n11349) );
  MUX2_X1 U13912 ( .A(n11349), .B(n11348), .S(n15519), .Z(n11350) );
  OAI21_X1 U13913 ( .B1(n11927), .B2(n12613), .A(n11350), .ZN(P3_U3453) );
  AND2_X1 U13914 ( .A1(n12973), .A2(n12853), .ZN(n11352) );
  OR2_X1 U13915 ( .A1(n12973), .A2(n12853), .ZN(n11351) );
  NAND2_X1 U13916 ( .A1(n11354), .A2(n13068), .ZN(n11356) );
  AOI22_X1 U13917 ( .A1(n11382), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n15283), 
        .B2(n11381), .ZN(n11355) );
  INV_X1 U13918 ( .A(n13196), .ZN(n12767) );
  XNOR2_X1 U13919 ( .A(n13460), .B(n12767), .ZN(n13448) );
  NAND2_X1 U13920 ( .A1(n13460), .A2(n12767), .ZN(n11357) );
  NAND2_X1 U13921 ( .A1(n11358), .A2(n13068), .ZN(n11360) );
  AOI22_X1 U13922 ( .A1(n15300), .A2(n11381), .B1(n11382), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n11359) );
  INV_X1 U13923 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n12760) );
  INV_X1 U13924 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11361) );
  OAI21_X1 U13925 ( .B1(n11363), .B2(n12760), .A(n11361), .ZN(n11364) );
  NAND2_X1 U13926 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n11362) );
  AND2_X1 U13927 ( .A1(n11364), .A2(n11374), .ZN(n13434) );
  NAND2_X1 U13928 ( .A1(n13434), .A2(n11502), .ZN(n11366) );
  AOI22_X1 U13929 ( .A1(n9306), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n6551), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n11365) );
  OAI211_X1 U13930 ( .C1(n11513), .C2(n11043), .A(n11366), .B(n11365), .ZN(
        n13195) );
  INV_X1 U13931 ( .A(n13195), .ZN(n12986) );
  NAND2_X1 U13932 ( .A1(n13438), .A2(n12986), .ZN(n11367) );
  OR2_X1 U13933 ( .A1(n11369), .A2(n13082), .ZN(n11371) );
  AOI22_X1 U13934 ( .A1(n11382), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n11381), 
        .B2(n13234), .ZN(n11370) );
  INV_X1 U13935 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n11378) );
  NAND2_X1 U13936 ( .A1(n11374), .A2(n11373), .ZN(n11375) );
  NAND2_X1 U13937 ( .A1(n11386), .A2(n11375), .ZN(n13417) );
  OR2_X1 U13938 ( .A1(n13417), .A2(n11492), .ZN(n11377) );
  AOI22_X1 U13939 ( .A1(n13072), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9306), 
        .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n11376) );
  OAI211_X1 U13940 ( .C1(n6549), .C2(n11378), .A(n11377), .B(n11376), .ZN(
        n13194) );
  INV_X1 U13941 ( .A(n13194), .ZN(n12718) );
  XNOR2_X1 U13942 ( .A(n13549), .B(n12718), .ZN(n13409) );
  OR2_X1 U13943 ( .A1(n13549), .A2(n12718), .ZN(n11379) );
  NAND2_X1 U13944 ( .A1(n11380), .A2(n13068), .ZN(n11384) );
  AOI22_X1 U13945 ( .A1(n11382), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11381), 
        .B2(n6984), .ZN(n11383) );
  INV_X1 U13946 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U13947 ( .A1(n11386), .A2(n11385), .ZN(n11387) );
  NAND2_X1 U13948 ( .A1(n11398), .A2(n11387), .ZN(n13398) );
  AOI22_X1 U13949 ( .A1(n13072), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n7659), 
        .B2(P2_REG0_REG_19__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U13950 ( .A1(n6551), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n11388) );
  OAI211_X1 U13951 ( .C1(n13398), .C2(n11492), .A(n11389), .B(n11388), .ZN(
        n13193) );
  INV_X1 U13952 ( .A(n13193), .ZN(n13119) );
  NAND2_X1 U13953 ( .A1(n13543), .A2(n13119), .ZN(n11390) );
  OR2_X1 U13954 ( .A1(n13543), .A2(n13119), .ZN(n11391) );
  NAND2_X1 U13955 ( .A1(n11392), .A2(n11391), .ZN(n13378) );
  OR2_X1 U13956 ( .A1(n11393), .A2(n13082), .ZN(n11396) );
  OR2_X1 U13957 ( .A1(n13083), .A2(n11394), .ZN(n11395) );
  INV_X1 U13958 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13796) );
  NAND2_X1 U13959 ( .A1(n11398), .A2(n13796), .ZN(n11399) );
  NAND2_X1 U13960 ( .A1(n11423), .A2(n11399), .ZN(n13384) );
  OR2_X1 U13961 ( .A1(n13384), .A2(n11492), .ZN(n11404) );
  INV_X1 U13962 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U13963 ( .A1(n6551), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n11401) );
  NAND2_X1 U13964 ( .A1(n13072), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n11400) );
  OAI211_X1 U13965 ( .C1(n9296), .C2(n13797), .A(n11401), .B(n11400), .ZN(
        n11402) );
  INV_X1 U13966 ( .A(n11402), .ZN(n11403) );
  NAND2_X1 U13967 ( .A1(n11404), .A2(n11403), .ZN(n13192) );
  XNOR2_X1 U13968 ( .A(n13537), .B(n13192), .ZN(n13388) );
  NAND2_X1 U13969 ( .A1(n13378), .A2(n13388), .ZN(n11406) );
  INV_X1 U13970 ( .A(n13537), .ZN(n13387) );
  NAND2_X1 U13971 ( .A1(n13387), .A2(n13192), .ZN(n11405) );
  NAND2_X1 U13972 ( .A1(n11407), .A2(n13068), .ZN(n11410) );
  OR2_X1 U13973 ( .A1(n13083), .A2(n11408), .ZN(n11409) );
  XNOR2_X1 U13974 ( .A(n11423), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n13371) );
  NAND2_X1 U13975 ( .A1(n13371), .A2(n11502), .ZN(n11415) );
  INV_X1 U13976 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13800) );
  NAND2_X1 U13977 ( .A1(n6551), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n11412) );
  NAND2_X1 U13978 ( .A1(n13072), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n11411) );
  OAI211_X1 U13979 ( .C1(n9296), .C2(n13800), .A(n11412), .B(n11411), .ZN(
        n11413) );
  INV_X1 U13980 ( .A(n11413), .ZN(n11414) );
  NAND2_X1 U13981 ( .A1(n11415), .A2(n11414), .ZN(n13191) );
  INV_X1 U13982 ( .A(n13191), .ZN(n12807) );
  NOR2_X1 U13983 ( .A1(n13367), .A2(n12807), .ZN(n11416) );
  NAND2_X1 U13984 ( .A1(n13367), .A2(n12807), .ZN(n11417) );
  NAND2_X1 U13985 ( .A1(n11418), .A2(n13068), .ZN(n11420) );
  OR2_X1 U13986 ( .A1(n13083), .A2(n13738), .ZN(n11419) );
  NAND2_X2 U13987 ( .A1(n11420), .A2(n11419), .ZN(n13526) );
  INV_X1 U13988 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12745) );
  INV_X1 U13989 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n11421) );
  OAI21_X1 U13990 ( .B1(n11423), .B2(n12745), .A(n11421), .ZN(n11424) );
  NAND2_X1 U13991 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n11422) );
  NAND2_X1 U13992 ( .A1(n11424), .A2(n11437), .ZN(n13356) );
  OR2_X1 U13993 ( .A1(n13356), .A2(n11492), .ZN(n11430) );
  INV_X1 U13994 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n11427) );
  NAND2_X1 U13995 ( .A1(n6551), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n11426) );
  NAND2_X1 U13996 ( .A1(n9306), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n11425) );
  OAI211_X1 U13997 ( .C1(n11427), .C2(n11513), .A(n11426), .B(n11425), .ZN(
        n11428) );
  INV_X1 U13998 ( .A(n11428), .ZN(n11429) );
  NAND2_X1 U13999 ( .A1(n11430), .A2(n11429), .ZN(n13190) );
  INV_X1 U14000 ( .A(n13190), .ZN(n11431) );
  AND2_X1 U14001 ( .A1(n13526), .A2(n11431), .ZN(n11432) );
  INV_X1 U14002 ( .A(n13526), .ZN(n13361) );
  NAND2_X1 U14003 ( .A1(n11433), .A2(n13068), .ZN(n11436) );
  OR2_X1 U14004 ( .A1(n13083), .A2(n11434), .ZN(n11435) );
  INV_X1 U14005 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12711) );
  NAND2_X1 U14006 ( .A1(n11437), .A2(n12711), .ZN(n11438) );
  NAND2_X1 U14007 ( .A1(n11456), .A2(n11438), .ZN(n12710) );
  INV_X1 U14008 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U14009 ( .A1(n7659), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n11440) );
  NAND2_X1 U14010 ( .A1(n6551), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n11439) );
  OAI211_X1 U14011 ( .C1(n11513), .C2(n11441), .A(n11440), .B(n11439), .ZN(
        n11442) );
  INV_X1 U14012 ( .A(n11442), .ZN(n11443) );
  OAI21_X1 U14013 ( .B1(n12710), .B2(n11492), .A(n11443), .ZN(n13189) );
  INV_X1 U14014 ( .A(n13189), .ZN(n12809) );
  INV_X1 U14015 ( .A(n13520), .ZN(n13340) );
  NAND2_X1 U14016 ( .A1(n11444), .A2(n13068), .ZN(n11446) );
  OR2_X1 U14017 ( .A1(n13083), .A2(n13906), .ZN(n11445) );
  XNOR2_X1 U14018 ( .A(n11456), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n13327) );
  NAND2_X1 U14019 ( .A1(n13327), .A2(n11502), .ZN(n11451) );
  INV_X1 U14020 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13330) );
  NAND2_X1 U14021 ( .A1(n6551), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U14022 ( .A1(n9306), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n11447) );
  OAI211_X1 U14023 ( .C1(n13330), .C2(n11513), .A(n11448), .B(n11447), .ZN(
        n11449) );
  INV_X1 U14024 ( .A(n11449), .ZN(n11450) );
  NAND2_X1 U14025 ( .A1(n11451), .A2(n11450), .ZN(n13188) );
  INV_X1 U14026 ( .A(n13188), .ZN(n11452) );
  XNOR2_X1 U14027 ( .A(n13332), .B(n11452), .ZN(n13320) );
  INV_X1 U14028 ( .A(n13320), .ZN(n13322) );
  NAND2_X1 U14029 ( .A1(n13332), .A2(n11452), .ZN(n11453) );
  NAND2_X1 U14030 ( .A1(n13901), .A2(n13068), .ZN(n11455) );
  OR2_X1 U14031 ( .A1(n13083), .A2(n13903), .ZN(n11454) );
  INV_X1 U14032 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12779) );
  INV_X1 U14033 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12752) );
  OAI21_X1 U14034 ( .B1(n11456), .B2(n12779), .A(n12752), .ZN(n11457) );
  AND2_X1 U14035 ( .A1(n11467), .A2(n11457), .ZN(n13312) );
  NAND2_X1 U14036 ( .A1(n13312), .A2(n11502), .ZN(n11462) );
  INV_X1 U14037 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13701) );
  NAND2_X1 U14038 ( .A1(n13072), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n11459) );
  NAND2_X1 U14039 ( .A1(n6551), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n11458) );
  OAI211_X1 U14040 ( .C1(n9296), .C2(n13701), .A(n11459), .B(n11458), .ZN(
        n11460) );
  INV_X1 U14041 ( .A(n11460), .ZN(n11461) );
  NAND2_X1 U14042 ( .A1(n11462), .A2(n11461), .ZN(n13187) );
  XNOR2_X1 U14043 ( .A(n13314), .B(n13187), .ZN(n13308) );
  NAND2_X1 U14044 ( .A1(n13309), .A2(n13308), .ZN(n11464) );
  INV_X1 U14045 ( .A(n13187), .ZN(n13043) );
  NAND2_X1 U14046 ( .A1(n13314), .A2(n13043), .ZN(n11463) );
  NAND2_X1 U14047 ( .A1(n11464), .A2(n11463), .ZN(n13298) );
  NAND2_X1 U14048 ( .A1(n13898), .A2(n13068), .ZN(n11466) );
  OR2_X1 U14049 ( .A1(n13083), .A2(n13899), .ZN(n11465) );
  INV_X1 U14050 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13662) );
  NAND2_X1 U14051 ( .A1(n11467), .A2(n13662), .ZN(n11468) );
  NAND2_X1 U14052 ( .A1(n13300), .A2(n11502), .ZN(n11474) );
  INV_X1 U14053 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U14054 ( .A1(n7659), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14055 ( .A1(n6551), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n11469) );
  OAI211_X1 U14056 ( .C1(n11471), .C2(n11513), .A(n11470), .B(n11469), .ZN(
        n11472) );
  INV_X1 U14057 ( .A(n11472), .ZN(n11473) );
  NAND2_X1 U14058 ( .A1(n11474), .A2(n11473), .ZN(n13186) );
  INV_X1 U14059 ( .A(n13186), .ZN(n11538) );
  OR2_X1 U14060 ( .A1(n13303), .A2(n11538), .ZN(n13118) );
  NAND2_X1 U14061 ( .A1(n13298), .A2(n13118), .ZN(n11475) );
  NAND2_X1 U14062 ( .A1(n13303), .A2(n11538), .ZN(n13117) );
  OR2_X1 U14063 ( .A1(n6565), .A2(n13897), .ZN(n11476) );
  XNOR2_X1 U14064 ( .A(n11489), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13290) );
  NAND2_X1 U14065 ( .A1(n13290), .A2(n11502), .ZN(n11482) );
  INV_X1 U14066 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n11479) );
  NAND2_X1 U14067 ( .A1(n9306), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n11478) );
  NAND2_X1 U14068 ( .A1(n6551), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n11477) );
  OAI211_X1 U14069 ( .C1(n11479), .C2(n11513), .A(n11478), .B(n11477), .ZN(
        n11480) );
  INV_X1 U14070 ( .A(n11480), .ZN(n11481) );
  NAND2_X1 U14071 ( .A1(n11482), .A2(n11481), .ZN(n13185) );
  INV_X1 U14072 ( .A(n13185), .ZN(n11499) );
  XNOR2_X1 U14073 ( .A(n13493), .B(n11499), .ZN(n13147) );
  NAND2_X1 U14074 ( .A1(n11483), .A2(n13068), .ZN(n11486) );
  OR2_X1 U14075 ( .A1(n13083), .A2(n11484), .ZN(n11485) );
  INV_X1 U14076 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12689) );
  INV_X1 U14077 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11487) );
  OAI21_X1 U14078 ( .B1(n11489), .B2(n12689), .A(n11487), .ZN(n11491) );
  NAND2_X1 U14079 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n11488) );
  NOR2_X1 U14080 ( .A1(n11489), .A2(n11488), .ZN(n11518) );
  INV_X1 U14081 ( .A(n11518), .ZN(n11490) );
  NAND2_X1 U14082 ( .A1(n11491), .A2(n11490), .ZN(n13271) );
  OR2_X1 U14083 ( .A1(n13271), .A2(n11492), .ZN(n11497) );
  INV_X1 U14084 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13275) );
  NAND2_X1 U14085 ( .A1(n6551), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U14086 ( .A1(n9306), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n11493) );
  OAI211_X1 U14087 ( .C1(n13275), .C2(n11513), .A(n11494), .B(n11493), .ZN(
        n11495) );
  INV_X1 U14088 ( .A(n11495), .ZN(n11496) );
  NAND2_X1 U14089 ( .A1(n11497), .A2(n11496), .ZN(n13184) );
  INV_X1 U14090 ( .A(n13184), .ZN(n11540) );
  NAND2_X1 U14091 ( .A1(n13490), .A2(n11540), .ZN(n11498) );
  NAND2_X1 U14092 ( .A1(n11500), .A2(n11498), .ZN(n13148) );
  NAND2_X1 U14093 ( .A1(n13493), .A2(n11499), .ZN(n13266) );
  OR2_X1 U14094 ( .A1(n6565), .A2(n13886), .ZN(n11501) );
  NAND2_X1 U14095 ( .A1(n11518), .A2(n11502), .ZN(n11508) );
  INV_X1 U14096 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n11505) );
  NAND2_X1 U14097 ( .A1(n6551), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n11504) );
  NAND2_X1 U14098 ( .A1(n7659), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n11503) );
  OAI211_X1 U14099 ( .C1(n11505), .C2(n11513), .A(n11504), .B(n11503), .ZN(
        n11506) );
  INV_X1 U14100 ( .A(n11506), .ZN(n11507) );
  NAND2_X1 U14101 ( .A1(n11508), .A2(n11507), .ZN(n13183) );
  NAND2_X1 U14102 ( .A1(n13184), .A2(n13167), .ZN(n11515) );
  AOI21_X1 U14103 ( .B1(n13169), .B2(P2_B_REG_SCAN_IN), .A(n12808), .ZN(n13252) );
  INV_X1 U14104 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13258) );
  NAND2_X1 U14105 ( .A1(n6551), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n11512) );
  NAND2_X1 U14106 ( .A1(n7659), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11511) );
  OAI211_X1 U14107 ( .C1(n11513), .C2(n13258), .A(n11512), .B(n11511), .ZN(
        n13182) );
  NAND2_X1 U14108 ( .A1(n13252), .A2(n13182), .ZN(n11514) );
  INV_X1 U14109 ( .A(n13438), .ZN(n13555) );
  AND2_X2 U14110 ( .A1(n13457), .A2(n13555), .ZN(n13433) );
  INV_X1 U14111 ( .A(n13549), .ZN(n13421) );
  NAND2_X1 U14112 ( .A1(n13433), .A2(n13421), .ZN(n13414) );
  NAND2_X1 U14113 ( .A1(n13387), .A2(n13396), .ZN(n13381) );
  NAND2_X1 U14114 ( .A1(n13513), .A2(n13337), .ZN(n13326) );
  OR2_X2 U14115 ( .A1(n13326), .A2(n13314), .ZN(n13311) );
  INV_X1 U14116 ( .A(n13490), .ZN(n13276) );
  AOI211_X1 U14117 ( .C1(n13484), .C2(n13273), .A(n13562), .B(n13257), .ZN(
        n13483) );
  INV_X1 U14118 ( .A(n13484), .ZN(n11520) );
  AOI22_X1 U14119 ( .A1(n15320), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n11518), 
        .B2(n15318), .ZN(n11519) );
  OAI21_X1 U14120 ( .B1(n11520), .B2(n13420), .A(n11519), .ZN(n11541) );
  OR2_X1 U14121 ( .A1(n12973), .A2(n13197), .ZN(n11521) );
  INV_X1 U14122 ( .A(n13448), .ZN(n13444) );
  NAND2_X1 U14123 ( .A1(n13460), .A2(n13196), .ZN(n11523) );
  XNOR2_X1 U14124 ( .A(n13438), .B(n12986), .ZN(n13430) );
  OR2_X1 U14125 ( .A1(n13549), .A2(n13194), .ZN(n11524) );
  NAND2_X1 U14126 ( .A1(n13422), .A2(n11524), .ZN(n13393) );
  NAND2_X1 U14127 ( .A1(n13543), .A2(n13193), .ZN(n11525) );
  NAND2_X1 U14128 ( .A1(n13393), .A2(n11525), .ZN(n11527) );
  OR2_X1 U14129 ( .A1(n13543), .A2(n13193), .ZN(n11526) );
  NOR2_X1 U14130 ( .A1(n13537), .A2(n13192), .ZN(n11528) );
  NAND2_X1 U14131 ( .A1(n13537), .A2(n13192), .ZN(n11529) );
  AND2_X1 U14132 ( .A1(n13367), .A2(n13191), .ZN(n11530) );
  NAND2_X1 U14133 ( .A1(n13526), .A2(n13190), .ZN(n11531) );
  OR2_X1 U14134 ( .A1(n13520), .A2(n13189), .ZN(n11532) );
  NAND2_X1 U14135 ( .A1(n13336), .A2(n11532), .ZN(n11534) );
  NAND2_X1 U14136 ( .A1(n13520), .A2(n13189), .ZN(n11533) );
  NAND2_X1 U14137 ( .A1(n11534), .A2(n11533), .ZN(n13321) );
  NAND2_X1 U14138 ( .A1(n13332), .A2(n13188), .ZN(n11535) );
  AND2_X1 U14139 ( .A1(n13314), .A2(n13187), .ZN(n11536) );
  OR2_X1 U14140 ( .A1(n13314), .A2(n13187), .ZN(n11537) );
  NOR2_X1 U14141 ( .A1(n13303), .A2(n13186), .ZN(n11539) );
  XNOR2_X1 U14142 ( .A(n11543), .B(n11542), .ZN(n15469) );
  NAND2_X1 U14143 ( .A1(n11997), .A2(n15508), .ZN(n15470) );
  NOR2_X1 U14144 ( .A1(n15470), .A2(n11544), .ZN(n11551) );
  OAI21_X1 U14145 ( .B1(n11546), .B2(n11542), .A(n11545), .ZN(n11549) );
  OAI22_X1 U14146 ( .A1(n11547), .A2(n12406), .B1(n8837), .B2(n12408), .ZN(
        n11548) );
  AOI21_X1 U14147 ( .B1(n11549), .B2(n12474), .A(n11548), .ZN(n11550) );
  OAI21_X1 U14148 ( .B1(n11601), .B2(n15469), .A(n11550), .ZN(n15471) );
  AOI211_X1 U14149 ( .C1(n12485), .C2(P3_REG3_REG_2__SCAN_IN), .A(n11551), .B(
        n15471), .ZN(n11552) );
  MUX2_X1 U14150 ( .A(n11553), .B(n11552), .S(n12490), .Z(n11554) );
  OAI21_X1 U14151 ( .B1(n15469), .B2(n12299), .A(n11554), .ZN(P3_U3231) );
  AOI21_X1 U14152 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n12485), .A(n11555), .ZN(
        n11556) );
  MUX2_X1 U14153 ( .A(n11557), .B(n11556), .S(n12490), .Z(n11558) );
  OAI21_X1 U14154 ( .B1(n11559), .B2(n12488), .A(n11558), .ZN(P3_U3233) );
  XNOR2_X1 U14155 ( .A(n14442), .B(n14639), .ZN(n11560) );
  NOR2_X1 U14156 ( .A1(n11560), .A2(n14589), .ZN(n14638) );
  NAND2_X1 U14157 ( .A1(n14315), .A2(n15059), .ZN(n11563) );
  NAND2_X1 U14158 ( .A1(n14317), .A2(n14554), .ZN(n11562) );
  INV_X1 U14159 ( .A(n14641), .ZN(n11566) );
  AOI21_X1 U14160 ( .B1(n14638), .B2(n14617), .A(n11566), .ZN(n11574) );
  OAI22_X1 U14161 ( .A1(n15104), .A2(n11567), .B1(n11804), .B2(n15091), .ZN(
        n11572) );
  OAI21_X1 U14162 ( .B1(n11570), .B2(n11569), .A(n11568), .ZN(n14642) );
  NOR2_X1 U14163 ( .A1(n14642), .A2(n14623), .ZN(n11571) );
  AOI211_X1 U14164 ( .C1(n15075), .C2(n14639), .A(n11572), .B(n11571), .ZN(
        n11573) );
  OAI21_X1 U14165 ( .B1(n11574), .B2(n15106), .A(n11573), .ZN(P1_U3265) );
  INV_X1 U14166 ( .A(n11811), .ZN(n11576) );
  OAI22_X1 U14167 ( .A1(n11576), .A2(n12387), .B1(n12490), .B2(n11575), .ZN(
        n11579) );
  NOR2_X1 U14168 ( .A1(n11577), .A2(n12486), .ZN(n11578) );
  OAI21_X1 U14169 ( .B1(n11581), .B2(n12493), .A(n11580), .ZN(P3_U3205) );
  INV_X1 U14170 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n11602) );
  NAND2_X1 U14171 ( .A1(n11582), .A2(n11983), .ZN(n11583) );
  AND2_X1 U14172 ( .A1(n12304), .A2(n11586), .ZN(n11585) );
  INV_X1 U14173 ( .A(n11586), .ZN(n11588) );
  NOR2_X1 U14174 ( .A1(n11588), .A2(n11587), .ZN(n11589) );
  NOR2_X1 U14175 ( .A1(n11590), .A2(n11589), .ZN(n11598) );
  AND2_X1 U14176 ( .A1(n12304), .A2(n11592), .ZN(n11591) );
  NAND2_X1 U14177 ( .A1(n12305), .A2(n11591), .ZN(n11596) );
  INV_X1 U14178 ( .A(n11592), .ZN(n11594) );
  OR2_X1 U14179 ( .A1(n11594), .A2(n11593), .ZN(n11595) );
  NAND2_X1 U14180 ( .A1(n11596), .A2(n11595), .ZN(n11597) );
  OAI21_X1 U14181 ( .B1(n11598), .B2(n11983), .A(n11597), .ZN(n11600) );
  OAI22_X1 U14182 ( .A1(n11666), .A2(n12408), .B1(n11860), .B2(n12406), .ZN(
        n11599) );
  OAI21_X1 U14183 ( .B1(n11671), .B2(n12556), .A(n11603), .ZN(P3_U3486) );
  INV_X1 U14184 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n11605) );
  MUX2_X1 U14185 ( .A(n11605), .B(n11604), .S(n15519), .Z(n11606) );
  OAI21_X1 U14186 ( .B1(n11671), .B2(n12613), .A(n11606), .ZN(P3_U3454) );
  NAND2_X1 U14187 ( .A1(n11607), .A2(n12490), .ZN(n11612) );
  INV_X1 U14188 ( .A(n11668), .ZN(n11609) );
  OAI22_X1 U14189 ( .A1(n11609), .A2(n12387), .B1(n12490), .B2(n11608), .ZN(
        n11610) );
  AOI21_X1 U14190 ( .B1(n11622), .B2(n12438), .A(n11610), .ZN(n11611) );
  OAI211_X1 U14191 ( .C1(n11613), .C2(n12299), .A(n11612), .B(n11611), .ZN(
        P3_U3206) );
  INV_X1 U14192 ( .A(n11614), .ZN(n11619) );
  NAND2_X1 U14193 ( .A1(n11615), .A2(n12485), .ZN(n12285) );
  NAND2_X1 U14194 ( .A1(n12486), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n11616) );
  OAI211_X1 U14195 ( .C1(n11617), .C2(n12488), .A(n12285), .B(n11616), .ZN(
        n11618) );
  AOI21_X1 U14196 ( .B1(n11619), .B2(n12490), .A(n11618), .ZN(n11620) );
  OAI21_X1 U14197 ( .B1(n11621), .B2(n12493), .A(n11620), .ZN(P3_U3204) );
  XNOR2_X1 U14198 ( .A(n11622), .B(n11655), .ZN(n11815) );
  NOR2_X1 U14199 ( .A1(n11815), .A2(n12169), .ZN(n11809) );
  AOI21_X1 U14200 ( .B1(n12169), .B2(n11815), .A(n11809), .ZN(n11663) );
  XNOR2_X1 U14201 ( .A(n12589), .B(n11655), .ZN(n11637) );
  XNOR2_X1 U14202 ( .A(n12605), .B(n11655), .ZN(n11626) );
  INV_X1 U14203 ( .A(n11626), .ZN(n11627) );
  XNOR2_X1 U14204 ( .A(n11626), .B(n11625), .ZN(n11824) );
  XOR2_X1 U14205 ( .A(n11655), .B(n12543), .Z(n11928) );
  OAI21_X1 U14206 ( .B1(n11930), .B2(n11829), .A(n11628), .ZN(n11865) );
  XNOR2_X1 U14207 ( .A(n12539), .B(n11655), .ZN(n11629) );
  XNOR2_X1 U14208 ( .A(n11629), .B(n12452), .ZN(n11864) );
  INV_X1 U14209 ( .A(n11629), .ZN(n11630) );
  XNOR2_X1 U14210 ( .A(n12535), .B(n11655), .ZN(n11631) );
  XNOR2_X1 U14211 ( .A(n11631), .B(n12405), .ZN(n11872) );
  XNOR2_X1 U14212 ( .A(n12598), .B(n11655), .ZN(n11632) );
  XNOR2_X1 U14213 ( .A(n11632), .B(n12422), .ZN(n11908) );
  INV_X1 U14214 ( .A(n11632), .ZN(n11633) );
  XNOR2_X1 U14215 ( .A(n12390), .B(n11655), .ZN(n11634) );
  XNOR2_X1 U14216 ( .A(n11634), .B(n12407), .ZN(n11841) );
  XNOR2_X1 U14217 ( .A(n12104), .B(n11655), .ZN(n11636) );
  XNOR2_X1 U14218 ( .A(n11636), .B(n12381), .ZN(n11891) );
  INV_X1 U14219 ( .A(n11634), .ZN(n11635) );
  NAND2_X1 U14220 ( .A1(n11635), .A2(n12407), .ZN(n11888) );
  XNOR2_X1 U14221 ( .A(n11637), .B(n12372), .ZN(n11847) );
  NAND2_X1 U14222 ( .A1(n11636), .A2(n12172), .ZN(n11848) );
  XNOR2_X1 U14223 ( .A(n11905), .B(n11655), .ZN(n11639) );
  NOR2_X1 U14224 ( .A1(n11638), .A2(n11639), .ZN(n11641) );
  XNOR2_X1 U14225 ( .A(n12338), .B(n11655), .ZN(n11643) );
  INV_X1 U14226 ( .A(n11642), .ZN(n11646) );
  INV_X1 U14227 ( .A(n11643), .ZN(n11645) );
  XNOR2_X1 U14228 ( .A(n11878), .B(n11807), .ZN(n11647) );
  NAND2_X1 U14229 ( .A1(n11647), .A2(n12335), .ZN(n11856) );
  INV_X1 U14230 ( .A(n11647), .ZN(n11648) );
  NAND2_X1 U14231 ( .A1(n11648), .A2(n12170), .ZN(n11649) );
  XNOR2_X1 U14232 ( .A(n11650), .B(n11807), .ZN(n11651) );
  NAND2_X1 U14233 ( .A1(n11651), .A2(n6554), .ZN(n11915) );
  INV_X1 U14234 ( .A(n11651), .ZN(n11652) );
  NAND2_X1 U14235 ( .A1(n11652), .A2(n12321), .ZN(n11653) );
  NAND2_X1 U14236 ( .A1(n11915), .A2(n11653), .ZN(n11855) );
  INV_X1 U14237 ( .A(n11855), .ZN(n11654) );
  XNOR2_X1 U14238 ( .A(n12295), .B(n11655), .ZN(n11658) );
  NOR2_X1 U14239 ( .A1(n11658), .A2(n12306), .ZN(n11657) );
  INV_X1 U14240 ( .A(n11657), .ZN(n11656) );
  AND2_X1 U14241 ( .A1(n11915), .A2(n11656), .ZN(n11661) );
  AOI21_X1 U14242 ( .B1(n12306), .B2(n11658), .A(n11657), .ZN(n11919) );
  OR2_X1 U14243 ( .A1(n11657), .A2(n11919), .ZN(n11659) );
  INV_X1 U14244 ( .A(n11659), .ZN(n11660) );
  OAI21_X1 U14245 ( .B1(n11663), .B2(n11662), .A(n11822), .ZN(n11664) );
  NAND2_X1 U14246 ( .A1(n11664), .A2(n11920), .ZN(n11670) );
  AOI22_X1 U14247 ( .A1(n12306), .A2(n11931), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11665) );
  OAI21_X1 U14248 ( .B1(n11666), .B2(n11933), .A(n11665), .ZN(n11667) );
  AOI21_X1 U14249 ( .B1(n11668), .B2(n11938), .A(n11667), .ZN(n11669) );
  OAI211_X1 U14250 ( .C1(n11671), .C2(n11935), .A(n11670), .B(n11669), .ZN(
        P3_U3154) );
  INV_X1 U14251 ( .A(n11674), .ZN(n11677) );
  INV_X1 U14252 ( .A(n11675), .ZN(n11676) );
  NAND2_X1 U14253 ( .A1(n11677), .A2(n11676), .ZN(n11678) );
  NAND2_X1 U14254 ( .A1(n14952), .A2(n11783), .ZN(n11681) );
  OR2_X1 U14255 ( .A1(n11683), .A2(n11798), .ZN(n11680) );
  NAND2_X1 U14256 ( .A1(n11681), .A2(n11680), .ZN(n11682) );
  XNOR2_X1 U14257 ( .A(n11682), .B(n11765), .ZN(n11686) );
  NOR2_X1 U14258 ( .A1(n11683), .A2(n11797), .ZN(n11684) );
  AOI21_X1 U14259 ( .B1(n14952), .B2(n10307), .A(n11684), .ZN(n11685) );
  NAND2_X1 U14260 ( .A1(n11686), .A2(n11685), .ZN(n11688) );
  OAI21_X1 U14261 ( .B1(n11686), .B2(n11685), .A(n11688), .ZN(n13921) );
  AOI22_X1 U14262 ( .A1(n14944), .A2(n11783), .B1(n10307), .B2(n14324), .ZN(
        n11689) );
  OAI22_X1 U14263 ( .A1(n14068), .A2(n11798), .B1(n11690), .B2(n11797), .ZN(
        n14063) );
  INV_X1 U14264 ( .A(n14063), .ZN(n11691) );
  NAND2_X1 U14265 ( .A1(n14714), .A2(n11783), .ZN(n11694) );
  NAND2_X1 U14266 ( .A1(n14323), .A2(n10307), .ZN(n11693) );
  NAND2_X1 U14267 ( .A1(n11694), .A2(n11693), .ZN(n11695) );
  XNOR2_X1 U14268 ( .A(n11695), .B(n11795), .ZN(n11699) );
  NAND2_X1 U14269 ( .A1(n14714), .A2(n10307), .ZN(n11697) );
  NAND2_X1 U14270 ( .A1(n14323), .A2(n11787), .ZN(n11696) );
  NAND2_X1 U14271 ( .A1(n11697), .A2(n11696), .ZN(n11698) );
  NOR2_X1 U14272 ( .A1(n11699), .A2(n11698), .ZN(n14000) );
  AOI21_X1 U14273 ( .B1(n11699), .B2(n11698), .A(n14000), .ZN(n13990) );
  INV_X1 U14274 ( .A(n14000), .ZN(n11700) );
  NAND2_X1 U14275 ( .A1(n14710), .A2(n11783), .ZN(n11702) );
  NAND2_X1 U14276 ( .A1(n14322), .A2(n10307), .ZN(n11701) );
  NAND2_X1 U14277 ( .A1(n11702), .A2(n11701), .ZN(n11703) );
  XNOR2_X1 U14278 ( .A(n11703), .B(n11765), .ZN(n11705) );
  AND2_X1 U14279 ( .A1(n14322), .A2(n11787), .ZN(n11704) );
  AOI21_X1 U14280 ( .B1(n14710), .B2(n10307), .A(n11704), .ZN(n11706) );
  NAND2_X1 U14281 ( .A1(n11705), .A2(n11706), .ZN(n11710) );
  INV_X1 U14282 ( .A(n11705), .ZN(n11708) );
  INV_X1 U14283 ( .A(n11706), .ZN(n11707) );
  NAND2_X1 U14284 ( .A1(n11708), .A2(n11707), .ZN(n11709) );
  AND2_X1 U14285 ( .A1(n11710), .A2(n11709), .ZN(n13999) );
  NAND2_X1 U14286 ( .A1(n14002), .A2(n11710), .ZN(n14042) );
  OAI22_X1 U14287 ( .A1(n14198), .A2(n11798), .B1(n14609), .B2(n11797), .ZN(
        n11716) );
  OAI22_X1 U14288 ( .A1(n14198), .A2(n11794), .B1(n14609), .B2(n11798), .ZN(
        n11711) );
  XNOR2_X1 U14289 ( .A(n11711), .B(n11795), .ZN(n11715) );
  XOR2_X1 U14290 ( .A(n11716), .B(n11715), .Z(n14043) );
  NAND2_X1 U14291 ( .A1(n14042), .A2(n14043), .ZN(n13948) );
  NOR2_X1 U14292 ( .A1(n11712), .A2(n11797), .ZN(n11713) );
  AOI21_X1 U14293 ( .B1(n14581), .B2(n10307), .A(n11713), .ZN(n11719) );
  AOI22_X1 U14294 ( .A1(n14581), .A2(n11783), .B1(n10307), .B2(n14555), .ZN(
        n11714) );
  XNOR2_X1 U14295 ( .A(n11714), .B(n11795), .ZN(n11720) );
  XOR2_X1 U14296 ( .A(n11719), .B(n11720), .Z(n13951) );
  INV_X1 U14297 ( .A(n11715), .ZN(n11718) );
  INV_X1 U14298 ( .A(n11716), .ZN(n11717) );
  NAND2_X1 U14299 ( .A1(n11718), .A2(n11717), .ZN(n13949) );
  OR2_X1 U14300 ( .A1(n11720), .A2(n11719), .ZN(n11721) );
  AND2_X1 U14301 ( .A1(n14577), .A2(n11787), .ZN(n11722) );
  AOI21_X1 U14302 ( .B1(n14688), .B2(n10307), .A(n11722), .ZN(n11725) );
  AOI22_X1 U14303 ( .A1(n14688), .A2(n11783), .B1(n10307), .B2(n14577), .ZN(
        n11723) );
  XNOR2_X1 U14304 ( .A(n11723), .B(n11795), .ZN(n11724) );
  XOR2_X1 U14305 ( .A(n11725), .B(n11724), .Z(n14021) );
  INV_X1 U14306 ( .A(n11724), .ZN(n11727) );
  INV_X1 U14307 ( .A(n11725), .ZN(n11726) );
  NAND2_X1 U14308 ( .A1(n11727), .A2(n11726), .ZN(n11728) );
  NAND2_X1 U14309 ( .A1(n14682), .A2(n11783), .ZN(n11731) );
  NAND2_X1 U14310 ( .A1(n14553), .A2(n10307), .ZN(n11730) );
  NAND2_X1 U14311 ( .A1(n11731), .A2(n11730), .ZN(n11732) );
  XNOR2_X1 U14312 ( .A(n11732), .B(n11765), .ZN(n11735) );
  AND2_X1 U14313 ( .A1(n14553), .A2(n11787), .ZN(n11733) );
  AOI21_X1 U14314 ( .B1(n14682), .B2(n10307), .A(n11733), .ZN(n11734) );
  NAND2_X1 U14315 ( .A1(n11735), .A2(n11734), .ZN(n14030) );
  OAI21_X1 U14316 ( .B1(n11735), .B2(n11734), .A(n14030), .ZN(n13970) );
  INV_X1 U14317 ( .A(n13970), .ZN(n11736) );
  OAI22_X1 U14318 ( .A1(n14676), .A2(n11794), .B1(n14216), .B2(n11798), .ZN(
        n11737) );
  XNOR2_X1 U14319 ( .A(n11737), .B(n11765), .ZN(n11739) );
  NOR2_X1 U14320 ( .A1(n14216), .A2(n11797), .ZN(n11738) );
  AOI21_X1 U14321 ( .B1(n14528), .B2(n10307), .A(n11738), .ZN(n11740) );
  NAND2_X1 U14322 ( .A1(n11739), .A2(n11740), .ZN(n13935) );
  INV_X1 U14323 ( .A(n11739), .ZN(n11742) );
  INV_X1 U14324 ( .A(n11740), .ZN(n11741) );
  NAND2_X1 U14325 ( .A1(n11742), .A2(n11741), .ZN(n11743) );
  AND2_X1 U14326 ( .A1(n13935), .A2(n11743), .ZN(n14031) );
  NAND2_X1 U14327 ( .A1(n14668), .A2(n11783), .ZN(n11746) );
  NAND2_X1 U14328 ( .A1(n14320), .A2(n10307), .ZN(n11745) );
  NAND2_X1 U14329 ( .A1(n11746), .A2(n11745), .ZN(n11747) );
  XNOR2_X1 U14330 ( .A(n11747), .B(n11765), .ZN(n11749) );
  AND2_X1 U14331 ( .A1(n11787), .A2(n14320), .ZN(n11748) );
  AOI21_X1 U14332 ( .B1(n14668), .B2(n10307), .A(n11748), .ZN(n11750) );
  NAND2_X1 U14333 ( .A1(n11749), .A2(n11750), .ZN(n14016) );
  INV_X1 U14334 ( .A(n11749), .ZN(n11752) );
  INV_X1 U14335 ( .A(n11750), .ZN(n11751) );
  NAND2_X1 U14336 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  NAND2_X1 U14337 ( .A1(n14664), .A2(n11783), .ZN(n11755) );
  NAND2_X1 U14338 ( .A1(n14512), .A2(n10307), .ZN(n11754) );
  NAND2_X1 U14339 ( .A1(n11755), .A2(n11754), .ZN(n11756) );
  XNOR2_X1 U14340 ( .A(n11756), .B(n11765), .ZN(n11758) );
  AND2_X1 U14341 ( .A1(n11787), .A2(n14512), .ZN(n11757) );
  AOI21_X1 U14342 ( .B1(n14664), .B2(n10307), .A(n11757), .ZN(n11759) );
  NAND2_X1 U14343 ( .A1(n11758), .A2(n11759), .ZN(n13982) );
  INV_X1 U14344 ( .A(n11758), .ZN(n11761) );
  INV_X1 U14345 ( .A(n11759), .ZN(n11760) );
  NAND2_X1 U14346 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  NAND2_X1 U14347 ( .A1(n14659), .A2(n11783), .ZN(n11764) );
  NAND2_X1 U14348 ( .A1(n14319), .A2(n10307), .ZN(n11763) );
  NAND2_X1 U14349 ( .A1(n11764), .A2(n11763), .ZN(n11766) );
  XNOR2_X1 U14350 ( .A(n11766), .B(n11765), .ZN(n11768) );
  AND2_X1 U14351 ( .A1(n11787), .A2(n14319), .ZN(n11767) );
  AOI21_X1 U14352 ( .B1(n14659), .B2(n10307), .A(n11767), .ZN(n11769) );
  NAND2_X1 U14353 ( .A1(n11768), .A2(n11769), .ZN(n11774) );
  INV_X1 U14354 ( .A(n11768), .ZN(n11771) );
  INV_X1 U14355 ( .A(n11769), .ZN(n11770) );
  NAND2_X1 U14356 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  NAND2_X1 U14357 ( .A1(n14652), .A2(n11783), .ZN(n11776) );
  NAND2_X1 U14358 ( .A1(n14318), .A2(n10307), .ZN(n11775) );
  NAND2_X1 U14359 ( .A1(n11776), .A2(n11775), .ZN(n11777) );
  XNOR2_X1 U14360 ( .A(n11777), .B(n11795), .ZN(n11781) );
  NAND2_X1 U14361 ( .A1(n14652), .A2(n10307), .ZN(n11779) );
  NAND2_X1 U14362 ( .A1(n11787), .A2(n14318), .ZN(n11778) );
  NAND2_X1 U14363 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  NOR2_X1 U14364 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  AOI21_X1 U14365 ( .B1(n11781), .B2(n11780), .A(n11782), .ZN(n14051) );
  NAND2_X1 U14366 ( .A1(n14644), .A2(n11783), .ZN(n11785) );
  NAND2_X1 U14367 ( .A1(n14317), .A2(n10307), .ZN(n11784) );
  NAND2_X1 U14368 ( .A1(n11785), .A2(n11784), .ZN(n11786) );
  XNOR2_X1 U14369 ( .A(n11786), .B(n11795), .ZN(n11791) );
  NAND2_X1 U14370 ( .A1(n14644), .A2(n10307), .ZN(n11789) );
  NAND2_X1 U14371 ( .A1(n11787), .A2(n14317), .ZN(n11788) );
  NAND2_X1 U14372 ( .A1(n11789), .A2(n11788), .ZN(n11790) );
  NOR2_X1 U14373 ( .A1(n11791), .A2(n11790), .ZN(n11792) );
  AOI21_X1 U14374 ( .B1(n11791), .B2(n11790), .A(n11792), .ZN(n13914) );
  INV_X1 U14375 ( .A(n11792), .ZN(n11793) );
  OAI22_X1 U14376 ( .A1(n14098), .A2(n11794), .B1(n14097), .B2(n11798), .ZN(
        n11796) );
  XNOR2_X1 U14377 ( .A(n11796), .B(n11795), .ZN(n11800) );
  OAI22_X1 U14378 ( .A1(n14098), .A2(n11798), .B1(n14097), .B2(n11797), .ZN(
        n11799) );
  XNOR2_X1 U14379 ( .A(n11800), .B(n11799), .ZN(n11801) );
  AOI22_X1 U14380 ( .A1(n14064), .A2(n14317), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11803) );
  NAND2_X1 U14381 ( .A1(n14023), .A2(n14315), .ZN(n11802) );
  OAI211_X1 U14382 ( .C1(n14026), .C2(n11804), .A(n11803), .B(n11802), .ZN(
        n11805) );
  AOI21_X1 U14383 ( .B1(n14639), .B2(n9398), .A(n11805), .ZN(n11806) );
  XNOR2_X1 U14384 ( .A(n11984), .B(n11807), .ZN(n11816) );
  INV_X1 U14385 ( .A(n11816), .ZN(n11808) );
  NAND2_X1 U14386 ( .A1(n11808), .A2(n11920), .ZN(n11823) );
  INV_X1 U14387 ( .A(n11809), .ZN(n11810) );
  NAND4_X1 U14388 ( .A1(n11822), .A2(n11920), .A3(n11816), .A4(n11810), .ZN(
        n11821) );
  AOI22_X1 U14389 ( .A1(n12169), .A2(n11931), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11813) );
  NAND2_X1 U14390 ( .A1(n11811), .A2(n11938), .ZN(n11812) );
  OAI211_X1 U14391 ( .C1(n11814), .C2(n11933), .A(n11813), .B(n11812), .ZN(
        n11818) );
  NOR4_X1 U14392 ( .A1(n11816), .A2(n11940), .A3(n12169), .A4(n11815), .ZN(
        n11817) );
  AOI211_X1 U14393 ( .C1(n11819), .C2(n11904), .A(n11818), .B(n11817), .ZN(
        n11820) );
  OAI211_X1 U14394 ( .C1(n11823), .C2(n11822), .A(n11821), .B(n11820), .ZN(
        P3_U3160) );
  AOI211_X1 U14395 ( .C1(n11825), .C2(n11824), .A(n11940), .B(n6700), .ZN(
        n11826) );
  INV_X1 U14396 ( .A(n11826), .ZN(n11832) );
  NAND2_X1 U14397 ( .A1(n12464), .A2(n11931), .ZN(n11828) );
  OAI211_X1 U14398 ( .C1(n11829), .C2(n11933), .A(n11828), .B(n11827), .ZN(
        n11830) );
  AOI21_X1 U14399 ( .B1(n12467), .B2(n11938), .A(n11830), .ZN(n11831) );
  OAI211_X1 U14400 ( .C1(n11935), .C2(n12605), .A(n11832), .B(n11831), .ZN(
        P3_U3155) );
  AOI21_X1 U14401 ( .B1(n12320), .B2(n11834), .A(n11833), .ZN(n11839) );
  AOI22_X1 U14402 ( .A1(n12171), .A2(n11931), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11836) );
  NAND2_X1 U14403 ( .A1(n11938), .A2(n12339), .ZN(n11835) );
  OAI211_X1 U14404 ( .C1(n12335), .C2(n11933), .A(n11836), .B(n11835), .ZN(
        n11837) );
  AOI21_X1 U14405 ( .B1(n12338), .B2(n11904), .A(n11837), .ZN(n11838) );
  OAI21_X1 U14406 ( .B1(n11839), .B2(n11940), .A(n11838), .ZN(P3_U3156) );
  OAI21_X1 U14407 ( .B1(n11841), .B2(n11840), .A(n11889), .ZN(n11842) );
  NAND2_X1 U14408 ( .A1(n11842), .A2(n11920), .ZN(n11846) );
  AND2_X1 U14409 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12269) );
  AOI21_X1 U14410 ( .B1(n12172), .B2(n11893), .A(n12269), .ZN(n11843) );
  OAI21_X1 U14411 ( .B1(n12382), .B2(n11895), .A(n11843), .ZN(n11844) );
  AOI21_X1 U14412 ( .B1(n12386), .B2(n11938), .A(n11844), .ZN(n11845) );
  OAI211_X1 U14413 ( .C1(n12527), .C2(n11935), .A(n11846), .B(n11845), .ZN(
        P3_U3159) );
  AOI21_X1 U14414 ( .B1(n11890), .B2(n11848), .A(n11847), .ZN(n11849) );
  OAI21_X1 U14415 ( .B1(n11850), .B2(n11849), .A(n11920), .ZN(n11854) );
  AOI22_X1 U14416 ( .A1(n12172), .A2(n11931), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11851) );
  OAI21_X1 U14417 ( .B1(n12360), .B2(n11933), .A(n11851), .ZN(n11852) );
  AOI21_X1 U14418 ( .B1(n12361), .B2(n11938), .A(n11852), .ZN(n11853) );
  OAI211_X1 U14419 ( .C1(n12589), .C2(n11935), .A(n11854), .B(n11853), .ZN(
        P3_U3163) );
  AND3_X1 U14420 ( .A1(n11879), .A2(n11856), .A3(n11855), .ZN(n11857) );
  OAI21_X1 U14421 ( .B1(n11858), .B2(n11857), .A(n11920), .ZN(n11863) );
  AOI22_X1 U14422 ( .A1(n12170), .A2(n11931), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11859) );
  OAI21_X1 U14423 ( .B1(n11860), .B2(n11933), .A(n11859), .ZN(n11861) );
  AOI21_X1 U14424 ( .B1(n12309), .B2(n11938), .A(n11861), .ZN(n11862) );
  OAI211_X1 U14425 ( .C1(n12573), .C2(n11935), .A(n11863), .B(n11862), .ZN(
        P3_U3165) );
  XNOR2_X1 U14426 ( .A(n11865), .B(n11864), .ZN(n11870) );
  NAND2_X1 U14427 ( .A1(n11931), .A2(n12463), .ZN(n11866) );
  NAND2_X1 U14428 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12219)
         );
  OAI211_X1 U14429 ( .C1(n12405), .C2(n11933), .A(n11866), .B(n12219), .ZN(
        n11868) );
  NOR2_X1 U14430 ( .A1(n12539), .A2(n11935), .ZN(n11867) );
  AOI211_X1 U14431 ( .C1(n12437), .C2(n11938), .A(n11868), .B(n11867), .ZN(
        n11869) );
  OAI21_X1 U14432 ( .B1(n11870), .B2(n11940), .A(n11869), .ZN(P3_U3166) );
  XOR2_X1 U14433 ( .A(n11872), .B(n11871), .Z(n11873) );
  NAND2_X1 U14434 ( .A1(n11873), .A2(n11920), .ZN(n11877) );
  NAND2_X1 U14435 ( .A1(n11931), .A2(n12452), .ZN(n11874) );
  NAND2_X1 U14436 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14908)
         );
  OAI211_X1 U14437 ( .C1(n12382), .C2(n11933), .A(n11874), .B(n14908), .ZN(
        n11875) );
  AOI21_X1 U14438 ( .B1(n11938), .B2(n12417), .A(n11875), .ZN(n11876) );
  OAI211_X1 U14439 ( .C1(n11935), .C2(n12535), .A(n11877), .B(n11876), .ZN(
        P3_U3168) );
  INV_X1 U14440 ( .A(n11878), .ZN(n12577) );
  INV_X1 U14441 ( .A(n11879), .ZN(n11883) );
  NOR3_X1 U14442 ( .A1(n11881), .A2(n11833), .A3(n11880), .ZN(n11882) );
  OAI21_X1 U14443 ( .B1(n11883), .B2(n11882), .A(n11920), .ZN(n11887) );
  AOI22_X1 U14444 ( .A1(n12321), .A2(n11893), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11884) );
  OAI21_X1 U14445 ( .B1(n12349), .B2(n11895), .A(n11884), .ZN(n11885) );
  AOI21_X1 U14446 ( .B1(n12324), .B2(n11938), .A(n11885), .ZN(n11886) );
  OAI211_X1 U14447 ( .C1(n12577), .C2(n11935), .A(n11887), .B(n11886), .ZN(
        P3_U3169) );
  AND2_X1 U14448 ( .A1(n11889), .A2(n11888), .ZN(n11892) );
  OAI211_X1 U14449 ( .C1(n11892), .C2(n11891), .A(n11920), .B(n11890), .ZN(
        n11898) );
  AOI22_X1 U14450 ( .A1(n11893), .A2(n12372), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11894) );
  OAI21_X1 U14451 ( .B1(n12407), .B2(n11895), .A(n11894), .ZN(n11896) );
  AOI21_X1 U14452 ( .B1(n12375), .B2(n11938), .A(n11896), .ZN(n11897) );
  OAI211_X1 U14453 ( .C1(n12593), .C2(n11935), .A(n11898), .B(n11897), .ZN(
        P3_U3173) );
  AOI21_X1 U14454 ( .B1(n12171), .B2(n11900), .A(n11899), .ZN(n11907) );
  NAND2_X1 U14455 ( .A1(n11938), .A2(n12350), .ZN(n11902) );
  AOI22_X1 U14456 ( .A1(n11931), .A2(n12372), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11901) );
  OAI211_X1 U14457 ( .C1(n12349), .C2(n11933), .A(n11902), .B(n11901), .ZN(
        n11903) );
  AOI21_X1 U14458 ( .B1(n11905), .B2(n11904), .A(n11903), .ZN(n11906) );
  OAI21_X1 U14459 ( .B1(n11907), .B2(n11940), .A(n11906), .ZN(P3_U3175) );
  XNOR2_X1 U14460 ( .A(n11909), .B(n11908), .ZN(n11914) );
  NAND2_X1 U14461 ( .A1(n11931), .A2(n12434), .ZN(n11910) );
  NAND2_X1 U14462 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12246)
         );
  OAI211_X1 U14463 ( .C1(n12407), .C2(n11933), .A(n11910), .B(n12246), .ZN(
        n11912) );
  NOR2_X1 U14464 ( .A1(n12598), .A2(n11935), .ZN(n11911) );
  AOI211_X1 U14465 ( .C1(n12409), .C2(n11938), .A(n11912), .B(n11911), .ZN(
        n11913) );
  OAI21_X1 U14466 ( .B1(n11914), .B2(n11940), .A(n11913), .ZN(P3_U3178) );
  NAND2_X1 U14467 ( .A1(n11916), .A2(n11915), .ZN(n11918) );
  NAND2_X1 U14468 ( .A1(n11918), .A2(n11919), .ZN(n11917) );
  OAI21_X1 U14469 ( .B1(n11919), .B2(n11918), .A(n11917), .ZN(n11921) );
  NAND2_X1 U14470 ( .A1(n11921), .A2(n11920), .ZN(n11926) );
  AOI22_X1 U14471 ( .A1(n12321), .A2(n11931), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11922) );
  OAI21_X1 U14472 ( .B1(n11923), .B2(n11933), .A(n11922), .ZN(n11924) );
  AOI21_X1 U14473 ( .B1(n12291), .B2(n11938), .A(n11924), .ZN(n11925) );
  OAI211_X1 U14474 ( .C1(n11927), .C2(n11935), .A(n11926), .B(n11925), .ZN(
        P3_U3180) );
  XNOR2_X1 U14475 ( .A(n11928), .B(n12463), .ZN(n11929) );
  XNOR2_X1 U14476 ( .A(n11930), .B(n11929), .ZN(n11941) );
  NAND2_X1 U14477 ( .A1(n11931), .A2(n12478), .ZN(n11932) );
  NAND2_X1 U14478 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12188)
         );
  OAI211_X1 U14479 ( .C1(n11934), .C2(n11933), .A(n11932), .B(n12188), .ZN(
        n11937) );
  NOR2_X1 U14480 ( .A1(n12543), .A2(n11935), .ZN(n11936) );
  AOI211_X1 U14481 ( .C1(n12447), .C2(n11938), .A(n11937), .B(n11936), .ZN(
        n11939) );
  OAI21_X1 U14482 ( .B1(n11941), .B2(n11940), .A(n11939), .ZN(P3_U3181) );
  INV_X1 U14483 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14742) );
  AND2_X1 U14484 ( .A1(n14742), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11942) );
  OAI22_X1 U14485 ( .A1(n11943), .A2(n11942), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n14742), .ZN(n11945) );
  XNOR2_X1 U14486 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11944) );
  XNOR2_X1 U14487 ( .A(n11945), .B(n11944), .ZN(n12618) );
  NAND2_X1 U14488 ( .A1(n12618), .A2(n11948), .ZN(n11947) );
  INV_X1 U14489 ( .A(SI_31_), .ZN(n12624) );
  OR2_X1 U14490 ( .A1(n11951), .A2(n12624), .ZN(n11946) );
  INV_X1 U14491 ( .A(n12563), .ZN(n12287) );
  NAND2_X1 U14492 ( .A1(n11949), .A2(n11948), .ZN(n11953) );
  OR2_X1 U14493 ( .A1(n8518), .A2(n11950), .ZN(n11952) );
  NAND2_X1 U14494 ( .A1(n11953), .A2(n11952), .ZN(n11957) );
  INV_X1 U14495 ( .A(n11958), .ZN(n12167) );
  AOI22_X1 U14496 ( .A1(n12563), .A2(n12284), .B1(n12569), .B2(n12167), .ZN(
        n12146) );
  NAND2_X1 U14497 ( .A1(n11955), .A2(n11954), .ZN(n11960) );
  OR2_X1 U14498 ( .A1(n12563), .A2(n12284), .ZN(n12145) );
  AOI21_X1 U14499 ( .B1(n11958), .B2(n11957), .A(n11956), .ZN(n11959) );
  OAI211_X1 U14500 ( .C1(n12569), .C2(n11961), .A(n11960), .B(n12144), .ZN(
        n11962) );
  OAI21_X1 U14501 ( .B1(n12287), .B2(n12146), .A(n11962), .ZN(n11963) );
  XNOR2_X1 U14502 ( .A(n11963), .B(n12268), .ZN(n12158) );
  INV_X1 U14503 ( .A(n12334), .ZN(n12329) );
  NAND2_X1 U14504 ( .A1(n12113), .A2(n12117), .ZN(n12345) );
  AND2_X1 U14505 ( .A1(n11965), .A2(n11964), .ZN(n12357) );
  INV_X1 U14506 ( .A(n12357), .ZN(n12355) );
  NOR4_X1 U14507 ( .A1(n11968), .A2(n6966), .A3(n11967), .A4(n11966), .ZN(
        n11970) );
  NAND4_X1 U14508 ( .A1(n11970), .A2(n11969), .A3(n12012), .A4(n12038), .ZN(
        n11973) );
  INV_X1 U14509 ( .A(n12050), .ZN(n12045) );
  NAND4_X1 U14510 ( .A1(n12027), .A2(n12008), .A3(n11971), .A4(n12032), .ZN(
        n11972) );
  NOR4_X1 U14511 ( .A1(n11973), .A2(n7607), .A3(n12045), .A4(n11972), .ZN(
        n11974) );
  INV_X1 U14512 ( .A(n12476), .ZN(n12472) );
  NAND4_X1 U14513 ( .A1(n11974), .A2(n12445), .A3(n12065), .A4(n12472), .ZN(
        n11975) );
  NOR4_X1 U14514 ( .A1(n12398), .A2(n11975), .A3(n12420), .A4(n12432), .ZN(
        n11976) );
  INV_X1 U14515 ( .A(n12370), .ZN(n12090) );
  NAND4_X1 U14516 ( .A1(n12355), .A2(n12392), .A3(n11976), .A4(n12090), .ZN(
        n11977) );
  NOR4_X1 U14517 ( .A1(n12318), .A2(n12329), .A3(n12345), .A4(n11977), .ZN(
        n11978) );
  NAND3_X1 U14518 ( .A1(n12132), .A2(n11978), .A3(n12301), .ZN(n11979) );
  NOR4_X1 U14519 ( .A1(n12141), .A2(n11984), .A3(n11983), .A4(n11979), .ZN(
        n11980) );
  NAND3_X1 U14520 ( .A1(n12144), .A2(n12146), .A3(n11980), .ZN(n11981) );
  XOR2_X1 U14521 ( .A(n12268), .B(n11981), .Z(n12154) );
  INV_X1 U14522 ( .A(n11982), .ZN(n11985) );
  OR2_X1 U14523 ( .A1(n11984), .A2(n11983), .ZN(n12134) );
  NOR2_X1 U14524 ( .A1(n12134), .A2(n12103), .ZN(n12138) );
  AOI21_X1 U14525 ( .B1(n11986), .B2(n11985), .A(n12138), .ZN(n12143) );
  NAND3_X1 U14526 ( .A1(n11987), .A2(n12163), .A3(n11988), .ZN(n11993) );
  INV_X1 U14527 ( .A(n11988), .ZN(n11989) );
  OAI211_X1 U14528 ( .C1(n11989), .C2(n11990), .A(n12129), .B(n11996), .ZN(
        n11992) );
  AOI22_X1 U14529 ( .A1(n11993), .A2(n11992), .B1(n11991), .B2(n11990), .ZN(
        n11994) );
  NOR2_X1 U14530 ( .A1(n11994), .A2(n11542), .ZN(n12001) );
  MUX2_X1 U14531 ( .A(n11996), .B(n11995), .S(n12129), .Z(n12000) );
  OAI21_X1 U14532 ( .B1(n11998), .B2(n11997), .A(n12010), .ZN(n11999) );
  AOI22_X1 U14533 ( .A1(n12001), .A2(n12000), .B1(n12103), .B2(n11999), .ZN(
        n12007) );
  INV_X1 U14534 ( .A(n12002), .ZN(n12006) );
  INV_X1 U14535 ( .A(n12003), .ZN(n12004) );
  OAI21_X1 U14536 ( .B1(n12006), .B2(n12004), .A(n12129), .ZN(n12005) );
  OAI21_X1 U14537 ( .B1(n12007), .B2(n12006), .A(n12005), .ZN(n12009) );
  OAI211_X1 U14538 ( .C1(n12103), .C2(n12010), .A(n12009), .B(n12008), .ZN(
        n12013) );
  NAND2_X1 U14539 ( .A1(n12025), .A2(n12011), .ZN(n12014) );
  AOI22_X1 U14540 ( .A1(n12013), .A2(n12012), .B1(n12129), .B2(n12014), .ZN(
        n12023) );
  INV_X1 U14541 ( .A(n12015), .ZN(n15480) );
  NOR3_X1 U14542 ( .A1(n12014), .A2(n12103), .A3(n15480), .ZN(n12017) );
  NOR2_X1 U14543 ( .A1(n12015), .A2(n12129), .ZN(n12016) );
  MUX2_X1 U14544 ( .A(n12017), .B(n12016), .S(n12179), .Z(n12022) );
  INV_X1 U14545 ( .A(n12024), .ZN(n12020) );
  INV_X1 U14546 ( .A(n12018), .ZN(n12019) );
  NOR2_X1 U14547 ( .A1(n12020), .A2(n12019), .ZN(n12021) );
  OAI22_X1 U14548 ( .A1(n12023), .A2(n12022), .B1(n12021), .B2(n12129), .ZN(
        n12028) );
  MUX2_X1 U14549 ( .A(n12025), .B(n12024), .S(n12129), .Z(n12026) );
  NAND3_X1 U14550 ( .A1(n12028), .A2(n12027), .A3(n12026), .ZN(n12033) );
  NAND2_X1 U14551 ( .A1(n12177), .A2(n15496), .ZN(n12029) );
  MUX2_X1 U14552 ( .A(n12030), .B(n12029), .S(n12129), .Z(n12031) );
  NAND3_X1 U14553 ( .A1(n12033), .A2(n12032), .A3(n12031), .ZN(n12039) );
  INV_X1 U14554 ( .A(n12034), .ZN(n15502) );
  NAND2_X1 U14555 ( .A1(n12176), .A2(n15502), .ZN(n12036) );
  MUX2_X1 U14556 ( .A(n12036), .B(n12035), .S(n12129), .Z(n12037) );
  NAND3_X1 U14557 ( .A1(n12039), .A2(n12038), .A3(n12037), .ZN(n12043) );
  MUX2_X1 U14558 ( .A(n12041), .B(n12040), .S(n12129), .Z(n12042) );
  AOI21_X1 U14559 ( .B1(n12043), .B2(n12042), .A(n7346), .ZN(n12048) );
  INV_X1 U14560 ( .A(n12044), .ZN(n12046) );
  AOI211_X1 U14561 ( .C1(n12173), .C2(n6739), .A(n12054), .B(n12047), .ZN(
        n12053) );
  INV_X1 U14562 ( .A(n12048), .ZN(n12051) );
  NAND3_X1 U14563 ( .A1(n12051), .A2(n12050), .A3(n12049), .ZN(n12052) );
  MUX2_X1 U14564 ( .A(n12055), .B(n12054), .S(n12129), .Z(n12056) );
  NOR2_X1 U14565 ( .A1(n12056), .A2(n12476), .ZN(n12061) );
  INV_X1 U14566 ( .A(n12061), .ZN(n12066) );
  NAND2_X1 U14567 ( .A1(n12058), .A2(n12057), .ZN(n12060) );
  AOI21_X1 U14568 ( .B1(n12061), .B2(n12060), .A(n12059), .ZN(n12062) );
  MUX2_X1 U14569 ( .A(n12063), .B(n12062), .S(n12129), .Z(n12064) );
  MUX2_X1 U14570 ( .A(n12068), .B(n6681), .S(n12129), .Z(n12069) );
  AOI21_X1 U14571 ( .B1(n12070), .B2(n12069), .A(n12450), .ZN(n12073) );
  AOI21_X1 U14572 ( .B1(n12078), .B2(n12071), .A(n12103), .ZN(n12072) );
  OAI21_X1 U14573 ( .B1(n12073), .B2(n12072), .A(n12074), .ZN(n12081) );
  INV_X1 U14574 ( .A(n12074), .ZN(n12077) );
  INV_X1 U14575 ( .A(n12075), .ZN(n12076) );
  OAI21_X1 U14576 ( .B1(n12077), .B2(n12076), .A(n12103), .ZN(n12080) );
  INV_X1 U14577 ( .A(n12078), .ZN(n12079) );
  AOI22_X1 U14578 ( .A1(n12081), .A2(n12080), .B1(n12079), .B2(n12103), .ZN(
        n12085) );
  INV_X1 U14579 ( .A(n12082), .ZN(n12086) );
  NOR3_X1 U14580 ( .A1(n12086), .A2(n12083), .A3(n12129), .ZN(n12094) );
  INV_X1 U14581 ( .A(n12101), .ZN(n12087) );
  MUX2_X1 U14582 ( .A(n12087), .B(n12086), .S(n12129), .Z(n12088) );
  INV_X1 U14583 ( .A(n12088), .ZN(n12089) );
  AND2_X1 U14584 ( .A1(n12090), .A2(n12089), .ZN(n12098) );
  NAND3_X1 U14585 ( .A1(n12091), .A2(n12402), .A3(n12098), .ZN(n12112) );
  INV_X1 U14586 ( .A(n12096), .ZN(n12092) );
  NOR2_X1 U14587 ( .A1(n12092), .A2(n12103), .ZN(n12102) );
  INV_X1 U14588 ( .A(n12093), .ZN(n12097) );
  INV_X1 U14589 ( .A(n12094), .ZN(n12095) );
  AOI21_X1 U14590 ( .B1(n12097), .B2(n12096), .A(n12095), .ZN(n12100) );
  INV_X1 U14591 ( .A(n12098), .ZN(n12099) );
  AOI211_X1 U14592 ( .C1(n12102), .C2(n12101), .A(n12100), .B(n12099), .ZN(
        n12108) );
  NOR2_X1 U14593 ( .A1(n12381), .A2(n12129), .ZN(n12106) );
  NOR2_X1 U14594 ( .A1(n12172), .A2(n12103), .ZN(n12105) );
  MUX2_X1 U14595 ( .A(n12106), .B(n12105), .S(n12104), .Z(n12107) );
  NOR3_X1 U14596 ( .A1(n12108), .A2(n12357), .A3(n12107), .ZN(n12111) );
  MUX2_X1 U14597 ( .A(n12109), .B(n6678), .S(n12129), .Z(n12110) );
  NOR2_X1 U14598 ( .A1(n12116), .A2(n7612), .ZN(n12114) );
  AOI22_X1 U14599 ( .A1(n12114), .A2(n12334), .B1(n12349), .B2(n12338), .ZN(
        n12115) );
  OAI21_X1 U14600 ( .B1(n12115), .B2(n12318), .A(n12120), .ZN(n12126) );
  INV_X1 U14601 ( .A(n12116), .ZN(n12118) );
  NAND3_X1 U14602 ( .A1(n12118), .A2(n12334), .A3(n12117), .ZN(n12124) );
  INV_X1 U14603 ( .A(n12119), .ZN(n12122) );
  OAI21_X1 U14604 ( .B1(n12122), .B2(n12121), .A(n12120), .ZN(n12123) );
  OAI21_X1 U14605 ( .B1(n12124), .B2(n12318), .A(n12123), .ZN(n12125) );
  NAND2_X1 U14606 ( .A1(n12573), .A2(n12129), .ZN(n12128) );
  OAI211_X1 U14607 ( .C1(n12321), .C2(n12129), .A(n12128), .B(n12127), .ZN(
        n12130) );
  NAND2_X1 U14608 ( .A1(n12133), .A2(n12132), .ZN(n12139) );
  INV_X1 U14609 ( .A(n12134), .ZN(n12136) );
  NAND3_X1 U14610 ( .A1(n12139), .A2(n12136), .A3(n12135), .ZN(n12142) );
  INV_X1 U14611 ( .A(n12144), .ZN(n12148) );
  INV_X1 U14612 ( .A(n12145), .ZN(n12147) );
  OAI22_X1 U14613 ( .A1(n12149), .A2(n12148), .B1(n12147), .B2(n12146), .ZN(
        n12150) );
  MUX2_X1 U14614 ( .A(n12152), .B(n12151), .S(n12150), .Z(n12153) );
  OAI21_X1 U14615 ( .B1(n12155), .B2(n12154), .A(n12153), .ZN(n12156) );
  AOI21_X1 U14616 ( .B1(n12158), .B2(n12157), .A(n12156), .ZN(n12166) );
  NAND4_X1 U14617 ( .A1(n12480), .A2(n12161), .A3(n12160), .A4(n12159), .ZN(
        n12162) );
  OAI211_X1 U14618 ( .C1(n12163), .C2(n12165), .A(n12162), .B(P3_B_REG_SCAN_IN), .ZN(n12164) );
  OAI21_X1 U14619 ( .B1(n12166), .B2(n12165), .A(n12164), .ZN(P3_U3296) );
  MUX2_X1 U14620 ( .A(n12167), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12181), .Z(
        P3_U3521) );
  MUX2_X1 U14621 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12168), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14622 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12169), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14623 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12306), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14624 ( .A(n12321), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12181), .Z(
        P3_U3516) );
  MUX2_X1 U14625 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12170), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14626 ( .A(n12320), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12181), .Z(
        P3_U3514) );
  MUX2_X1 U14627 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12171), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14628 ( .A(n12372), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12181), .Z(
        P3_U3512) );
  MUX2_X1 U14629 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12172), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14630 ( .A(n12422), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12181), .Z(
        P3_U3509) );
  MUX2_X1 U14631 ( .A(n12434), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12181), .Z(
        P3_U3508) );
  MUX2_X1 U14632 ( .A(n12452), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12181), .Z(
        P3_U3507) );
  MUX2_X1 U14633 ( .A(n12463), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12181), .Z(
        P3_U3506) );
  MUX2_X1 U14634 ( .A(n12478), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12181), .Z(
        P3_U3505) );
  MUX2_X1 U14635 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12464), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14636 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12481), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14637 ( .A(n12173), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12181), .Z(
        P3_U3502) );
  MUX2_X1 U14638 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12174), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14639 ( .A(n12175), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12181), .Z(
        P3_U3500) );
  MUX2_X1 U14640 ( .A(n12176), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12181), .Z(
        P3_U3499) );
  MUX2_X1 U14641 ( .A(n12177), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12181), .Z(
        P3_U3498) );
  MUX2_X1 U14642 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12178), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14643 ( .A(n12179), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12181), .Z(
        P3_U3495) );
  MUX2_X1 U14644 ( .A(n12180), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12181), .Z(
        P3_U3493) );
  MUX2_X1 U14645 ( .A(n12182), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12181), .Z(
        P3_U3491) );
  INV_X1 U14646 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12197) );
  AOI21_X1 U14647 ( .B1(n12197), .B2(n12185), .A(n12208), .ZN(n12203) );
  OAI21_X1 U14648 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12187), .A(n12223), 
        .ZN(n12191) );
  INV_X1 U14649 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14854) );
  INV_X1 U14650 ( .A(n12222), .ZN(n12196) );
  NAND2_X1 U14651 ( .A1(n14907), .A2(n12196), .ZN(n12189) );
  OAI211_X1 U14652 ( .C1(n14854), .C2(n14910), .A(n12189), .B(n12188), .ZN(
        n12190) );
  AOI21_X1 U14653 ( .B1(n12191), .B2(n15461), .A(n12190), .ZN(n12202) );
  MUX2_X1 U14654 ( .A(n12193), .B(n12192), .S(n12275), .Z(n12194) );
  NAND2_X1 U14655 ( .A1(n12195), .A2(n12194), .ZN(n12214) );
  XNOR2_X1 U14656 ( .A(n12214), .B(n12196), .ZN(n12199) );
  MUX2_X1 U14657 ( .A(n12197), .B(n6753), .S(n12275), .Z(n12198) );
  NAND2_X1 U14658 ( .A1(n12199), .A2(n12198), .ZN(n12216) );
  OAI21_X1 U14659 ( .B1(n12199), .B2(n12198), .A(n12216), .ZN(n12200) );
  NAND2_X1 U14660 ( .A1(n12200), .A2(n12280), .ZN(n12201) );
  OAI211_X1 U14661 ( .C1(n12203), .C2(n15465), .A(n12202), .B(n12201), .ZN(
        P3_U3197) );
  INV_X1 U14662 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12204) );
  NAND2_X1 U14663 ( .A1(n12249), .A2(n12204), .ZN(n12206) );
  NAND2_X1 U14664 ( .A1(n12220), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12205) );
  AND2_X1 U14665 ( .A1(n12206), .A2(n12205), .ZN(n12211) );
  INV_X1 U14666 ( .A(n12232), .ZN(n12209) );
  AOI21_X1 U14667 ( .B1(n12211), .B2(n12210), .A(n12209), .ZN(n12230) );
  MUX2_X1 U14668 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12275), .Z(n12212) );
  NAND2_X1 U14669 ( .A1(n12212), .A2(n12249), .ZN(n12236) );
  INV_X1 U14670 ( .A(n12212), .ZN(n12213) );
  NAND2_X1 U14671 ( .A1(n12213), .A2(n12220), .ZN(n12238) );
  NAND2_X1 U14672 ( .A1(n12236), .A2(n12238), .ZN(n12217) );
  OR2_X1 U14673 ( .A1(n12214), .A2(n12222), .ZN(n12215) );
  NAND2_X1 U14674 ( .A1(n12216), .A2(n12215), .ZN(n12237) );
  XOR2_X1 U14675 ( .A(n12217), .B(n12237), .Z(n12228) );
  NAND2_X1 U14676 ( .A1(n15458), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n12218) );
  OAI211_X1 U14677 ( .C1(n15452), .C2(n12249), .A(n12219), .B(n12218), .ZN(
        n12227) );
  XNOR2_X1 U14678 ( .A(n12220), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12247) );
  NAND2_X1 U14679 ( .A1(n12222), .A2(n12221), .ZN(n12224) );
  XOR2_X1 U14680 ( .A(n12247), .B(n12248), .Z(n12225) );
  NOR2_X1 U14681 ( .A1(n12225), .A2(n12258), .ZN(n12226) );
  AOI211_X1 U14682 ( .C1(n12228), .C2(n12280), .A(n12227), .B(n12226), .ZN(
        n12229) );
  OAI21_X1 U14683 ( .B1(n12230), .B2(n15465), .A(n12229), .ZN(P3_U3198) );
  NAND2_X1 U14684 ( .A1(n12249), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12231) );
  INV_X1 U14685 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14903) );
  NAND2_X1 U14686 ( .A1(n12273), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12264) );
  OAI21_X1 U14687 ( .B1(n12273), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12264), 
        .ZN(n12234) );
  NAND2_X1 U14688 ( .A1(n12237), .A2(n12236), .ZN(n12239) );
  NAND2_X1 U14689 ( .A1(n12239), .A2(n12238), .ZN(n14914) );
  MUX2_X1 U14690 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12275), .Z(n12240) );
  XNOR2_X1 U14691 ( .A(n12240), .B(n12252), .ZN(n14915) );
  NAND2_X1 U14692 ( .A1(n12240), .A2(n12252), .ZN(n12241) );
  NAND2_X1 U14693 ( .A1(n14912), .A2(n12241), .ZN(n12274) );
  XNOR2_X1 U14694 ( .A(n12274), .B(n12267), .ZN(n12244) );
  INV_X1 U14695 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12242) );
  INV_X1 U14696 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12530) );
  MUX2_X1 U14697 ( .A(n12242), .B(n12530), .S(n12275), .Z(n12243) );
  NAND2_X1 U14698 ( .A1(n12244), .A2(n12243), .ZN(n12272) );
  OAI21_X1 U14699 ( .B1(n12244), .B2(n12243), .A(n12272), .ZN(n12262) );
  NAND2_X1 U14700 ( .A1(n15458), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12245) );
  OAI211_X1 U14701 ( .C1(n15452), .C2(n12273), .A(n12246), .B(n12245), .ZN(
        n12261) );
  NAND2_X1 U14702 ( .A1(n12249), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12250) );
  NAND2_X1 U14703 ( .A1(n12253), .A2(n12252), .ZN(n12257) );
  XNOR2_X1 U14704 ( .A(n12253), .B(n14906), .ZN(n14905) );
  XNOR2_X1 U14705 ( .A(n12267), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12255) );
  INV_X1 U14706 ( .A(n12255), .ZN(n12256) );
  NAND3_X1 U14707 ( .A1(n12257), .A2(n14904), .A3(n12256), .ZN(n12259) );
  AOI21_X1 U14708 ( .B1(n12266), .B2(n12259), .A(n12258), .ZN(n12260) );
  AOI211_X1 U14709 ( .C1(n12280), .C2(n12262), .A(n12261), .B(n12260), .ZN(
        n12263) );
  XNOR2_X1 U14710 ( .A(n12268), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12277) );
  XNOR2_X1 U14711 ( .A(n12268), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12276) );
  NAND2_X1 U14712 ( .A1(n14907), .A2(n12268), .ZN(n12271) );
  AOI21_X1 U14713 ( .B1(n15458), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n12269), 
        .ZN(n12270) );
  OAI21_X1 U14714 ( .B1(n12274), .B2(n12273), .A(n12272), .ZN(n12279) );
  MUX2_X1 U14715 ( .A(n12277), .B(n12276), .S(n12275), .Z(n12278) );
  XNOR2_X1 U14716 ( .A(n12279), .B(n12278), .ZN(n12281) );
  NAND2_X1 U14717 ( .A1(n12281), .A2(n12280), .ZN(n12282) );
  AOI21_X1 U14718 ( .B1(n12285), .B2(n12495), .A(n12486), .ZN(n12288) );
  AOI21_X1 U14719 ( .B1(n12486), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12288), 
        .ZN(n12286) );
  OAI21_X1 U14720 ( .B1(n12287), .B2(n12488), .A(n12286), .ZN(P3_U3202) );
  AOI21_X1 U14721 ( .B1(n12486), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12288), 
        .ZN(n12289) );
  OAI21_X1 U14722 ( .B1(n12569), .B2(n12488), .A(n12289), .ZN(P3_U3203) );
  NAND2_X1 U14723 ( .A1(n12290), .A2(n12490), .ZN(n12297) );
  INV_X1 U14724 ( .A(n12291), .ZN(n12293) );
  OAI22_X1 U14725 ( .A1(n12293), .A2(n12387), .B1(n12490), .B2(n12292), .ZN(
        n12294) );
  AOI21_X1 U14726 ( .B1(n12295), .B2(n12438), .A(n12294), .ZN(n12296) );
  OAI211_X1 U14727 ( .C1(n12299), .C2(n12298), .A(n12297), .B(n12296), .ZN(
        P3_U3207) );
  OAI21_X1 U14728 ( .B1(n12302), .B2(n12301), .A(n12300), .ZN(n12502) );
  INV_X1 U14729 ( .A(n12502), .ZN(n12313) );
  OAI211_X1 U14730 ( .C1(n12305), .C2(n12304), .A(n12303), .B(n12474), .ZN(
        n12308) );
  NAND2_X1 U14731 ( .A1(n12306), .A2(n12479), .ZN(n12307) );
  OAI211_X1 U14732 ( .C1(n12335), .C2(n12406), .A(n12308), .B(n12307), .ZN(
        n12501) );
  AOI22_X1 U14733 ( .A1(n12309), .A2(n12485), .B1(n12486), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12310) );
  OAI21_X1 U14734 ( .B1(n12573), .B2(n12488), .A(n12310), .ZN(n12311) );
  AOI21_X1 U14735 ( .B1(n12501), .B2(n12490), .A(n12311), .ZN(n12312) );
  OAI21_X1 U14736 ( .B1(n12313), .B2(n12493), .A(n12312), .ZN(P3_U3208) );
  OAI21_X1 U14737 ( .B1(n12316), .B2(n12315), .A(n12314), .ZN(n12506) );
  INV_X1 U14738 ( .A(n12506), .ZN(n12328) );
  OAI211_X1 U14739 ( .C1(n12319), .C2(n12318), .A(n12317), .B(n12474), .ZN(
        n12323) );
  AOI22_X1 U14740 ( .A1(n12321), .A2(n12479), .B1(n12480), .B2(n12320), .ZN(
        n12322) );
  NAND2_X1 U14741 ( .A1(n12323), .A2(n12322), .ZN(n12505) );
  AOI22_X1 U14742 ( .A1(n12485), .A2(n12324), .B1(n12486), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12325) );
  OAI21_X1 U14743 ( .B1(n12577), .B2(n12488), .A(n12325), .ZN(n12326) );
  AOI21_X1 U14744 ( .B1(n12505), .B2(n12490), .A(n12326), .ZN(n12327) );
  OAI21_X1 U14745 ( .B1(n12328), .B2(n12493), .A(n12327), .ZN(P3_U3209) );
  XNOR2_X1 U14746 ( .A(n12330), .B(n12329), .ZN(n12509) );
  INV_X1 U14747 ( .A(n12509), .ZN(n12343) );
  INV_X1 U14748 ( .A(n12331), .ZN(n12332) );
  AOI211_X1 U14749 ( .C1(n12334), .C2(n12333), .A(n12404), .B(n12332), .ZN(
        n12337) );
  OAI22_X1 U14750 ( .A1(n12335), .A2(n12408), .B1(n12360), .B2(n12406), .ZN(
        n12336) );
  OR2_X1 U14751 ( .A1(n12337), .A2(n12336), .ZN(n12508) );
  INV_X1 U14752 ( .A(n12338), .ZN(n12581) );
  AOI22_X1 U14753 ( .A1(n12486), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12485), 
        .B2(n12339), .ZN(n12340) );
  OAI21_X1 U14754 ( .B1(n12581), .B2(n12488), .A(n12340), .ZN(n12341) );
  AOI21_X1 U14755 ( .B1(n12508), .B2(n12490), .A(n12341), .ZN(n12342) );
  OAI21_X1 U14756 ( .B1(n12493), .B2(n12343), .A(n12342), .ZN(P3_U3210) );
  XNOR2_X1 U14757 ( .A(n12344), .B(n12345), .ZN(n12513) );
  INV_X1 U14758 ( .A(n12513), .ZN(n12354) );
  XNOR2_X1 U14759 ( .A(n12346), .B(n12345), .ZN(n12347) );
  OAI222_X1 U14760 ( .A1(n12408), .A2(n12349), .B1(n12406), .B2(n12348), .C1(
        n12347), .C2(n12404), .ZN(n12512) );
  AOI22_X1 U14761 ( .A1(n12486), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12485), 
        .B2(n12350), .ZN(n12351) );
  OAI21_X1 U14762 ( .B1(n12585), .B2(n12488), .A(n12351), .ZN(n12352) );
  AOI21_X1 U14763 ( .B1(n12512), .B2(n12490), .A(n12352), .ZN(n12353) );
  OAI21_X1 U14764 ( .B1(n12493), .B2(n12354), .A(n12353), .ZN(P3_U3211) );
  XNOR2_X1 U14765 ( .A(n12356), .B(n12355), .ZN(n12517) );
  INV_X1 U14766 ( .A(n12517), .ZN(n12365) );
  XNOR2_X1 U14767 ( .A(n12358), .B(n12357), .ZN(n12359) );
  OAI222_X1 U14768 ( .A1(n12408), .A2(n12360), .B1(n12406), .B2(n12381), .C1(
        n12404), .C2(n12359), .ZN(n12516) );
  AOI22_X1 U14769 ( .A1(n12486), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12485), 
        .B2(n12361), .ZN(n12362) );
  OAI21_X1 U14770 ( .B1(n12589), .B2(n12488), .A(n12362), .ZN(n12363) );
  AOI21_X1 U14771 ( .B1(n12516), .B2(n12490), .A(n12363), .ZN(n12364) );
  OAI21_X1 U14772 ( .B1(n12493), .B2(n12365), .A(n12364), .ZN(P3_U3212) );
  AOI21_X1 U14773 ( .B1(n12370), .B2(n12368), .A(n12367), .ZN(n12521) );
  INV_X1 U14774 ( .A(n12521), .ZN(n12379) );
  OAI211_X1 U14775 ( .C1(n12371), .C2(n12370), .A(n12369), .B(n12474), .ZN(
        n12374) );
  NAND2_X1 U14776 ( .A1(n12372), .A2(n12479), .ZN(n12373) );
  OAI211_X1 U14777 ( .C1(n12407), .C2(n12406), .A(n12374), .B(n12373), .ZN(
        n12520) );
  AOI22_X1 U14778 ( .A1(n12486), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n12485), 
        .B2(n12375), .ZN(n12376) );
  OAI21_X1 U14779 ( .B1(n12593), .B2(n12488), .A(n12376), .ZN(n12377) );
  AOI21_X1 U14780 ( .B1(n12520), .B2(n12490), .A(n12377), .ZN(n12378) );
  OAI21_X1 U14781 ( .B1(n12493), .B2(n12379), .A(n12378), .ZN(P3_U3213) );
  AOI21_X1 U14782 ( .B1(n12380), .B2(n12392), .A(n12404), .ZN(n12385) );
  OAI22_X1 U14783 ( .A1(n12382), .A2(n12406), .B1(n12381), .B2(n12408), .ZN(
        n12383) );
  AOI21_X1 U14784 ( .B1(n12385), .B2(n12384), .A(n12383), .ZN(n12526) );
  INV_X1 U14785 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13744) );
  INV_X1 U14786 ( .A(n12386), .ZN(n12388) );
  OAI22_X1 U14787 ( .A1(n12490), .A2(n13744), .B1(n12388), .B2(n12387), .ZN(
        n12389) );
  AOI21_X1 U14788 ( .B1(n12390), .B2(n12438), .A(n12389), .ZN(n12395) );
  OAI21_X1 U14789 ( .B1(n12393), .B2(n12392), .A(n12391), .ZN(n12524) );
  NAND2_X1 U14790 ( .A1(n12524), .A2(n12457), .ZN(n12394) );
  OAI211_X1 U14791 ( .C1(n12526), .C2(n12486), .A(n12395), .B(n12394), .ZN(
        P3_U3214) );
  AOI21_X1 U14792 ( .B1(n12398), .B2(n12397), .A(n12396), .ZN(n12529) );
  INV_X1 U14793 ( .A(n12529), .ZN(n12413) );
  INV_X1 U14794 ( .A(n12399), .ZN(n12400) );
  AOI21_X1 U14795 ( .B1(n12402), .B2(n12401), .A(n12400), .ZN(n12403) );
  OAI222_X1 U14796 ( .A1(n12408), .A2(n12407), .B1(n12406), .B2(n12405), .C1(
        n12404), .C2(n12403), .ZN(n12528) );
  AOI22_X1 U14797 ( .A1(n12486), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n12485), 
        .B2(n12409), .ZN(n12410) );
  OAI21_X1 U14798 ( .B1(n12598), .B2(n12488), .A(n12410), .ZN(n12411) );
  AOI21_X1 U14799 ( .B1(n12528), .B2(n12490), .A(n12411), .ZN(n12412) );
  OAI21_X1 U14800 ( .B1(n12493), .B2(n12413), .A(n12412), .ZN(P3_U3215) );
  OAI21_X1 U14801 ( .B1(n12416), .B2(n12415), .A(n12414), .ZN(n12532) );
  AOI22_X1 U14802 ( .A1(n12486), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12485), 
        .B2(n12417), .ZN(n12418) );
  OAI21_X1 U14803 ( .B1(n12535), .B2(n12488), .A(n12418), .ZN(n12426) );
  OAI211_X1 U14804 ( .C1(n12421), .C2(n12420), .A(n12419), .B(n12474), .ZN(
        n12424) );
  AOI22_X1 U14805 ( .A1(n12480), .A2(n12452), .B1(n12422), .B2(n12479), .ZN(
        n12423) );
  NOR2_X1 U14806 ( .A1(n12534), .A2(n12486), .ZN(n12425) );
  AOI211_X1 U14807 ( .C1(n12457), .C2(n12532), .A(n12426), .B(n12425), .ZN(
        n12427) );
  INV_X1 U14808 ( .A(n12427), .ZN(P3_U3216) );
  OAI21_X1 U14809 ( .B1(n12430), .B2(n12429), .A(n12428), .ZN(n12536) );
  OAI211_X1 U14810 ( .C1(n12433), .C2(n12432), .A(n12431), .B(n12474), .ZN(
        n12436) );
  AOI22_X1 U14811 ( .A1(n12480), .A2(n12463), .B1(n12434), .B2(n12479), .ZN(
        n12435) );
  AOI22_X1 U14812 ( .A1(n12486), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12485), 
        .B2(n12437), .ZN(n12441) );
  NAND2_X1 U14813 ( .A1(n12439), .A2(n12438), .ZN(n12440) );
  OAI211_X1 U14814 ( .C1(n12538), .C2(n12486), .A(n12441), .B(n12440), .ZN(
        n12442) );
  AOI21_X1 U14815 ( .B1(n12457), .B2(n12536), .A(n12442), .ZN(n12443) );
  INV_X1 U14816 ( .A(n12443), .ZN(P3_U3217) );
  OAI21_X1 U14817 ( .B1(n12446), .B2(n12445), .A(n12444), .ZN(n12540) );
  AOI22_X1 U14818 ( .A1(n12486), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12485), 
        .B2(n12447), .ZN(n12448) );
  OAI21_X1 U14819 ( .B1(n12543), .B2(n12488), .A(n12448), .ZN(n12456) );
  OAI211_X1 U14820 ( .C1(n12451), .C2(n12450), .A(n12449), .B(n12474), .ZN(
        n12454) );
  AOI22_X1 U14821 ( .A1(n12480), .A2(n12478), .B1(n12452), .B2(n12479), .ZN(
        n12453) );
  NOR2_X1 U14822 ( .A1(n12542), .A2(n12486), .ZN(n12455) );
  AOI211_X1 U14823 ( .C1(n12457), .C2(n12540), .A(n12456), .B(n12455), .ZN(
        n12458) );
  INV_X1 U14824 ( .A(n12458), .ZN(P3_U3218) );
  XNOR2_X1 U14825 ( .A(n12459), .B(n12461), .ZN(n12545) );
  INV_X1 U14826 ( .A(n12545), .ZN(n12471) );
  OAI211_X1 U14827 ( .C1(n12462), .C2(n12461), .A(n12460), .B(n12474), .ZN(
        n12466) );
  AOI22_X1 U14828 ( .A1(n12464), .A2(n12480), .B1(n12479), .B2(n12463), .ZN(
        n12465) );
  NAND2_X1 U14829 ( .A1(n12466), .A2(n12465), .ZN(n12544) );
  AOI22_X1 U14830 ( .A1(n12486), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n12485), 
        .B2(n12467), .ZN(n12468) );
  OAI21_X1 U14831 ( .B1(n12605), .B2(n12488), .A(n12468), .ZN(n12469) );
  AOI21_X1 U14832 ( .B1(n12544), .B2(n12490), .A(n12469), .ZN(n12470) );
  OAI21_X1 U14833 ( .B1(n12471), .B2(n12493), .A(n12470), .ZN(P3_U3219) );
  XNOR2_X1 U14834 ( .A(n12473), .B(n12472), .ZN(n12549) );
  INV_X1 U14835 ( .A(n12549), .ZN(n12492) );
  OAI211_X1 U14836 ( .C1(n12477), .C2(n12476), .A(n12475), .B(n12474), .ZN(
        n12483) );
  AOI22_X1 U14837 ( .A1(n12481), .A2(n12480), .B1(n12479), .B2(n12478), .ZN(
        n12482) );
  NAND2_X1 U14838 ( .A1(n12483), .A2(n12482), .ZN(n12548) );
  AOI22_X1 U14839 ( .A1(n12486), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n12485), 
        .B2(n12484), .ZN(n12487) );
  OAI21_X1 U14840 ( .B1(n12609), .B2(n12488), .A(n12487), .ZN(n12489) );
  AOI21_X1 U14841 ( .B1(n12548), .B2(n12490), .A(n12489), .ZN(n12491) );
  OAI21_X1 U14842 ( .B1(n12493), .B2(n12492), .A(n12491), .ZN(P3_U3220) );
  INV_X1 U14843 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12497) );
  NAND2_X1 U14844 ( .A1(n12563), .A2(n12494), .ZN(n12496) );
  INV_X1 U14845 ( .A(n12495), .ZN(n12564) );
  NAND2_X1 U14846 ( .A1(n12564), .A2(n15540), .ZN(n12499) );
  OAI211_X1 U14847 ( .C1(n15540), .C2(n12497), .A(n12496), .B(n12499), .ZN(
        P3_U3490) );
  NAND2_X1 U14848 ( .A1(n15538), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12498) );
  OAI211_X1 U14849 ( .C1(n12569), .C2(n12556), .A(n12499), .B(n12498), .ZN(
        P3_U3489) );
  INV_X1 U14850 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12503) );
  AOI21_X1 U14851 ( .B1(n15518), .B2(n12502), .A(n12501), .ZN(n12570) );
  MUX2_X1 U14852 ( .A(n12503), .B(n12570), .S(n15540), .Z(n12504) );
  OAI21_X1 U14853 ( .B1(n12573), .B2(n12556), .A(n12504), .ZN(P3_U3484) );
  INV_X1 U14854 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13740) );
  AOI21_X1 U14855 ( .B1(n15518), .B2(n12506), .A(n12505), .ZN(n12574) );
  MUX2_X1 U14856 ( .A(n13740), .B(n12574), .S(n15540), .Z(n12507) );
  OAI21_X1 U14857 ( .B1(n12577), .B2(n12556), .A(n12507), .ZN(P3_U3483) );
  INV_X1 U14858 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12510) );
  AOI21_X1 U14859 ( .B1(n12509), .B2(n15518), .A(n12508), .ZN(n12578) );
  MUX2_X1 U14860 ( .A(n12510), .B(n12578), .S(n15540), .Z(n12511) );
  OAI21_X1 U14861 ( .B1(n12581), .B2(n12556), .A(n12511), .ZN(P3_U3482) );
  INV_X1 U14862 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12514) );
  AOI21_X1 U14863 ( .B1(n12513), .B2(n15518), .A(n12512), .ZN(n12582) );
  MUX2_X1 U14864 ( .A(n12514), .B(n12582), .S(n15540), .Z(n12515) );
  OAI21_X1 U14865 ( .B1(n12585), .B2(n12556), .A(n12515), .ZN(P3_U3481) );
  INV_X1 U14866 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12518) );
  AOI21_X1 U14867 ( .B1(n12517), .B2(n15518), .A(n12516), .ZN(n12586) );
  MUX2_X1 U14868 ( .A(n12518), .B(n12586), .S(n15540), .Z(n12519) );
  OAI21_X1 U14869 ( .B1(n12589), .B2(n12556), .A(n12519), .ZN(P3_U3480) );
  INV_X1 U14870 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12522) );
  AOI21_X1 U14871 ( .B1(n12521), .B2(n15518), .A(n12520), .ZN(n12590) );
  MUX2_X1 U14872 ( .A(n12522), .B(n12590), .S(n15540), .Z(n12523) );
  OAI21_X1 U14873 ( .B1(n12593), .B2(n12556), .A(n12523), .ZN(P3_U3479) );
  NAND2_X1 U14874 ( .A1(n12524), .A2(n15518), .ZN(n12525) );
  OAI211_X1 U14875 ( .C1(n12527), .C2(n15515), .A(n12526), .B(n12525), .ZN(
        n12594) );
  MUX2_X1 U14876 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12594), .S(n15540), .Z(
        P3_U3478) );
  AOI21_X1 U14877 ( .B1(n12529), .B2(n15518), .A(n12528), .ZN(n12595) );
  MUX2_X1 U14878 ( .A(n12530), .B(n12595), .S(n15540), .Z(n12531) );
  OAI21_X1 U14879 ( .B1(n12598), .B2(n12556), .A(n12531), .ZN(P3_U3477) );
  NAND2_X1 U14880 ( .A1(n12532), .A2(n15518), .ZN(n12533) );
  OAI211_X1 U14881 ( .C1(n12535), .C2(n15515), .A(n12534), .B(n12533), .ZN(
        n12599) );
  MUX2_X1 U14882 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12599), .S(n15540), .Z(
        P3_U3476) );
  NAND2_X1 U14883 ( .A1(n12536), .A2(n15518), .ZN(n12537) );
  OAI211_X1 U14884 ( .C1(n12539), .C2(n15515), .A(n12538), .B(n12537), .ZN(
        n12600) );
  MUX2_X1 U14885 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12600), .S(n15540), .Z(
        P3_U3475) );
  NAND2_X1 U14886 ( .A1(n12540), .A2(n15518), .ZN(n12541) );
  OAI211_X1 U14887 ( .C1(n12543), .C2(n15515), .A(n12542), .B(n12541), .ZN(
        n12601) );
  MUX2_X1 U14888 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n12601), .S(n15540), .Z(
        P3_U3474) );
  INV_X1 U14889 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12546) );
  AOI21_X1 U14890 ( .B1(n15518), .B2(n12545), .A(n12544), .ZN(n12602) );
  MUX2_X1 U14891 ( .A(n12546), .B(n12602), .S(n15540), .Z(n12547) );
  OAI21_X1 U14892 ( .B1(n12556), .B2(n12605), .A(n12547), .ZN(P3_U3473) );
  INV_X1 U14893 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12550) );
  AOI21_X1 U14894 ( .B1(n12549), .B2(n15518), .A(n12548), .ZN(n12606) );
  MUX2_X1 U14895 ( .A(n12550), .B(n12606), .S(n15540), .Z(n12551) );
  OAI21_X1 U14896 ( .B1(n12556), .B2(n12609), .A(n12551), .ZN(P3_U3472) );
  AOI21_X1 U14897 ( .B1(n15518), .B2(n12553), .A(n12552), .ZN(n12610) );
  MUX2_X1 U14898 ( .A(n12554), .B(n12610), .S(n15540), .Z(n12555) );
  OAI21_X1 U14899 ( .B1(n12614), .B2(n12556), .A(n12555), .ZN(P3_U3471) );
  NAND2_X1 U14900 ( .A1(n12557), .A2(n15518), .ZN(n12559) );
  AND3_X1 U14901 ( .A1(n12560), .A2(n12559), .A3(n12558), .ZN(n15467) );
  INV_X1 U14902 ( .A(n15467), .ZN(n12561) );
  MUX2_X1 U14903 ( .A(P3_REG1_REG_1__SCAN_IN), .B(n12561), .S(n15540), .Z(
        P3_U3460) );
  INV_X1 U14904 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12566) );
  INV_X1 U14905 ( .A(n12613), .ZN(n12562) );
  NAND2_X1 U14906 ( .A1(n12563), .A2(n12562), .ZN(n12565) );
  NAND2_X1 U14907 ( .A1(n12564), .A2(n15519), .ZN(n12568) );
  OAI211_X1 U14908 ( .C1(n15519), .C2(n12566), .A(n12565), .B(n12568), .ZN(
        P3_U3458) );
  NAND2_X1 U14909 ( .A1(n15521), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12567) );
  OAI211_X1 U14910 ( .C1(n12569), .C2(n12613), .A(n12568), .B(n12567), .ZN(
        P3_U3457) );
  INV_X1 U14911 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12571) );
  MUX2_X1 U14912 ( .A(n12571), .B(n12570), .S(n15519), .Z(n12572) );
  OAI21_X1 U14913 ( .B1(n12573), .B2(n12613), .A(n12572), .ZN(P3_U3452) );
  INV_X1 U14914 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12575) );
  MUX2_X1 U14915 ( .A(n12575), .B(n12574), .S(n15519), .Z(n12576) );
  OAI21_X1 U14916 ( .B1(n12577), .B2(n12613), .A(n12576), .ZN(P3_U3451) );
  MUX2_X1 U14917 ( .A(n12579), .B(n12578), .S(n15519), .Z(n12580) );
  OAI21_X1 U14918 ( .B1(n12581), .B2(n12613), .A(n12580), .ZN(P3_U3450) );
  INV_X1 U14919 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12583) );
  MUX2_X1 U14920 ( .A(n12583), .B(n12582), .S(n15519), .Z(n12584) );
  OAI21_X1 U14921 ( .B1(n12585), .B2(n12613), .A(n12584), .ZN(P3_U3449) );
  INV_X1 U14922 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12587) );
  MUX2_X1 U14923 ( .A(n12587), .B(n12586), .S(n15519), .Z(n12588) );
  OAI21_X1 U14924 ( .B1(n12589), .B2(n12613), .A(n12588), .ZN(P3_U3448) );
  INV_X1 U14925 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12591) );
  MUX2_X1 U14926 ( .A(n12591), .B(n12590), .S(n15519), .Z(n12592) );
  OAI21_X1 U14927 ( .B1(n12593), .B2(n12613), .A(n12592), .ZN(P3_U3447) );
  MUX2_X1 U14928 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n12594), .S(n15519), .Z(
        P3_U3446) );
  INV_X1 U14929 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12596) );
  MUX2_X1 U14930 ( .A(n12596), .B(n12595), .S(n15519), .Z(n12597) );
  OAI21_X1 U14931 ( .B1(n12598), .B2(n12613), .A(n12597), .ZN(P3_U3444) );
  MUX2_X1 U14932 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12599), .S(n15519), .Z(
        P3_U3441) );
  MUX2_X1 U14933 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n12600), .S(n15519), .Z(
        P3_U3438) );
  MUX2_X1 U14934 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n12601), .S(n15519), .Z(
        P3_U3435) );
  INV_X1 U14935 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12603) );
  MUX2_X1 U14936 ( .A(n12603), .B(n12602), .S(n15519), .Z(n12604) );
  OAI21_X1 U14937 ( .B1(n12613), .B2(n12605), .A(n12604), .ZN(P3_U3432) );
  INV_X1 U14938 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12607) );
  MUX2_X1 U14939 ( .A(n12607), .B(n12606), .S(n15519), .Z(n12608) );
  OAI21_X1 U14940 ( .B1(n12613), .B2(n12609), .A(n12608), .ZN(P3_U3429) );
  INV_X1 U14941 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n12611) );
  MUX2_X1 U14942 ( .A(n12611), .B(n12610), .S(n15519), .Z(n12612) );
  OAI21_X1 U14943 ( .B1(n12614), .B2(n12613), .A(n12612), .ZN(P3_U3426) );
  MUX2_X1 U14944 ( .A(n12616), .B(P3_D_REG_0__SCAN_IN), .S(n12615), .Z(
        P3_U3376) );
  NAND2_X1 U14945 ( .A1(n12618), .A2(n12617), .ZN(n12622) );
  OR4_X1 U14946 ( .A1(n12620), .A2(P3_IR_REG_30__SCAN_IN), .A3(n12619), .A4(
        P3_U3151), .ZN(n12621) );
  OAI211_X1 U14947 ( .C1(n12624), .C2(n12623), .A(n12622), .B(n12621), .ZN(
        P3_U3264) );
  INV_X1 U14948 ( .A(n12625), .ZN(n12626) );
  OAI222_X1 U14949 ( .A1(n12623), .A2(n12630), .B1(P3_U3151), .B2(n12628), 
        .C1(n12627), .C2(n12626), .ZN(P3_U3266) );
  INV_X1 U14950 ( .A(n12631), .ZN(n12632) );
  AOI21_X1 U14951 ( .B1(n12834), .B2(n12632), .A(n12854), .ZN(n12637) );
  NOR3_X1 U14952 ( .A1(n12852), .A2(n12634), .A3(n12633), .ZN(n12636) );
  OAI21_X1 U14953 ( .B1(n12637), .B2(n12636), .A(n12635), .ZN(n12641) );
  AOI22_X1 U14954 ( .A1(n15402), .A2(n12831), .B1(n12862), .B2(n12638), .ZN(
        n12640) );
  NAND2_X1 U14955 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13228) );
  NAND2_X1 U14956 ( .A1(n12838), .A2(n15401), .ZN(n12639) );
  NAND4_X1 U14957 ( .A1(n12641), .A2(n12640), .A3(n13228), .A4(n12639), .ZN(
        P2_U3185) );
  NAND2_X1 U14958 ( .A1(n13190), .A2(n9845), .ZN(n12675) );
  INV_X1 U14959 ( .A(n12675), .ZN(n12815) );
  XNOR2_X1 U14960 ( .A(n13526), .B(n12667), .ZN(n12676) );
  INV_X1 U14961 ( .A(n12676), .ZN(n12813) );
  XNOR2_X1 U14962 ( .A(n13577), .B(n12684), .ZN(n12644) );
  NAND2_X1 U14963 ( .A1(n9845), .A2(n13198), .ZN(n12645) );
  XNOR2_X1 U14964 ( .A(n12644), .B(n12645), .ZN(n12704) );
  AND2_X1 U14965 ( .A1(n12704), .A2(n12642), .ZN(n12643) );
  INV_X1 U14966 ( .A(n12644), .ZN(n12646) );
  NAND2_X1 U14967 ( .A1(n12646), .A2(n12645), .ZN(n12647) );
  NAND2_X1 U14968 ( .A1(n12700), .A2(n12647), .ZN(n12649) );
  XNOR2_X1 U14969 ( .A(n12973), .B(n12667), .ZN(n12648) );
  OR2_X1 U14970 ( .A1(n12649), .A2(n12648), .ZN(n12650) );
  XNOR2_X1 U14971 ( .A(n13460), .B(n12684), .ZN(n12769) );
  NAND2_X1 U14972 ( .A1(n9845), .A2(n13196), .ZN(n12651) );
  XNOR2_X1 U14973 ( .A(n12769), .B(n12651), .ZN(n12757) );
  INV_X1 U14974 ( .A(n12769), .ZN(n12652) );
  NAND2_X1 U14975 ( .A1(n12652), .A2(n12651), .ZN(n12653) );
  XNOR2_X1 U14976 ( .A(n13438), .B(n12684), .ZN(n12654) );
  NAND2_X1 U14977 ( .A1(n13195), .A2(n9845), .ZN(n12655) );
  XNOR2_X1 U14978 ( .A(n12654), .B(n12655), .ZN(n12770) );
  INV_X1 U14979 ( .A(n12654), .ZN(n12656) );
  NAND2_X1 U14980 ( .A1(n12656), .A2(n12655), .ZN(n12657) );
  XNOR2_X1 U14981 ( .A(n13549), .B(n12732), .ZN(n12658) );
  AND2_X1 U14982 ( .A1(n13194), .A2(n9845), .ZN(n12659) );
  NAND2_X1 U14983 ( .A1(n12658), .A2(n12659), .ZN(n12662) );
  INV_X1 U14984 ( .A(n12658), .ZN(n12716) );
  INV_X1 U14985 ( .A(n12659), .ZN(n12660) );
  NAND2_X1 U14986 ( .A1(n12716), .A2(n12660), .ZN(n12661) );
  NAND2_X1 U14987 ( .A1(n12662), .A2(n12661), .ZN(n12827) );
  XNOR2_X1 U14988 ( .A(n13543), .B(n12732), .ZN(n12664) );
  NAND2_X1 U14989 ( .A1(n13193), .A2(n9845), .ZN(n12665) );
  XNOR2_X1 U14990 ( .A(n12664), .B(n12665), .ZN(n12725) );
  AND2_X1 U14991 ( .A1(n12725), .A2(n12662), .ZN(n12663) );
  INV_X1 U14992 ( .A(n12664), .ZN(n12666) );
  XNOR2_X1 U14993 ( .A(n13537), .B(n12667), .ZN(n12668) );
  NAND2_X1 U14994 ( .A1(n13192), .A2(n9845), .ZN(n12669) );
  AND2_X1 U14995 ( .A1(n12668), .A2(n12669), .ZN(n12797) );
  INV_X1 U14996 ( .A(n12668), .ZN(n12671) );
  INV_X1 U14997 ( .A(n12669), .ZN(n12670) );
  NAND2_X1 U14998 ( .A1(n12671), .A2(n12670), .ZN(n12798) );
  XNOR2_X1 U14999 ( .A(n13367), .B(n12684), .ZN(n12674) );
  NAND2_X1 U15000 ( .A1(n13191), .A2(n9845), .ZN(n12672) );
  XNOR2_X1 U15001 ( .A(n12674), .B(n12672), .ZN(n12743) );
  NAND2_X1 U15002 ( .A1(n12744), .A2(n12743), .ZN(n12812) );
  INV_X1 U15003 ( .A(n12672), .ZN(n12673) );
  NAND2_X1 U15004 ( .A1(n12674), .A2(n12673), .ZN(n12811) );
  XNOR2_X1 U15005 ( .A(n13520), .B(n12732), .ZN(n12678) );
  NOR2_X1 U15006 ( .A1(n12809), .A2(n12677), .ZN(n12706) );
  XNOR2_X1 U15007 ( .A(n13513), .B(n12732), .ZN(n12680) );
  NAND2_X1 U15008 ( .A1(n13188), .A2(n9845), .ZN(n12679) );
  XNOR2_X1 U15009 ( .A(n12680), .B(n12679), .ZN(n12777) );
  XNOR2_X1 U15010 ( .A(n13314), .B(n12684), .ZN(n12682) );
  NAND2_X1 U15011 ( .A1(n13187), .A2(n9845), .ZN(n12681) );
  XNOR2_X1 U15012 ( .A(n12682), .B(n12681), .ZN(n12750) );
  INV_X1 U15013 ( .A(n12681), .ZN(n12683) );
  AOI22_X1 U15014 ( .A1(n12751), .A2(n12750), .B1(n12683), .B2(n12682), .ZN(
        n12845) );
  AND2_X1 U15015 ( .A1(n13186), .A2(n9845), .ZN(n12686) );
  XNOR2_X1 U15016 ( .A(n13303), .B(n12684), .ZN(n12685) );
  NOR2_X1 U15017 ( .A1(n12685), .A2(n12686), .ZN(n12687) );
  AOI21_X1 U15018 ( .B1(n12686), .B2(n12685), .A(n12687), .ZN(n12844) );
  NAND2_X1 U15019 ( .A1(n12845), .A2(n12844), .ZN(n12843) );
  INV_X1 U15020 ( .A(n12687), .ZN(n12688) );
  NAND2_X1 U15021 ( .A1(n12843), .A2(n12688), .ZN(n12731) );
  NAND2_X1 U15022 ( .A1(n13185), .A2(n9845), .ZN(n12728) );
  XNOR2_X1 U15023 ( .A(n13493), .B(n12732), .ZN(n12727) );
  XOR2_X1 U15024 ( .A(n12728), .B(n12727), .Z(n12730) );
  XNOR2_X1 U15025 ( .A(n12731), .B(n12730), .ZN(n12693) );
  AOI22_X1 U15026 ( .A1(n13184), .A2(n12848), .B1(n13167), .B2(n13186), .ZN(
        n13285) );
  OAI22_X1 U15027 ( .A1(n13285), .A2(n12860), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12689), .ZN(n12690) );
  AOI21_X1 U15028 ( .B1(n13290), .B2(n12862), .A(n12690), .ZN(n12692) );
  NAND2_X1 U15029 ( .A1(n13493), .A2(n12831), .ZN(n12691) );
  OAI211_X1 U15030 ( .C1(n12693), .C2(n12854), .A(n12692), .B(n12691), .ZN(
        P2_U3186) );
  NOR3_X1 U15031 ( .A1(n12695), .A2(n12694), .A3(n12852), .ZN(n12696) );
  AOI21_X1 U15032 ( .B1(n6691), .B2(n12846), .A(n12696), .ZN(n12705) );
  NAND2_X1 U15033 ( .A1(n12838), .A2(n12697), .ZN(n12698) );
  NAND2_X1 U15034 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15265)
         );
  OAI211_X1 U15035 ( .C1(n12825), .C2(n12699), .A(n12698), .B(n15265), .ZN(
        n12702) );
  NOR2_X1 U15036 ( .A1(n12700), .A2(n12854), .ZN(n12701) );
  AOI211_X1 U15037 ( .C1(n13577), .C2(n12831), .A(n12702), .B(n12701), .ZN(
        n12703) );
  OAI21_X1 U15038 ( .B1(n12705), .B2(n12704), .A(n12703), .ZN(P2_U3187) );
  NAND2_X1 U15039 ( .A1(n12818), .A2(n13189), .ZN(n12709) );
  OR2_X1 U15040 ( .A1(n12854), .A2(n12706), .ZN(n12708) );
  MUX2_X1 U15041 ( .A(n12709), .B(n12708), .S(n12707), .Z(n12714) );
  INV_X1 U15042 ( .A(n12710), .ZN(n13338) );
  AOI22_X1 U15043 ( .A1(n13188), .A2(n12848), .B1(n13167), .B2(n13190), .ZN(
        n13344) );
  OAI22_X1 U15044 ( .A1(n12860), .A2(n13344), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12711), .ZN(n12712) );
  AOI21_X1 U15045 ( .B1(n13338), .B2(n12862), .A(n12712), .ZN(n12713) );
  OAI211_X1 U15046 ( .C1(n13340), .C2(n12866), .A(n12714), .B(n12713), .ZN(
        P2_U3188) );
  INV_X1 U15047 ( .A(n12715), .ZN(n12826) );
  NOR3_X1 U15048 ( .A1(n12716), .A2(n12718), .A3(n12852), .ZN(n12717) );
  AOI21_X1 U15049 ( .B1(n12826), .B2(n12846), .A(n12717), .ZN(n12726) );
  INV_X1 U15050 ( .A(n13192), .ZN(n12719) );
  OAI22_X1 U15051 ( .A1(n12719), .A2(n12808), .B1(n12718), .B2(n12806), .ZN(
        n13542) );
  AOI22_X1 U15052 ( .A1(n12838), .A2(n13542), .B1(P2_REG3_REG_19__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12720) );
  OAI21_X1 U15053 ( .B1(n13398), .B2(n12825), .A(n12720), .ZN(n12723) );
  NOR2_X1 U15054 ( .A1(n12721), .A2(n12854), .ZN(n12722) );
  AOI211_X1 U15055 ( .C1(n13543), .C2(n12831), .A(n12723), .B(n12722), .ZN(
        n12724) );
  OAI21_X1 U15056 ( .B1(n12726), .B2(n12725), .A(n12724), .ZN(P2_U3191) );
  INV_X1 U15057 ( .A(n12727), .ZN(n12729) );
  OAI22_X1 U15058 ( .A1(n12731), .A2(n12730), .B1(n12729), .B2(n12728), .ZN(
        n12736) );
  NAND2_X1 U15059 ( .A1(n13184), .A2(n9845), .ZN(n12733) );
  XNOR2_X1 U15060 ( .A(n12733), .B(n12732), .ZN(n12734) );
  XNOR2_X1 U15061 ( .A(n13490), .B(n12734), .ZN(n12735) );
  XNOR2_X1 U15062 ( .A(n12736), .B(n12735), .ZN(n12742) );
  NAND2_X1 U15063 ( .A1(n13185), .A2(n13167), .ZN(n12738) );
  NAND2_X1 U15064 ( .A1(n13183), .A2(n12848), .ZN(n12737) );
  NAND2_X1 U15065 ( .A1(n12738), .A2(n12737), .ZN(n13267) );
  AOI22_X1 U15066 ( .A1(n13267), .A2(n12838), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12739) );
  OAI21_X1 U15067 ( .B1(n13271), .B2(n12825), .A(n12739), .ZN(n12740) );
  AOI21_X1 U15068 ( .B1(n13490), .B2(n12831), .A(n12740), .ZN(n12741) );
  OAI21_X1 U15069 ( .B1(n12742), .B2(n12854), .A(n12741), .ZN(P2_U3192) );
  XNOR2_X1 U15070 ( .A(n12744), .B(n12743), .ZN(n12749) );
  AOI22_X1 U15071 ( .A1(n13190), .A2(n12848), .B1(n13167), .B2(n13192), .ZN(
        n13530) );
  OAI22_X1 U15072 ( .A1(n12860), .A2(n13530), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12745), .ZN(n12746) );
  AOI21_X1 U15073 ( .B1(n13371), .B2(n12862), .A(n12746), .ZN(n12748) );
  NAND2_X1 U15074 ( .A1(n13367), .A2(n12831), .ZN(n12747) );
  OAI211_X1 U15075 ( .C1(n12749), .C2(n12854), .A(n12748), .B(n12747), .ZN(
        P2_U3195) );
  XNOR2_X1 U15076 ( .A(n12751), .B(n12750), .ZN(n12756) );
  AOI22_X1 U15077 ( .A1(n13186), .A2(n12848), .B1(n13167), .B2(n13188), .ZN(
        n13504) );
  OAI22_X1 U15078 ( .A1(n13504), .A2(n12860), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12752), .ZN(n12753) );
  AOI21_X1 U15079 ( .B1(n13312), .B2(n12862), .A(n12753), .ZN(n12755) );
  NAND2_X1 U15080 ( .A1(n13314), .A2(n12831), .ZN(n12754) );
  OAI211_X1 U15081 ( .C1(n12756), .C2(n12854), .A(n12755), .B(n12754), .ZN(
        P2_U3197) );
  OAI21_X1 U15082 ( .B1(n12758), .B2(n12757), .A(n12766), .ZN(n12759) );
  NAND2_X1 U15083 ( .A1(n12759), .A2(n12846), .ZN(n12763) );
  AOI22_X1 U15084 ( .A1(n13195), .A2(n12848), .B1(n13167), .B2(n13197), .ZN(
        n13453) );
  OAI22_X1 U15085 ( .A1(n12860), .A2(n13453), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12760), .ZN(n12761) );
  AOI21_X1 U15086 ( .B1(n13458), .B2(n12862), .A(n12761), .ZN(n12762) );
  OAI211_X1 U15087 ( .C1(n13561), .C2(n12866), .A(n12763), .B(n12762), .ZN(
        P2_U3198) );
  INV_X1 U15088 ( .A(n13434), .ZN(n12765) );
  AOI22_X1 U15089 ( .A1(n13194), .A2(n12848), .B1(n13167), .B2(n13196), .ZN(
        n13553) );
  INV_X1 U15090 ( .A(n13553), .ZN(n13435) );
  AOI22_X1 U15091 ( .A1(n12838), .A2(n13435), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12764) );
  OAI21_X1 U15092 ( .B1(n12765), .B2(n12825), .A(n12764), .ZN(n12774) );
  INV_X1 U15093 ( .A(n12766), .ZN(n12772) );
  NOR2_X1 U15094 ( .A1(n12852), .A2(n12767), .ZN(n12768) );
  AOI21_X1 U15095 ( .B1(n12769), .B2(n12846), .A(n12768), .ZN(n12771) );
  NOR3_X1 U15096 ( .A1(n12772), .A2(n12771), .A3(n12770), .ZN(n12773) );
  AOI211_X1 U15097 ( .C1(n13438), .C2(n12831), .A(n12774), .B(n12773), .ZN(
        n12775) );
  OAI21_X1 U15098 ( .B1(n12776), .B2(n12854), .A(n12775), .ZN(P2_U3200) );
  XNOR2_X1 U15099 ( .A(n12778), .B(n12777), .ZN(n12783) );
  AOI22_X1 U15100 ( .A1(n13187), .A2(n12848), .B1(n13167), .B2(n13189), .ZN(
        n13511) );
  OAI22_X1 U15101 ( .A1(n13511), .A2(n12860), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12779), .ZN(n12781) );
  NOR2_X1 U15102 ( .A1(n13513), .A2(n12866), .ZN(n12780) );
  AOI211_X1 U15103 ( .C1(n12862), .C2(n13327), .A(n12781), .B(n12780), .ZN(
        n12782) );
  OAI21_X1 U15104 ( .B1(n12783), .B2(n12854), .A(n12782), .ZN(P2_U3201) );
  OAI21_X1 U15105 ( .B1(n12790), .B2(n12785), .A(n12784), .ZN(n12786) );
  NAND2_X1 U15106 ( .A1(n12786), .A2(n12846), .ZN(n12796) );
  AOI22_X1 U15107 ( .A1(n12838), .A2(n12787), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12795) );
  INV_X1 U15108 ( .A(n12788), .ZN(n12789) );
  AOI22_X1 U15109 ( .A1(n12900), .A2(n12831), .B1(n12862), .B2(n12789), .ZN(
        n12794) );
  INV_X1 U15110 ( .A(n12790), .ZN(n12792) );
  NAND4_X1 U15111 ( .A1(n12818), .A2(n12792), .A3(n12791), .A4(n13210), .ZN(
        n12793) );
  NAND4_X1 U15112 ( .A1(n12796), .A2(n12795), .A3(n12794), .A4(n12793), .ZN(
        P2_U3202) );
  INV_X1 U15113 ( .A(n12797), .ZN(n12799) );
  NAND2_X1 U15114 ( .A1(n12799), .A2(n12798), .ZN(n12800) );
  XNOR2_X1 U15115 ( .A(n12801), .B(n12800), .ZN(n12805) );
  OAI22_X1 U15116 ( .A1(n12807), .A2(n12808), .B1(n13119), .B2(n12806), .ZN(
        n13379) );
  AOI22_X1 U15117 ( .A1(n12838), .A2(n13379), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12802) );
  OAI21_X1 U15118 ( .B1(n13384), .B2(n12825), .A(n12802), .ZN(n12803) );
  AOI21_X1 U15119 ( .B1(n13537), .B2(n12831), .A(n12803), .ZN(n12804) );
  OAI21_X1 U15120 ( .B1(n12805), .B2(n12854), .A(n12804), .ZN(P2_U3205) );
  OAI22_X1 U15121 ( .A1(n12809), .A2(n12808), .B1(n12807), .B2(n12806), .ZN(
        n13525) );
  AOI22_X1 U15122 ( .A1(n13525), .A2(n12838), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12810) );
  OAI21_X1 U15123 ( .B1(n13356), .B2(n12825), .A(n12810), .ZN(n12817) );
  NAND2_X1 U15124 ( .A1(n12812), .A2(n12811), .ZN(n12814) );
  XNOR2_X1 U15125 ( .A(n12814), .B(n12813), .ZN(n12819) );
  NOR3_X1 U15126 ( .A1(n12819), .A2(n12815), .A3(n12854), .ZN(n12816) );
  AOI211_X1 U15127 ( .C1(n13526), .C2(n12831), .A(n12817), .B(n12816), .ZN(
        n12821) );
  NAND3_X1 U15128 ( .A1(n12819), .A2(n12818), .A3(n13190), .ZN(n12820) );
  NAND2_X1 U15129 ( .A1(n12821), .A2(n12820), .ZN(P2_U3207) );
  NAND2_X1 U15130 ( .A1(n13193), .A2(n12848), .ZN(n12823) );
  NAND2_X1 U15131 ( .A1(n13195), .A2(n13167), .ZN(n12822) );
  NAND2_X1 U15132 ( .A1(n12823), .A2(n12822), .ZN(n13411) );
  AOI22_X1 U15133 ( .A1(n12838), .A2(n13411), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12824) );
  OAI21_X1 U15134 ( .B1(n13417), .B2(n12825), .A(n12824), .ZN(n12830) );
  AOI211_X1 U15135 ( .C1(n12828), .C2(n12827), .A(n12854), .B(n12826), .ZN(
        n12829) );
  AOI211_X1 U15136 ( .C1(n13549), .C2(n12831), .A(n12830), .B(n12829), .ZN(
        n12832) );
  INV_X1 U15137 ( .A(n12832), .ZN(P2_U3210) );
  NAND2_X1 U15138 ( .A1(n12835), .A2(n12834), .ZN(n12842) );
  AOI22_X1 U15139 ( .A1(n15393), .A2(n12831), .B1(n12862), .B2(n12836), .ZN(
        n12840) );
  NAND2_X1 U15140 ( .A1(n12838), .A2(n12837), .ZN(n12839) );
  NAND4_X1 U15141 ( .A1(n12842), .A2(n12841), .A3(n12840), .A4(n12839), .ZN(
        P2_U3211) );
  OAI21_X1 U15142 ( .B1(n12845), .B2(n12844), .A(n12843), .ZN(n12847) );
  NAND2_X1 U15143 ( .A1(n12847), .A2(n12846), .ZN(n12851) );
  AOI22_X1 U15144 ( .A1(n13185), .A2(n12848), .B1(n13167), .B2(n13187), .ZN(
        n13498) );
  OAI22_X1 U15145 ( .A1(n13498), .A2(n12860), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13662), .ZN(n12849) );
  AOI21_X1 U15146 ( .B1(n13300), .B2(n12862), .A(n12849), .ZN(n12850) );
  OAI211_X1 U15147 ( .C1(n7234), .C2(n12866), .A(n12851), .B(n12850), .ZN(
        P2_U3212) );
  OAI22_X1 U15148 ( .A1(n12855), .A2(n12854), .B1(n12853), .B2(n12852), .ZN(
        n12857) );
  NAND2_X1 U15149 ( .A1(n12857), .A2(n12856), .ZN(n12865) );
  INV_X1 U15150 ( .A(n12858), .ZN(n12863) );
  OAI22_X1 U15151 ( .A1(n12860), .A2(n13567), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12859), .ZN(n12861) );
  AOI21_X1 U15152 ( .B1(n12863), .B2(n12862), .A(n12861), .ZN(n12864) );
  OAI211_X1 U15153 ( .C1(n13568), .C2(n12866), .A(n12865), .B(n12864), .ZN(
        P2_U3213) );
  NAND2_X1 U15154 ( .A1(n12961), .A2(n13470), .ZN(n12870) );
  NAND2_X1 U15155 ( .A1(n12871), .A2(n12878), .ZN(n12873) );
  NAND2_X1 U15156 ( .A1(n12873), .A2(n12872), .ZN(n12875) );
  NAND2_X1 U15157 ( .A1(n12875), .A2(n12874), .ZN(n12877) );
  NAND2_X1 U15158 ( .A1(n13036), .A2(n13470), .ZN(n12880) );
  NAND2_X1 U15159 ( .A1(n13212), .A2(n12961), .ZN(n12879) );
  NAND2_X1 U15160 ( .A1(n12880), .A2(n12879), .ZN(n12881) );
  NAND2_X1 U15161 ( .A1(n12883), .A2(n12882), .ZN(n12884) );
  NAND2_X1 U15162 ( .A1(n12961), .A2(n13211), .ZN(n12887) );
  NAND2_X1 U15163 ( .A1(n13036), .A2(n12888), .ZN(n12886) );
  AOI22_X1 U15164 ( .A1(n13211), .A2(n13036), .B1(n12947), .B2(n12888), .ZN(
        n12889) );
  NAND2_X1 U15165 ( .A1(n13210), .A2(n13036), .ZN(n12894) );
  INV_X1 U15166 ( .A(n13036), .ZN(n12947) );
  NAND2_X1 U15167 ( .A1(n12947), .A2(n15370), .ZN(n12893) );
  NAND2_X1 U15168 ( .A1(n12894), .A2(n12893), .ZN(n12896) );
  AOI22_X1 U15169 ( .A1(n13210), .A2(n13098), .B1(n13036), .B2(n15370), .ZN(
        n12895) );
  NAND2_X1 U15170 ( .A1(n13209), .A2(n12947), .ZN(n12899) );
  NAND2_X1 U15171 ( .A1(n12878), .A2(n12900), .ZN(n12898) );
  NAND2_X1 U15172 ( .A1(n12899), .A2(n12898), .ZN(n12902) );
  AOI22_X1 U15173 ( .A1(n13209), .A2(n12878), .B1(n13098), .B2(n12900), .ZN(
        n12901) );
  NAND2_X1 U15174 ( .A1(n15385), .A2(n12947), .ZN(n12904) );
  NAND2_X1 U15175 ( .A1(n13208), .A2(n12878), .ZN(n12903) );
  NAND2_X1 U15176 ( .A1(n12904), .A2(n12903), .ZN(n12906) );
  AOI22_X1 U15177 ( .A1(n15385), .A2(n12878), .B1(n13208), .B2(n13098), .ZN(
        n12905) );
  NOR2_X1 U15178 ( .A1(n12907), .A2(n12906), .ZN(n12908) );
  NAND2_X1 U15179 ( .A1(n15393), .A2(n13036), .ZN(n12911) );
  NAND2_X1 U15180 ( .A1(n13207), .A2(n12947), .ZN(n12910) );
  NAND2_X1 U15181 ( .A1(n12911), .A2(n12910), .ZN(n12913) );
  AOI22_X1 U15182 ( .A1(n15393), .A2(n13098), .B1(n13036), .B2(n13207), .ZN(
        n12912) );
  NAND2_X1 U15183 ( .A1(n15402), .A2(n12947), .ZN(n12916) );
  NAND2_X1 U15184 ( .A1(n13206), .A2(n12878), .ZN(n12915) );
  NAND2_X1 U15185 ( .A1(n12916), .A2(n12915), .ZN(n12921) );
  NAND2_X1 U15186 ( .A1(n15402), .A2(n13036), .ZN(n12917) );
  OAI21_X1 U15187 ( .B1(n12918), .B2(n13036), .A(n12917), .ZN(n12919) );
  NAND2_X1 U15188 ( .A1(n12924), .A2(n13036), .ZN(n12923) );
  NAND2_X1 U15189 ( .A1(n13205), .A2(n12947), .ZN(n12922) );
  NAND2_X1 U15190 ( .A1(n12923), .A2(n12922), .ZN(n12926) );
  AOI22_X1 U15191 ( .A1(n12924), .A2(n13098), .B1(n13036), .B2(n13205), .ZN(
        n12925) );
  NAND2_X1 U15192 ( .A1(n15412), .A2(n13098), .ZN(n12928) );
  NAND2_X1 U15193 ( .A1(n13203), .A2(n13036), .ZN(n12927) );
  NAND2_X1 U15194 ( .A1(n12928), .A2(n12927), .ZN(n12933) );
  NAND2_X1 U15195 ( .A1(n12934), .A2(n12933), .ZN(n12932) );
  NAND2_X1 U15196 ( .A1(n15412), .A2(n12878), .ZN(n12929) );
  OAI21_X1 U15197 ( .B1(n12930), .B2(n13036), .A(n12929), .ZN(n12931) );
  NAND2_X1 U15198 ( .A1(n12932), .A2(n12931), .ZN(n12935) );
  NAND2_X1 U15199 ( .A1(n15420), .A2(n12878), .ZN(n12937) );
  NAND2_X1 U15200 ( .A1(n13202), .A2(n12947), .ZN(n12936) );
  AOI22_X1 U15201 ( .A1(n15420), .A2(n13098), .B1(n13036), .B2(n13202), .ZN(
        n12938) );
  NAND2_X1 U15202 ( .A1(n12941), .A2(n12947), .ZN(n12940) );
  NAND2_X1 U15203 ( .A1(n13201), .A2(n13036), .ZN(n12939) );
  AOI22_X1 U15204 ( .A1(n12941), .A2(n12878), .B1(n13201), .B2(n12947), .ZN(
        n12942) );
  INV_X1 U15205 ( .A(n12942), .ZN(n12943) );
  NAND2_X1 U15206 ( .A1(n13855), .A2(n13036), .ZN(n12946) );
  NAND2_X1 U15207 ( .A1(n13200), .A2(n12947), .ZN(n12945) );
  NAND2_X1 U15208 ( .A1(n13855), .A2(n12947), .ZN(n12948) );
  OAI21_X1 U15209 ( .B1(n12949), .B2(n12961), .A(n12948), .ZN(n12950) );
  NAND2_X1 U15210 ( .A1(n13582), .A2(n13098), .ZN(n12952) );
  NAND2_X1 U15211 ( .A1(n13199), .A2(n13036), .ZN(n12951) );
  NAND2_X1 U15212 ( .A1(n12952), .A2(n12951), .ZN(n12954) );
  AOI22_X1 U15213 ( .A1(n13582), .A2(n12878), .B1(n13199), .B2(n13098), .ZN(
        n12953) );
  NOR2_X1 U15214 ( .A1(n12955), .A2(n12954), .ZN(n12956) );
  NAND2_X1 U15215 ( .A1(n13577), .A2(n13036), .ZN(n12959) );
  NAND2_X1 U15216 ( .A1(n13198), .A2(n12947), .ZN(n12958) );
  NAND2_X1 U15217 ( .A1(n12959), .A2(n12958), .ZN(n12964) );
  NAND2_X1 U15218 ( .A1(n13577), .A2(n12947), .ZN(n12960) );
  OAI21_X1 U15219 ( .B1(n12962), .B2(n12961), .A(n12960), .ZN(n12963) );
  AND2_X1 U15220 ( .A1(n13195), .A2(n13036), .ZN(n12966) );
  AOI21_X1 U15221 ( .B1(n13438), .B2(n13098), .A(n12966), .ZN(n12989) );
  NAND2_X1 U15222 ( .A1(n13438), .A2(n13036), .ZN(n12968) );
  NAND2_X1 U15223 ( .A1(n13195), .A2(n13098), .ZN(n12967) );
  NAND2_X1 U15224 ( .A1(n12968), .A2(n12967), .ZN(n12987) );
  AND2_X1 U15225 ( .A1(n13196), .A2(n13036), .ZN(n12969) );
  AOI21_X1 U15226 ( .B1(n13460), .B2(n13098), .A(n12969), .ZN(n12983) );
  NAND2_X1 U15227 ( .A1(n13460), .A2(n13036), .ZN(n12971) );
  NAND2_X1 U15228 ( .A1(n13196), .A2(n13098), .ZN(n12970) );
  NAND2_X1 U15229 ( .A1(n12971), .A2(n12970), .ZN(n12982) );
  AOI22_X1 U15230 ( .A1(n12989), .A2(n12987), .B1(n12983), .B2(n12982), .ZN(
        n12978) );
  AND2_X1 U15231 ( .A1(n13197), .A2(n13036), .ZN(n12972) );
  AOI21_X1 U15232 ( .B1(n12973), .B2(n13098), .A(n12972), .ZN(n12980) );
  NAND2_X1 U15233 ( .A1(n12973), .A2(n13036), .ZN(n12975) );
  NAND2_X1 U15234 ( .A1(n13197), .A2(n13098), .ZN(n12974) );
  NAND2_X1 U15235 ( .A1(n12975), .A2(n12974), .ZN(n12979) );
  NAND2_X1 U15236 ( .A1(n12980), .A2(n12979), .ZN(n12976) );
  INV_X1 U15237 ( .A(n12978), .ZN(n12981) );
  OR3_X1 U15238 ( .A1(n12981), .A2(n12980), .A3(n12979), .ZN(n12995) );
  INV_X1 U15239 ( .A(n12982), .ZN(n12985) );
  INV_X1 U15240 ( .A(n12983), .ZN(n12984) );
  NAND2_X1 U15241 ( .A1(n12985), .A2(n12984), .ZN(n12988) );
  NAND3_X1 U15242 ( .A1(n12988), .A2(n12986), .A3(n13555), .ZN(n12993) );
  INV_X1 U15243 ( .A(n12987), .ZN(n12992) );
  INV_X1 U15244 ( .A(n12988), .ZN(n12991) );
  INV_X1 U15245 ( .A(n12989), .ZN(n12990) );
  AOI22_X1 U15246 ( .A1(n12993), .A2(n12992), .B1(n12991), .B2(n12990), .ZN(
        n12994) );
  AND2_X1 U15247 ( .A1(n13194), .A2(n13098), .ZN(n12996) );
  AOI21_X1 U15248 ( .B1(n13549), .B2(n12878), .A(n12996), .ZN(n13000) );
  NAND2_X1 U15249 ( .A1(n13549), .A2(n13098), .ZN(n12998) );
  NAND2_X1 U15250 ( .A1(n13194), .A2(n13036), .ZN(n12997) );
  NAND2_X1 U15251 ( .A1(n12998), .A2(n12997), .ZN(n12999) );
  NAND2_X1 U15252 ( .A1(n13001), .A2(n13000), .ZN(n13002) );
  NAND2_X1 U15253 ( .A1(n13543), .A2(n13098), .ZN(n13005) );
  NAND2_X1 U15254 ( .A1(n13193), .A2(n13036), .ZN(n13004) );
  AOI22_X1 U15255 ( .A1(n13543), .A2(n12878), .B1(n13193), .B2(n12947), .ZN(
        n13006) );
  NAND2_X1 U15256 ( .A1(n13537), .A2(n13036), .ZN(n13008) );
  NAND2_X1 U15257 ( .A1(n13192), .A2(n12947), .ZN(n13007) );
  NAND2_X1 U15258 ( .A1(n13008), .A2(n13007), .ZN(n13010) );
  AOI22_X1 U15259 ( .A1(n13537), .A2(n13098), .B1(n13036), .B2(n13192), .ZN(
        n13009) );
  NAND2_X1 U15260 ( .A1(n13367), .A2(n13098), .ZN(n13013) );
  NAND2_X1 U15261 ( .A1(n13191), .A2(n13036), .ZN(n13012) );
  NAND2_X1 U15262 ( .A1(n13013), .A2(n13012), .ZN(n13015) );
  AOI22_X1 U15263 ( .A1(n13367), .A2(n12878), .B1(n13191), .B2(n13098), .ZN(
        n13014) );
  NOR2_X1 U15264 ( .A1(n13016), .A2(n13015), .ZN(n13017) );
  NAND2_X1 U15265 ( .A1(n13526), .A2(n13036), .ZN(n13020) );
  NAND2_X1 U15266 ( .A1(n13190), .A2(n13098), .ZN(n13019) );
  NAND2_X1 U15267 ( .A1(n13020), .A2(n13019), .ZN(n13022) );
  AOI22_X1 U15268 ( .A1(n13526), .A2(n13098), .B1(n13036), .B2(n13190), .ZN(
        n13021) );
  NAND2_X1 U15269 ( .A1(n13520), .A2(n12961), .ZN(n13025) );
  NAND2_X1 U15270 ( .A1(n13189), .A2(n12878), .ZN(n13024) );
  NAND2_X1 U15271 ( .A1(n13025), .A2(n13024), .ZN(n13031) );
  NAND2_X1 U15272 ( .A1(n13520), .A2(n13036), .ZN(n13027) );
  NAND2_X1 U15273 ( .A1(n13189), .A2(n13098), .ZN(n13026) );
  NAND2_X1 U15274 ( .A1(n13027), .A2(n13026), .ZN(n13028) );
  NAND2_X1 U15275 ( .A1(n13029), .A2(n13028), .ZN(n13035) );
  INV_X1 U15276 ( .A(n13030), .ZN(n13033) );
  INV_X1 U15277 ( .A(n13031), .ZN(n13032) );
  NAND2_X1 U15278 ( .A1(n13033), .A2(n13032), .ZN(n13034) );
  NAND2_X1 U15279 ( .A1(n13332), .A2(n13036), .ZN(n13038) );
  NAND2_X1 U15280 ( .A1(n13188), .A2(n13098), .ZN(n13037) );
  AOI22_X1 U15281 ( .A1(n13332), .A2(n12947), .B1(n13036), .B2(n13188), .ZN(
        n13039) );
  NAND2_X1 U15282 ( .A1(n13314), .A2(n13098), .ZN(n13041) );
  NAND2_X1 U15283 ( .A1(n13187), .A2(n12878), .ZN(n13040) );
  NAND2_X1 U15284 ( .A1(n13041), .A2(n13040), .ZN(n13045) );
  NAND2_X1 U15285 ( .A1(n13314), .A2(n13036), .ZN(n13042) );
  INV_X1 U15286 ( .A(n13044), .ZN(n13047) );
  NAND2_X1 U15287 ( .A1(n13303), .A2(n12878), .ZN(n13050) );
  NAND2_X1 U15288 ( .A1(n13186), .A2(n13098), .ZN(n13049) );
  NAND2_X1 U15289 ( .A1(n13050), .A2(n13049), .ZN(n13052) );
  AOI22_X1 U15290 ( .A1(n13303), .A2(n13098), .B1(n12878), .B2(n13186), .ZN(
        n13051) );
  NAND2_X1 U15291 ( .A1(n13493), .A2(n13098), .ZN(n13055) );
  NAND2_X1 U15292 ( .A1(n13185), .A2(n13036), .ZN(n13054) );
  NAND2_X1 U15293 ( .A1(n13055), .A2(n13054), .ZN(n13100) );
  INV_X1 U15294 ( .A(n13056), .ZN(n13057) );
  NOR2_X1 U15295 ( .A1(n13057), .A2(SI_29_), .ZN(n13058) );
  MUX2_X1 U15296 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n13064), .Z(n13061) );
  NAND2_X1 U15297 ( .A1(n13061), .A2(SI_30_), .ZN(n13063) );
  OAI21_X1 U15298 ( .B1(SI_30_), .B2(n13061), .A(n13063), .ZN(n13078) );
  INV_X1 U15299 ( .A(n13078), .ZN(n13062) );
  NAND2_X1 U15300 ( .A1(n13077), .A2(n13062), .ZN(n13081) );
  NAND2_X1 U15301 ( .A1(n13081), .A2(n13063), .ZN(n13067) );
  MUX2_X1 U15302 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n13064), .Z(n13065) );
  XNOR2_X1 U15303 ( .A(n13065), .B(SI_31_), .ZN(n13066) );
  NAND2_X1 U15304 ( .A1(n14088), .A2(n13068), .ZN(n13071) );
  INV_X1 U15305 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13069) );
  OR2_X1 U15306 ( .A1(n6565), .A2(n13069), .ZN(n13070) );
  INV_X1 U15307 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13683) );
  NAND2_X1 U15308 ( .A1(n13072), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U15309 ( .A1(n9306), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n13073) );
  OAI211_X1 U15310 ( .C1(n6549), .C2(n13683), .A(n13074), .B(n13073), .ZN(
        n13251) );
  INV_X1 U15311 ( .A(n13251), .ZN(n13075) );
  NAND2_X1 U15312 ( .A1(n13253), .A2(n13075), .ZN(n13113) );
  OR2_X1 U15313 ( .A1(n13253), .A2(n13075), .ZN(n13076) );
  INV_X1 U15314 ( .A(n13077), .ZN(n13079) );
  NAND2_X1 U15315 ( .A1(n13079), .A2(n13078), .ZN(n13080) );
  OR2_X1 U15316 ( .A1(n13083), .A2(n13884), .ZN(n13084) );
  AND2_X1 U15317 ( .A1(n13182), .A2(n12878), .ZN(n13086) );
  AOI21_X1 U15318 ( .B1(n13261), .B2(n12961), .A(n13086), .ZN(n13107) );
  NAND2_X1 U15319 ( .A1(n13261), .A2(n13036), .ZN(n13090) );
  NAND2_X1 U15320 ( .A1(n13251), .A2(n13098), .ZN(n13087) );
  NAND2_X1 U15321 ( .A1(n13172), .A2(n15314), .ZN(n13159) );
  NAND4_X1 U15322 ( .A1(n10346), .A2(n13087), .A3(n13163), .A4(n13159), .ZN(
        n13088) );
  NAND2_X1 U15323 ( .A1(n13088), .A2(n13182), .ZN(n13089) );
  NAND2_X1 U15324 ( .A1(n13090), .A2(n13089), .ZN(n13106) );
  AND2_X1 U15325 ( .A1(n13183), .A2(n13036), .ZN(n13091) );
  AOI21_X1 U15326 ( .B1(n13484), .B2(n12961), .A(n13091), .ZN(n13104) );
  NAND2_X1 U15327 ( .A1(n13484), .A2(n12878), .ZN(n13093) );
  NAND2_X1 U15328 ( .A1(n13183), .A2(n13098), .ZN(n13092) );
  NAND2_X1 U15329 ( .A1(n13093), .A2(n13092), .ZN(n13103) );
  AND2_X1 U15330 ( .A1(n13184), .A2(n13036), .ZN(n13094) );
  AOI21_X1 U15331 ( .B1(n13490), .B2(n12961), .A(n13094), .ZN(n13102) );
  NAND2_X1 U15332 ( .A1(n13490), .A2(n13036), .ZN(n13096) );
  NAND2_X1 U15333 ( .A1(n13184), .A2(n13098), .ZN(n13095) );
  NAND2_X1 U15334 ( .A1(n13096), .A2(n13095), .ZN(n13101) );
  NAND2_X1 U15335 ( .A1(n13102), .A2(n13101), .ZN(n13097) );
  AOI22_X1 U15336 ( .A1(n13493), .A2(n12878), .B1(n13185), .B2(n13098), .ZN(
        n13099) );
  OAI22_X1 U15337 ( .A1(n13104), .A2(n13103), .B1(n13102), .B2(n13101), .ZN(
        n13105) );
  OR2_X1 U15338 ( .A1(n13116), .A2(n13105), .ZN(n13110) );
  INV_X1 U15339 ( .A(n13106), .ZN(n13109) );
  INV_X1 U15340 ( .A(n13107), .ZN(n13108) );
  AOI22_X1 U15341 ( .A1(n13111), .A2(n13110), .B1(n13109), .B2(n13108), .ZN(
        n13115) );
  NAND2_X1 U15342 ( .A1(n13036), .A2(n13251), .ZN(n13112) );
  OAI22_X1 U15343 ( .A1(n13113), .A2(n13036), .B1(n13112), .B2(n13253), .ZN(
        n13114) );
  XNOR2_X1 U15344 ( .A(n13261), .B(n13182), .ZN(n13152) );
  XNOR2_X1 U15345 ( .A(n13543), .B(n13119), .ZN(n13404) );
  NOR2_X1 U15346 ( .A1(n15362), .A2(n6561), .ZN(n13123) );
  NAND4_X1 U15347 ( .A1(n13123), .A2(n13122), .A3(n13121), .A4(n6954), .ZN(
        n13126) );
  NOR3_X1 U15348 ( .A1(n13126), .A2(n13125), .A3(n13124), .ZN(n13129) );
  NAND4_X1 U15349 ( .A1(n13130), .A2(n13129), .A3(n13128), .A4(n13127), .ZN(
        n13131) );
  NOR2_X1 U15350 ( .A1(n13132), .A2(n13131), .ZN(n13135) );
  NAND4_X1 U15351 ( .A1(n13136), .A2(n13135), .A3(n13134), .A4(n13133), .ZN(
        n13137) );
  OR4_X1 U15352 ( .A1(n13430), .A2(n13448), .A3(n13138), .A4(n13137), .ZN(
        n13139) );
  OR4_X1 U15353 ( .A1(n13409), .A2(n13141), .A3(n13140), .A4(n13139), .ZN(
        n13142) );
  NOR2_X1 U15354 ( .A1(n13404), .A2(n13142), .ZN(n13143) );
  XNOR2_X1 U15355 ( .A(n13367), .B(n13191), .ZN(n13365) );
  NAND4_X1 U15356 ( .A1(n13352), .A2(n13143), .A3(n13365), .A4(n13388), .ZN(
        n13144) );
  NOR2_X1 U15357 ( .A1(n13320), .A2(n13144), .ZN(n13145) );
  XNOR2_X1 U15358 ( .A(n13520), .B(n13189), .ZN(n13342) );
  NAND4_X1 U15359 ( .A1(n13297), .A2(n13145), .A3(n13308), .A4(n13342), .ZN(
        n13146) );
  NOR3_X1 U15360 ( .A1(n13148), .A2(n13147), .A3(n13146), .ZN(n13150) );
  NAND3_X1 U15361 ( .A1(n10346), .A2(n13157), .A3(n6984), .ZN(n13158) );
  OAI211_X1 U15362 ( .C1(n13173), .C2(n13174), .A(n13159), .B(n13158), .ZN(
        n13160) );
  NAND2_X1 U15363 ( .A1(n13160), .A2(n13177), .ZN(n13161) );
  NAND2_X1 U15364 ( .A1(n10346), .A2(n13244), .ZN(n13162) );
  OAI211_X1 U15365 ( .C1(n13172), .C2(n13164), .A(n13163), .B(n13162), .ZN(
        n13165) );
  NAND4_X1 U15366 ( .A1(n15358), .A2(n13169), .A3(n13168), .A4(n13167), .ZN(
        n13170) );
  OAI211_X1 U15367 ( .C1(n13172), .C2(n13171), .A(n13170), .B(P2_B_REG_SCAN_IN), .ZN(n13180) );
  INV_X1 U15368 ( .A(n13173), .ZN(n13178) );
  INV_X1 U15369 ( .A(n15314), .ZN(n13176) );
  INV_X1 U15370 ( .A(n13174), .ZN(n13175) );
  NAND4_X1 U15371 ( .A1(n13178), .A2(n13177), .A3(n13176), .A4(n13175), .ZN(
        n13179) );
  INV_X2 U15372 ( .A(P2_U3947), .ZN(n13204) );
  MUX2_X1 U15373 ( .A(n13251), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13204), .Z(
        P2_U3562) );
  MUX2_X1 U15374 ( .A(n13182), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13204), .Z(
        P2_U3561) );
  MUX2_X1 U15375 ( .A(n13183), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13204), .Z(
        P2_U3560) );
  MUX2_X1 U15376 ( .A(n13184), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13204), .Z(
        P2_U3559) );
  MUX2_X1 U15377 ( .A(n13185), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13204), .Z(
        P2_U3558) );
  MUX2_X1 U15378 ( .A(n13186), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13204), .Z(
        P2_U3557) );
  MUX2_X1 U15379 ( .A(n13187), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13204), .Z(
        P2_U3556) );
  MUX2_X1 U15380 ( .A(n13188), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13204), .Z(
        P2_U3555) );
  MUX2_X1 U15381 ( .A(n13189), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13204), .Z(
        P2_U3554) );
  MUX2_X1 U15382 ( .A(n13190), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13204), .Z(
        P2_U3553) );
  MUX2_X1 U15383 ( .A(n13191), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13204), .Z(
        P2_U3552) );
  MUX2_X1 U15384 ( .A(n13192), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13204), .Z(
        P2_U3551) );
  MUX2_X1 U15385 ( .A(n13193), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13204), .Z(
        P2_U3550) );
  MUX2_X1 U15386 ( .A(n13194), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13204), .Z(
        P2_U3549) );
  MUX2_X1 U15387 ( .A(n13195), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13204), .Z(
        P2_U3548) );
  MUX2_X1 U15388 ( .A(n13196), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13204), .Z(
        P2_U3547) );
  MUX2_X1 U15389 ( .A(n13197), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13204), .Z(
        P2_U3546) );
  MUX2_X1 U15390 ( .A(n13198), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13204), .Z(
        P2_U3545) );
  MUX2_X1 U15391 ( .A(n13199), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13204), .Z(
        P2_U3544) );
  MUX2_X1 U15392 ( .A(n13200), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13204), .Z(
        P2_U3543) );
  MUX2_X1 U15393 ( .A(n13201), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13204), .Z(
        P2_U3542) );
  MUX2_X1 U15394 ( .A(n13202), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13204), .Z(
        P2_U3541) );
  MUX2_X1 U15395 ( .A(n13203), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13204), .Z(
        P2_U3540) );
  MUX2_X1 U15396 ( .A(n13205), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13204), .Z(
        P2_U3539) );
  MUX2_X1 U15397 ( .A(n13206), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13204), .Z(
        P2_U3538) );
  MUX2_X1 U15398 ( .A(n13207), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13204), .Z(
        P2_U3537) );
  MUX2_X1 U15399 ( .A(n13208), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13204), .Z(
        P2_U3536) );
  MUX2_X1 U15400 ( .A(n13209), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13204), .Z(
        P2_U3535) );
  MUX2_X1 U15401 ( .A(n13210), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13204), .Z(
        P2_U3534) );
  MUX2_X1 U15402 ( .A(n13211), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13204), .Z(
        P2_U3533) );
  MUX2_X1 U15403 ( .A(n13212), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13204), .Z(
        P2_U3532) );
  MUX2_X1 U15404 ( .A(n9847), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13204), .Z(
        P2_U3531) );
  INV_X1 U15405 ( .A(n13213), .ZN(n13218) );
  NOR3_X1 U15406 ( .A1(n13216), .A2(n13215), .A3(n13214), .ZN(n13217) );
  NOR3_X1 U15407 ( .A1(n13218), .A2(n13217), .A3(n15242), .ZN(n13219) );
  AOI21_X1 U15408 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(n15294), .A(n13219), .ZN(
        n13229) );
  NAND2_X1 U15409 ( .A1(n15299), .A2(n13220), .ZN(n13227) );
  MUX2_X1 U15410 ( .A(n9236), .B(P2_REG1_REG_7__SCAN_IN), .S(n13220), .Z(
        n13221) );
  NAND3_X1 U15411 ( .A1(n13223), .A2(n13222), .A3(n13221), .ZN(n13224) );
  NAND3_X1 U15412 ( .A1(n15302), .A2(n13225), .A3(n13224), .ZN(n13226) );
  NAND4_X1 U15413 ( .A1(n13229), .A2(n13228), .A3(n13227), .A4(n13226), .ZN(
        P2_U3221) );
  NOR2_X1 U15414 ( .A1(n13234), .A2(n13230), .ZN(n13231) );
  INV_X1 U15415 ( .A(n13243), .ZN(n13241) );
  INV_X1 U15416 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13238) );
  NAND2_X1 U15417 ( .A1(n13234), .A2(n13233), .ZN(n13236) );
  NAND2_X1 U15418 ( .A1(n13236), .A2(n13235), .ZN(n13237) );
  XNOR2_X1 U15419 ( .A(n13238), .B(n13237), .ZN(n13242) );
  OAI21_X1 U15420 ( .B1(n13242), .B2(n13239), .A(n15273), .ZN(n13240) );
  AOI21_X1 U15421 ( .B1(n13241), .B2(n15296), .A(n13240), .ZN(n13246) );
  AOI22_X1 U15422 ( .A1(n13243), .A2(n15296), .B1(n15302), .B2(n13242), .ZN(
        n13245) );
  MUX2_X1 U15423 ( .A(n13246), .B(n13245), .S(n13244), .Z(n13248) );
  NAND2_X1 U15424 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n13247)
         );
  OAI211_X1 U15425 ( .C1(n7766), .C2(n13249), .A(n13248), .B(n13247), .ZN(
        P2_U3233) );
  NAND2_X1 U15426 ( .A1(n13482), .A2(n13257), .ZN(n13256) );
  XOR2_X1 U15427 ( .A(n13256), .B(n13253), .Z(n13250) );
  NAND2_X1 U15428 ( .A1(n13250), .A2(n13431), .ZN(n13478) );
  NAND2_X1 U15429 ( .A1(n13252), .A2(n13251), .ZN(n13480) );
  NOR2_X1 U15430 ( .A1(n15320), .A2(n13480), .ZN(n13259) );
  INV_X1 U15431 ( .A(n13253), .ZN(n13479) );
  NOR2_X1 U15432 ( .A1(n13479), .A2(n13420), .ZN(n13254) );
  AOI211_X1 U15433 ( .C1(n15320), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13259), 
        .B(n13254), .ZN(n13255) );
  OAI21_X1 U15434 ( .B1(n13478), .B2(n13440), .A(n13255), .ZN(P2_U3234) );
  OAI211_X1 U15435 ( .C1(n13482), .C2(n13257), .A(n13256), .B(n13431), .ZN(
        n13481) );
  NOR2_X1 U15436 ( .A1(n13472), .A2(n13258), .ZN(n13260) );
  AOI211_X1 U15437 ( .C1(n13261), .C2(n13471), .A(n13260), .B(n13259), .ZN(
        n13262) );
  OAI21_X1 U15438 ( .B1(n13481), .B2(n13440), .A(n13262), .ZN(P2_U3235) );
  XNOR2_X1 U15439 ( .A(n13263), .B(n13265), .ZN(n13491) );
  NAND2_X1 U15440 ( .A1(n13264), .A2(n15409), .ZN(n13270) );
  AOI21_X1 U15441 ( .B1(n13281), .B2(n13266), .A(n13265), .ZN(n13269) );
  INV_X1 U15442 ( .A(n13267), .ZN(n13268) );
  NOR2_X1 U15443 ( .A1(n13271), .A2(n13397), .ZN(n13272) );
  OAI21_X1 U15444 ( .B1(n13488), .B2(n13272), .A(n13472), .ZN(n13279) );
  INV_X1 U15445 ( .A(n13288), .ZN(n13274) );
  AOI211_X1 U15446 ( .C1(n13490), .C2(n13274), .A(n13562), .B(n7231), .ZN(
        n13489) );
  OAI22_X1 U15447 ( .A1(n13276), .A2(n13420), .B1(n13472), .B2(n13275), .ZN(
        n13277) );
  AOI21_X1 U15448 ( .B1(n13489), .B2(n13467), .A(n13277), .ZN(n13278) );
  OAI211_X1 U15449 ( .C1(n13465), .C2(n13491), .A(n13279), .B(n13278), .ZN(
        P2_U3237) );
  XNOR2_X1 U15450 ( .A(n13280), .B(n13282), .ZN(n13492) );
  INV_X1 U15451 ( .A(n13492), .ZN(n13295) );
  OAI21_X1 U15452 ( .B1(n13283), .B2(n13282), .A(n13281), .ZN(n13284) );
  NAND2_X1 U15453 ( .A1(n13284), .A2(n15409), .ZN(n13286) );
  NAND2_X1 U15454 ( .A1(n13286), .A2(n13285), .ZN(n13496) );
  NAND2_X1 U15455 ( .A1(n13493), .A2(n6600), .ZN(n13287) );
  NAND2_X1 U15456 ( .A1(n13287), .A2(n13431), .ZN(n13289) );
  OR2_X1 U15457 ( .A1(n13289), .A2(n13288), .ZN(n13494) );
  AOI22_X1 U15458 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(n15320), .B1(n13290), 
        .B2(n15318), .ZN(n13292) );
  NAND2_X1 U15459 ( .A1(n13493), .A2(n13471), .ZN(n13291) );
  OAI211_X1 U15460 ( .C1(n13494), .C2(n13440), .A(n13292), .B(n13291), .ZN(
        n13293) );
  AOI21_X1 U15461 ( .B1(n13496), .B2(n13472), .A(n13293), .ZN(n13294) );
  OAI21_X1 U15462 ( .B1(n13295), .B2(n13465), .A(n13294), .ZN(P2_U3238) );
  XNOR2_X1 U15463 ( .A(n13296), .B(n13297), .ZN(n13503) );
  XNOR2_X1 U15464 ( .A(n13298), .B(n13297), .ZN(n13501) );
  AOI21_X1 U15465 ( .B1(n13303), .B2(n13311), .A(n13562), .ZN(n13299) );
  NAND2_X1 U15466 ( .A1(n13299), .A2(n6600), .ZN(n13499) );
  AOI22_X1 U15467 ( .A1(n15320), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13300), 
        .B2(n15318), .ZN(n13301) );
  OAI21_X1 U15468 ( .B1(n13498), .B2(n15320), .A(n13301), .ZN(n13302) );
  AOI21_X1 U15469 ( .B1(n13303), .B2(n13471), .A(n13302), .ZN(n13304) );
  OAI21_X1 U15470 ( .B1(n13499), .B2(n13440), .A(n13304), .ZN(n13305) );
  AOI21_X1 U15471 ( .B1(n13501), .B2(n13406), .A(n13305), .ZN(n13306) );
  OAI21_X1 U15472 ( .B1(n13503), .B2(n13465), .A(n13306), .ZN(P2_U3239) );
  XOR2_X1 U15473 ( .A(n13307), .B(n13308), .Z(n13510) );
  XNOR2_X1 U15474 ( .A(n13309), .B(n13308), .ZN(n13508) );
  NAND2_X1 U15475 ( .A1(n13326), .A2(n13314), .ZN(n13310) );
  NAND3_X1 U15476 ( .A1(n13311), .A2(n13431), .A3(n13310), .ZN(n13505) );
  INV_X1 U15477 ( .A(n13312), .ZN(n13313) );
  OAI22_X1 U15478 ( .A1(n13504), .A2(n15320), .B1(n13313), .B2(n13397), .ZN(
        n13316) );
  INV_X1 U15479 ( .A(n13314), .ZN(n13506) );
  NOR2_X1 U15480 ( .A1(n13506), .A2(n13420), .ZN(n13315) );
  AOI211_X1 U15481 ( .C1(n15320), .C2(P2_REG2_REG_25__SCAN_IN), .A(n13316), 
        .B(n13315), .ZN(n13317) );
  OAI21_X1 U15482 ( .B1(n13440), .B2(n13505), .A(n13317), .ZN(n13318) );
  AOI21_X1 U15483 ( .B1(n13508), .B2(n13406), .A(n13318), .ZN(n13319) );
  OAI21_X1 U15484 ( .B1(n13510), .B2(n13465), .A(n13319), .ZN(P2_U3240) );
  XNOR2_X1 U15485 ( .A(n13321), .B(n13320), .ZN(n13517) );
  XNOR2_X1 U15486 ( .A(n13323), .B(n13322), .ZN(n13515) );
  AOI21_X1 U15487 ( .B1(n13332), .B2(n13324), .A(n13562), .ZN(n13325) );
  NAND2_X1 U15488 ( .A1(n13326), .A2(n13325), .ZN(n13512) );
  INV_X1 U15489 ( .A(n13511), .ZN(n13328) );
  AOI22_X1 U15490 ( .A1(n13328), .A2(n13472), .B1(n13327), .B2(n15318), .ZN(
        n13329) );
  OAI21_X1 U15491 ( .B1(n13330), .B2(n13472), .A(n13329), .ZN(n13331) );
  AOI21_X1 U15492 ( .B1(n13332), .B2(n13471), .A(n13331), .ZN(n13333) );
  OAI21_X1 U15493 ( .B1(n13512), .B2(n13440), .A(n13333), .ZN(n13334) );
  AOI21_X1 U15494 ( .B1(n13515), .B2(n13406), .A(n13334), .ZN(n13335) );
  OAI21_X1 U15495 ( .B1(n13517), .B2(n13465), .A(n13335), .ZN(P2_U3241) );
  XOR2_X1 U15496 ( .A(n13336), .B(n13342), .Z(n13522) );
  AOI211_X1 U15497 ( .C1(n13520), .C2(n13355), .A(n13562), .B(n13337), .ZN(
        n13519) );
  AOI22_X1 U15498 ( .A1(n15320), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13338), 
        .B2(n15318), .ZN(n13339) );
  OAI21_X1 U15499 ( .B1(n13340), .B2(n13420), .A(n13339), .ZN(n13341) );
  AOI21_X1 U15500 ( .B1(n13519), .B2(n13467), .A(n13341), .ZN(n13347) );
  XNOR2_X1 U15501 ( .A(n13343), .B(n13342), .ZN(n13345) );
  OAI21_X1 U15502 ( .B1(n13345), .B2(n13575), .A(n13344), .ZN(n13518) );
  NAND2_X1 U15503 ( .A1(n13518), .A2(n13472), .ZN(n13346) );
  OAI211_X1 U15504 ( .C1(n13522), .C2(n13465), .A(n13347), .B(n13346), .ZN(
        P2_U3242) );
  XOR2_X1 U15505 ( .A(n13352), .B(n13348), .Z(n13529) );
  INV_X1 U15506 ( .A(n13349), .ZN(n13350) );
  AOI21_X1 U15507 ( .B1(n13352), .B2(n13351), .A(n13350), .ZN(n13523) );
  INV_X1 U15508 ( .A(n13370), .ZN(n13353) );
  AOI21_X1 U15509 ( .B1(n13526), .B2(n13353), .A(n13562), .ZN(n13354) );
  AND2_X1 U15510 ( .A1(n13355), .A2(n13354), .ZN(n13524) );
  NAND2_X1 U15511 ( .A1(n13524), .A2(n13467), .ZN(n13360) );
  INV_X1 U15512 ( .A(n13525), .ZN(n13357) );
  OAI22_X1 U15513 ( .A1(n13357), .A2(n15320), .B1(n13356), .B2(n13397), .ZN(
        n13358) );
  AOI21_X1 U15514 ( .B1(P2_REG2_REG_22__SCAN_IN), .B2(n15320), .A(n13358), 
        .ZN(n13359) );
  OAI211_X1 U15515 ( .C1(n13361), .C2(n13420), .A(n13360), .B(n13359), .ZN(
        n13362) );
  AOI21_X1 U15516 ( .B1(n13523), .B2(n13469), .A(n13362), .ZN(n13363) );
  OAI21_X1 U15517 ( .B1(n13529), .B2(n13443), .A(n13363), .ZN(P2_U3243) );
  XNOR2_X1 U15518 ( .A(n13364), .B(n13365), .ZN(n13535) );
  XNOR2_X1 U15519 ( .A(n13366), .B(n13365), .ZN(n13533) );
  NAND2_X1 U15520 ( .A1(n13367), .A2(n13381), .ZN(n13368) );
  NAND2_X1 U15521 ( .A1(n13368), .A2(n13431), .ZN(n13369) );
  NOR2_X1 U15522 ( .A1(n13370), .A2(n13369), .ZN(n13532) );
  NAND2_X1 U15523 ( .A1(n13532), .A2(n13467), .ZN(n13375) );
  INV_X1 U15524 ( .A(n13371), .ZN(n13372) );
  OAI22_X1 U15525 ( .A1(n15320), .A2(n13530), .B1(n13372), .B2(n13397), .ZN(
        n13373) );
  AOI21_X1 U15526 ( .B1(P2_REG2_REG_21__SCAN_IN), .B2(n15320), .A(n13373), 
        .ZN(n13374) );
  OAI211_X1 U15527 ( .C1(n7433), .C2(n13420), .A(n13375), .B(n13374), .ZN(
        n13376) );
  AOI21_X1 U15528 ( .B1(n13533), .B2(n13469), .A(n13376), .ZN(n13377) );
  OAI21_X1 U15529 ( .B1(n13443), .B2(n13535), .A(n13377), .ZN(P2_U3244) );
  XOR2_X1 U15530 ( .A(n13378), .B(n13388), .Z(n13380) );
  AOI21_X1 U15531 ( .B1(n13380), .B2(n15409), .A(n13379), .ZN(n13539) );
  INV_X1 U15532 ( .A(n13396), .ZN(n13383) );
  INV_X1 U15533 ( .A(n13381), .ZN(n13382) );
  AOI211_X1 U15534 ( .C1(n13537), .C2(n13383), .A(n13562), .B(n13382), .ZN(
        n13536) );
  INV_X1 U15535 ( .A(n13384), .ZN(n13385) );
  AOI22_X1 U15536 ( .A1(n15320), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13385), 
        .B2(n15318), .ZN(n13386) );
  OAI21_X1 U15537 ( .B1(n13387), .B2(n13420), .A(n13386), .ZN(n13391) );
  XNOR2_X1 U15538 ( .A(n13389), .B(n13388), .ZN(n13540) );
  NOR2_X1 U15539 ( .A1(n13540), .A2(n13465), .ZN(n13390) );
  AOI211_X1 U15540 ( .C1(n13536), .C2(n13467), .A(n13391), .B(n13390), .ZN(
        n13392) );
  OAI21_X1 U15541 ( .B1(n15320), .B2(n13539), .A(n13392), .ZN(P2_U3245) );
  XOR2_X1 U15542 ( .A(n13393), .B(n13404), .Z(n13547) );
  NAND2_X1 U15543 ( .A1(n13543), .A2(n13414), .ZN(n13394) );
  NAND2_X1 U15544 ( .A1(n13394), .A2(n13431), .ZN(n13395) );
  NOR2_X1 U15545 ( .A1(n13396), .A2(n13395), .ZN(n13541) );
  INV_X1 U15546 ( .A(n13543), .ZN(n13402) );
  INV_X1 U15547 ( .A(n13542), .ZN(n13399) );
  OAI22_X1 U15548 ( .A1(n15320), .A2(n13399), .B1(n13398), .B2(n13397), .ZN(
        n13400) );
  AOI21_X1 U15549 ( .B1(P2_REG2_REG_19__SCAN_IN), .B2(n15320), .A(n13400), 
        .ZN(n13401) );
  OAI21_X1 U15550 ( .B1(n13402), .B2(n13420), .A(n13401), .ZN(n13403) );
  AOI21_X1 U15551 ( .B1(n13541), .B2(n13467), .A(n13403), .ZN(n13408) );
  XNOR2_X1 U15552 ( .A(n13405), .B(n13404), .ZN(n13544) );
  NAND2_X1 U15553 ( .A1(n13544), .A2(n13406), .ZN(n13407) );
  OAI211_X1 U15554 ( .C1(n13547), .C2(n13465), .A(n13408), .B(n13407), .ZN(
        P2_U3246) );
  AOI21_X1 U15555 ( .B1(n13410), .B2(n13409), .A(n13575), .ZN(n13413) );
  AOI21_X1 U15556 ( .B1(n13413), .B2(n13412), .A(n13411), .ZN(n13551) );
  INV_X1 U15557 ( .A(n13433), .ZN(n13416) );
  INV_X1 U15558 ( .A(n13414), .ZN(n13415) );
  AOI211_X1 U15559 ( .C1(n13549), .C2(n13416), .A(n13562), .B(n13415), .ZN(
        n13548) );
  INV_X1 U15560 ( .A(n13417), .ZN(n13418) );
  AOI22_X1 U15561 ( .A1(n15320), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13418), 
        .B2(n15318), .ZN(n13419) );
  OAI21_X1 U15562 ( .B1(n13421), .B2(n13420), .A(n13419), .ZN(n13426) );
  INV_X1 U15563 ( .A(n13422), .ZN(n13423) );
  AOI21_X1 U15564 ( .B1(n7160), .B2(n13424), .A(n13423), .ZN(n13552) );
  NOR2_X1 U15565 ( .A1(n13552), .A2(n13465), .ZN(n13425) );
  AOI211_X1 U15566 ( .C1(n13548), .C2(n13467), .A(n13426), .B(n13425), .ZN(
        n13427) );
  OAI21_X1 U15567 ( .B1(n15320), .B2(n13551), .A(n13427), .ZN(P2_U3247) );
  XNOR2_X1 U15568 ( .A(n13428), .B(n13430), .ZN(n13559) );
  XOR2_X1 U15569 ( .A(n13430), .B(n13429), .Z(n13557) );
  OAI21_X1 U15570 ( .B1(n13457), .B2(n13555), .A(n13431), .ZN(n13432) );
  OR2_X1 U15571 ( .A1(n13433), .A2(n13432), .ZN(n13554) );
  AOI22_X1 U15572 ( .A1(n13472), .A2(n13435), .B1(n13434), .B2(n15318), .ZN(
        n13436) );
  OAI21_X1 U15573 ( .B1(n11043), .B2(n13472), .A(n13436), .ZN(n13437) );
  AOI21_X1 U15574 ( .B1(n13438), .B2(n13471), .A(n13437), .ZN(n13439) );
  OAI21_X1 U15575 ( .B1(n13554), .B2(n13440), .A(n13439), .ZN(n13441) );
  AOI21_X1 U15576 ( .B1(n13557), .B2(n13469), .A(n13441), .ZN(n13442) );
  OAI21_X1 U15577 ( .B1(n13559), .B2(n13443), .A(n13442), .ZN(P2_U3248) );
  NAND2_X1 U15578 ( .A1(n13445), .A2(n13444), .ZN(n13446) );
  NAND2_X1 U15579 ( .A1(n13447), .A2(n13446), .ZN(n13560) );
  NAND2_X1 U15580 ( .A1(n13449), .A2(n13448), .ZN(n13450) );
  NAND2_X1 U15581 ( .A1(n13451), .A2(n13450), .ZN(n13452) );
  NAND2_X1 U15582 ( .A1(n13452), .A2(n15409), .ZN(n13454) );
  NAND2_X1 U15583 ( .A1(n13454), .A2(n13453), .ZN(n13566) );
  NOR2_X1 U15584 ( .A1(n13455), .A2(n13561), .ZN(n13456) );
  AOI22_X1 U15585 ( .A1(n13460), .A2(n13459), .B1(n13458), .B2(n15318), .ZN(
        n13461) );
  OAI21_X1 U15586 ( .B1(n13563), .B2(n9845), .A(n13461), .ZN(n13462) );
  OAI21_X1 U15587 ( .B1(n13566), .B2(n13462), .A(n13472), .ZN(n13464) );
  NAND2_X1 U15588 ( .A1(n15320), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13463) );
  OAI211_X1 U15589 ( .C1(n13560), .C2(n13465), .A(n13464), .B(n13463), .ZN(
        P2_U3249) );
  AOI22_X1 U15590 ( .A1(n13469), .A2(n13468), .B1(n13467), .B2(n13466), .ZN(
        n13477) );
  AOI22_X1 U15591 ( .A1(n13471), .A2(n13470), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n15318), .ZN(n13476) );
  MUX2_X1 U15592 ( .A(n13474), .B(n13473), .S(n13472), .Z(n13475) );
  NAND3_X1 U15593 ( .A1(n13477), .A2(n13476), .A3(n13475), .ZN(P2_U3264) );
  OAI211_X1 U15594 ( .C1(n13479), .C2(n15379), .A(n13478), .B(n13480), .ZN(
        n13860) );
  MUX2_X1 U15595 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13860), .S(n15443), .Z(
        P2_U3530) );
  OAI211_X1 U15596 ( .C1(n13482), .C2(n15379), .A(n13481), .B(n13480), .ZN(
        n13861) );
  MUX2_X1 U15597 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13861), .S(n15443), .Z(
        P2_U3529) );
  AOI21_X1 U15598 ( .B1(n15421), .B2(n13484), .A(n13483), .ZN(n13485) );
  MUX2_X1 U15599 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13862), .S(n15443), .Z(
        P2_U3528) );
  MUX2_X1 U15600 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13863), .S(n15443), .Z(
        P2_U3527) );
  AND2_X1 U15601 ( .A1(n13492), .A2(n13571), .ZN(n13497) );
  OAI21_X1 U15602 ( .B1(n7235), .B2(n15379), .A(n13494), .ZN(n13495) );
  MUX2_X1 U15603 ( .A(n13864), .B(P2_REG1_REG_27__SCAN_IN), .S(n15441), .Z(
        P2_U3526) );
  OAI211_X1 U15604 ( .C1(n7234), .C2(n15379), .A(n13499), .B(n13498), .ZN(
        n13500) );
  AOI21_X1 U15605 ( .B1(n13501), .B2(n15409), .A(n13500), .ZN(n13502) );
  OAI21_X1 U15606 ( .B1(n15405), .B2(n13503), .A(n13502), .ZN(n13865) );
  MUX2_X1 U15607 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13865), .S(n15443), .Z(
        P2_U3525) );
  OAI211_X1 U15608 ( .C1(n13506), .C2(n15379), .A(n13505), .B(n13504), .ZN(
        n13507) );
  AOI21_X1 U15609 ( .B1(n13508), .B2(n15409), .A(n13507), .ZN(n13509) );
  OAI21_X1 U15610 ( .B1(n13510), .B2(n15405), .A(n13509), .ZN(n13866) );
  MUX2_X1 U15611 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13866), .S(n15443), .Z(
        P2_U3524) );
  OAI211_X1 U15612 ( .C1(n13513), .C2(n15379), .A(n13512), .B(n13511), .ZN(
        n13514) );
  AOI21_X1 U15613 ( .B1(n13515), .B2(n15409), .A(n13514), .ZN(n13516) );
  OAI21_X1 U15614 ( .B1(n15405), .B2(n13517), .A(n13516), .ZN(n13867) );
  MUX2_X1 U15615 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13867), .S(n15443), .Z(
        P2_U3523) );
  AOI211_X1 U15616 ( .C1(n15421), .C2(n13520), .A(n13519), .B(n13518), .ZN(
        n13521) );
  OAI21_X1 U15617 ( .B1(n15405), .B2(n13522), .A(n13521), .ZN(n13868) );
  MUX2_X1 U15618 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13868), .S(n15443), .Z(
        P2_U3522) );
  NAND2_X1 U15619 ( .A1(n13523), .A2(n13571), .ZN(n13528) );
  AOI211_X1 U15620 ( .C1(n15421), .C2(n13526), .A(n13525), .B(n13524), .ZN(
        n13527) );
  OAI211_X1 U15621 ( .C1(n13575), .C2(n13529), .A(n13528), .B(n13527), .ZN(
        n13869) );
  MUX2_X1 U15622 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13869), .S(n15443), .Z(
        P2_U3521) );
  OAI21_X1 U15623 ( .B1(n7433), .B2(n15379), .A(n13530), .ZN(n13531) );
  AOI211_X1 U15624 ( .C1(n13533), .C2(n13571), .A(n13532), .B(n13531), .ZN(
        n13534) );
  OAI21_X1 U15625 ( .B1(n13575), .B2(n13535), .A(n13534), .ZN(n13870) );
  MUX2_X1 U15626 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13870), .S(n15443), .Z(
        P2_U3520) );
  AOI21_X1 U15627 ( .B1(n15421), .B2(n13537), .A(n13536), .ZN(n13538) );
  OAI211_X1 U15628 ( .C1(n15405), .C2(n13540), .A(n13539), .B(n13538), .ZN(
        n13871) );
  MUX2_X1 U15629 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13871), .S(n15443), .Z(
        P2_U3519) );
  AOI211_X1 U15630 ( .C1(n15421), .C2(n13543), .A(n13542), .B(n13541), .ZN(
        n13546) );
  NAND2_X1 U15631 ( .A1(n13544), .A2(n15409), .ZN(n13545) );
  OAI211_X1 U15632 ( .C1(n13547), .C2(n15405), .A(n13546), .B(n13545), .ZN(
        n13872) );
  MUX2_X1 U15633 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13872), .S(n15443), .Z(
        P2_U3518) );
  AOI21_X1 U15634 ( .B1(n15421), .B2(n13549), .A(n13548), .ZN(n13550) );
  OAI211_X1 U15635 ( .C1(n13552), .C2(n15405), .A(n13551), .B(n13550), .ZN(
        n13873) );
  MUX2_X1 U15636 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13873), .S(n15443), .Z(
        P2_U3517) );
  OAI211_X1 U15637 ( .C1(n13555), .C2(n15379), .A(n13554), .B(n13553), .ZN(
        n13556) );
  AOI21_X1 U15638 ( .B1(n13557), .B2(n13571), .A(n13556), .ZN(n13558) );
  OAI21_X1 U15639 ( .B1(n13575), .B2(n13559), .A(n13558), .ZN(n13874) );
  MUX2_X1 U15640 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13874), .S(n15443), .Z(
        P2_U3516) );
  NOR2_X1 U15641 ( .A1(n13560), .A2(n15405), .ZN(n13565) );
  OAI22_X1 U15642 ( .A1(n13563), .A2(n13562), .B1(n13561), .B2(n15379), .ZN(
        n13564) );
  MUX2_X1 U15643 ( .A(n13875), .B(P2_REG1_REG_16__SCAN_IN), .S(n15441), .Z(
        P2_U3515) );
  OAI21_X1 U15644 ( .B1(n13568), .B2(n15379), .A(n13567), .ZN(n13569) );
  AOI211_X1 U15645 ( .C1(n13572), .C2(n13571), .A(n13570), .B(n13569), .ZN(
        n13573) );
  OAI21_X1 U15646 ( .B1(n13575), .B2(n13574), .A(n13573), .ZN(n13876) );
  MUX2_X1 U15647 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13876), .S(n15443), .Z(
        P2_U3514) );
  AOI21_X1 U15648 ( .B1(n15421), .B2(n13577), .A(n13576), .ZN(n13578) );
  OAI211_X1 U15649 ( .C1(n15405), .C2(n13580), .A(n13579), .B(n13578), .ZN(
        n13877) );
  MUX2_X1 U15650 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13877), .S(n15443), .Z(
        P2_U3513) );
  AOI21_X1 U15651 ( .B1(n15421), .B2(n13582), .A(n13581), .ZN(n13583) );
  OAI211_X1 U15652 ( .C1(n15405), .C2(n13585), .A(n13584), .B(n13583), .ZN(
        n13878) );
  MUX2_X1 U15653 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13878), .S(n15443), .Z(
        n13852) );
  INV_X1 U15654 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15112) );
  AOI22_X1 U15655 ( .A1(n13801), .A2(keyinput56), .B1(keyinput110), .B2(n15112), .ZN(n13586) );
  OAI221_X1 U15656 ( .B1(n13801), .B2(keyinput56), .C1(n15112), .C2(
        keyinput110), .A(n13586), .ZN(n13595) );
  INV_X1 U15657 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14776) );
  AOI22_X1 U15658 ( .A1(n13588), .A2(keyinput65), .B1(keyinput63), .B2(n14776), 
        .ZN(n13587) );
  OAI221_X1 U15659 ( .B1(n13588), .B2(keyinput65), .C1(n14776), .C2(keyinput63), .A(n13587), .ZN(n13594) );
  INV_X1 U15660 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U15661 ( .A1(n15128), .A2(keyinput37), .B1(keyinput79), .B2(n10763), 
        .ZN(n13589) );
  OAI221_X1 U15662 ( .B1(n15128), .B2(keyinput37), .C1(n10763), .C2(keyinput79), .A(n13589), .ZN(n13593) );
  INV_X1 U15663 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14364) );
  AOI22_X1 U15664 ( .A1(n13591), .A2(keyinput104), .B1(keyinput39), .B2(n14364), .ZN(n13590) );
  OAI221_X1 U15665 ( .B1(n13591), .B2(keyinput104), .C1(n14364), .C2(
        keyinput39), .A(n13590), .ZN(n13592) );
  NOR4_X1 U15666 ( .A1(n13595), .A2(n13594), .A3(n13593), .A4(n13592), .ZN(
        n13625) );
  INV_X1 U15667 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15346) );
  AOI22_X1 U15668 ( .A1(n13597), .A2(keyinput48), .B1(keyinput8), .B2(n15346), 
        .ZN(n13596) );
  OAI221_X1 U15669 ( .B1(n13597), .B2(keyinput48), .C1(n15346), .C2(keyinput8), 
        .A(n13596), .ZN(n13604) );
  INV_X1 U15670 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15132) );
  AOI22_X1 U15671 ( .A1(n15341), .A2(keyinput66), .B1(keyinput16), .B2(n15132), 
        .ZN(n13598) );
  OAI221_X1 U15672 ( .B1(n15341), .B2(keyinput66), .C1(n15132), .C2(keyinput16), .A(n13598), .ZN(n13603) );
  INV_X1 U15673 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15133) );
  AOI22_X1 U15674 ( .A1(n15439), .A2(keyinput53), .B1(keyinput68), .B2(n15133), 
        .ZN(n13599) );
  OAI221_X1 U15675 ( .B1(n15439), .B2(keyinput53), .C1(n15133), .C2(keyinput68), .A(n13599), .ZN(n13602) );
  AOI22_X1 U15676 ( .A1(n15446), .A2(keyinput107), .B1(keyinput76), .B2(n7879), 
        .ZN(n13600) );
  OAI221_X1 U15677 ( .B1(n15446), .B2(keyinput107), .C1(n7879), .C2(keyinput76), .A(n13600), .ZN(n13601) );
  NOR4_X1 U15678 ( .A1(n13604), .A2(n13603), .A3(n13602), .A4(n13601), .ZN(
        n13624) );
  AOI22_X1 U15679 ( .A1(n13606), .A2(keyinput92), .B1(n15526), .B2(keyinput29), 
        .ZN(n13605) );
  OAI221_X1 U15680 ( .B1(n13606), .B2(keyinput92), .C1(n15526), .C2(keyinput29), .A(n13605), .ZN(n13614) );
  AOI22_X1 U15681 ( .A1(n13792), .A2(keyinput103), .B1(keyinput81), .B2(n13608), .ZN(n13607) );
  OAI221_X1 U15682 ( .B1(n13792), .B2(keyinput103), .C1(n13608), .C2(
        keyinput81), .A(n13607), .ZN(n13613) );
  INV_X1 U15683 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15119) );
  AOI22_X1 U15684 ( .A1(n13810), .A2(keyinput99), .B1(n15119), .B2(keyinput42), 
        .ZN(n13609) );
  OAI221_X1 U15685 ( .B1(n13810), .B2(keyinput99), .C1(n15119), .C2(keyinput42), .A(n13609), .ZN(n13612) );
  INV_X1 U15686 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n13610) );
  XNOR2_X1 U15687 ( .A(n13610), .B(keyinput80), .ZN(n13611) );
  NOR4_X1 U15688 ( .A1(n13614), .A2(n13613), .A3(n13612), .A4(n13611), .ZN(
        n13623) );
  INV_X1 U15689 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n13835) );
  AOI22_X1 U15690 ( .A1(n13835), .A2(keyinput31), .B1(keyinput64), .B2(n7993), 
        .ZN(n13615) );
  OAI221_X1 U15691 ( .B1(n13835), .B2(keyinput31), .C1(n7993), .C2(keyinput64), 
        .A(n13615), .ZN(n13621) );
  AOI22_X1 U15692 ( .A1(n9557), .A2(keyinput24), .B1(n9384), .B2(keyinput126), 
        .ZN(n13616) );
  OAI221_X1 U15693 ( .B1(n9557), .B2(keyinput24), .C1(n9384), .C2(keyinput126), 
        .A(n13616), .ZN(n13620) );
  XNOR2_X1 U15694 ( .A(n13617), .B(keyinput15), .ZN(n13619) );
  XNOR2_X1 U15695 ( .A(n15356), .B(keyinput30), .ZN(n13618) );
  NOR4_X1 U15696 ( .A1(n13621), .A2(n13620), .A3(n13619), .A4(n13618), .ZN(
        n13622) );
  NAND4_X1 U15697 ( .A1(n13625), .A2(n13624), .A3(n13623), .A4(n13622), .ZN(
        n13725) );
  INV_X1 U15698 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15130) );
  INV_X1 U15699 ( .A(keyinput46), .ZN(n13627) );
  AOI22_X1 U15700 ( .A1(n15130), .A2(keyinput38), .B1(P3_ADDR_REG_11__SCAN_IN), 
        .B2(n13627), .ZN(n13626) );
  OAI221_X1 U15701 ( .B1(n15130), .B2(keyinput38), .C1(n13627), .C2(
        P3_ADDR_REG_11__SCAN_IN), .A(n13626), .ZN(n13639) );
  INV_X1 U15702 ( .A(keyinput59), .ZN(n13629) );
  AOI22_X1 U15703 ( .A1(n13630), .A2(keyinput13), .B1(P3_DATAO_REG_31__SCAN_IN), .B2(n13629), .ZN(n13628) );
  OAI221_X1 U15704 ( .B1(n13630), .B2(keyinput13), .C1(n13629), .C2(
        P3_DATAO_REG_31__SCAN_IN), .A(n13628), .ZN(n13638) );
  INV_X1 U15705 ( .A(keyinput86), .ZN(n13632) );
  AOI22_X1 U15706 ( .A1(n13820), .A2(keyinput47), .B1(P1_ADDR_REG_12__SCAN_IN), 
        .B2(n13632), .ZN(n13631) );
  OAI221_X1 U15707 ( .B1(n13820), .B2(keyinput47), .C1(n13632), .C2(
        P1_ADDR_REG_12__SCAN_IN), .A(n13631), .ZN(n13637) );
  INV_X1 U15708 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n13635) );
  INV_X1 U15709 ( .A(keyinput111), .ZN(n13634) );
  AOI22_X1 U15710 ( .A1(n13635), .A2(keyinput27), .B1(P2_ADDR_REG_15__SCAN_IN), 
        .B2(n13634), .ZN(n13633) );
  OAI221_X1 U15711 ( .B1(n13635), .B2(keyinput27), .C1(n13634), .C2(
        P2_ADDR_REG_15__SCAN_IN), .A(n13633), .ZN(n13636) );
  NOR4_X1 U15712 ( .A1(n13639), .A2(n13638), .A3(n13637), .A4(n13636), .ZN(
        n13676) );
  AOI22_X1 U15713 ( .A1(n14806), .A2(keyinput2), .B1(n8008), .B2(keyinput82), 
        .ZN(n13640) );
  OAI221_X1 U15714 ( .B1(n14806), .B2(keyinput2), .C1(n8008), .C2(keyinput82), 
        .A(n13640), .ZN(n13651) );
  AOI22_X1 U15715 ( .A1(n14897), .A2(keyinput74), .B1(n13642), .B2(keyinput54), 
        .ZN(n13641) );
  OAI221_X1 U15716 ( .B1(n14897), .B2(keyinput74), .C1(n13642), .C2(keyinput54), .A(n13641), .ZN(n13650) );
  AOI22_X1 U15717 ( .A1(n13645), .A2(keyinput72), .B1(n13644), .B2(keyinput23), 
        .ZN(n13643) );
  OAI221_X1 U15718 ( .B1(n13645), .B2(keyinput72), .C1(n13644), .C2(keyinput23), .A(n13643), .ZN(n13649) );
  INV_X1 U15719 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15328) );
  INV_X1 U15720 ( .A(keyinput6), .ZN(n13647) );
  AOI22_X1 U15721 ( .A1(n15328), .A2(keyinput96), .B1(P3_DATAO_REG_3__SCAN_IN), 
        .B2(n13647), .ZN(n13646) );
  OAI221_X1 U15722 ( .B1(n15328), .B2(keyinput96), .C1(n13647), .C2(
        P3_DATAO_REG_3__SCAN_IN), .A(n13646), .ZN(n13648) );
  NOR4_X1 U15723 ( .A1(n13651), .A2(n13650), .A3(n13649), .A4(n13648), .ZN(
        n13675) );
  INV_X1 U15724 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14872) );
  AOI22_X1 U15725 ( .A1(n14872), .A2(keyinput1), .B1(n11427), .B2(keyinput124), 
        .ZN(n13652) );
  OAI221_X1 U15726 ( .B1(n14872), .B2(keyinput1), .C1(n11427), .C2(keyinput124), .A(n13652), .ZN(n13659) );
  INV_X1 U15727 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15126) );
  XNOR2_X1 U15728 ( .A(n15126), .B(keyinput112), .ZN(n13658) );
  XOR2_X1 U15729 ( .A(n8229), .B(keyinput88), .Z(n13656) );
  INV_X1 U15730 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15520) );
  XOR2_X1 U15731 ( .A(n15520), .B(keyinput51), .Z(n13655) );
  XNOR2_X1 U15732 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput84), .ZN(n13654) );
  XNOR2_X1 U15733 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput85), .ZN(n13653) );
  NAND4_X1 U15734 ( .A1(n13656), .A2(n13655), .A3(n13654), .A4(n13653), .ZN(
        n13657) );
  NOR3_X1 U15735 ( .A1(n13659), .A2(n13658), .A3(n13657), .ZN(n13674) );
  INV_X1 U15736 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U15737 ( .A1(n13662), .A2(keyinput20), .B1(keyinput95), .B2(n13661), 
        .ZN(n13660) );
  OAI221_X1 U15738 ( .B1(n13662), .B2(keyinput20), .C1(n13661), .C2(keyinput95), .A(n13660), .ZN(n13667) );
  AOI22_X1 U15739 ( .A1(n13783), .A2(keyinput71), .B1(n13782), .B2(keyinput36), 
        .ZN(n13663) );
  OAI221_X1 U15740 ( .B1(n13783), .B2(keyinput71), .C1(n13782), .C2(keyinput36), .A(n13663), .ZN(n13666) );
  XNOR2_X1 U15741 ( .A(keyinput123), .B(n7697), .ZN(n13665) );
  XNOR2_X1 U15742 ( .A(keyinput105), .B(n11207), .ZN(n13664) );
  OR4_X1 U15743 ( .A1(n13667), .A2(n13666), .A3(n13665), .A4(n13664), .ZN(
        n13672) );
  INV_X1 U15744 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13793) );
  INV_X1 U15745 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13795) );
  AOI22_X1 U15746 ( .A1(n13793), .A2(keyinput0), .B1(n13795), .B2(keyinput7), 
        .ZN(n13668) );
  OAI221_X1 U15747 ( .B1(n13793), .B2(keyinput0), .C1(n13795), .C2(keyinput7), 
        .A(n13668), .ZN(n13671) );
  AOI22_X1 U15748 ( .A1(n14760), .A2(keyinput22), .B1(n7766), .B2(keyinput108), 
        .ZN(n13669) );
  OAI221_X1 U15749 ( .B1(n14760), .B2(keyinput22), .C1(n7766), .C2(keyinput108), .A(n13669), .ZN(n13670) );
  NOR3_X1 U15750 ( .A1(n13672), .A2(n13671), .A3(n13670), .ZN(n13673) );
  NAND4_X1 U15751 ( .A1(n13676), .A2(n13675), .A3(n13674), .A4(n13673), .ZN(
        n13724) );
  XOR2_X1 U15752 ( .A(keyinput28), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n13679) );
  INV_X1 U15753 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15123) );
  AOI22_X1 U15754 ( .A1(n9564), .A2(keyinput113), .B1(n15123), .B2(keyinput57), 
        .ZN(n13677) );
  OAI221_X1 U15755 ( .B1(n9564), .B2(keyinput113), .C1(n15123), .C2(keyinput57), .A(n13677), .ZN(n13678) );
  AOI211_X1 U15756 ( .C1(n9218), .C2(keyinput34), .A(n13679), .B(n13678), .ZN(
        n13680) );
  OAI21_X1 U15757 ( .B1(n9218), .B2(keyinput34), .A(n13680), .ZN(n13723) );
  AOI22_X1 U15758 ( .A1(n8423), .A2(keyinput17), .B1(keyinput70), .B2(n10604), 
        .ZN(n13681) );
  OAI221_X1 U15759 ( .B1(n8423), .B2(keyinput17), .C1(n10604), .C2(keyinput70), 
        .A(n13681), .ZN(n13706) );
  INV_X1 U15760 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15111) );
  AOI22_X1 U15761 ( .A1(n15111), .A2(keyinput125), .B1(keyinput102), .B2(
        n13683), .ZN(n13682) );
  OAI221_X1 U15762 ( .B1(n15111), .B2(keyinput125), .C1(n13683), .C2(
        keyinput102), .A(n13682), .ZN(n13699) );
  XNOR2_X1 U15763 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput45), .ZN(n13687) );
  XNOR2_X1 U15764 ( .A(P2_REG0_REG_19__SCAN_IN), .B(keyinput33), .ZN(n13686)
         );
  XNOR2_X1 U15765 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput100), .ZN(n13685) );
  XNOR2_X1 U15766 ( .A(SI_16_), .B(keyinput106), .ZN(n13684) );
  NAND4_X1 U15767 ( .A1(n13687), .A2(n13686), .A3(n13685), .A4(n13684), .ZN(
        n13698) );
  XNOR2_X1 U15768 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput75), .ZN(n13691) );
  XNOR2_X1 U15769 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput62), .ZN(n13690) );
  XNOR2_X1 U15770 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput73), .ZN(n13689) );
  XNOR2_X1 U15771 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput55), .ZN(n13688) );
  NAND4_X1 U15772 ( .A1(n13691), .A2(n13690), .A3(n13689), .A4(n13688), .ZN(
        n13697) );
  XNOR2_X1 U15773 ( .A(P3_REG1_REG_1__SCAN_IN), .B(keyinput61), .ZN(n13695) );
  XNOR2_X1 U15774 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput97), .ZN(n13694) );
  XNOR2_X1 U15775 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput25), .ZN(n13693) );
  XNOR2_X1 U15776 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput4), .ZN(n13692) );
  NAND4_X1 U15777 ( .A1(n13695), .A2(n13694), .A3(n13693), .A4(n13692), .ZN(
        n13696) );
  OR4_X1 U15778 ( .A1(n13699), .A2(n13698), .A3(n13697), .A4(n13696), .ZN(
        n13705) );
  AOI22_X1 U15779 ( .A1(n13701), .A2(keyinput118), .B1(n13776), .B2(
        keyinput115), .ZN(n13700) );
  OAI221_X1 U15780 ( .B1(n13701), .B2(keyinput118), .C1(n13776), .C2(
        keyinput115), .A(n13700), .ZN(n13704) );
  INV_X1 U15781 ( .A(keyinput78), .ZN(n13702) );
  XNOR2_X1 U15782 ( .A(n13702), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n13703) );
  NOR4_X1 U15783 ( .A1(n13706), .A2(n13705), .A3(n13704), .A4(n13703), .ZN(
        n13721) );
  XNOR2_X1 U15784 ( .A(n15342), .B(keyinput52), .ZN(n13717) );
  XNOR2_X1 U15785 ( .A(SI_2_), .B(keyinput9), .ZN(n13710) );
  XNOR2_X1 U15786 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput19), .ZN(n13709) );
  XNOR2_X1 U15787 ( .A(P1_REG3_REG_28__SCAN_IN), .B(keyinput114), .ZN(n13708)
         );
  XNOR2_X1 U15788 ( .A(P2_REG0_REG_21__SCAN_IN), .B(keyinput127), .ZN(n13707)
         );
  NAND4_X1 U15789 ( .A1(n13710), .A2(n13709), .A3(n13708), .A4(n13707), .ZN(
        n13716) );
  XNOR2_X1 U15790 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput40), .ZN(n13714) );
  XNOR2_X1 U15791 ( .A(P3_IR_REG_22__SCAN_IN), .B(keyinput83), .ZN(n13713) );
  XNOR2_X1 U15792 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput5), .ZN(n13712) );
  XNOR2_X1 U15793 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput119), .ZN(n13711) );
  NAND4_X1 U15794 ( .A1(n13714), .A2(n13713), .A3(n13712), .A4(n13711), .ZN(
        n13715) );
  NOR3_X1 U15795 ( .A1(n13717), .A2(n13716), .A3(n13715), .ZN(n13720) );
  INV_X1 U15796 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15125) );
  XOR2_X1 U15797 ( .A(keyinput117), .B(n15125), .Z(n13719) );
  XOR2_X1 U15798 ( .A(keyinput122), .B(n14791), .Z(n13718) );
  NAND4_X1 U15799 ( .A1(n13721), .A2(n13720), .A3(n13719), .A4(n13718), .ZN(
        n13722) );
  NOR4_X1 U15800 ( .A1(n13725), .A2(n13724), .A3(n13723), .A4(n13722), .ZN(
        n13775) );
  AOI22_X1 U15801 ( .A1(n13794), .A2(keyinput12), .B1(keyinput91), .B2(n13727), 
        .ZN(n13726) );
  OAI221_X1 U15802 ( .B1(n13794), .B2(keyinput12), .C1(n13727), .C2(keyinput91), .A(n13726), .ZN(n13736) );
  INV_X1 U15803 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U15804 ( .A1(n15322), .A2(keyinput69), .B1(keyinput21), .B2(n9763), 
        .ZN(n13728) );
  OAI221_X1 U15805 ( .B1(n15322), .B2(keyinput69), .C1(n9763), .C2(keyinput21), 
        .A(n13728), .ZN(n13735) );
  AOI22_X1 U15806 ( .A1(n15348), .A2(keyinput121), .B1(keyinput58), .B2(n13730), .ZN(n13729) );
  OAI221_X1 U15807 ( .B1(n15348), .B2(keyinput121), .C1(n13730), .C2(
        keyinput58), .A(n13729), .ZN(n13734) );
  AOI22_X1 U15808 ( .A1(n13732), .A2(keyinput93), .B1(n9584), .B2(keyinput67), 
        .ZN(n13731) );
  OAI221_X1 U15809 ( .B1(n13732), .B2(keyinput93), .C1(n9584), .C2(keyinput67), 
        .A(n13731), .ZN(n13733) );
  NOR4_X1 U15810 ( .A1(n13736), .A2(n13735), .A3(n13734), .A4(n13733), .ZN(
        n13774) );
  INV_X1 U15811 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14080) );
  AOI22_X1 U15812 ( .A1(n13738), .A2(keyinput18), .B1(keyinput94), .B2(n14080), 
        .ZN(n13737) );
  OAI221_X1 U15813 ( .B1(n13738), .B2(keyinput18), .C1(n14080), .C2(keyinput94), .A(n13737), .ZN(n13748) );
  INV_X1 U15814 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U15815 ( .A1(n15129), .A2(keyinput90), .B1(n13740), .B2(keyinput87), 
        .ZN(n13739) );
  OAI221_X1 U15816 ( .B1(n15129), .B2(keyinput90), .C1(n13740), .C2(keyinput87), .A(n13739), .ZN(n13747) );
  AOI22_X1 U15817 ( .A1(n13973), .A2(keyinput43), .B1(keyinput116), .B2(n13742), .ZN(n13741) );
  AOI22_X1 U15818 ( .A1(n13744), .A2(keyinput11), .B1(keyinput32), .B2(n11035), 
        .ZN(n13743) );
  OAI221_X1 U15819 ( .B1(n13744), .B2(keyinput11), .C1(n11035), .C2(keyinput32), .A(n13743), .ZN(n13745) );
  NOR4_X1 U15820 ( .A1(n13748), .A2(n13747), .A3(n13746), .A4(n13745), .ZN(
        n13772) );
  AOI22_X1 U15821 ( .A1(n13797), .A2(keyinput3), .B1(n8419), .B2(keyinput109), 
        .ZN(n13749) );
  OAI221_X1 U15822 ( .B1(n13797), .B2(keyinput3), .C1(n8419), .C2(keyinput109), 
        .A(n13749), .ZN(n13757) );
  INV_X1 U15823 ( .A(keyinput41), .ZN(n13751) );
  AOI22_X1 U15824 ( .A1(n14750), .A2(keyinput44), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n13751), .ZN(n13750) );
  OAI221_X1 U15825 ( .B1(n14750), .B2(keyinput44), .C1(n13751), .C2(
        P1_ADDR_REG_15__SCAN_IN), .A(n13750), .ZN(n13756) );
  INV_X1 U15826 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15338) );
  AOI22_X1 U15827 ( .A1(n15338), .A2(keyinput98), .B1(keyinput50), .B2(n13796), 
        .ZN(n13752) );
  OAI221_X1 U15828 ( .B1(n15338), .B2(keyinput98), .C1(n13796), .C2(keyinput50), .A(n13752), .ZN(n13755) );
  INV_X1 U15829 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13815) );
  AOI22_X1 U15830 ( .A1(n15345), .A2(keyinput77), .B1(keyinput35), .B2(n13815), 
        .ZN(n13753) );
  OAI221_X1 U15831 ( .B1(n15345), .B2(keyinput77), .C1(n13815), .C2(keyinput35), .A(n13753), .ZN(n13754) );
  NOR4_X1 U15832 ( .A1(n13757), .A2(n13756), .A3(n13755), .A4(n13754), .ZN(
        n13771) );
  INV_X1 U15833 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n13759) );
  AOI22_X1 U15834 ( .A1(n13759), .A2(keyinput120), .B1(keyinput101), .B2(n9562), .ZN(n13758) );
  OAI221_X1 U15835 ( .B1(n13759), .B2(keyinput120), .C1(n9562), .C2(
        keyinput101), .A(n13758), .ZN(n13769) );
  INV_X1 U15836 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n13824) );
  AOI22_X1 U15837 ( .A1(n13761), .A2(keyinput10), .B1(n13824), .B2(keyinput26), 
        .ZN(n13760) );
  OAI221_X1 U15838 ( .B1(n13761), .B2(keyinput10), .C1(n13824), .C2(keyinput26), .A(n13760), .ZN(n13768) );
  AOI22_X1 U15839 ( .A1(n13763), .A2(keyinput14), .B1(keyinput60), .B2(n13829), 
        .ZN(n13762) );
  OAI221_X1 U15840 ( .B1(n13763), .B2(keyinput14), .C1(n13829), .C2(keyinput60), .A(n13762), .ZN(n13767) );
  INV_X1 U15841 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n13825) );
  INV_X1 U15842 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n13765) );
  AOI22_X1 U15843 ( .A1(n13825), .A2(keyinput89), .B1(n13765), .B2(keyinput49), 
        .ZN(n13764) );
  OAI221_X1 U15844 ( .B1(n13825), .B2(keyinput89), .C1(n13765), .C2(keyinput49), .A(n13764), .ZN(n13766) );
  NOR4_X1 U15845 ( .A1(n13769), .A2(n13768), .A3(n13767), .A4(n13766), .ZN(
        n13770) );
  AND3_X1 U15846 ( .A1(n13772), .A2(n13771), .A3(n13770), .ZN(n13773) );
  NAND3_X1 U15847 ( .A1(n13775), .A2(n13774), .A3(n13773), .ZN(n13850) );
  NOR4_X1 U15848 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .A3(P3_DATAO_REG_30__SCAN_IN), .A4(n13776), .ZN(n13777) );
  NAND3_X1 U15849 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), 
        .A3(n13777), .ZN(n13791) );
  NAND4_X1 U15850 ( .A1(P1_REG0_REG_30__SCAN_IN), .A2(P3_DATAO_REG_1__SCAN_IN), 
        .A3(n13778), .A4(n9564), .ZN(n13779) );
  NOR3_X1 U15851 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_REG0_REG_10__SCAN_IN), 
        .A3(n13779), .ZN(n13789) );
  NAND4_X1 U15852 ( .A1(P3_REG1_REG_24__SCAN_IN), .A2(P1_DATAO_REG_22__SCAN_IN), .A3(P1_D_REG_9__SCAN_IN), .A4(n14080), .ZN(n13787) );
  INV_X1 U15853 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13780) );
  NAND4_X1 U15854 ( .A1(P2_REG1_REG_2__SCAN_IN), .A2(P2_REG1_REG_1__SCAN_IN), 
        .A3(n13780), .A4(n15439), .ZN(n13781) );
  NOR2_X1 U15855 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(n13781), .ZN(n13784) );
  NAND4_X1 U15856 ( .A1(n13784), .A2(P1_D_REG_5__SCAN_IN), .A3(n13783), .A4(
        n13782), .ZN(n13786) );
  NAND4_X1 U15857 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P2_REG1_REG_31__SCAN_IN), 
        .A3(P1_ADDR_REG_13__SCAN_IN), .A4(P2_ADDR_REG_8__SCAN_IN), .ZN(n13785)
         );
  NOR3_X1 U15858 ( .A1(n13787), .A2(n13786), .A3(n13785), .ZN(n13788) );
  NAND4_X1 U15859 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_REG1_REG_4__SCAN_IN), 
        .A3(n13789), .A4(n13788), .ZN(n13790) );
  NOR4_X1 U15860 ( .A1(P2_REG0_REG_25__SCAN_IN), .A2(n13792), .A3(n13791), 
        .A4(n13790), .ZN(n13848) );
  NAND4_X1 U15861 ( .A1(SI_15_), .A2(n13795), .A3(n13794), .A4(n13793), .ZN(
        n13809) );
  NAND4_X1 U15862 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_REG2_REG_9__SCAN_IN), 
        .A3(P1_REG3_REG_17__SCAN_IN), .A4(P1_REG0_REG_0__SCAN_IN), .ZN(n13808)
         );
  NOR4_X1 U15863 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P2_DATAO_REG_26__SCAN_IN), 
        .A3(P1_ADDR_REG_15__SCAN_IN), .A4(n13796), .ZN(n13798) );
  NAND4_X1 U15864 ( .A1(n13799), .A2(P3_ADDR_REG_10__SCAN_IN), .A3(n13798), 
        .A4(n13797), .ZN(n13807) );
  NOR4_X1 U15865 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(SI_18_), .A3(
        P1_REG3_REG_28__SCAN_IN), .A4(P1_REG2_REG_1__SCAN_IN), .ZN(n13805) );
  NOR4_X1 U15866 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P1_REG1_REG_24__SCAN_IN), 
        .A3(P1_REG2_REG_4__SCAN_IN), .A4(n13800), .ZN(n13804) );
  NOR4_X1 U15867 ( .A1(n15112), .A2(n13801), .A3(n15130), .A4(
        P1_REG2_REG_23__SCAN_IN), .ZN(n13803) );
  NOR4_X1 U15868 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(P3_DATAO_REG_31__SCAN_IN), 
        .A3(P3_ADDR_REG_11__SCAN_IN), .A4(n9557), .ZN(n13802) );
  NAND4_X1 U15869 ( .A1(n13805), .A2(n13804), .A3(n13803), .A4(n13802), .ZN(
        n13806) );
  NOR4_X1 U15870 ( .A1(n13809), .A2(n13808), .A3(n13807), .A4(n13806), .ZN(
        n13847) );
  NAND4_X1 U15871 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .A3(n15119), .A4(n13810), .ZN(n13812) );
  NAND4_X1 U15872 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n13811) );
  OR3_X1 U15873 ( .A1(n13812), .A2(n13811), .A3(P3_DATAO_REG_21__SCAN_IN), 
        .ZN(n13819) );
  NAND4_X1 U15874 ( .A1(P3_REG1_REG_1__SCAN_IN), .A2(P1_REG1_REG_16__SCAN_IN), 
        .A3(P3_DATAO_REG_3__SCAN_IN), .A4(n7697), .ZN(n13818) );
  INV_X1 U15875 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n13813) );
  NAND4_X1 U15876 ( .A1(n13814), .A2(n13813), .A3(P2_IR_REG_18__SCAN_IN), .A4(
        P2_IR_REG_9__SCAN_IN), .ZN(n13817) );
  NAND4_X1 U15877 ( .A1(n13815), .A2(P2_REG2_REG_13__SCAN_IN), .A3(
        P2_REG3_REG_13__SCAN_IN), .A4(P2_REG1_REG_10__SCAN_IN), .ZN(n13816) );
  NOR4_X1 U15878 ( .A1(n13819), .A2(n13818), .A3(n13817), .A4(n13816), .ZN(
        n13845) );
  NAND4_X1 U15879 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG0_REG_26__SCAN_IN), 
        .A3(P1_REG2_REG_13__SCAN_IN), .A4(n15520), .ZN(n13823) );
  NAND4_X1 U15880 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(n13821), .A3(n14897), 
        .A4(n13820), .ZN(n13822) );
  NOR2_X1 U15881 ( .A1(n13823), .A2(n13822), .ZN(n13826) );
  NAND4_X1 U15882 ( .A1(n13826), .A2(n14806), .A3(n13825), .A4(n13824), .ZN(
        n13827) );
  NOR2_X1 U15883 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(n13827), .ZN(n13828) );
  NAND4_X1 U15884 ( .A1(n13828), .A2(P1_ADDR_REG_8__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n13834) );
  NAND4_X1 U15885 ( .A1(n13830), .A2(n13829), .A3(n14352), .A4(
        P1_REG2_REG_12__SCAN_IN), .ZN(n13833) );
  NAND4_X1 U15886 ( .A1(n13831), .A2(P2_DATAO_REG_28__SCAN_IN), .A3(
        P2_DATAO_REG_6__SCAN_IN), .A4(P3_IR_REG_10__SCAN_IN), .ZN(n13832) );
  NOR3_X1 U15887 ( .A1(n13834), .A2(n13833), .A3(n13832), .ZN(n13840) );
  NAND4_X1 U15888 ( .A1(n8423), .A2(n10604), .A3(n13835), .A4(n7993), .ZN(
        n13837) );
  NAND4_X1 U15889 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .A3(P2_ADDR_REG_2__SCAN_IN), .A4(n14760), .ZN(n13836) );
  NOR2_X1 U15890 ( .A1(n13837), .A2(n13836), .ZN(n13839) );
  AND4_X1 U15891 ( .A1(n13840), .A2(n13839), .A3(n15356), .A4(n13838), .ZN(
        n13844) );
  INV_X1 U15892 ( .A(n13841), .ZN(n13842) );
  AND4_X1 U15893 ( .A1(n13845), .A2(n13844), .A3(n13843), .A4(n13842), .ZN(
        n13846) );
  NAND3_X1 U15894 ( .A1(n13848), .A2(n13847), .A3(n13846), .ZN(n13849) );
  XNOR2_X1 U15895 ( .A(n13850), .B(n13849), .ZN(n13851) );
  XNOR2_X1 U15896 ( .A(n13852), .B(n13851), .ZN(P2_U3512) );
  AOI211_X1 U15897 ( .C1(n15421), .C2(n13855), .A(n13854), .B(n13853), .ZN(
        n13858) );
  NAND2_X1 U15898 ( .A1(n13856), .A2(n15409), .ZN(n13857) );
  OAI211_X1 U15899 ( .C1(n13859), .C2(n15405), .A(n13858), .B(n13857), .ZN(
        n13879) );
  MUX2_X1 U15900 ( .A(n13879), .B(P2_REG1_REG_12__SCAN_IN), .S(n15441), .Z(
        P2_U3511) );
  MUX2_X1 U15901 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13860), .S(n15431), .Z(
        P2_U3498) );
  MUX2_X1 U15902 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13861), .S(n15431), .Z(
        P2_U3497) );
  MUX2_X1 U15903 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13862), .S(n15431), .Z(
        P2_U3496) );
  MUX2_X1 U15904 ( .A(n13864), .B(P2_REG0_REG_27__SCAN_IN), .S(n15429), .Z(
        P2_U3494) );
  MUX2_X1 U15905 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13865), .S(n15431), .Z(
        P2_U3493) );
  MUX2_X1 U15906 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13866), .S(n15431), .Z(
        P2_U3492) );
  MUX2_X1 U15907 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13867), .S(n15431), .Z(
        P2_U3491) );
  MUX2_X1 U15908 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13868), .S(n15431), .Z(
        P2_U3490) );
  MUX2_X1 U15909 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13869), .S(n15431), .Z(
        P2_U3489) );
  MUX2_X1 U15910 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13870), .S(n15431), .Z(
        P2_U3488) );
  MUX2_X1 U15911 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13871), .S(n15431), .Z(
        P2_U3487) );
  MUX2_X1 U15912 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13872), .S(n15431), .Z(
        P2_U3486) );
  MUX2_X1 U15913 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13873), .S(n15431), .Z(
        P2_U3484) );
  MUX2_X1 U15914 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13874), .S(n15431), .Z(
        P2_U3481) );
  MUX2_X1 U15915 ( .A(n13875), .B(P2_REG0_REG_16__SCAN_IN), .S(n15429), .Z(
        P2_U3478) );
  MUX2_X1 U15916 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13876), .S(n15431), .Z(
        P2_U3475) );
  MUX2_X1 U15917 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13877), .S(n15431), .Z(
        P2_U3472) );
  MUX2_X1 U15918 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13878), .S(n15431), .Z(
        P2_U3469) );
  MUX2_X1 U15919 ( .A(n13879), .B(P2_REG0_REG_12__SCAN_IN), .S(n15429), .Z(
        P2_U3466) );
  INV_X1 U15920 ( .A(n14088), .ZN(n14741) );
  NOR4_X1 U15921 ( .A1(n13880), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13881), .A4(
        P2_U3088), .ZN(n13882) );
  AOI21_X1 U15922 ( .B1(n13890), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13882), 
        .ZN(n13883) );
  OAI21_X1 U15923 ( .B1(n14741), .B2(n13908), .A(n13883), .ZN(P2_U3296) );
  OAI222_X1 U15924 ( .A1(n13908), .A2(n14744), .B1(P2_U3088), .B2(n9285), .C1(
        n13884), .C2(n13905), .ZN(P2_U3297) );
  INV_X1 U15925 ( .A(n13885), .ZN(n14747) );
  OAI222_X1 U15926 ( .A1(n13908), .A2(n14747), .B1(P2_U3088), .B2(n13887), 
        .C1(n13886), .C2(n13905), .ZN(P2_U3298) );
  AOI21_X1 U15927 ( .B1(n13890), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13889), 
        .ZN(n13891) );
  OAI21_X1 U15928 ( .B1(n13892), .B2(n13908), .A(n13891), .ZN(P2_U3299) );
  NAND2_X1 U15929 ( .A1(n13894), .A2(n13893), .ZN(n13896) );
  OAI211_X1 U15930 ( .C1(n13905), .C2(n13897), .A(n13896), .B(n13895), .ZN(
        P2_U3300) );
  INV_X1 U15931 ( .A(n13898), .ZN(n14749) );
  OAI222_X1 U15932 ( .A1(n13900), .A2(P2_U3088), .B1(n13908), .B2(n14749), 
        .C1(n13899), .C2(n13905), .ZN(P2_U3301) );
  INV_X1 U15933 ( .A(n13901), .ZN(n14752) );
  OAI222_X1 U15934 ( .A1(n13905), .A2(n13903), .B1(n13908), .B2(n14752), .C1(
        n13902), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15935 ( .A(n13904), .ZN(n13909) );
  OAI222_X1 U15936 ( .A1(n13909), .A2(P2_U3088), .B1(n13908), .B2(n13907), 
        .C1(n13906), .C2(n13905), .ZN(P2_U3303) );
  INV_X1 U15937 ( .A(n13910), .ZN(n13912) );
  MUX2_X1 U15938 ( .A(n13912), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15939 ( .A(n14026), .ZN(n14071) );
  INV_X1 U15940 ( .A(n13915), .ZN(n14445) );
  AOI22_X1 U15941 ( .A1(n14316), .A2(n15059), .B1(n14554), .B2(n14318), .ZN(
        n14439) );
  INV_X1 U15942 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13916) );
  OAI22_X1 U15943 ( .A1(n14439), .A2(n14055), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13916), .ZN(n13917) );
  AOI21_X1 U15944 ( .B1(n14071), .B2(n14445), .A(n13917), .ZN(n13918) );
  AOI21_X1 U15945 ( .B1(n13921), .B2(n13920), .A(n6901), .ZN(n13929) );
  INV_X1 U15946 ( .A(n14064), .ZN(n13955) );
  NAND2_X1 U15947 ( .A1(n14071), .A2(n13922), .ZN(n13925) );
  AOI21_X1 U15948 ( .B1(n14023), .B2(n14324), .A(n13923), .ZN(n13924) );
  OAI211_X1 U15949 ( .C1(n13926), .C2(n13955), .A(n13925), .B(n13924), .ZN(
        n13927) );
  AOI21_X1 U15950 ( .B1(n14952), .B2(n9398), .A(n13927), .ZN(n13928) );
  OAI21_X1 U15951 ( .B1(n13929), .B2(n14074), .A(n13928), .ZN(P1_U3215) );
  AOI22_X1 U15952 ( .A1(n14023), .A2(n14512), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13931) );
  NAND2_X1 U15953 ( .A1(n14064), .A2(n6940), .ZN(n13930) );
  OAI211_X1 U15954 ( .C1(n14026), .C2(n14516), .A(n13931), .B(n13930), .ZN(
        n13938) );
  NAND3_X1 U15955 ( .A1(n13933), .A2(n13935), .A3(n7641), .ZN(n13936) );
  AOI21_X1 U15956 ( .B1(n13932), .B2(n13936), .A(n14074), .ZN(n13937) );
  AOI211_X1 U15957 ( .C1(n14668), .C2(n9398), .A(n13938), .B(n13937), .ZN(
        n13939) );
  INV_X1 U15958 ( .A(n13939), .ZN(P1_U3216) );
  OAI211_X1 U15959 ( .C1(n13942), .C2(n13941), .A(n13940), .B(n14052), .ZN(
        n13947) );
  AOI22_X1 U15960 ( .A1(n14116), .A2(n9398), .B1(n14064), .B2(n14336), .ZN(
        n13946) );
  NOR2_X1 U15961 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13943), .ZN(n14366) );
  NOR2_X1 U15962 ( .A1(n14026), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13944) );
  AOI211_X1 U15963 ( .C1(n14023), .C2(n14334), .A(n14366), .B(n13944), .ZN(
        n13945) );
  NAND3_X1 U15964 ( .A1(n13947), .A2(n13946), .A3(n13945), .ZN(P1_U3218) );
  INV_X1 U15965 ( .A(n14581), .ZN(n14698) );
  AND2_X1 U15966 ( .A1(n13948), .A2(n13949), .ZN(n13952) );
  OAI211_X1 U15967 ( .C1(n13952), .C2(n13951), .A(n14052), .B(n13950), .ZN(
        n13959) );
  NAND2_X1 U15968 ( .A1(n14577), .A2(n14023), .ZN(n13954) );
  OAI211_X1 U15969 ( .C1(n13955), .C2(n14609), .A(n13954), .B(n13953), .ZN(
        n13956) );
  AOI21_X1 U15970 ( .B1(n13957), .B2(n14071), .A(n13956), .ZN(n13958) );
  OAI211_X1 U15971 ( .C1(n14698), .C2(n14067), .A(n13959), .B(n13958), .ZN(
        P1_U3219) );
  NOR2_X1 U15972 ( .A1(n13961), .A2(n13960), .ZN(n13963) );
  OAI21_X1 U15973 ( .B1(n13963), .B2(n13962), .A(n14052), .ZN(n13968) );
  AOI22_X1 U15974 ( .A1(n14023), .A2(n14336), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n13964), .ZN(n13967) );
  AOI22_X1 U15975 ( .A1(n13965), .A2(n9398), .B1(n14064), .B2(n14338), .ZN(
        n13966) );
  NAND3_X1 U15976 ( .A1(n13968), .A2(n13967), .A3(n13966), .ZN(P1_U3222) );
  INV_X1 U15977 ( .A(n13969), .ZN(n14033) );
  AOI21_X1 U15978 ( .B1(n13971), .B2(n13970), .A(n14033), .ZN(n13977) );
  NOR2_X1 U15979 ( .A1(n14026), .A2(n14538), .ZN(n13975) );
  NOR2_X1 U15980 ( .A1(n14216), .A2(n14608), .ZN(n13972) );
  AOI21_X1 U15981 ( .B1(n14577), .B2(n14554), .A(n13972), .ZN(n14534) );
  OAI22_X1 U15982 ( .A1(n14534), .A2(n14055), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13973), .ZN(n13974) );
  AOI211_X1 U15983 ( .C1(n14682), .C2(n9398), .A(n13975), .B(n13974), .ZN(
        n13976) );
  OAI21_X1 U15984 ( .B1(n13977), .B2(n14074), .A(n13976), .ZN(P1_U3223) );
  AOI22_X1 U15985 ( .A1(n14023), .A2(n14318), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13979) );
  NAND2_X1 U15986 ( .A1(n14064), .A2(n14512), .ZN(n13978) );
  OAI211_X1 U15987 ( .C1(n14026), .C2(n14479), .A(n13979), .B(n13978), .ZN(
        n13986) );
  NAND3_X1 U15988 ( .A1(n13980), .A2(n13982), .A3(n7646), .ZN(n13983) );
  AOI21_X1 U15989 ( .B1(n13984), .B2(n13983), .A(n14074), .ZN(n13985) );
  INV_X1 U15990 ( .A(n13987), .ZN(P1_U3225) );
  OAI21_X1 U15991 ( .B1(n13990), .B2(n13989), .A(n13988), .ZN(n13991) );
  NAND2_X1 U15992 ( .A1(n13991), .A2(n14052), .ZN(n13998) );
  NOR2_X1 U15993 ( .A1(n14026), .A2(n13992), .ZN(n13996) );
  OAI21_X1 U15994 ( .B1(n14066), .B2(n13994), .A(n13993), .ZN(n13995) );
  AOI211_X1 U15995 ( .C1(n14064), .C2(n14324), .A(n13996), .B(n13995), .ZN(
        n13997) );
  OAI211_X1 U15996 ( .C1(n7633), .C2(n14067), .A(n13998), .B(n13997), .ZN(
        P1_U3226) );
  INV_X1 U15997 ( .A(n14710), .ZN(n14011) );
  INV_X1 U15998 ( .A(n13988), .ZN(n14001) );
  NOR3_X1 U15999 ( .A1(n14001), .A2(n14000), .A3(n13999), .ZN(n14004) );
  INV_X1 U16000 ( .A(n14002), .ZN(n14003) );
  OAI21_X1 U16001 ( .B1(n14004), .B2(n14003), .A(n14052), .ZN(n14010) );
  NAND2_X1 U16002 ( .A1(n14023), .A2(n14321), .ZN(n14006) );
  NAND2_X1 U16003 ( .A1(n14006), .A2(n14005), .ZN(n14008) );
  NOR2_X1 U16004 ( .A1(n14026), .A2(n14619), .ZN(n14007) );
  AOI211_X1 U16005 ( .C1(n14064), .C2(n14323), .A(n14008), .B(n14007), .ZN(
        n14009) );
  OAI211_X1 U16006 ( .C1(n14011), .C2(n14067), .A(n14010), .B(n14009), .ZN(
        P1_U3228) );
  AOI22_X1 U16007 ( .A1(n14023), .A2(n14319), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14013) );
  NAND2_X1 U16008 ( .A1(n14064), .A2(n14320), .ZN(n14012) );
  OAI211_X1 U16009 ( .C1(n14026), .C2(n14498), .A(n14013), .B(n14012), .ZN(
        n14019) );
  INV_X1 U16010 ( .A(n14014), .ZN(n14015) );
  NAND3_X1 U16011 ( .A1(n13932), .A2(n14016), .A3(n14015), .ZN(n14017) );
  AOI21_X1 U16012 ( .B1(n13980), .B2(n14017), .A(n14074), .ZN(n14018) );
  AOI211_X1 U16013 ( .C1(n14664), .C2(n9398), .A(n14019), .B(n14018), .ZN(
        n14020) );
  INV_X1 U16014 ( .A(n14020), .ZN(P1_U3229) );
  XNOR2_X1 U16015 ( .A(n14022), .B(n14021), .ZN(n14029) );
  AOI22_X1 U16016 ( .A1(n14553), .A2(n14023), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14025) );
  NAND2_X1 U16017 ( .A1(n14555), .A2(n14064), .ZN(n14024) );
  OAI211_X1 U16018 ( .C1(n14026), .C2(n14559), .A(n14025), .B(n14024), .ZN(
        n14027) );
  AOI21_X1 U16019 ( .B1(n14688), .B2(n9398), .A(n14027), .ZN(n14028) );
  OAI21_X1 U16020 ( .B1(n14029), .B2(n14074), .A(n14028), .ZN(P1_U3233) );
  INV_X1 U16021 ( .A(n14030), .ZN(n14032) );
  NOR3_X1 U16022 ( .A1(n14033), .A2(n14032), .A3(n14031), .ZN(n14035) );
  INV_X1 U16023 ( .A(n13933), .ZN(n14034) );
  OAI21_X1 U16024 ( .B1(n14035), .B2(n14034), .A(n14052), .ZN(n14041) );
  INV_X1 U16025 ( .A(n14036), .ZN(n14525) );
  AND2_X1 U16026 ( .A1(n14320), .A2(n15059), .ZN(n14037) );
  AOI21_X1 U16027 ( .B1(n14553), .B2(n14554), .A(n14037), .ZN(n14674) );
  INV_X1 U16028 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14038) );
  OAI22_X1 U16029 ( .A1(n14674), .A2(n14055), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14038), .ZN(n14039) );
  AOI21_X1 U16030 ( .B1(n14525), .B2(n14071), .A(n14039), .ZN(n14040) );
  OAI211_X1 U16031 ( .C1(n14067), .C2(n14676), .A(n14041), .B(n14040), .ZN(
        P1_U3235) );
  OAI21_X1 U16032 ( .B1(n14043), .B2(n14042), .A(n13948), .ZN(n14044) );
  NAND2_X1 U16033 ( .A1(n14044), .A2(n14052), .ZN(n14048) );
  INV_X1 U16034 ( .A(n14045), .ZN(n14595) );
  AOI22_X1 U16035 ( .A1(n14555), .A2(n15059), .B1(n14554), .B2(n14322), .ZN(
        n14594) );
  NAND2_X1 U16036 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15045)
         );
  OAI21_X1 U16037 ( .B1(n14594), .B2(n14055), .A(n15045), .ZN(n14046) );
  AOI21_X1 U16038 ( .B1(n14595), .B2(n14071), .A(n14046), .ZN(n14047) );
  OAI211_X1 U16039 ( .C1(n14198), .C2(n14067), .A(n14048), .B(n14047), .ZN(
        P1_U3238) );
  OAI21_X1 U16040 ( .B1(n14051), .B2(n14050), .A(n14049), .ZN(n14053) );
  NAND2_X1 U16041 ( .A1(n14053), .A2(n14052), .ZN(n14059) );
  INV_X1 U16042 ( .A(n14460), .ZN(n14057) );
  AOI22_X1 U16043 ( .A1(n14554), .A2(n14319), .B1(n14317), .B2(n15059), .ZN(
        n14649) );
  INV_X1 U16044 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14054) );
  OAI22_X1 U16045 ( .A1(n14055), .A2(n14649), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14054), .ZN(n14056) );
  AOI21_X1 U16046 ( .B1(n14071), .B2(n14057), .A(n14056), .ZN(n14058) );
  OAI211_X1 U16047 ( .C1(n14463), .C2(n14067), .A(n14059), .B(n14058), .ZN(
        P1_U3240) );
  INV_X1 U16048 ( .A(n14060), .ZN(n14061) );
  AOI21_X1 U16049 ( .B1(n14063), .B2(n14062), .A(n14061), .ZN(n14075) );
  NAND2_X1 U16050 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15031)
         );
  NAND2_X1 U16051 ( .A1(n14064), .A2(n14325), .ZN(n14065) );
  OAI211_X1 U16052 ( .C1(n14066), .C2(n14607), .A(n15031), .B(n14065), .ZN(
        n14070) );
  NOR2_X1 U16053 ( .A1(n14068), .A2(n14067), .ZN(n14069) );
  AOI211_X1 U16054 ( .C1(n14072), .C2(n14071), .A(n14070), .B(n14069), .ZN(
        n14073) );
  OAI21_X1 U16055 ( .B1(n14075), .B2(n14074), .A(n14073), .ZN(P1_U3241) );
  NAND2_X1 U16056 ( .A1(n14076), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n14079) );
  NAND2_X1 U16057 ( .A1(n14077), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n14078) );
  OAI211_X1 U16058 ( .C1(n14081), .C2(n14080), .A(n14079), .B(n14078), .ZN(
        n14418) );
  NAND2_X1 U16059 ( .A1(n8306), .A2(n14598), .ZN(n14082) );
  NOR2_X1 U16060 ( .A1(n14418), .A2(n14123), .ZN(n14090) );
  AND2_X1 U16061 ( .A1(n14418), .A2(n14206), .ZN(n14089) );
  MUX2_X1 U16062 ( .A(n14090), .B(n14089), .S(n14633), .Z(n14304) );
  NAND2_X1 U16063 ( .A1(n14092), .A2(n14091), .ZN(n14093) );
  NAND2_X1 U16064 ( .A1(n14094), .A2(n14093), .ZN(n14095) );
  INV_X1 U16065 ( .A(n14095), .ZN(n14096) );
  NOR2_X1 U16066 ( .A1(n14096), .A2(n14302), .ZN(n14303) );
  MUX2_X1 U16067 ( .A(n14098), .B(n14097), .S(n14252), .Z(n14241) );
  MUX2_X1 U16068 ( .A(n14327), .B(n14885), .S(n14155), .Z(n14164) );
  NAND2_X1 U16069 ( .A1(n14338), .A2(n14099), .ZN(n14100) );
  NAND2_X1 U16070 ( .A1(n14101), .A2(n14100), .ZN(n15138) );
  XNOR2_X1 U16071 ( .A(n14101), .B(n14123), .ZN(n14102) );
  OAI21_X1 U16072 ( .B1(n15138), .B2(n14103), .A(n14102), .ZN(n14105) );
  MUX2_X1 U16073 ( .A(n14106), .B(n14107), .S(n14155), .Z(n14104) );
  NAND2_X1 U16074 ( .A1(n14105), .A2(n14104), .ZN(n14109) );
  MUX2_X1 U16075 ( .A(n14107), .B(n14106), .S(n14155), .Z(n14108) );
  NAND3_X1 U16076 ( .A1(n14109), .A2(n14268), .A3(n14108), .ZN(n14115) );
  NAND2_X1 U16077 ( .A1(n14336), .A2(n14206), .ZN(n14113) );
  NAND2_X1 U16078 ( .A1(n14110), .A2(n14252), .ZN(n14112) );
  MUX2_X1 U16079 ( .A(n14113), .B(n14112), .S(n14111), .Z(n14114) );
  NAND3_X1 U16080 ( .A1(n14115), .A2(n14269), .A3(n14114), .ZN(n14121) );
  NAND2_X1 U16081 ( .A1(n14123), .A2(n14116), .ZN(n14119) );
  MUX2_X1 U16082 ( .A(n14119), .B(n14118), .S(n14335), .Z(n14120) );
  NAND2_X1 U16083 ( .A1(n14121), .A2(n14120), .ZN(n14127) );
  MUX2_X1 U16084 ( .A(n14122), .B(n15147), .S(n14155), .Z(n14126) );
  MUX2_X1 U16085 ( .A(n14334), .B(n14124), .S(n14206), .Z(n14125) );
  OAI21_X1 U16086 ( .B1(n14127), .B2(n14126), .A(n14125), .ZN(n14129) );
  NAND2_X1 U16087 ( .A1(n14127), .A2(n14126), .ZN(n14128) );
  MUX2_X1 U16088 ( .A(n15152), .B(n14333), .S(n14155), .Z(n14131) );
  MUX2_X1 U16089 ( .A(n14333), .B(n15152), .S(n14155), .Z(n14130) );
  MUX2_X1 U16090 ( .A(n14332), .B(n15160), .S(n14155), .Z(n14134) );
  MUX2_X1 U16091 ( .A(n14332), .B(n15160), .S(n14206), .Z(n14133) );
  MUX2_X1 U16092 ( .A(n14331), .B(n14135), .S(n14206), .Z(n14139) );
  NAND2_X1 U16093 ( .A1(n14138), .A2(n14139), .ZN(n14137) );
  MUX2_X1 U16094 ( .A(n14331), .B(n14135), .S(n14155), .Z(n14136) );
  NAND2_X1 U16095 ( .A1(n14137), .A2(n14136), .ZN(n14143) );
  INV_X1 U16096 ( .A(n14138), .ZN(n14141) );
  INV_X1 U16097 ( .A(n14139), .ZN(n14140) );
  NAND2_X1 U16098 ( .A1(n14141), .A2(n14140), .ZN(n14142) );
  NAND2_X1 U16099 ( .A1(n14143), .A2(n14142), .ZN(n14145) );
  MUX2_X1 U16100 ( .A(n14330), .B(n15089), .S(n14155), .Z(n14146) );
  MUX2_X1 U16101 ( .A(n14330), .B(n15089), .S(n14206), .Z(n14144) );
  INV_X1 U16102 ( .A(n14146), .ZN(n14147) );
  MUX2_X1 U16103 ( .A(n14329), .B(n15076), .S(n14206), .Z(n14150) );
  MUX2_X1 U16104 ( .A(n14329), .B(n15076), .S(n14155), .Z(n14148) );
  NAND2_X1 U16105 ( .A1(n14149), .A2(n14148), .ZN(n14152) );
  MUX2_X1 U16106 ( .A(n14328), .B(n15188), .S(n14155), .Z(n14154) );
  MUX2_X1 U16107 ( .A(n14328), .B(n15188), .S(n14206), .Z(n14153) );
  MUX2_X1 U16108 ( .A(n15058), .B(n14934), .S(n14206), .Z(n14158) );
  MUX2_X1 U16109 ( .A(n15058), .B(n14934), .S(n14155), .Z(n14156) );
  INV_X1 U16110 ( .A(n14158), .ZN(n14159) );
  MUX2_X1 U16111 ( .A(n14327), .B(n14885), .S(n14206), .Z(n14160) );
  NAND2_X1 U16112 ( .A1(n14161), .A2(n14160), .ZN(n14162) );
  OAI21_X1 U16113 ( .B1(n14164), .B2(n14163), .A(n14162), .ZN(n14168) );
  AND2_X1 U16114 ( .A1(n14173), .A2(n14165), .ZN(n14169) );
  AND2_X1 U16115 ( .A1(n14174), .A2(n14166), .ZN(n14170) );
  MUX2_X1 U16116 ( .A(n14326), .B(n14961), .S(n14206), .Z(n14175) );
  NOR2_X1 U16117 ( .A1(n14961), .A2(n14123), .ZN(n14176) );
  NOR2_X1 U16118 ( .A1(n14326), .A2(n14252), .ZN(n14172) );
  OR3_X1 U16119 ( .A1(n14175), .A2(n14176), .A3(n14172), .ZN(n14167) );
  NAND4_X1 U16120 ( .A1(n14168), .A2(n14169), .A3(n14170), .A4(n14167), .ZN(
        n14187) );
  INV_X1 U16121 ( .A(n14169), .ZN(n14183) );
  INV_X1 U16122 ( .A(n14170), .ZN(n14179) );
  OR2_X1 U16123 ( .A1(n14179), .A2(n14206), .ZN(n14171) );
  OAI21_X1 U16124 ( .B1(n14183), .B2(n14252), .A(n14171), .ZN(n14185) );
  NAND2_X1 U16125 ( .A1(n14175), .A2(n14172), .ZN(n14182) );
  MUX2_X1 U16126 ( .A(n14174), .B(n14173), .S(n14252), .Z(n14181) );
  INV_X1 U16127 ( .A(n14175), .ZN(n14178) );
  INV_X1 U16128 ( .A(n14176), .ZN(n14177) );
  OR3_X1 U16129 ( .A1(n14179), .A2(n14178), .A3(n14177), .ZN(n14180) );
  OAI211_X1 U16130 ( .C1(n14183), .C2(n14182), .A(n14181), .B(n14180), .ZN(
        n14184) );
  AOI21_X1 U16131 ( .B1(n14289), .B2(n14185), .A(n14184), .ZN(n14186) );
  NAND2_X1 U16132 ( .A1(n14187), .A2(n14186), .ZN(n14191) );
  MUX2_X1 U16133 ( .A(n14323), .B(n14714), .S(n14206), .Z(n14190) );
  NAND2_X1 U16134 ( .A1(n14191), .A2(n14190), .ZN(n14189) );
  MUX2_X1 U16135 ( .A(n14323), .B(n14714), .S(n14252), .Z(n14188) );
  NAND2_X1 U16136 ( .A1(n14189), .A2(n14188), .ZN(n14193) );
  OR2_X1 U16137 ( .A1(n14191), .A2(n14190), .ZN(n14192) );
  NAND2_X1 U16138 ( .A1(n14193), .A2(n14192), .ZN(n14197) );
  MUX2_X1 U16139 ( .A(n14322), .B(n14710), .S(n14252), .Z(n14194) );
  MUX2_X1 U16140 ( .A(n14609), .B(n14198), .S(n14252), .Z(n14199) );
  MUX2_X1 U16141 ( .A(n14203), .B(n14202), .S(n14206), .Z(n14204) );
  NAND2_X1 U16142 ( .A1(n14205), .A2(n14204), .ZN(n14210) );
  MUX2_X1 U16143 ( .A(n14577), .B(n14688), .S(n14206), .Z(n14207) );
  INV_X1 U16144 ( .A(n14207), .ZN(n14209) );
  MUX2_X1 U16145 ( .A(n14688), .B(n14577), .S(n14206), .Z(n14208) );
  OAI21_X1 U16146 ( .B1(n14210), .B2(n14209), .A(n14208), .ZN(n14212) );
  NAND2_X1 U16147 ( .A1(n14210), .A2(n14209), .ZN(n14211) );
  MUX2_X1 U16148 ( .A(n14553), .B(n14682), .S(n14252), .Z(n14214) );
  MUX2_X1 U16149 ( .A(n14682), .B(n14553), .S(n14252), .Z(n14213) );
  MUX2_X1 U16150 ( .A(n14676), .B(n14216), .S(n14252), .Z(n14215) );
  INV_X1 U16151 ( .A(n14215), .ZN(n14218) );
  MUX2_X1 U16152 ( .A(n14216), .B(n14676), .S(n14252), .Z(n14217) );
  AOI21_X1 U16153 ( .B1(n14219), .B2(n14218), .A(n14217), .ZN(n14220) );
  MUX2_X1 U16154 ( .A(n14668), .B(n14320), .S(n14206), .Z(n14222) );
  MUX2_X1 U16155 ( .A(n14668), .B(n14320), .S(n14252), .Z(n14221) );
  MUX2_X1 U16156 ( .A(n14664), .B(n14512), .S(n14252), .Z(n14224) );
  MUX2_X1 U16157 ( .A(n14512), .B(n14664), .S(n14252), .Z(n14223) );
  OR2_X1 U16158 ( .A1(n14225), .A2(n14224), .ZN(n14226) );
  NAND2_X1 U16159 ( .A1(n14227), .A2(n14226), .ZN(n14229) );
  MUX2_X1 U16160 ( .A(n14319), .B(n14659), .S(n14252), .Z(n14230) );
  MUX2_X1 U16161 ( .A(n14659), .B(n14319), .S(n14252), .Z(n14228) );
  INV_X1 U16162 ( .A(n14230), .ZN(n14231) );
  MUX2_X1 U16163 ( .A(n14652), .B(n14318), .S(n14252), .Z(n14234) );
  MUX2_X1 U16164 ( .A(n14652), .B(n14318), .S(n14123), .Z(n14232) );
  NAND2_X1 U16165 ( .A1(n14233), .A2(n14232), .ZN(n14236) );
  NAND2_X1 U16166 ( .A1(n14236), .A2(n14235), .ZN(n14237) );
  MUX2_X1 U16167 ( .A(n14317), .B(n14644), .S(n14252), .Z(n14238) );
  MUX2_X1 U16168 ( .A(n14644), .B(n14317), .S(n14252), .Z(n14239) );
  MUX2_X1 U16169 ( .A(n14316), .B(n14639), .S(n14252), .Z(n14240) );
  OR2_X1 U16170 ( .A1(n14744), .A2(n14242), .ZN(n14244) );
  OR2_X1 U16171 ( .A1(n7896), .A2(n14742), .ZN(n14243) );
  OAI21_X1 U16172 ( .B1(n14418), .B2(n14245), .A(n14314), .ZN(n14246) );
  INV_X1 U16173 ( .A(n14246), .ZN(n14247) );
  NAND2_X1 U16174 ( .A1(n14418), .A2(n14252), .ZN(n14250) );
  INV_X1 U16175 ( .A(n14314), .ZN(n14248) );
  AOI21_X1 U16176 ( .B1(n14250), .B2(n14249), .A(n14248), .ZN(n14251) );
  AOI21_X1 U16177 ( .B1(n14415), .B2(n14123), .A(n14251), .ZN(n14261) );
  MUX2_X1 U16178 ( .A(n14253), .B(n14315), .S(n14252), .Z(n14257) );
  INV_X1 U16179 ( .A(n14257), .ZN(n14254) );
  MUX2_X1 U16180 ( .A(n14315), .B(n14253), .S(n14252), .Z(n14256) );
  AOI22_X1 U16181 ( .A1(n14259), .A2(n14261), .B1(n14254), .B2(n14256), .ZN(
        n14255) );
  INV_X1 U16182 ( .A(n14256), .ZN(n14258) );
  NAND2_X1 U16183 ( .A1(n14258), .A2(n14257), .ZN(n14260) );
  INV_X1 U16184 ( .A(n14260), .ZN(n14264) );
  INV_X1 U16185 ( .A(n14261), .ZN(n14263) );
  AOI21_X1 U16186 ( .B1(n14261), .B2(n14260), .A(n14259), .ZN(n14262) );
  AOI21_X1 U16187 ( .B1(n14264), .B2(n14263), .A(n14262), .ZN(n14265) );
  XNOR2_X1 U16188 ( .A(n14633), .B(n14418), .ZN(n14300) );
  AOI21_X1 U16189 ( .B1(n14266), .B2(n14265), .A(n14300), .ZN(n14267) );
  XNOR2_X1 U16190 ( .A(n14415), .B(n14314), .ZN(n14297) );
  INV_X1 U16191 ( .A(n15138), .ZN(n14270) );
  NAND4_X1 U16192 ( .A1(n14271), .A2(n14270), .A3(n14269), .A4(n14268), .ZN(
        n14274) );
  NOR3_X1 U16193 ( .A1(n14274), .A2(n14273), .A3(n14272), .ZN(n14277) );
  NAND4_X1 U16194 ( .A1(n14278), .A2(n14277), .A3(n14276), .A4(n14275), .ZN(
        n14279) );
  OR4_X1 U16195 ( .A1(n14281), .A2(n15056), .A3(n14280), .A4(n14279), .ZN(
        n14282) );
  NOR2_X1 U16196 ( .A1(n14283), .A2(n14282), .ZN(n14286) );
  NAND4_X1 U16197 ( .A1(n14602), .A2(n14286), .A3(n14285), .A4(n14284), .ZN(
        n14287) );
  OR4_X1 U16198 ( .A1(n14591), .A2(n14289), .A3(n14288), .A4(n14287), .ZN(
        n14290) );
  NOR2_X1 U16199 ( .A1(n14291), .A2(n14290), .ZN(n14292) );
  NAND4_X1 U16200 ( .A1(n14520), .A2(n14292), .A3(n14565), .A4(n14545), .ZN(
        n14293) );
  NOR2_X1 U16201 ( .A1(n14493), .A2(n14293), .ZN(n14294) );
  AND4_X1 U16202 ( .A1(n14455), .A2(n14294), .A3(n14471), .A4(n14509), .ZN(
        n14296) );
  NAND4_X1 U16203 ( .A1(n14297), .A2(n14296), .A3(n14450), .A4(n14295), .ZN(
        n14298) );
  NOR3_X1 U16204 ( .A1(n14300), .A2(n14299), .A3(n14298), .ZN(n14301) );
  XOR2_X1 U16205 ( .A(n14598), .B(n14301), .Z(n14307) );
  INV_X1 U16206 ( .A(n14302), .ZN(n14306) );
  AOI21_X1 U16207 ( .B1(n14304), .B2(n14303), .A(n14311), .ZN(n14305) );
  OAI21_X1 U16208 ( .B1(n14307), .B2(n14306), .A(n14305), .ZN(n14313) );
  NAND3_X1 U16209 ( .A1(n14309), .A2(n6559), .A3(n14554), .ZN(n14310) );
  OAI211_X1 U16210 ( .C1(n14756), .C2(n14311), .A(n14310), .B(P1_B_REG_SCAN_IN), .ZN(n14312) );
  MUX2_X1 U16211 ( .A(n14418), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14337), .Z(
        P1_U3591) );
  MUX2_X1 U16212 ( .A(n14314), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14337), .Z(
        P1_U3590) );
  MUX2_X1 U16213 ( .A(n14315), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14337), .Z(
        P1_U3589) );
  MUX2_X1 U16214 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14316), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16215 ( .A(n14317), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14337), .Z(
        P1_U3587) );
  MUX2_X1 U16216 ( .A(n14318), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14337), .Z(
        P1_U3586) );
  MUX2_X1 U16217 ( .A(n14319), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14337), .Z(
        P1_U3585) );
  MUX2_X1 U16218 ( .A(n14512), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14337), .Z(
        P1_U3584) );
  MUX2_X1 U16219 ( .A(n14320), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14337), .Z(
        P1_U3583) );
  MUX2_X1 U16220 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n6940), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16221 ( .A(n14553), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14337), .Z(
        P1_U3581) );
  MUX2_X1 U16222 ( .A(n14577), .B(P1_DATAO_REG_20__SCAN_IN), .S(n14337), .Z(
        P1_U3580) );
  MUX2_X1 U16223 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14555), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16224 ( .A(n14321), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14337), .Z(
        P1_U3578) );
  MUX2_X1 U16225 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14322), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16226 ( .A(n14323), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14337), .Z(
        P1_U3576) );
  MUX2_X1 U16227 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14324), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16228 ( .A(n14325), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14337), .Z(
        P1_U3574) );
  MUX2_X1 U16229 ( .A(n14326), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14337), .Z(
        P1_U3573) );
  MUX2_X1 U16230 ( .A(n14327), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14337), .Z(
        P1_U3572) );
  MUX2_X1 U16231 ( .A(n15058), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14337), .Z(
        P1_U3571) );
  MUX2_X1 U16232 ( .A(n14328), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14337), .Z(
        P1_U3570) );
  MUX2_X1 U16233 ( .A(n14329), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14337), .Z(
        P1_U3569) );
  MUX2_X1 U16234 ( .A(n14330), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14337), .Z(
        P1_U3568) );
  MUX2_X1 U16235 ( .A(n14331), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14337), .Z(
        P1_U3567) );
  MUX2_X1 U16236 ( .A(n14332), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14337), .Z(
        P1_U3566) );
  MUX2_X1 U16237 ( .A(n14333), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14337), .Z(
        P1_U3565) );
  MUX2_X1 U16238 ( .A(n14334), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14337), .Z(
        P1_U3564) );
  MUX2_X1 U16239 ( .A(n14335), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14337), .Z(
        P1_U3563) );
  MUX2_X1 U16240 ( .A(n14336), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14337), .Z(
        P1_U3562) );
  MUX2_X1 U16241 ( .A(n14624), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14337), .Z(
        P1_U3561) );
  MUX2_X1 U16242 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14338), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16243 ( .C1(n14341), .C2(n14340), .A(n15040), .B(n14339), .ZN(
        n14350) );
  MUX2_X1 U16244 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9013), .S(n14342), .Z(
        n14343) );
  OAI21_X1 U16245 ( .B1(n15000), .B2(n7503), .A(n14343), .ZN(n14344) );
  NAND3_X1 U16246 ( .A1(n15035), .A2(n14345), .A3(n14344), .ZN(n14349) );
  NAND2_X1 U16247 ( .A1(n15038), .A2(n14346), .ZN(n14348) );
  AOI22_X1 U16248 ( .A1(n15006), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14347) );
  NAND4_X1 U16249 ( .A1(n14350), .A2(n14349), .A3(n14348), .A4(n14347), .ZN(
        P1_U3244) );
  INV_X1 U16250 ( .A(n14351), .ZN(n14354) );
  OAI22_X1 U16251 ( .A1(n15047), .A2(n14761), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14352), .ZN(n14353) );
  AOI21_X1 U16252 ( .B1(n14354), .B2(n15038), .A(n14353), .ZN(n14362) );
  OAI211_X1 U16253 ( .C1(n14356), .C2(n14355), .A(n15035), .B(n14371), .ZN(
        n14361) );
  INV_X1 U16254 ( .A(n14376), .ZN(n14357) );
  OAI211_X1 U16255 ( .C1(n14359), .C2(n14358), .A(n15040), .B(n14357), .ZN(
        n14360) );
  NAND4_X1 U16256 ( .A1(n14363), .A2(n14362), .A3(n14361), .A4(n14360), .ZN(
        P1_U3245) );
  NOR2_X1 U16257 ( .A1(n15047), .A2(n14364), .ZN(n14365) );
  AOI211_X1 U16258 ( .C1(n15038), .C2(n14367), .A(n14366), .B(n14365), .ZN(
        n14381) );
  MUX2_X1 U16259 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9020), .S(n14368), .Z(
        n14369) );
  NAND3_X1 U16260 ( .A1(n14371), .A2(n14370), .A3(n14369), .ZN(n14372) );
  NAND3_X1 U16261 ( .A1(n15035), .A2(n14373), .A3(n14372), .ZN(n14380) );
  OR3_X1 U16262 ( .A1(n14376), .A2(n14375), .A3(n14374), .ZN(n14377) );
  NAND3_X1 U16263 ( .A1(n15040), .A2(n14378), .A3(n14377), .ZN(n14379) );
  NAND3_X1 U16264 ( .A1(n14381), .A2(n14380), .A3(n14379), .ZN(P1_U3246) );
  INV_X1 U16265 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14773) );
  NOR2_X1 U16266 ( .A1(n15047), .A2(n14773), .ZN(n14382) );
  AOI211_X1 U16267 ( .C1(n15038), .C2(n14391), .A(n14383), .B(n14382), .ZN(
        n14399) );
  INV_X1 U16268 ( .A(n14384), .ZN(n14386) );
  MUX2_X1 U16269 ( .A(n9157), .B(P1_REG2_REG_7__SCAN_IN), .S(n14391), .Z(
        n14385) );
  NAND2_X1 U16270 ( .A1(n14386), .A2(n14385), .ZN(n14388) );
  OAI211_X1 U16271 ( .C1(n14389), .C2(n14388), .A(n14387), .B(n15040), .ZN(
        n14398) );
  INV_X1 U16272 ( .A(n14390), .ZN(n14393) );
  MUX2_X1 U16273 ( .A(n15202), .B(P1_REG1_REG_7__SCAN_IN), .S(n14391), .Z(
        n14392) );
  NAND2_X1 U16274 ( .A1(n14393), .A2(n14392), .ZN(n14395) );
  OAI211_X1 U16275 ( .C1(n14396), .C2(n14395), .A(n14394), .B(n15035), .ZN(
        n14397) );
  NAND3_X1 U16276 ( .A1(n14399), .A2(n14398), .A3(n14397), .ZN(P1_U3250) );
  OAI21_X1 U16277 ( .B1(n14402), .B2(n14401), .A(n14400), .ZN(n14403) );
  NAND2_X1 U16278 ( .A1(n14403), .A2(n15035), .ZN(n14414) );
  INV_X1 U16279 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14831) );
  OAI21_X1 U16280 ( .B1(n15047), .B2(n14831), .A(n14404), .ZN(n14405) );
  AOI21_X1 U16281 ( .B1(n14406), .B2(n15038), .A(n14405), .ZN(n14413) );
  OR3_X1 U16282 ( .A1(n14409), .A2(n14408), .A3(n14407), .ZN(n14410) );
  NAND3_X1 U16283 ( .A1(n14411), .A2(n15040), .A3(n14410), .ZN(n14412) );
  NAND3_X1 U16284 ( .A1(n14414), .A2(n14413), .A3(n14412), .ZN(P1_U3254) );
  NAND2_X1 U16285 ( .A1(n14636), .A2(n14422), .ZN(n14421) );
  XNOR2_X1 U16286 ( .A(n14633), .B(n14421), .ZN(n14416) );
  NAND2_X1 U16287 ( .A1(n14416), .A2(n8988), .ZN(n14632) );
  NAND2_X1 U16288 ( .A1(n14418), .A2(n14417), .ZN(n14634) );
  NOR2_X1 U16289 ( .A1(n15106), .A2(n14634), .ZN(n14424) );
  NOR2_X1 U16290 ( .A1(n14633), .A2(n14541), .ZN(n14419) );
  AOI211_X1 U16291 ( .C1(n15106), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14424), 
        .B(n14419), .ZN(n14420) );
  OAI21_X1 U16292 ( .B1(n14632), .B2(n14583), .A(n14420), .ZN(P1_U3263) );
  OAI211_X1 U16293 ( .C1(n14636), .C2(n14422), .A(n14421), .B(n8988), .ZN(
        n14635) );
  NOR2_X1 U16294 ( .A1(n14636), .A2(n14541), .ZN(n14423) );
  AOI211_X1 U16295 ( .C1(n15106), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14424), 
        .B(n14423), .ZN(n14425) );
  OAI21_X1 U16296 ( .B1(n14583), .B2(n14635), .A(n14425), .ZN(P1_U3264) );
  INV_X1 U16297 ( .A(n14426), .ZN(n14428) );
  OAI21_X1 U16298 ( .B1(n14598), .B2(n14428), .A(n14427), .ZN(n14429) );
  NAND2_X1 U16299 ( .A1(n14429), .A2(n15104), .ZN(n14436) );
  OAI22_X1 U16300 ( .A1(n14431), .A2(n6716), .B1(n14430), .B2(n15091), .ZN(
        n14434) );
  NOR2_X1 U16301 ( .A1(n14432), .A2(n14541), .ZN(n14433) );
  AOI211_X1 U16302 ( .C1(n15106), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14434), 
        .B(n14433), .ZN(n14435) );
  OAI211_X1 U16303 ( .C1(n14437), .C2(n14623), .A(n14436), .B(n14435), .ZN(
        P1_U3356) );
  XNOR2_X1 U16304 ( .A(n14438), .B(n14450), .ZN(n14441) );
  INV_X1 U16305 ( .A(n14439), .ZN(n14440) );
  AOI21_X1 U16306 ( .B1(n14441), .B2(n15139), .A(n14440), .ZN(n14646) );
  INV_X1 U16307 ( .A(n14459), .ZN(n14444) );
  INV_X1 U16308 ( .A(n14442), .ZN(n14443) );
  AOI211_X1 U16309 ( .C1(n14644), .C2(n14444), .A(n14589), .B(n14443), .ZN(
        n14643) );
  AOI22_X1 U16310 ( .A1(n15106), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n15073), 
        .B2(n14445), .ZN(n14446) );
  OAI21_X1 U16311 ( .B1(n14447), .B2(n14541), .A(n14446), .ZN(n14451) );
  OAI21_X1 U16312 ( .B1(n14454), .B2(n14453), .A(n14452), .ZN(n14655) );
  XNOR2_X1 U16313 ( .A(n14456), .B(n14455), .ZN(n14648) );
  NAND2_X1 U16314 ( .A1(n14648), .A2(n14627), .ZN(n14466) );
  NAND2_X1 U16315 ( .A1(n14652), .A2(n14473), .ZN(n14457) );
  NAND2_X1 U16316 ( .A1(n14457), .A2(n8988), .ZN(n14458) );
  NOR2_X1 U16317 ( .A1(n14459), .A2(n14458), .ZN(n14650) );
  OAI22_X1 U16318 ( .A1(n15106), .A2(n14649), .B1(n14460), .B2(n15091), .ZN(
        n14461) );
  AOI21_X1 U16319 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n15106), .A(n14461), 
        .ZN(n14462) );
  OAI21_X1 U16320 ( .B1(n14463), .B2(n14541), .A(n14462), .ZN(n14464) );
  AOI21_X1 U16321 ( .B1(n14650), .B2(n15101), .A(n14464), .ZN(n14465) );
  OAI211_X1 U16322 ( .C1(n14655), .C2(n14623), .A(n14466), .B(n14465), .ZN(
        P1_U3267) );
  OAI21_X1 U16323 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(n14662) );
  OAI21_X1 U16324 ( .B1(n14472), .B2(n14471), .A(n14470), .ZN(n14656) );
  NAND2_X1 U16325 ( .A1(n14656), .A2(n14627), .ZN(n14485) );
  INV_X1 U16326 ( .A(n14496), .ZN(n14475) );
  INV_X1 U16327 ( .A(n14473), .ZN(n14474) );
  AOI211_X1 U16328 ( .C1(n14659), .C2(n14475), .A(n14589), .B(n14474), .ZN(
        n14657) );
  NAND2_X1 U16329 ( .A1(n14657), .A2(n14617), .ZN(n14478) );
  OAI22_X1 U16330 ( .A1(n14476), .A2(n14606), .B1(n8247), .B2(n14608), .ZN(
        n14658) );
  INV_X1 U16331 ( .A(n14658), .ZN(n14477) );
  OAI211_X1 U16332 ( .C1(n15091), .C2(n14479), .A(n14478), .B(n14477), .ZN(
        n14483) );
  OAI22_X1 U16333 ( .A1(n14481), .A2(n14541), .B1(n14480), .B2(n15104), .ZN(
        n14482) );
  AOI21_X1 U16334 ( .B1(n14483), .B2(n15104), .A(n14482), .ZN(n14484) );
  OAI211_X1 U16335 ( .C1(n14662), .C2(n14623), .A(n14485), .B(n14484), .ZN(
        P1_U3268) );
  AOI21_X1 U16336 ( .B1(n14488), .B2(n14487), .A(n14486), .ZN(n14667) );
  INV_X1 U16337 ( .A(n14667), .ZN(n14502) );
  OAI22_X1 U16338 ( .A1(n14490), .A2(n14606), .B1(n14489), .B2(n14608), .ZN(
        n14495) );
  AOI211_X1 U16339 ( .C1(n14493), .C2(n14492), .A(n15084), .B(n14491), .ZN(
        n14494) );
  AOI211_X1 U16340 ( .C1(n15167), .C2(n14502), .A(n14495), .B(n14494), .ZN(
        n14666) );
  AOI211_X1 U16341 ( .C1(n14664), .C2(n6572), .A(n14589), .B(n14496), .ZN(
        n14663) );
  NOR2_X1 U16342 ( .A1(n14497), .A2(n14541), .ZN(n14501) );
  OAI22_X1 U16343 ( .A1(n15104), .A2(n14499), .B1(n14498), .B2(n15091), .ZN(
        n14500) );
  AOI211_X1 U16344 ( .C1(n14663), .C2(n15101), .A(n14501), .B(n14500), .ZN(
        n14504) );
  NAND2_X1 U16345 ( .A1(n14502), .A2(n15081), .ZN(n14503) );
  OAI211_X1 U16346 ( .C1(n14666), .C2(n15106), .A(n14504), .B(n14503), .ZN(
        P1_U3269) );
  NAND2_X1 U16347 ( .A1(n14505), .A2(n14509), .ZN(n14506) );
  NAND2_X1 U16348 ( .A1(n14507), .A2(n14506), .ZN(n14671) );
  OAI21_X1 U16349 ( .B1(n14510), .B2(n14509), .A(n14508), .ZN(n14511) );
  NAND2_X1 U16350 ( .A1(n14511), .A2(n15139), .ZN(n14514) );
  AOI22_X1 U16351 ( .A1(n6940), .A2(n14554), .B1(n15059), .B2(n14512), .ZN(
        n14513) );
  NAND2_X1 U16352 ( .A1(n14514), .A2(n14513), .ZN(n14673) );
  AOI21_X1 U16353 ( .B1(n14668), .B2(n14524), .A(n14589), .ZN(n14515) );
  NAND2_X1 U16354 ( .A1(n14515), .A2(n6572), .ZN(n14669) );
  OAI22_X1 U16355 ( .A1(n14669), .A2(n14598), .B1(n15091), .B2(n14516), .ZN(
        n14517) );
  OAI21_X1 U16356 ( .B1(n14673), .B2(n14517), .A(n15104), .ZN(n14519) );
  AOI22_X1 U16357 ( .A1(n14668), .A2(n15075), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15106), .ZN(n14518) );
  OAI211_X1 U16358 ( .C1(n14671), .C2(n14623), .A(n14519), .B(n14518), .ZN(
        P1_U3270) );
  XNOR2_X1 U16359 ( .A(n14521), .B(n14520), .ZN(n14680) );
  XNOR2_X1 U16360 ( .A(n14523), .B(n14522), .ZN(n14678) );
  OAI211_X1 U16361 ( .C1(n14676), .C2(n14537), .A(n8988), .B(n14524), .ZN(
        n14675) );
  AOI22_X1 U16362 ( .A1(n15106), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14525), 
        .B2(n15073), .ZN(n14526) );
  OAI21_X1 U16363 ( .B1(n14674), .B2(n15106), .A(n14526), .ZN(n14527) );
  AOI21_X1 U16364 ( .B1(n14528), .B2(n15075), .A(n14527), .ZN(n14529) );
  OAI21_X1 U16365 ( .B1(n14675), .B2(n14583), .A(n14529), .ZN(n14530) );
  AOI21_X1 U16366 ( .B1(n14678), .B2(n15102), .A(n14530), .ZN(n14531) );
  OAI21_X1 U16367 ( .B1(n14680), .B2(n14532), .A(n14531), .ZN(P1_U3271) );
  XOR2_X1 U16368 ( .A(n14533), .B(n14545), .Z(n14536) );
  INV_X1 U16369 ( .A(n14534), .ZN(n14535) );
  AOI21_X1 U16370 ( .B1(n14536), .B2(n15139), .A(n14535), .ZN(n14684) );
  AOI211_X1 U16371 ( .C1(n14682), .C2(n14562), .A(n14589), .B(n14537), .ZN(
        n14681) );
  INV_X1 U16372 ( .A(n14538), .ZN(n14539) );
  AOI22_X1 U16373 ( .A1(n14539), .A2(n15073), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15106), .ZN(n14540) );
  OAI21_X1 U16374 ( .B1(n6812), .B2(n14541), .A(n14540), .ZN(n14547) );
  INV_X1 U16375 ( .A(n14542), .ZN(n14543) );
  AOI21_X1 U16376 ( .B1(n14545), .B2(n14544), .A(n14543), .ZN(n14685) );
  NOR2_X1 U16377 ( .A1(n14685), .A2(n14623), .ZN(n14546) );
  AOI211_X1 U16378 ( .C1(n14681), .C2(n15101), .A(n14547), .B(n14546), .ZN(
        n14548) );
  OAI21_X1 U16379 ( .B1(n15106), .B2(n14684), .A(n14548), .ZN(P1_U3272) );
  NAND2_X1 U16380 ( .A1(n14550), .A2(n14549), .ZN(n14551) );
  NAND3_X1 U16381 ( .A1(n14552), .A2(n15139), .A3(n14551), .ZN(n14557) );
  AOI22_X1 U16382 ( .A1(n14555), .A2(n14554), .B1(n14553), .B2(n15059), .ZN(
        n14556) );
  NAND2_X1 U16383 ( .A1(n14557), .A2(n14556), .ZN(n14693) );
  INV_X1 U16384 ( .A(n14693), .ZN(n14569) );
  INV_X1 U16385 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14558) );
  OAI22_X1 U16386 ( .A1(n14559), .A2(n15091), .B1(n14558), .B2(n15104), .ZN(
        n14564) );
  INV_X1 U16387 ( .A(n14575), .ZN(n14560) );
  AOI21_X1 U16388 ( .B1(n14688), .B2(n14560), .A(n14589), .ZN(n14561) );
  NAND2_X1 U16389 ( .A1(n14562), .A2(n14561), .ZN(n14689) );
  NOR2_X1 U16390 ( .A1(n14689), .A2(n14583), .ZN(n14563) );
  AOI211_X1 U16391 ( .C1(n15075), .C2(n14688), .A(n14564), .B(n14563), .ZN(
        n14568) );
  NAND2_X1 U16392 ( .A1(n14566), .A2(n14565), .ZN(n14686) );
  NAND3_X1 U16393 ( .A1(n14687), .A2(n14686), .A3(n15102), .ZN(n14567) );
  OAI211_X1 U16394 ( .C1(n14569), .C2(n15106), .A(n14568), .B(n14567), .ZN(
        P1_U3273) );
  XNOR2_X1 U16395 ( .A(n14570), .B(n14572), .ZN(n14702) );
  OAI21_X1 U16396 ( .B1(n14573), .B2(n14572), .A(n14571), .ZN(n14700) );
  AND2_X1 U16397 ( .A1(n14581), .A2(n14587), .ZN(n14574) );
  OR3_X1 U16398 ( .A1(n14575), .A2(n14574), .A3(n14589), .ZN(n14697) );
  NOR2_X1 U16399 ( .A1(n14609), .A2(n14606), .ZN(n14576) );
  AOI21_X1 U16400 ( .B1(n14577), .B2(n15059), .A(n14576), .ZN(n14696) );
  OAI21_X1 U16401 ( .B1(n14578), .B2(n15091), .A(n14696), .ZN(n14579) );
  MUX2_X1 U16402 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14579), .S(n15104), .Z(
        n14580) );
  AOI21_X1 U16403 ( .B1(n14581), .B2(n15075), .A(n14580), .ZN(n14582) );
  OAI21_X1 U16404 ( .B1(n14697), .B2(n14583), .A(n14582), .ZN(n14584) );
  AOI21_X1 U16405 ( .B1(n14700), .B2(n14627), .A(n14584), .ZN(n14585) );
  OAI21_X1 U16406 ( .B1(n14702), .B2(n14623), .A(n14585), .ZN(P1_U3274) );
  XNOR2_X1 U16407 ( .A(n14586), .B(n14591), .ZN(n14708) );
  INV_X1 U16408 ( .A(n14616), .ZN(n14590) );
  INV_X1 U16409 ( .A(n14587), .ZN(n14588) );
  AOI211_X1 U16410 ( .C1(n14705), .C2(n14590), .A(n14589), .B(n14588), .ZN(
        n14703) );
  INV_X1 U16411 ( .A(n14703), .ZN(n14597) );
  XNOR2_X1 U16412 ( .A(n14592), .B(n14591), .ZN(n14593) );
  NAND2_X1 U16413 ( .A1(n14593), .A2(n15139), .ZN(n14707) );
  INV_X1 U16414 ( .A(n14594), .ZN(n14704) );
  AOI21_X1 U16415 ( .B1(n14595), .B2(n15073), .A(n14704), .ZN(n14596) );
  OAI211_X1 U16416 ( .C1(n14598), .C2(n14597), .A(n14707), .B(n14596), .ZN(
        n14599) );
  NAND2_X1 U16417 ( .A1(n14599), .A2(n15104), .ZN(n14601) );
  AOI22_X1 U16418 ( .A1(n14705), .A2(n15075), .B1(n15106), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n14600) );
  OAI211_X1 U16419 ( .C1(n14623), .C2(n14708), .A(n14601), .B(n14600), .ZN(
        P1_U3275) );
  XNOR2_X1 U16420 ( .A(n14603), .B(n14602), .ZN(n14713) );
  AOI21_X1 U16421 ( .B1(n14605), .B2(n14604), .A(n15084), .ZN(n14612) );
  OAI22_X1 U16422 ( .A1(n14609), .A2(n14608), .B1(n14607), .B2(n14606), .ZN(
        n14610) );
  AOI21_X1 U16423 ( .B1(n14612), .B2(n14611), .A(n14610), .ZN(n14712) );
  NAND2_X1 U16424 ( .A1(n14613), .A2(n14710), .ZN(n14614) );
  NAND2_X1 U16425 ( .A1(n14614), .A2(n8988), .ZN(n14615) );
  NOR2_X1 U16426 ( .A1(n14616), .A2(n14615), .ZN(n14709) );
  NAND2_X1 U16427 ( .A1(n14709), .A2(n14617), .ZN(n14618) );
  OAI211_X1 U16428 ( .C1(n15091), .C2(n14619), .A(n14712), .B(n14618), .ZN(
        n14620) );
  NAND2_X1 U16429 ( .A1(n14620), .A2(n15104), .ZN(n14622) );
  AOI22_X1 U16430 ( .A1(n14710), .A2(n15075), .B1(n15106), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n14621) );
  OAI211_X1 U16431 ( .C1(n14713), .C2(n14623), .A(n14622), .B(n14621), .ZN(
        P1_U3276) );
  NAND2_X1 U16432 ( .A1(n14624), .A2(n15059), .ZN(n15143) );
  OAI22_X1 U16433 ( .A1(n15106), .A2(n15143), .B1(n14625), .B2(n15091), .ZN(
        n14626) );
  AOI21_X1 U16434 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n15106), .A(n14626), .ZN(
        n14631) );
  OAI21_X1 U16435 ( .B1(n15102), .B2(n14627), .A(n15138), .ZN(n14630) );
  OAI21_X1 U16436 ( .B1(n14628), .B2(n15075), .A(n15141), .ZN(n14629) );
  NAND3_X1 U16437 ( .A1(n14631), .A2(n14630), .A3(n14629), .ZN(P1_U3293) );
  OAI211_X1 U16438 ( .C1(n15191), .C2(n14633), .A(n14632), .B(n14634), .ZN(
        n14719) );
  MUX2_X1 U16439 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14719), .S(n15209), .Z(
        P1_U3559) );
  OAI211_X1 U16440 ( .C1(n15191), .C2(n14636), .A(n14635), .B(n14634), .ZN(
        n14720) );
  MUX2_X1 U16441 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14720), .S(n15209), .Z(
        P1_U3558) );
  MUX2_X1 U16442 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14637), .S(n15209), .Z(
        P1_U3557) );
  AOI21_X1 U16443 ( .B1(n14639), .B2(n15159), .A(n14638), .ZN(n14640) );
  MUX2_X1 U16444 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14721), .S(n15209), .Z(
        P1_U3556) );
  AOI21_X1 U16445 ( .B1(n14644), .B2(n15159), .A(n14643), .ZN(n14645) );
  OAI211_X1 U16446 ( .C1(n14647), .C2(n14964), .A(n14646), .B(n14645), .ZN(
        n14722) );
  MUX2_X1 U16447 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14722), .S(n15209), .Z(
        P1_U3555) );
  NAND2_X1 U16448 ( .A1(n14648), .A2(n15139), .ZN(n14654) );
  INV_X1 U16449 ( .A(n14649), .ZN(n14651) );
  AOI211_X1 U16450 ( .C1(n14652), .C2(n15159), .A(n14651), .B(n14650), .ZN(
        n14653) );
  OAI211_X1 U16451 ( .C1(n14964), .C2(n14655), .A(n14654), .B(n14653), .ZN(
        n14723) );
  MUX2_X1 U16452 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14723), .S(n15209), .Z(
        P1_U3554) );
  NAND2_X1 U16453 ( .A1(n14656), .A2(n15139), .ZN(n14661) );
  AOI211_X1 U16454 ( .C1(n14659), .C2(n15159), .A(n14658), .B(n14657), .ZN(
        n14660) );
  OAI211_X1 U16455 ( .C1(n14964), .C2(n14662), .A(n14661), .B(n14660), .ZN(
        n14724) );
  MUX2_X1 U16456 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14724), .S(n15209), .Z(
        P1_U3553) );
  AOI21_X1 U16457 ( .B1(n14664), .B2(n15159), .A(n14663), .ZN(n14665) );
  OAI211_X1 U16458 ( .C1(n14667), .C2(n15163), .A(n14666), .B(n14665), .ZN(
        n14725) );
  MUX2_X1 U16459 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14725), .S(n15209), .Z(
        P1_U3552) );
  NAND2_X1 U16460 ( .A1(n14668), .A2(n15159), .ZN(n14670) );
  OAI211_X1 U16461 ( .C1(n14671), .C2(n14964), .A(n14670), .B(n14669), .ZN(
        n14672) );
  MUX2_X1 U16462 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14726), .S(n15209), .Z(
        P1_U3551) );
  OAI211_X1 U16463 ( .C1(n15191), .C2(n14676), .A(n14675), .B(n14674), .ZN(
        n14677) );
  AOI21_X1 U16464 ( .B1(n14678), .B2(n15195), .A(n14677), .ZN(n14679) );
  OAI21_X1 U16465 ( .B1(n14680), .B2(n15084), .A(n14679), .ZN(n14727) );
  MUX2_X1 U16466 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14727), .S(n15209), .Z(
        P1_U3550) );
  AOI21_X1 U16467 ( .B1(n14682), .B2(n15159), .A(n14681), .ZN(n14683) );
  OAI211_X1 U16468 ( .C1(n14964), .C2(n14685), .A(n14684), .B(n14683), .ZN(
        n14728) );
  MUX2_X1 U16469 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14728), .S(n15209), .Z(
        P1_U3549) );
  NAND3_X1 U16470 ( .A1(n14687), .A2(n14686), .A3(n15195), .ZN(n14691) );
  NAND2_X1 U16471 ( .A1(n14688), .A2(n15159), .ZN(n14690) );
  NAND3_X1 U16472 ( .A1(n14691), .A2(n14690), .A3(n14689), .ZN(n14692) );
  NOR2_X1 U16473 ( .A1(n14693), .A2(n14692), .ZN(n14729) );
  MUX2_X1 U16474 ( .A(n14694), .B(n14729), .S(n15209), .Z(n14695) );
  INV_X1 U16475 ( .A(n14695), .ZN(P1_U3548) );
  OAI211_X1 U16476 ( .C1(n14698), .C2(n15191), .A(n14697), .B(n14696), .ZN(
        n14699) );
  AOI21_X1 U16477 ( .B1(n14700), .B2(n15139), .A(n14699), .ZN(n14701) );
  OAI21_X1 U16478 ( .B1(n14964), .B2(n14702), .A(n14701), .ZN(n14732) );
  MUX2_X1 U16479 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14732), .S(n15209), .Z(
        P1_U3547) );
  AOI211_X1 U16480 ( .C1(n14705), .C2(n15159), .A(n14704), .B(n14703), .ZN(
        n14706) );
  OAI211_X1 U16481 ( .C1(n14964), .C2(n14708), .A(n14707), .B(n14706), .ZN(
        n14733) );
  MUX2_X1 U16482 ( .A(n14733), .B(P1_REG1_REG_18__SCAN_IN), .S(n15206), .Z(
        P1_U3546) );
  AOI21_X1 U16483 ( .B1(n14710), .B2(n15159), .A(n14709), .ZN(n14711) );
  OAI211_X1 U16484 ( .C1(n14964), .C2(n14713), .A(n14712), .B(n14711), .ZN(
        n14734) );
  MUX2_X1 U16485 ( .A(n14734), .B(P1_REG1_REG_17__SCAN_IN), .S(n15206), .Z(
        P1_U3545) );
  AOI22_X1 U16486 ( .A1(n14715), .A2(n8988), .B1(n14714), .B2(n15159), .ZN(
        n14716) );
  OAI211_X1 U16487 ( .C1(n14964), .C2(n14718), .A(n14717), .B(n14716), .ZN(
        n14735) );
  MUX2_X1 U16488 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14735), .S(n15209), .Z(
        P1_U3544) );
  MUX2_X1 U16489 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14719), .S(n15197), .Z(
        P1_U3527) );
  MUX2_X1 U16490 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14720), .S(n15197), .Z(
        P1_U3526) );
  MUX2_X1 U16491 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14721), .S(n15197), .Z(
        P1_U3524) );
  MUX2_X1 U16492 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14722), .S(n15197), .Z(
        P1_U3523) );
  MUX2_X1 U16493 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14723), .S(n15197), .Z(
        P1_U3522) );
  MUX2_X1 U16494 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14724), .S(n15197), .Z(
        P1_U3521) );
  MUX2_X1 U16495 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14725), .S(n15197), .Z(
        P1_U3520) );
  MUX2_X1 U16496 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14726), .S(n15197), .Z(
        P1_U3519) );
  MUX2_X1 U16497 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14727), .S(n15197), .Z(
        P1_U3518) );
  MUX2_X1 U16498 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14728), .S(n15197), .Z(
        P1_U3517) );
  INV_X1 U16499 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14730) );
  MUX2_X1 U16500 ( .A(n14730), .B(n14729), .S(n15197), .Z(n14731) );
  INV_X1 U16501 ( .A(n14731), .ZN(P1_U3516) );
  MUX2_X1 U16502 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14732), .S(n15197), .Z(
        P1_U3515) );
  MUX2_X1 U16503 ( .A(n14733), .B(P1_REG0_REG_18__SCAN_IN), .S(n15196), .Z(
        P1_U3513) );
  MUX2_X1 U16504 ( .A(n14734), .B(P1_REG0_REG_17__SCAN_IN), .S(n15196), .Z(
        P1_U3510) );
  MUX2_X1 U16505 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14735), .S(n15197), .Z(
        P1_U3507) );
  NOR4_X1 U16506 ( .A1(n14737), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14736), .A4(
        P1_U3086), .ZN(n14738) );
  AOI21_X1 U16507 ( .B1(n14739), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14738), 
        .ZN(n14740) );
  OAI21_X1 U16508 ( .B1(n14741), .B2(n14753), .A(n14740), .ZN(P1_U3324) );
  OAI222_X1 U16509 ( .A1(n14753), .A2(n14744), .B1(P1_U3086), .B2(n14743), 
        .C1(n14742), .C2(n14755), .ZN(P1_U3325) );
  OAI222_X1 U16510 ( .A1(n14753), .A2(n14747), .B1(P1_U3086), .B2(n14746), 
        .C1(n14745), .C2(n14755), .ZN(P1_U3326) );
  OAI222_X1 U16511 ( .A1(n14755), .A2(n14750), .B1(n14753), .B2(n14749), .C1(
        n14748), .C2(P1_U3086), .ZN(P1_U3329) );
  OAI222_X1 U16512 ( .A1(n14755), .A2(n14754), .B1(n14753), .B2(n14752), .C1(
        P1_U3086), .C2(n14751), .ZN(P1_U3330) );
  MUX2_X1 U16513 ( .A(n14757), .B(n14756), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16514 ( .A(n14758), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16515 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14782) );
  NOR2_X1 U16516 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n14776), .ZN(n14779) );
  NAND2_X1 U16517 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n14791), .ZN(n14790) );
  OAI21_X1 U16518 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(n14760), .A(n14759), .ZN(
        n14789) );
  XOR2_X1 U16519 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14787) );
  INV_X1 U16520 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14762) );
  NOR2_X1 U16521 ( .A1(n14763), .A2(n14762), .ZN(n14765) );
  INV_X1 U16522 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14768) );
  NOR2_X1 U16523 ( .A1(n14767), .A2(n14768), .ZN(n14770) );
  AND2_X1 U16524 ( .A1(n14806), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14771) );
  NOR2_X1 U16525 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14772), .ZN(n14775) );
  XNOR2_X1 U16526 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14772), .ZN(n14810) );
  INV_X1 U16527 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14777) );
  AOI22_X1 U16528 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P3_ADDR_REG_8__SCAN_IN), 
        .B1(n14777), .B2(n14776), .ZN(n14783) );
  XOR2_X1 U16529 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n14780), .Z(n14817) );
  NAND2_X1 U16530 ( .A1(n14818), .A2(n14817), .ZN(n14781) );
  XOR2_X1 U16531 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n14823) );
  XOR2_X1 U16532 ( .A(n14824), .B(n14823), .Z(n14822) );
  XOR2_X1 U16533 ( .A(n14784), .B(n14783), .Z(n14814) );
  NAND2_X1 U16534 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14786), .ZN(n14802) );
  XNOR2_X1 U16535 ( .A(n14788), .B(n14787), .ZN(n14870) );
  XNOR2_X1 U16536 ( .A(n14790), .B(n14789), .ZN(n14793) );
  NAND2_X1 U16537 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14793), .ZN(n14795) );
  OAI21_X1 U16538 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n14791), .A(n14790), .ZN(
        n14792) );
  INV_X1 U16539 ( .A(n14792), .ZN(n15544) );
  NOR2_X1 U16540 ( .A1(n9371), .A2(n15544), .ZN(n15551) );
  NAND2_X1 U16541 ( .A1(n15551), .A2(n15550), .ZN(n14794) );
  NAND2_X1 U16542 ( .A1(n14870), .A2(n14871), .ZN(n14796) );
  NOR2_X1 U16543 ( .A1(n14870), .A2(n14871), .ZN(n14869) );
  XNOR2_X1 U16544 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14797), .ZN(n14799) );
  NOR2_X1 U16545 ( .A1(n14798), .A2(n14799), .ZN(n15548) );
  NOR2_X1 U16546 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15547), .ZN(n14800) );
  NAND2_X1 U16547 ( .A1(n15542), .A2(n15541), .ZN(n14801) );
  NAND2_X1 U16548 ( .A1(n14804), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14809) );
  NOR2_X1 U16549 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n14806), .ZN(n14805) );
  AOI21_X1 U16550 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n14806), .A(n14805), .ZN(
        n14808) );
  XOR2_X1 U16551 ( .A(n14808), .B(n14807), .Z(n14874) );
  NAND2_X1 U16552 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14811), .ZN(n14812) );
  XNOR2_X1 U16553 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14810), .ZN(n15546) );
  NOR2_X1 U16554 ( .A1(n14814), .A2(n14813), .ZN(n14816) );
  XNOR2_X1 U16555 ( .A(n14818), .B(n14817), .ZN(n14820) );
  XNOR2_X1 U16556 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n14827) );
  INV_X1 U16557 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14826) );
  XNOR2_X1 U16558 ( .A(n14827), .B(n14830), .ZN(n14979) );
  XNOR2_X1 U16559 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n14832) );
  INV_X1 U16560 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14828) );
  NAND2_X1 U16561 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n14828), .ZN(n14829) );
  XOR2_X1 U16562 ( .A(n14832), .B(n14835), .Z(n14984) );
  NAND2_X1 U16563 ( .A1(n14983), .A2(n14984), .ZN(n14833) );
  AND2_X1 U16564 ( .A1(n14834), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n14836) );
  XOR2_X1 U16565 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .Z(n14837) );
  XOR2_X1 U16566 ( .A(n14842), .B(n14837), .Z(n14838) );
  NOR2_X1 U16567 ( .A1(n14839), .A2(n14838), .ZN(n14987) );
  INV_X1 U16568 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14843) );
  INV_X1 U16569 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14840) );
  NAND2_X1 U16570 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14840), .ZN(n14841) );
  XOR2_X1 U16571 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n14844) );
  XOR2_X1 U16572 ( .A(n14850), .B(n14844), .Z(n14845) );
  XNOR2_X1 U16573 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14851) );
  INV_X1 U16574 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14847) );
  NAND2_X1 U16575 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n14847), .ZN(n14849) );
  XOR2_X1 U16576 ( .A(n14851), .B(n14856), .Z(n14853) );
  NAND2_X1 U16577 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14854), .ZN(n14855) );
  INV_X1 U16578 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15033) );
  AOI22_X1 U16579 ( .A1(n14856), .A2(n14855), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n15033), .ZN(n14857) );
  XOR2_X1 U16580 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n14857), .Z(n14858) );
  XNOR2_X1 U16581 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n14858), .ZN(n14997) );
  NOR2_X1 U16582 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14857), .ZN(n14860) );
  XNOR2_X1 U16583 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14863), .ZN(n14864) );
  XOR2_X1 U16584 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14864), .Z(n14861) );
  NOR2_X1 U16585 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14863), .ZN(n14866) );
  INV_X1 U16586 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14911) );
  NOR2_X1 U16587 ( .A1(n14911), .A2(n14864), .ZN(n14865) );
  NOR2_X1 U16588 ( .A1(n14866), .A2(n14865), .ZN(n14895) );
  XOR2_X1 U16589 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14894) );
  XNOR2_X1 U16590 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14893), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16591 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14867) );
  OAI21_X1 U16592 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14867), 
        .ZN(U28) );
  AOI21_X1 U16593 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14868) );
  OAI21_X1 U16594 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14868), 
        .ZN(U29) );
  AOI21_X1 U16595 ( .B1(n14871), .B2(n14870), .A(n14869), .ZN(n14873) );
  XNOR2_X1 U16596 ( .A(n14873), .B(n14872), .ZN(SUB_1596_U61) );
  XOR2_X1 U16597 ( .A(n14875), .B(n14874), .Z(SUB_1596_U57) );
  XNOR2_X1 U16598 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14876), .ZN(SUB_1596_U55)
         );
  NOR2_X1 U16599 ( .A1(n14878), .A2(n14877), .ZN(n14879) );
  XOR2_X1 U16600 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14879), .Z(SUB_1596_U54) );
  NOR2_X1 U16601 ( .A1(n14881), .A2(n14880), .ZN(n14882) );
  XOR2_X1 U16602 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14882), .Z(SUB_1596_U70)
         );
  INV_X1 U16603 ( .A(n14887), .ZN(n14889) );
  AOI211_X1 U16604 ( .C1(n14885), .C2(n15159), .A(n14884), .B(n14883), .ZN(
        n14886) );
  OAI21_X1 U16605 ( .B1(n15163), .B2(n14887), .A(n14886), .ZN(n14888) );
  AOI21_X1 U16606 ( .B1(n15167), .B2(n14889), .A(n14888), .ZN(n14891) );
  INV_X1 U16607 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14890) );
  AOI22_X1 U16608 ( .A1(n15197), .A2(n14891), .B1(n14890), .B2(n15196), .ZN(
        P1_U3495) );
  AOI22_X1 U16609 ( .A1(n15209), .A2(n14891), .B1(n9409), .B2(n15206), .ZN(
        P1_U3540) );
  XNOR2_X1 U16610 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14892), .ZN(SUB_1596_U63)
         );
  INV_X1 U16611 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15048) );
  NOR2_X1 U16612 ( .A1(n14895), .A2(n14894), .ZN(n14896) );
  AOI21_X1 U16613 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n15048), .A(n14896), 
        .ZN(n14900) );
  XNOR2_X1 U16614 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14898) );
  XNOR2_X1 U16615 ( .A(n14898), .B(n14897), .ZN(n14899) );
  AOI21_X1 U16616 ( .B1(n14903), .B2(n14902), .A(n14901), .ZN(n14920) );
  OAI21_X1 U16617 ( .B1(n14905), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14904), 
        .ZN(n14918) );
  NAND2_X1 U16618 ( .A1(n14907), .A2(n14906), .ZN(n14909) );
  OAI211_X1 U16619 ( .C1(n14911), .C2(n14910), .A(n14909), .B(n14908), .ZN(
        n14917) );
  INV_X1 U16620 ( .A(n14912), .ZN(n14913) );
  AOI211_X1 U16621 ( .C1(n14915), .C2(n14914), .A(n15454), .B(n14913), .ZN(
        n14916) );
  AOI211_X1 U16622 ( .C1(n15461), .C2(n14918), .A(n14917), .B(n14916), .ZN(
        n14919) );
  OAI21_X1 U16623 ( .B1(n14920), .B2(n15465), .A(n14919), .ZN(P3_U3199) );
  OAI21_X1 U16624 ( .B1(n15515), .B2(n6739), .A(n14921), .ZN(n14922) );
  AOI21_X1 U16625 ( .B1(n15518), .B2(n14923), .A(n14922), .ZN(n14925) );
  INV_X1 U16626 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14924) );
  AOI22_X1 U16627 ( .A1(n15540), .A2(n14925), .B1(n14924), .B2(n15538), .ZN(
        P3_U3470) );
  INV_X1 U16628 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14926) );
  AOI22_X1 U16629 ( .A1(n15521), .A2(n14926), .B1(n14925), .B2(n15519), .ZN(
        P3_U3423) );
  INV_X1 U16630 ( .A(n14927), .ZN(n14928) );
  AOI21_X1 U16631 ( .B1(n14928), .B2(n14935), .A(n15084), .ZN(n14931) );
  AOI21_X1 U16632 ( .B1(n14931), .B2(n14930), .A(n14929), .ZN(n14968) );
  INV_X1 U16633 ( .A(n14932), .ZN(n14933) );
  AOI222_X1 U16634 ( .A1(n14934), .A2(n15075), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n15106), .C1(n15073), .C2(n14933), .ZN(n14941) );
  XNOR2_X1 U16635 ( .A(n14936), .B(n14935), .ZN(n14971) );
  OAI211_X1 U16636 ( .C1(n14969), .C2(n14938), .A(n8988), .B(n14937), .ZN(
        n14967) );
  INV_X1 U16637 ( .A(n14967), .ZN(n14939) );
  AOI22_X1 U16638 ( .A1(n14971), .A2(n15102), .B1(n15101), .B2(n14939), .ZN(
        n14940) );
  OAI211_X1 U16639 ( .C1(n15106), .C2(n14968), .A(n14941), .B(n14940), .ZN(
        P1_U3282) );
  AOI211_X1 U16640 ( .C1(n14944), .C2(n15159), .A(n14943), .B(n14942), .ZN(
        n14945) );
  OAI21_X1 U16641 ( .B1(n14946), .B2(n14964), .A(n14945), .ZN(n14947) );
  AOI21_X1 U16642 ( .B1(n14948), .B2(n15139), .A(n14947), .ZN(n14973) );
  AOI22_X1 U16643 ( .A1(n15209), .A2(n14973), .B1(n8111), .B2(n15206), .ZN(
        P1_U3543) );
  NAND3_X1 U16644 ( .A1(n14950), .A2(n14949), .A3(n15195), .ZN(n14955) );
  AOI21_X1 U16645 ( .B1(n14952), .B2(n15159), .A(n14951), .ZN(n14954) );
  NAND3_X1 U16646 ( .A1(n14955), .A2(n14954), .A3(n14953), .ZN(n14956) );
  AOI21_X1 U16647 ( .B1(n14957), .B2(n15139), .A(n14956), .ZN(n14974) );
  AOI22_X1 U16648 ( .A1(n15209), .A2(n14974), .B1(n8082), .B2(n15206), .ZN(
        P1_U3542) );
  INV_X1 U16649 ( .A(n14958), .ZN(n14960) );
  AOI211_X1 U16650 ( .C1(n14961), .C2(n15159), .A(n14960), .B(n14959), .ZN(
        n14963) );
  OAI211_X1 U16651 ( .C1(n14965), .C2(n14964), .A(n14963), .B(n14962), .ZN(
        n14966) );
  INV_X1 U16652 ( .A(n14966), .ZN(n14975) );
  AOI22_X1 U16653 ( .A1(n15209), .A2(n14975), .B1(n9557), .B2(n15206), .ZN(
        P1_U3541) );
  OAI211_X1 U16654 ( .C1(n14969), .C2(n15191), .A(n14968), .B(n14967), .ZN(
        n14970) );
  AOI21_X1 U16655 ( .B1(n14971), .B2(n15195), .A(n14970), .ZN(n14977) );
  AOI22_X1 U16656 ( .A1(n15209), .A2(n14977), .B1(n8033), .B2(n15206), .ZN(
        P1_U3539) );
  INV_X1 U16657 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U16658 ( .A1(n15197), .A2(n14973), .B1(n14972), .B2(n15196), .ZN(
        P1_U3504) );
  AOI22_X1 U16659 ( .A1(n15197), .A2(n14974), .B1(n8083), .B2(n15196), .ZN(
        P1_U3501) );
  AOI22_X1 U16660 ( .A1(n15197), .A2(n14975), .B1(n8067), .B2(n15196), .ZN(
        P1_U3498) );
  INV_X1 U16661 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14976) );
  AOI22_X1 U16662 ( .A1(n15197), .A2(n14977), .B1(n14976), .B2(n15196), .ZN(
        P1_U3492) );
  AOI21_X1 U16663 ( .B1(n14980), .B2(n14979), .A(n14978), .ZN(n14981) );
  XNOR2_X1 U16664 ( .A(n14981), .B(n9492), .ZN(SUB_1596_U69) );
  AOI21_X1 U16665 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n14985) );
  XNOR2_X1 U16666 ( .A(n14985), .B(n9519), .ZN(SUB_1596_U68) );
  NOR2_X1 U16667 ( .A1(n14987), .A2(n14986), .ZN(n14988) );
  XOR2_X1 U16668 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14988), .Z(SUB_1596_U67)
         );
  NOR2_X1 U16669 ( .A1(n14990), .A2(n14989), .ZN(n14991) );
  XOR2_X1 U16670 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n14991), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16671 ( .A1(n14993), .A2(n14992), .ZN(n14994) );
  XOR2_X1 U16672 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14994), .Z(SUB_1596_U65)
         );
  OAI21_X1 U16673 ( .B1(n14997), .B2(n14996), .A(n14995), .ZN(n14998) );
  XNOR2_X1 U16674 ( .A(n14998), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  AOI21_X1 U16675 ( .B1(n6560), .B2(n15000), .A(n14999), .ZN(n15002) );
  XNOR2_X1 U16676 ( .A(n15002), .B(P1_IR_REG_0__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U16677 ( .A1(n15006), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15003) );
  OAI21_X1 U16678 ( .B1(n15005), .B2(n15004), .A(n15003), .ZN(P1_U3243) );
  NAND2_X1 U16679 ( .A1(n15006), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n15007) );
  OAI211_X1 U16680 ( .C1(n15029), .C2(n15009), .A(n15008), .B(n15007), .ZN(
        n15010) );
  INV_X1 U16681 ( .A(n15010), .ZN(n15019) );
  OAI211_X1 U16682 ( .C1(n15013), .C2(n15012), .A(n15011), .B(n15035), .ZN(
        n15018) );
  OAI211_X1 U16683 ( .C1(n15016), .C2(n15015), .A(n15014), .B(n15040), .ZN(
        n15017) );
  NAND3_X1 U16684 ( .A1(n15019), .A2(n15018), .A3(n15017), .ZN(P1_U3256) );
  AOI21_X1 U16685 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n15021), .A(n15020), 
        .ZN(n15026) );
  AOI21_X1 U16686 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n15023), .A(n15022), 
        .ZN(n15024) );
  OAI222_X1 U16687 ( .A1(n15029), .A2(n15028), .B1(n15027), .B2(n15026), .C1(
        n15025), .C2(n15024), .ZN(n15030) );
  INV_X1 U16688 ( .A(n15030), .ZN(n15032) );
  OAI211_X1 U16689 ( .C1(n15033), .C2(n15047), .A(n15032), .B(n15031), .ZN(
        P1_U3258) );
  OAI211_X1 U16690 ( .C1(n15036), .C2(P1_REG1_REG_18__SCAN_IN), .A(n15035), 
        .B(n15034), .ZN(n15044) );
  NAND2_X1 U16691 ( .A1(n15038), .A2(n15037), .ZN(n15043) );
  OAI211_X1 U16692 ( .C1(n15041), .C2(P1_REG2_REG_18__SCAN_IN), .A(n15040), 
        .B(n15039), .ZN(n15042) );
  AND3_X1 U16693 ( .A1(n15044), .A2(n15043), .A3(n15042), .ZN(n15046) );
  OAI211_X1 U16694 ( .C1(n15048), .C2(n15047), .A(n15046), .B(n15045), .ZN(
        P1_U3261) );
  AOI21_X1 U16695 ( .B1(n15049), .B2(n15056), .A(n15084), .ZN(n15053) );
  INV_X1 U16696 ( .A(n15050), .ZN(n15051) );
  AOI21_X1 U16697 ( .B1(n15053), .B2(n15052), .A(n15051), .ZN(n15190) );
  INV_X1 U16698 ( .A(n15054), .ZN(n15055) );
  AOI222_X1 U16699 ( .A1(n15188), .A2(n15075), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n15106), .C1(n15055), .C2(n15073), .ZN(n15063) );
  XNOR2_X1 U16700 ( .A(n15057), .B(n15056), .ZN(n15194) );
  XOR2_X1 U16701 ( .A(n15078), .B(n15188), .Z(n15060) );
  AOI22_X1 U16702 ( .A1(n15060), .A2(n8988), .B1(n15059), .B2(n15058), .ZN(
        n15189) );
  INV_X1 U16703 ( .A(n15189), .ZN(n15061) );
  AOI22_X1 U16704 ( .A1(n15194), .A2(n15102), .B1(n15101), .B2(n15061), .ZN(
        n15062) );
  OAI211_X1 U16705 ( .C1(n15106), .C2(n15190), .A(n15063), .B(n15062), .ZN(
        P1_U3283) );
  OAI21_X1 U16706 ( .B1(n15065), .B2(n15066), .A(n15064), .ZN(n15071) );
  XNOR2_X1 U16707 ( .A(n15067), .B(n15066), .ZN(n15077) );
  NOR2_X1 U16708 ( .A1(n15077), .A2(n15068), .ZN(n15069) );
  AOI211_X1 U16709 ( .C1(n15139), .C2(n15071), .A(n15070), .B(n15069), .ZN(
        n15182) );
  INV_X1 U16710 ( .A(n15072), .ZN(n15074) );
  AOI222_X1 U16711 ( .A1(n15076), .A2(n15075), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n15106), .C1(n15074), .C2(n15073), .ZN(n15083) );
  INV_X1 U16712 ( .A(n15077), .ZN(n15185) );
  INV_X1 U16713 ( .A(n15098), .ZN(n15079) );
  OAI211_X1 U16714 ( .C1(n15079), .C2(n15181), .A(n8988), .B(n15078), .ZN(
        n15180) );
  INV_X1 U16715 ( .A(n15180), .ZN(n15080) );
  AOI22_X1 U16716 ( .A1(n15185), .A2(n15081), .B1(n15101), .B2(n15080), .ZN(
        n15082) );
  OAI211_X1 U16717 ( .C1(n15106), .C2(n15182), .A(n15083), .B(n15082), .ZN(
        P1_U3284) );
  AOI21_X1 U16718 ( .B1(n15085), .B2(n15095), .A(n15084), .ZN(n15088) );
  AOI21_X1 U16719 ( .B1(n15088), .B2(n15087), .A(n15086), .ZN(n15175) );
  INV_X1 U16720 ( .A(n15175), .ZN(n15094) );
  INV_X1 U16721 ( .A(n15089), .ZN(n15176) );
  OAI22_X1 U16722 ( .A1(n15176), .A2(n15092), .B1(n15091), .B2(n15090), .ZN(
        n15093) );
  NOR2_X1 U16723 ( .A1(n15094), .A2(n15093), .ZN(n15105) );
  XNOR2_X1 U16724 ( .A(n15096), .B(n15095), .ZN(n15178) );
  INV_X1 U16725 ( .A(n15097), .ZN(n15099) );
  OAI211_X1 U16726 ( .C1(n15099), .C2(n15176), .A(n8988), .B(n15098), .ZN(
        n15174) );
  INV_X1 U16727 ( .A(n15174), .ZN(n15100) );
  AOI22_X1 U16728 ( .A1(n15178), .A2(n15102), .B1(n15101), .B2(n15100), .ZN(
        n15103) );
  OAI221_X1 U16729 ( .B1(n15106), .B2(n15105), .C1(n15104), .C2(n7979), .A(
        n15103), .ZN(P1_U3285) );
  INV_X1 U16730 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15107) );
  NOR2_X1 U16731 ( .A1(n15137), .A2(n15107), .ZN(P1_U3294) );
  INV_X1 U16732 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15108) );
  NOR2_X1 U16733 ( .A1(n15137), .A2(n15108), .ZN(P1_U3295) );
  INV_X1 U16734 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15109) );
  NOR2_X1 U16735 ( .A1(n15137), .A2(n15109), .ZN(P1_U3296) );
  INV_X1 U16736 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15110) );
  NOR2_X1 U16737 ( .A1(n15137), .A2(n15110), .ZN(P1_U3297) );
  NOR2_X1 U16738 ( .A1(n15137), .A2(n15111), .ZN(P1_U3298) );
  NOR2_X1 U16739 ( .A1(n15137), .A2(n15112), .ZN(P1_U3299) );
  INV_X1 U16740 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15113) );
  NOR2_X1 U16741 ( .A1(n15137), .A2(n15113), .ZN(P1_U3300) );
  INV_X1 U16742 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15114) );
  NOR2_X1 U16743 ( .A1(n15137), .A2(n15114), .ZN(P1_U3301) );
  INV_X1 U16744 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15115) );
  NOR2_X1 U16745 ( .A1(n15137), .A2(n15115), .ZN(P1_U3302) );
  INV_X1 U16746 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15116) );
  NOR2_X1 U16747 ( .A1(n15137), .A2(n15116), .ZN(P1_U3303) );
  INV_X1 U16748 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15117) );
  NOR2_X1 U16749 ( .A1(n15137), .A2(n15117), .ZN(P1_U3304) );
  INV_X1 U16750 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15118) );
  NOR2_X1 U16751 ( .A1(n15137), .A2(n15118), .ZN(P1_U3305) );
  NOR2_X1 U16752 ( .A1(n15137), .A2(n15119), .ZN(P1_U3306) );
  INV_X1 U16753 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15120) );
  NOR2_X1 U16754 ( .A1(n15137), .A2(n15120), .ZN(P1_U3307) );
  INV_X1 U16755 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15121) );
  NOR2_X1 U16756 ( .A1(n15137), .A2(n15121), .ZN(P1_U3308) );
  INV_X1 U16757 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15122) );
  NOR2_X1 U16758 ( .A1(n15137), .A2(n15122), .ZN(P1_U3309) );
  NOR2_X1 U16759 ( .A1(n15137), .A2(n15123), .ZN(P1_U3310) );
  INV_X1 U16760 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15124) );
  NOR2_X1 U16761 ( .A1(n15137), .A2(n15124), .ZN(P1_U3311) );
  NOR2_X1 U16762 ( .A1(n15137), .A2(n15125), .ZN(P1_U3312) );
  NOR2_X1 U16763 ( .A1(n15137), .A2(n15126), .ZN(P1_U3313) );
  INV_X1 U16764 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U16765 ( .A1(n15137), .A2(n15127), .ZN(P1_U3314) );
  NOR2_X1 U16766 ( .A1(n15137), .A2(n15128), .ZN(P1_U3315) );
  NOR2_X1 U16767 ( .A1(n15137), .A2(n15129), .ZN(P1_U3316) );
  NOR2_X1 U16768 ( .A1(n15137), .A2(n15130), .ZN(P1_U3317) );
  INV_X1 U16769 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15131) );
  NOR2_X1 U16770 ( .A1(n15137), .A2(n15131), .ZN(P1_U3318) );
  NOR2_X1 U16771 ( .A1(n15137), .A2(n15132), .ZN(P1_U3319) );
  NOR2_X1 U16772 ( .A1(n15137), .A2(n15133), .ZN(P1_U3320) );
  INV_X1 U16773 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15134) );
  NOR2_X1 U16774 ( .A1(n15137), .A2(n15134), .ZN(P1_U3321) );
  INV_X1 U16775 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15135) );
  NOR2_X1 U16776 ( .A1(n15137), .A2(n15135), .ZN(P1_U3322) );
  INV_X1 U16777 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15136) );
  NOR2_X1 U16778 ( .A1(n15137), .A2(n15136), .ZN(P1_U3323) );
  OAI21_X1 U16779 ( .B1(n15195), .B2(n15139), .A(n15138), .ZN(n15144) );
  NAND3_X1 U16780 ( .A1(n15141), .A2(n15140), .A3(n8306), .ZN(n15142) );
  AND3_X1 U16781 ( .A1(n15144), .A2(n15143), .A3(n15142), .ZN(n15198) );
  AOI22_X1 U16782 ( .A1(n15197), .A2(n15198), .B1(n7879), .B2(n15196), .ZN(
        P1_U3459) );
  OAI211_X1 U16783 ( .C1(n15147), .C2(n15191), .A(n15146), .B(n15145), .ZN(
        n15148) );
  AOI21_X1 U16784 ( .B1(n15149), .B2(n15195), .A(n15148), .ZN(n15199) );
  INV_X1 U16785 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15150) );
  AOI22_X1 U16786 ( .A1(n15197), .A2(n15199), .B1(n15150), .B2(n15196), .ZN(
        P1_U3471) );
  AOI21_X1 U16787 ( .B1(n15152), .B2(n15159), .A(n15151), .ZN(n15153) );
  OAI211_X1 U16788 ( .C1(n15155), .C2(n15163), .A(n15154), .B(n15153), .ZN(
        n15156) );
  INV_X1 U16789 ( .A(n15156), .ZN(n15200) );
  INV_X1 U16790 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15157) );
  AOI22_X1 U16791 ( .A1(n15197), .A2(n15200), .B1(n15157), .B2(n15196), .ZN(
        P1_U3474) );
  INV_X1 U16792 ( .A(n15164), .ZN(n15166) );
  AOI21_X1 U16793 ( .B1(n15160), .B2(n15159), .A(n15158), .ZN(n15161) );
  OAI211_X1 U16794 ( .C1(n15164), .C2(n15163), .A(n15162), .B(n15161), .ZN(
        n15165) );
  AOI21_X1 U16795 ( .B1(n15167), .B2(n15166), .A(n15165), .ZN(n15201) );
  INV_X1 U16796 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15168) );
  AOI22_X1 U16797 ( .A1(n15197), .A2(n15201), .B1(n15168), .B2(n15196), .ZN(
        P1_U3477) );
  OAI211_X1 U16798 ( .C1(n15171), .C2(n15191), .A(n15170), .B(n15169), .ZN(
        n15172) );
  AOI21_X1 U16799 ( .B1(n15173), .B2(n15195), .A(n15172), .ZN(n15203) );
  AOI22_X1 U16800 ( .A1(n15197), .A2(n15203), .B1(n7962), .B2(n15196), .ZN(
        P1_U3480) );
  OAI211_X1 U16801 ( .C1(n15176), .C2(n15191), .A(n15175), .B(n15174), .ZN(
        n15177) );
  AOI21_X1 U16802 ( .B1(n15178), .B2(n15195), .A(n15177), .ZN(n15204) );
  INV_X1 U16803 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15179) );
  AOI22_X1 U16804 ( .A1(n15197), .A2(n15204), .B1(n15179), .B2(n15196), .ZN(
        P1_U3483) );
  OAI21_X1 U16805 ( .B1(n15181), .B2(n15191), .A(n15180), .ZN(n15184) );
  INV_X1 U16806 ( .A(n15182), .ZN(n15183) );
  AOI211_X1 U16807 ( .C1(n15186), .C2(n15185), .A(n15184), .B(n15183), .ZN(
        n15205) );
  INV_X1 U16808 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15187) );
  AOI22_X1 U16809 ( .A1(n15197), .A2(n15205), .B1(n15187), .B2(n15196), .ZN(
        P1_U3486) );
  INV_X1 U16810 ( .A(n15188), .ZN(n15192) );
  OAI211_X1 U16811 ( .C1(n15192), .C2(n15191), .A(n15190), .B(n15189), .ZN(
        n15193) );
  AOI21_X1 U16812 ( .B1(n15195), .B2(n15194), .A(n15193), .ZN(n15208) );
  AOI22_X1 U16813 ( .A1(n15197), .A2(n15208), .B1(n8008), .B2(n15196), .ZN(
        P1_U3489) );
  AOI22_X1 U16814 ( .A1(n15209), .A2(n15198), .B1(n15000), .B2(n15206), .ZN(
        P1_U3528) );
  AOI22_X1 U16815 ( .A1(n15209), .A2(n15199), .B1(n7917), .B2(n15206), .ZN(
        P1_U3532) );
  AOI22_X1 U16816 ( .A1(n15209), .A2(n15200), .B1(n7933), .B2(n15206), .ZN(
        P1_U3533) );
  AOI22_X1 U16817 ( .A1(n15209), .A2(n15201), .B1(n9149), .B2(n15206), .ZN(
        P1_U3534) );
  AOI22_X1 U16818 ( .A1(n15209), .A2(n15203), .B1(n15202), .B2(n15206), .ZN(
        P1_U3535) );
  AOI22_X1 U16819 ( .A1(n15209), .A2(n15204), .B1(n9148), .B2(n15206), .ZN(
        P1_U3536) );
  AOI22_X1 U16820 ( .A1(n15209), .A2(n15205), .B1(n7993), .B2(n15206), .ZN(
        P1_U3537) );
  AOI22_X1 U16821 ( .A1(n15209), .A2(n15208), .B1(n15207), .B2(n15206), .ZN(
        P1_U3538) );
  NOR2_X1 U16822 ( .A1(n15294), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI21_X1 U16823 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15210), .ZN(n15221) );
  NOR2_X1 U16824 ( .A1(n15211), .A2(n9364), .ZN(n15214) );
  OAI211_X1 U16825 ( .C1(n15214), .C2(n15213), .A(n15296), .B(n15212), .ZN(
        n15220) );
  NAND2_X1 U16826 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15294), .ZN(n15219) );
  OAI211_X1 U16827 ( .C1(n15217), .C2(n15216), .A(n15302), .B(n15215), .ZN(
        n15218) );
  NAND4_X1 U16828 ( .A1(n15221), .A2(n15220), .A3(n15219), .A4(n15218), .ZN(
        P2_U3215) );
  INV_X1 U16829 ( .A(n15222), .ZN(n15223) );
  OAI21_X1 U16830 ( .B1(n15273), .B2(n15224), .A(n15223), .ZN(n15225) );
  AOI21_X1 U16831 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15294), .A(n15225), .ZN(
        n15235) );
  OAI211_X1 U16832 ( .C1(n15228), .C2(n15227), .A(n15302), .B(n15226), .ZN(
        n15234) );
  AOI211_X1 U16833 ( .C1(n15231), .C2(n15230), .A(n15229), .B(n15242), .ZN(
        n15232) );
  INV_X1 U16834 ( .A(n15232), .ZN(n15233) );
  NAND3_X1 U16835 ( .A1(n15235), .A2(n15234), .A3(n15233), .ZN(P2_U3217) );
  OAI21_X1 U16836 ( .B1(n15237), .B2(n15236), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15238) );
  OAI21_X1 U16837 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15238), .ZN(n15250) );
  OAI211_X1 U16838 ( .C1(n15241), .C2(n15240), .A(n15302), .B(n15239), .ZN(
        n15249) );
  NAND2_X1 U16839 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15294), .ZN(n15248) );
  AOI211_X1 U16840 ( .C1(n15245), .C2(n15244), .A(n15243), .B(n15242), .ZN(
        n15246) );
  INV_X1 U16841 ( .A(n15246), .ZN(n15247) );
  NAND4_X1 U16842 ( .A1(n15250), .A2(n15249), .A3(n15248), .A4(n15247), .ZN(
        P2_U3218) );
  AOI22_X1 U16843 ( .A1(n15294), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n15261) );
  OAI211_X1 U16844 ( .C1(n15253), .C2(n15252), .A(n15251), .B(n15296), .ZN(
        n15260) );
  OAI211_X1 U16845 ( .C1(n15256), .C2(n15255), .A(n15254), .B(n15302), .ZN(
        n15259) );
  NAND2_X1 U16846 ( .A1(n15299), .A2(n15257), .ZN(n15258) );
  NAND4_X1 U16847 ( .A1(n15261), .A2(n15260), .A3(n15259), .A4(n15258), .ZN(
        P2_U3227) );
  OAI211_X1 U16848 ( .C1(n15263), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15296), 
        .B(n15262), .ZN(n15264) );
  NAND2_X1 U16849 ( .A1(n15265), .A2(n15264), .ZN(n15266) );
  AOI21_X1 U16850 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(n15294), .A(n15266), 
        .ZN(n15271) );
  OAI211_X1 U16851 ( .C1(n15269), .C2(n15268), .A(n15302), .B(n15267), .ZN(
        n15270) );
  OAI211_X1 U16852 ( .C1(n15273), .C2(n15272), .A(n15271), .B(n15270), .ZN(
        P2_U3228) );
  AOI22_X1 U16853 ( .A1(n15294), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15282) );
  NAND2_X1 U16854 ( .A1(n15299), .A2(n15274), .ZN(n15281) );
  XOR2_X1 U16855 ( .A(P2_REG2_REG_15__SCAN_IN), .B(n15275), .Z(n15276) );
  NAND2_X1 U16856 ( .A1(n15276), .A2(n15296), .ZN(n15280) );
  XNOR2_X1 U16857 ( .A(n15277), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n15278) );
  NAND2_X1 U16858 ( .A1(n15302), .A2(n15278), .ZN(n15279) );
  NAND4_X1 U16859 ( .A1(n15282), .A2(n15281), .A3(n15280), .A4(n15279), .ZN(
        P2_U3229) );
  AOI22_X1 U16860 ( .A1(n15294), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n15293) );
  NAND2_X1 U16861 ( .A1(n15299), .A2(n15283), .ZN(n15292) );
  OAI211_X1 U16862 ( .C1(n15286), .C2(n15285), .A(n15296), .B(n15284), .ZN(
        n15291) );
  OAI211_X1 U16863 ( .C1(n15289), .C2(n15288), .A(n15302), .B(n15287), .ZN(
        n15290) );
  NAND4_X1 U16864 ( .A1(n15293), .A2(n15292), .A3(n15291), .A4(n15290), .ZN(
        P2_U3230) );
  AOI22_X1 U16865 ( .A1(n15294), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n15308) );
  OAI211_X1 U16866 ( .C1(n15298), .C2(n15297), .A(n15296), .B(n15295), .ZN(
        n15307) );
  NAND2_X1 U16867 ( .A1(n15300), .A2(n15299), .ZN(n15306) );
  OAI211_X1 U16868 ( .C1(n15304), .C2(n15303), .A(n15302), .B(n15301), .ZN(
        n15305) );
  NAND4_X1 U16869 ( .A1(n15308), .A2(n15307), .A3(n15306), .A4(n15305), .ZN(
        P2_U3231) );
  OAI21_X1 U16870 ( .B1(n15428), .B2(n15409), .A(n15362), .ZN(n15311) );
  INV_X1 U16871 ( .A(n15309), .ZN(n15310) );
  NAND2_X1 U16872 ( .A1(n15311), .A2(n15310), .ZN(n15360) );
  INV_X1 U16873 ( .A(n15362), .ZN(n15316) );
  NAND2_X1 U16874 ( .A1(n15313), .A2(n15312), .ZN(n15359) );
  OAI22_X1 U16875 ( .A1(n15316), .A2(n15315), .B1(n15314), .B2(n15359), .ZN(
        n15317) );
  AOI211_X1 U16876 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n15318), .A(n15360), .B(
        n15317), .ZN(n15319) );
  AOI22_X1 U16877 ( .A1(n15320), .A2(n9364), .B1(n15319), .B2(n13472), .ZN(
        P2_U3265) );
  NOR2_X1 U16878 ( .A1(n15353), .A2(n15322), .ZN(P2_U3266) );
  INV_X1 U16879 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15323) );
  NOR2_X1 U16880 ( .A1(n15353), .A2(n15323), .ZN(P2_U3267) );
  INV_X1 U16881 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15324) );
  NOR2_X1 U16882 ( .A1(n15353), .A2(n15324), .ZN(P2_U3268) );
  INV_X1 U16883 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15325) );
  NOR2_X1 U16884 ( .A1(n15353), .A2(n15325), .ZN(P2_U3269) );
  INV_X1 U16885 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15326) );
  NOR2_X1 U16886 ( .A1(n15336), .A2(n15326), .ZN(P2_U3270) );
  INV_X1 U16887 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15327) );
  NOR2_X1 U16888 ( .A1(n15336), .A2(n15327), .ZN(P2_U3271) );
  NOR2_X1 U16889 ( .A1(n15336), .A2(n15328), .ZN(P2_U3272) );
  INV_X1 U16890 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15329) );
  NOR2_X1 U16891 ( .A1(n15336), .A2(n15329), .ZN(P2_U3273) );
  INV_X1 U16892 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15330) );
  NOR2_X1 U16893 ( .A1(n15336), .A2(n15330), .ZN(P2_U3274) );
  INV_X1 U16894 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15331) );
  NOR2_X1 U16895 ( .A1(n15336), .A2(n15331), .ZN(P2_U3275) );
  INV_X1 U16896 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15332) );
  NOR2_X1 U16897 ( .A1(n15336), .A2(n15332), .ZN(P2_U3276) );
  INV_X1 U16898 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U16899 ( .A1(n15336), .A2(n15333), .ZN(P2_U3277) );
  INV_X1 U16900 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15334) );
  NOR2_X1 U16901 ( .A1(n15336), .A2(n15334), .ZN(P2_U3278) );
  INV_X1 U16902 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U16903 ( .A1(n15336), .A2(n15335), .ZN(P2_U3279) );
  INV_X1 U16904 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15337) );
  NOR2_X1 U16905 ( .A1(n15353), .A2(n15337), .ZN(P2_U3280) );
  NOR2_X1 U16906 ( .A1(n15353), .A2(n15338), .ZN(P2_U3281) );
  INV_X1 U16907 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15339) );
  NOR2_X1 U16908 ( .A1(n15353), .A2(n15339), .ZN(P2_U3282) );
  INV_X1 U16909 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15340) );
  NOR2_X1 U16910 ( .A1(n15353), .A2(n15340), .ZN(P2_U3283) );
  NOR2_X1 U16911 ( .A1(n15353), .A2(n15341), .ZN(P2_U3284) );
  NOR2_X1 U16912 ( .A1(n15353), .A2(n15342), .ZN(P2_U3285) );
  INV_X1 U16913 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15343) );
  NOR2_X1 U16914 ( .A1(n15353), .A2(n15343), .ZN(P2_U3286) );
  INV_X1 U16915 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15344) );
  NOR2_X1 U16916 ( .A1(n15353), .A2(n15344), .ZN(P2_U3287) );
  NOR2_X1 U16917 ( .A1(n15353), .A2(n15345), .ZN(P2_U3288) );
  NOR2_X1 U16918 ( .A1(n15353), .A2(n15346), .ZN(P2_U3289) );
  INV_X1 U16919 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15347) );
  NOR2_X1 U16920 ( .A1(n15353), .A2(n15347), .ZN(P2_U3290) );
  NOR2_X1 U16921 ( .A1(n15353), .A2(n15348), .ZN(P2_U3291) );
  INV_X1 U16922 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U16923 ( .A1(n15353), .A2(n15349), .ZN(P2_U3292) );
  INV_X1 U16924 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15350) );
  NOR2_X1 U16925 ( .A1(n15353), .A2(n15350), .ZN(P2_U3293) );
  INV_X1 U16926 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15351) );
  NOR2_X1 U16927 ( .A1(n15353), .A2(n15351), .ZN(P2_U3294) );
  INV_X1 U16928 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15352) );
  NOR2_X1 U16929 ( .A1(n15353), .A2(n15352), .ZN(P2_U3295) );
  MUX2_X1 U16930 ( .A(P2_D_REG_0__SCAN_IN), .B(n15354), .S(n15353), .Z(
        P2_U3416) );
  AOI22_X1 U16931 ( .A1(n15358), .A2(n15357), .B1(n15356), .B2(n15355), .ZN(
        P2_U3417) );
  INV_X1 U16932 ( .A(n15359), .ZN(n15361) );
  AOI211_X1 U16933 ( .C1(n15363), .C2(n15362), .A(n15361), .B(n15360), .ZN(
        n15433) );
  AOI22_X1 U16934 ( .A1(n15431), .A2(n15433), .B1(n15364), .B2(n15429), .ZN(
        P2_U3430) );
  INV_X1 U16935 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U16936 ( .A1(n15431), .A2(n15366), .B1(n15365), .B2(n15429), .ZN(
        P2_U3433) );
  INV_X1 U16937 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15367) );
  AOI22_X1 U16938 ( .A1(n15431), .A2(n15368), .B1(n15367), .B2(n15429), .ZN(
        P2_U3436) );
  AOI21_X1 U16939 ( .B1(n15421), .B2(n15370), .A(n15369), .ZN(n15371) );
  OAI211_X1 U16940 ( .C1(n15405), .C2(n15373), .A(n15372), .B(n15371), .ZN(
        n15374) );
  INV_X1 U16941 ( .A(n15374), .ZN(n15434) );
  INV_X1 U16942 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15375) );
  AOI22_X1 U16943 ( .A1(n15431), .A2(n15434), .B1(n15375), .B2(n15429), .ZN(
        P2_U3439) );
  INV_X1 U16944 ( .A(n15376), .ZN(n15383) );
  NOR2_X1 U16945 ( .A1(n15376), .A2(n15423), .ZN(n15382) );
  OAI211_X1 U16946 ( .C1(n15380), .C2(n15379), .A(n15378), .B(n15377), .ZN(
        n15381) );
  AOI211_X1 U16947 ( .C1(n15428), .C2(n15383), .A(n15382), .B(n15381), .ZN(
        n15435) );
  INV_X1 U16948 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15384) );
  AOI22_X1 U16949 ( .A1(n15431), .A2(n15435), .B1(n15384), .B2(n15429), .ZN(
        P2_U3442) );
  AND2_X1 U16950 ( .A1(n15385), .A2(n15421), .ZN(n15386) );
  NOR2_X1 U16951 ( .A1(n15387), .A2(n15386), .ZN(n15390) );
  OR2_X1 U16952 ( .A1(n15388), .A2(n15405), .ZN(n15389) );
  AND3_X1 U16953 ( .A1(n15391), .A2(n15390), .A3(n15389), .ZN(n15436) );
  INV_X1 U16954 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15392) );
  AOI22_X1 U16955 ( .A1(n15431), .A2(n15436), .B1(n15392), .B2(n15429), .ZN(
        P2_U3445) );
  AND2_X1 U16956 ( .A1(n15393), .A2(n15421), .ZN(n15394) );
  NOR2_X1 U16957 ( .A1(n15395), .A2(n15394), .ZN(n15398) );
  OR2_X1 U16958 ( .A1(n15396), .A2(n15405), .ZN(n15397) );
  AND3_X1 U16959 ( .A1(n15399), .A2(n15398), .A3(n15397), .ZN(n15437) );
  INV_X1 U16960 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15400) );
  AOI22_X1 U16961 ( .A1(n15431), .A2(n15437), .B1(n15400), .B2(n15429), .ZN(
        P2_U3448) );
  AOI21_X1 U16962 ( .B1(n15402), .B2(n15421), .A(n15401), .ZN(n15404) );
  OAI211_X1 U16963 ( .C1(n15406), .C2(n15405), .A(n15404), .B(n15403), .ZN(
        n15407) );
  AOI21_X1 U16964 ( .B1(n15409), .B2(n15408), .A(n15407), .ZN(n15438) );
  INV_X1 U16965 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U16966 ( .A1(n15431), .A2(n15438), .B1(n15410), .B2(n15429), .ZN(
        P2_U3451) );
  INV_X1 U16967 ( .A(n15414), .ZN(n15417) );
  AOI21_X1 U16968 ( .B1(n15421), .B2(n15412), .A(n15411), .ZN(n15413) );
  OAI21_X1 U16969 ( .B1(n15414), .B2(n15423), .A(n15413), .ZN(n15415) );
  AOI211_X1 U16970 ( .C1(n15428), .C2(n15417), .A(n15416), .B(n15415), .ZN(
        n15440) );
  INV_X1 U16971 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U16972 ( .A1(n15431), .A2(n15440), .B1(n15418), .B2(n15429), .ZN(
        P2_U3457) );
  INV_X1 U16973 ( .A(n15424), .ZN(n15427) );
  AOI21_X1 U16974 ( .B1(n15421), .B2(n15420), .A(n15419), .ZN(n15422) );
  OAI21_X1 U16975 ( .B1(n15424), .B2(n15423), .A(n15422), .ZN(n15425) );
  AOI211_X1 U16976 ( .C1(n15428), .C2(n15427), .A(n15426), .B(n15425), .ZN(
        n15442) );
  INV_X1 U16977 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15430) );
  AOI22_X1 U16978 ( .A1(n15431), .A2(n15442), .B1(n15430), .B2(n15429), .ZN(
        P2_U3460) );
  INV_X1 U16979 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15432) );
  AOI22_X1 U16980 ( .A1(n15443), .A2(n15433), .B1(n15432), .B2(n15441), .ZN(
        P2_U3499) );
  AOI22_X1 U16981 ( .A1(n15443), .A2(n15434), .B1(n9223), .B2(n15441), .ZN(
        P2_U3502) );
  AOI22_X1 U16982 ( .A1(n15443), .A2(n15435), .B1(n9231), .B2(n15441), .ZN(
        P2_U3503) );
  AOI22_X1 U16983 ( .A1(n15443), .A2(n15436), .B1(n9233), .B2(n15441), .ZN(
        P2_U3504) );
  AOI22_X1 U16984 ( .A1(n15443), .A2(n15437), .B1(n9235), .B2(n15441), .ZN(
        P2_U3505) );
  AOI22_X1 U16985 ( .A1(n15443), .A2(n15438), .B1(n9236), .B2(n15441), .ZN(
        P2_U3506) );
  AOI22_X1 U16986 ( .A1(n15443), .A2(n15440), .B1(n15439), .B2(n15441), .ZN(
        P2_U3508) );
  AOI22_X1 U16987 ( .A1(n15443), .A2(n15442), .B1(n9384), .B2(n15441), .ZN(
        P2_U3509) );
  NOR2_X1 U16988 ( .A1(P3_U3897), .A2(n15458), .ZN(P3_U3150) );
  AOI21_X1 U16989 ( .B1(n15446), .B2(n15445), .A(n15444), .ZN(n15466) );
  INV_X1 U16990 ( .A(n15447), .ZN(n15449) );
  NAND2_X1 U16991 ( .A1(n15449), .A2(n15448), .ZN(n15450) );
  XNOR2_X1 U16992 ( .A(n15451), .B(n15450), .ZN(n15455) );
  OAI22_X1 U16993 ( .A1(n15455), .A2(n15454), .B1(n15453), .B2(n15452), .ZN(
        n15456) );
  AOI211_X1 U16994 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15458), .A(n15457), .B(
        n15456), .ZN(n15464) );
  OAI21_X1 U16995 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15460), .A(n15459), .ZN(
        n15462) );
  NAND2_X1 U16996 ( .A1(n15462), .A2(n15461), .ZN(n15463) );
  OAI211_X1 U16997 ( .C1(n15466), .C2(n15465), .A(n15464), .B(n15463), .ZN(
        P3_U3191) );
  AOI22_X1 U16998 ( .A1(n15521), .A2(n15468), .B1(n15467), .B2(n15519), .ZN(
        P3_U3393) );
  INV_X1 U16999 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15474) );
  INV_X1 U17000 ( .A(n15469), .ZN(n15473) );
  INV_X1 U17001 ( .A(n15470), .ZN(n15472) );
  AOI211_X1 U17002 ( .C1(n15473), .C2(n15509), .A(n15472), .B(n15471), .ZN(
        n15523) );
  AOI22_X1 U17003 ( .A1(n15521), .A2(n15474), .B1(n15523), .B2(n15519), .ZN(
        P3_U3396) );
  INV_X1 U17004 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15479) );
  OAI22_X1 U17005 ( .A1(n15476), .A2(n15497), .B1(n15515), .B2(n15475), .ZN(
        n15477) );
  NOR2_X1 U17006 ( .A1(n15478), .A2(n15477), .ZN(n15525) );
  AOI22_X1 U17007 ( .A1(n15521), .A2(n15479), .B1(n15525), .B2(n15519), .ZN(
        P3_U3399) );
  INV_X1 U17008 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15484) );
  OAI22_X1 U17009 ( .A1(n15481), .A2(n15497), .B1(n15515), .B2(n15480), .ZN(
        n15482) );
  NOR2_X1 U17010 ( .A1(n15483), .A2(n15482), .ZN(n15527) );
  AOI22_X1 U17011 ( .A1(n15521), .A2(n15484), .B1(n15527), .B2(n15519), .ZN(
        P3_U3402) );
  INV_X1 U17012 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15490) );
  INV_X1 U17013 ( .A(n15485), .ZN(n15487) );
  OAI22_X1 U17014 ( .A1(n15487), .A2(n15497), .B1(n15515), .B2(n15486), .ZN(
        n15488) );
  NOR2_X1 U17015 ( .A1(n15489), .A2(n15488), .ZN(n15529) );
  AOI22_X1 U17016 ( .A1(n15521), .A2(n15490), .B1(n15529), .B2(n15519), .ZN(
        P3_U3405) );
  INV_X1 U17017 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15495) );
  OAI22_X1 U17018 ( .A1(n15492), .A2(n15497), .B1(n15491), .B2(n15515), .ZN(
        n15493) );
  NOR2_X1 U17019 ( .A1(n15494), .A2(n15493), .ZN(n15531) );
  AOI22_X1 U17020 ( .A1(n15521), .A2(n15495), .B1(n15531), .B2(n15519), .ZN(
        P3_U3408) );
  INV_X1 U17021 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15501) );
  OAI22_X1 U17022 ( .A1(n15498), .A2(n15497), .B1(n15515), .B2(n15496), .ZN(
        n15499) );
  NOR2_X1 U17023 ( .A1(n15500), .A2(n15499), .ZN(n15533) );
  AOI22_X1 U17024 ( .A1(n15521), .A2(n15501), .B1(n15533), .B2(n15519), .ZN(
        P3_U3411) );
  INV_X1 U17025 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15506) );
  NOR2_X1 U17026 ( .A1(n15502), .A2(n15515), .ZN(n15504) );
  AOI211_X1 U17027 ( .C1(n15509), .C2(n15505), .A(n15504), .B(n15503), .ZN(
        n15535) );
  AOI22_X1 U17028 ( .A1(n15521), .A2(n15506), .B1(n15535), .B2(n15519), .ZN(
        P3_U3414) );
  AOI22_X1 U17029 ( .A1(n15510), .A2(n15509), .B1(n15508), .B2(n15507), .ZN(
        n15511) );
  AND2_X1 U17030 ( .A1(n15512), .A2(n15511), .ZN(n15537) );
  AOI22_X1 U17031 ( .A1(n15521), .A2(n7072), .B1(n15537), .B2(n15519), .ZN(
        P3_U3417) );
  OAI21_X1 U17032 ( .B1(n15515), .B2(n15514), .A(n15513), .ZN(n15516) );
  AOI21_X1 U17033 ( .B1(n15518), .B2(n15517), .A(n15516), .ZN(n15539) );
  AOI22_X1 U17034 ( .A1(n15521), .A2(n15520), .B1(n15539), .B2(n15519), .ZN(
        P3_U3420) );
  AOI22_X1 U17035 ( .A1(n15540), .A2(n15523), .B1(n15522), .B2(n15538), .ZN(
        P3_U3461) );
  INV_X1 U17036 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15524) );
  AOI22_X1 U17037 ( .A1(n15540), .A2(n15525), .B1(n15524), .B2(n15538), .ZN(
        P3_U3462) );
  AOI22_X1 U17038 ( .A1(n15540), .A2(n15527), .B1(n15526), .B2(n15538), .ZN(
        P3_U3463) );
  INV_X1 U17039 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15528) );
  AOI22_X1 U17040 ( .A1(n15540), .A2(n15529), .B1(n15528), .B2(n15538), .ZN(
        P3_U3464) );
  AOI22_X1 U17041 ( .A1(n15540), .A2(n15531), .B1(n15530), .B2(n15538), .ZN(
        P3_U3465) );
  INV_X1 U17042 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U17043 ( .A1(n15540), .A2(n15533), .B1(n15532), .B2(n15538), .ZN(
        P3_U3466) );
  AOI22_X1 U17044 ( .A1(n15540), .A2(n15535), .B1(n15534), .B2(n15538), .ZN(
        P3_U3467) );
  AOI22_X1 U17045 ( .A1(n15540), .A2(n15537), .B1(n15536), .B2(n15538), .ZN(
        P3_U3468) );
  AOI22_X1 U17046 ( .A1(n15540), .A2(n15539), .B1(n10604), .B2(n15538), .ZN(
        P3_U3469) );
  XOR2_X1 U17047 ( .A(n15542), .B(n15541), .Z(SUB_1596_U59) );
  XNOR2_X1 U17048 ( .A(n15543), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17049 ( .B1(n15544), .B2(n9371), .A(n15551), .ZN(SUB_1596_U53) );
  XOR2_X1 U17050 ( .A(n15545), .B(n15546), .Z(SUB_1596_U56) );
  NOR2_X1 U17051 ( .A1(n15548), .A2(n15547), .ZN(n15549) );
  XOR2_X1 U17052 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15549), .Z(SUB_1596_U60) );
  XOR2_X1 U17053 ( .A(n15551), .B(n15550), .Z(SUB_1596_U5) );
  CLKBUF_X2 U7305 ( .A(n14123), .Z(n14206) );
  CLKBUF_X3 U7390 ( .A(n8486), .Z(n6567) );
  INV_X4 U7392 ( .A(n12129), .ZN(n12103) );
  INV_X4 U7394 ( .A(n8312), .ZN(n14077) );
  INV_X2 U7479 ( .A(n14589), .ZN(n8988) );
endmodule

