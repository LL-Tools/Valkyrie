

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738;

  OAI21_X1 U3670 ( .B1(n4500), .B2(n3780), .A(n3778), .ZN(n6942) );
  AOI21_X1 U3671 ( .B1(n4041), .B2(n4049), .A(n4209), .ZN(n4057) );
  CLKBUF_X2 U3672 ( .A(n4970), .Z(n3673) );
  CLKBUF_X2 U3673 ( .A(n3676), .Z(n3666) );
  CLKBUF_X2 U3674 ( .A(n3944), .Z(n4979) );
  CLKBUF_X2 U3675 ( .A(n4115), .Z(n7224) );
  INV_X1 U3676 ( .A(n3662), .ZN(n3949) );
  AND2_X1 U3677 ( .A1(n3814), .A2(n5282), .ZN(n3665) );
  INV_X1 U3678 ( .A(n3909), .ZN(n3636) );
  INV_X2 U3679 ( .A(n3636), .ZN(n3637) );
  AND2_X1 U3680 ( .A1(n5133), .A2(n5282), .ZN(n3677) );
  NAND2_X1 U3681 ( .A1(n3989), .A2(n4017), .ZN(n4440) );
  CLKBUF_X2 U3682 ( .A(n4301), .Z(n4448) );
  NOR2_X1 U3683 ( .A1(n7313), .A2(n6513), .ZN(n6500) );
  NAND2_X1 U3684 ( .A1(n3954), .A2(n4503), .ZN(n3986) );
  NOR2_X1 U3685 ( .A1(n7317), .A2(n7585), .ZN(n7598) );
  OR2_X1 U3686 ( .A1(n7693), .A2(n7671), .ZN(n5167) );
  NAND2_X1 U3687 ( .A1(n3971), .A2(n3988), .ZN(n4330) );
  INV_X1 U3688 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7691) );
  INV_X1 U3689 ( .A(n4017), .ZN(n3669) );
  NAND4_X1 U3690 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3638)
         );
  AND2_X2 U3691 ( .A1(n5271), .A2(n3820), .ZN(n3944) );
  AND2_X1 U3692 ( .A1(n3814), .A2(n5282), .ZN(n3639) );
  AND2_X1 U3693 ( .A1(n3814), .A2(n5282), .ZN(n4977) );
  BUF_X1 U3694 ( .A(n3945), .Z(n3640) );
  BUF_X2 U3695 ( .A(n3945), .Z(n3641) );
  BUF_X4 U3696 ( .A(n3945), .Z(n3642) );
  AND2_X1 U3697 ( .A1(n3814), .A2(n5271), .ZN(n3643) );
  AND2_X2 U3698 ( .A1(n3814), .A2(n5271), .ZN(n3678) );
  AND2_X1 U3699 ( .A1(n3814), .A2(n5271), .ZN(n3909) );
  AND2_X1 U3700 ( .A1(n4725), .A2(n4724), .ZN(n6495) );
  INV_X1 U3701 ( .A(n6568), .ZN(n3645) );
  CLKBUF_X2 U3702 ( .A(n5366), .Z(n5411) );
  CLKBUF_X1 U3703 ( .A(n5090), .Z(n3667) );
  NAND2_X1 U3704 ( .A1(n4052), .A2(n4051), .ZN(n5552) );
  BUF_X1 U3705 ( .A(n5087), .Z(n3668) );
  AND3_X1 U3706 ( .A1(n3801), .A2(n3947), .A3(n3946), .ZN(n3969) );
  AND4_X1 U3707 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(n3878)
         );
  AND4_X1 U3708 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3899)
         );
  CLKBUF_X2 U3709 ( .A(n4971), .Z(n4908) );
  BUF_X2 U3710 ( .A(n4676), .Z(n4950) );
  BUF_X2 U3711 ( .A(n3927), .Z(n4972) );
  AND2_X2 U3713 ( .A1(n3820), .A2(n3819), .ZN(n3945) );
  INV_X2 U3714 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3804) );
  OR2_X1 U3715 ( .A1(n6953), .A2(n6952), .ZN(n6955) );
  AND2_X1 U3716 ( .A1(n5056), .A2(n5055), .ZN(n5057) );
  NOR2_X1 U3717 ( .A1(n6390), .A2(n7595), .ZN(n3748) );
  AOI21_X1 U3718 ( .B1(n6989), .B2(n3769), .A(n3767), .ZN(n3766) );
  OR2_X1 U3719 ( .A1(n6550), .A2(n7059), .ZN(n5056) );
  CLKBUF_X1 U3720 ( .A(n6437), .Z(n6438) );
  NAND2_X1 U3721 ( .A1(n4228), .A2(n4227), .ZN(n7060) );
  NAND2_X1 U3722 ( .A1(n6317), .A2(n4226), .ZN(n4228) );
  CLKBUF_X1 U3723 ( .A(n6532), .Z(n6533) );
  AND2_X2 U3724 ( .A1(n6532), .A2(n3789), .ZN(n6460) );
  OAI21_X1 U3725 ( .B1(n4235), .B2(n3768), .A(n4234), .ZN(n3767) );
  NOR2_X1 U3726 ( .A1(n3758), .A2(n3755), .ZN(n3754) );
  OR2_X1 U3727 ( .A1(n3649), .A2(n6170), .ZN(n3648) );
  XNOR2_X1 U3728 ( .A(n4451), .B(n5029), .ZN(n6381) );
  NOR2_X1 U3729 ( .A1(n4235), .A2(n3771), .ZN(n3769) );
  XNOR2_X1 U3730 ( .A(n4206), .B(n5865), .ZN(n5771) );
  AND2_X1 U3731 ( .A1(n7510), .A2(n5039), .ZN(n7570) );
  INV_X8 U3732 ( .A(n7031), .ZN(n7030) );
  NAND2_X1 U3733 ( .A1(n4205), .A2(n4204), .ZN(n4206) );
  INV_X4 U3734 ( .A(n7016), .ZN(n7031) );
  OR2_X1 U3735 ( .A1(n4561), .A2(n4210), .ZN(n4205) );
  NAND2_X1 U3736 ( .A1(n4541), .A2(n4540), .ZN(n5492) );
  AND2_X1 U3737 ( .A1(n3688), .A2(n4128), .ZN(n7388) );
  NOR2_X1 U3738 ( .A1(n5776), .A2(n7293), .ZN(n5930) );
  NAND2_X1 U3739 ( .A1(n4522), .A2(n4521), .ZN(n5194) );
  CLKBUF_X1 U3740 ( .A(n7520), .Z(n7610) );
  OR2_X1 U3741 ( .A1(n5182), .A2(n4520), .ZN(n5201) );
  AND2_X1 U3742 ( .A1(n6371), .A2(REIP_REG_3__SCAN_IN), .ZN(n6143) );
  NOR3_X1 U3743 ( .A1(n7501), .A2(n7506), .A3(n7507), .ZN(n6371) );
  AND2_X1 U3744 ( .A1(n5179), .A2(n5180), .ZN(n5182) );
  NAND2_X1 U3745 ( .A1(n4123), .A2(n4122), .ZN(n5297) );
  NAND2_X1 U3746 ( .A1(n5108), .A2(n5107), .ZN(n7425) );
  INV_X1 U3747 ( .A(n4090), .ZN(n4088) );
  AOI21_X1 U3748 ( .B1(n5087), .B2(n7691), .A(n4087), .ZN(n4090) );
  XNOR2_X1 U3749 ( .A(n5289), .B(n5287), .ZN(n5090) );
  AOI21_X1 U3750 ( .B1(n5552), .B2(n4508), .A(n7669), .ZN(n5115) );
  NAND2_X1 U3751 ( .A1(n4104), .A2(n4103), .ZN(n5289) );
  INV_X1 U3752 ( .A(n5167), .ZN(n3646) );
  NOR2_X1 U3753 ( .A1(n6165), .A2(n6164), .ZN(n6198) );
  NAND2_X1 U3754 ( .A1(n4293), .A2(n4292), .ZN(n7693) );
  OAI21_X1 U3755 ( .B1(n4291), .B2(n4289), .A(n3745), .ZN(n4293) );
  NAND2_X1 U3756 ( .A1(n4509), .A2(n7691), .ZN(n4047) );
  AND2_X1 U3757 ( .A1(n4740), .A2(n4739), .ZN(n6496) );
  NAND2_X1 U3758 ( .A1(n4110), .A2(n4109), .ZN(n5287) );
  NAND2_X1 U3759 ( .A1(n4462), .A2(n3679), .ZN(n4021) );
  NAND2_X1 U3760 ( .A1(n4260), .A2(n3743), .ZN(n4269) );
  INV_X1 U3761 ( .A(n4306), .ZN(n3971) );
  AND3_X1 U3762 ( .A1(n4024), .A2(n4020), .A3(n4019), .ZN(n4060) );
  NAND2_X1 U3763 ( .A1(n3966), .A2(n3967), .ZN(n5130) );
  NAND2_X1 U3764 ( .A1(n4440), .A2(n4448), .ZN(n5228) );
  CLKBUF_X2 U3765 ( .A(n3987), .Z(n3675) );
  NAND2_X1 U3766 ( .A1(n5191), .A2(n4448), .ZN(n4437) );
  NAND2_X1 U3767 ( .A1(n4256), .A2(n4073), .ZN(n4288) );
  AND2_X1 U3768 ( .A1(n3951), .A2(n4508), .ZN(n4295) );
  INV_X2 U3769 ( .A(n3969), .ZN(n4312) );
  INV_X1 U3770 ( .A(n4017), .ZN(n3922) );
  OR2_X1 U3771 ( .A1(n4016), .A2(n4015), .ZN(n4214) );
  AND4_X2 U3772 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3662)
         );
  NAND2_X2 U3773 ( .A1(n3839), .A2(n3838), .ZN(n5073) );
  AND4_X1 U3774 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3921)
         );
  AND4_X1 U3775 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  AND4_X1 U3776 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3876)
         );
  AND4_X1 U3777 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3947)
         );
  AND4_X1 U3778 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3828)
         );
  AND4_X1 U3779 ( .A1(n3847), .A2(n3846), .A3(n3845), .A4(n3844), .ZN(n3858)
         );
  AND4_X1 U3780 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3838)
         );
  AND4_X1 U3781 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3877)
         );
  AND4_X1 U3782 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3879)
         );
  AND4_X1 U3783 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3856)
         );
  AND4_X1 U3784 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3900)
         );
  AND4_X1 U3785 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3857)
         );
  AND4_X1 U3786 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3898)
         );
  AND4_X1 U3787 ( .A1(n3843), .A2(n3842), .A3(n3841), .A4(n3840), .ZN(n3859)
         );
  AND4_X1 U3788 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3920)
         );
  AND4_X1 U3789 ( .A1(n3832), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(n3839)
         );
  AND4_X1 U3790 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3825)
         );
  AND4_X1 U3791 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3919)
         );
  AND4_X1 U3792 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3826)
         );
  AND4_X1 U3793 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3827)
         );
  AND4_X1 U3794 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3918)
         );
  NAND2_X2 U3795 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7706), .ZN(n7334) );
  BUF_X2 U3796 ( .A(n3998), .Z(n4978) );
  NAND2_X2 U3797 ( .A1(n7706), .A2(n7702), .ZN(n7342) );
  BUF_X2 U3798 ( .A(n3936), .Z(n4955) );
  AND2_X2 U3799 ( .A1(n5274), .A2(n5144), .ZN(n4115) );
  AND2_X2 U3800 ( .A1(n3804), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5274)
         );
  AND2_X2 U3801 ( .A1(n5129), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3814)
         );
  AND2_X2 U3802 ( .A1(n3809), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5133)
         );
  INV_X2 U3803 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n7669) );
  AND2_X2 U3804 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5282) );
  AND2_X2 U3805 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5144) );
  NOR2_X2 U3806 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3819) );
  NOR2_X2 U3807 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3820) );
  NAND2_X1 U3808 ( .A1(n3696), .A2(n3650), .ZN(n3647) );
  AND2_X2 U3809 ( .A1(n3647), .A2(n3648), .ZN(n6214) );
  INV_X1 U3810 ( .A(n4219), .ZN(n3649) );
  AND2_X1 U3811 ( .A1(n4218), .A2(n4219), .ZN(n3650) );
  OAI21_X1 U3812 ( .B1(n5085), .B2(n4686), .A(n4850), .ZN(n4520) );
  AND2_X2 U3813 ( .A1(n3652), .A2(n4088), .ZN(n3651) );
  AND2_X2 U3814 ( .A1(n4063), .A2(n4062), .ZN(n3652) );
  NOR2_X2 U3815 ( .A1(n6351), .A2(n3653), .ZN(n6497) );
  NAND2_X1 U3816 ( .A1(n4724), .A2(n6496), .ZN(n3653) );
  AND2_X1 U3817 ( .A1(n6302), .A2(n3654), .ZN(n6336) );
  AND2_X1 U3818 ( .A1(n6304), .A2(n3655), .ZN(n3654) );
  INV_X1 U3819 ( .A(n6337), .ZN(n3655) );
  AND2_X1 U3820 ( .A1(n4017), .A2(n3965), .ZN(n5191) );
  AND2_X1 U3821 ( .A1(n3954), .A2(n3965), .ZN(n4294) );
  NAND2_X1 U3822 ( .A1(n6246), .A2(n3659), .ZN(n3656) );
  AND2_X2 U3823 ( .A1(n3656), .A2(n3657), .ZN(n6317) );
  OR2_X1 U3824 ( .A1(n3658), .A2(n3777), .ZN(n3657) );
  INV_X1 U3825 ( .A(n4225), .ZN(n3658) );
  AND2_X1 U3826 ( .A1(n6247), .A2(n4225), .ZN(n3659) );
  CLKBUF_X1 U3827 ( .A(n7399), .Z(n3660) );
  AND2_X1 U3828 ( .A1(n4064), .A2(n3772), .ZN(n3661) );
  NAND2_X2 U3829 ( .A1(n4022), .A2(n4021), .ZN(n4066) );
  NAND2_X1 U3830 ( .A1(n4150), .A2(n4149), .ZN(n4173) );
  AND2_X1 U3831 ( .A1(n3819), .A2(n5144), .ZN(n3663) );
  AND2_X2 U3832 ( .A1(n3819), .A2(n5144), .ZN(n3664) );
  AND2_X2 U3833 ( .A1(n5271), .A2(n5133), .ZN(n4970) );
  OAI21_X1 U3834 ( .B1(n4561), .B2(n4686), .A(n4560), .ZN(n5448) );
  OAI211_X2 U3835 ( .C1(n4068), .C2(n3781), .A(n3975), .B(n3775), .ZN(n4064)
         );
  AND2_X1 U3836 ( .A1(n5133), .A2(n5282), .ZN(n3676) );
  INV_X2 U3837 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3731) );
  OR2_X1 U3838 ( .A1(n5083), .A2(n4210), .ZN(n3688) );
  NAND2_X1 U3839 ( .A1(n3765), .A2(n5216), .ZN(n7382) );
  NAND2_X2 U3840 ( .A1(n4124), .A2(n3706), .ZN(n5085) );
  NAND2_X2 U3841 ( .A1(n3652), .A2(n4088), .ZN(n4124) );
  AND2_X1 U3842 ( .A1(n4503), .A2(n3952), .ZN(n4508) );
  AND3_X1 U3843 ( .A1(n3949), .A2(STATE2_REG_0__SCAN_IN), .A3(n4017), .ZN(
        n4275) );
  NAND2_X2 U3844 ( .A1(n6460), .A2(n6461), .ZN(n6448) );
  OAI21_X2 U3845 ( .B1(n7390), .B2(n4468), .A(n7388), .ZN(n3764) );
  NAND2_X2 U3846 ( .A1(n4101), .A2(n4100), .ZN(n7390) );
  NAND2_X1 U3847 ( .A1(n3662), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4256) );
  NOR2_X4 U3848 ( .A1(n6448), .A2(n6450), .ZN(n6437) );
  NAND2_X2 U3849 ( .A1(n3702), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4068) );
  OAI21_X2 U3850 ( .B1(n7060), .B2(n4230), .A(n4229), .ZN(n7052) );
  OAI21_X2 U3851 ( .B1(n4068), .B2(n3809), .A(n3977), .ZN(n4022) );
  OAI21_X2 U3852 ( .B1(n6989), .B2(n3689), .A(n3770), .ZN(n7024) );
  NAND2_X2 U3853 ( .A1(n7052), .A2(n4231), .ZN(n6989) );
  OAI22_X1 U3854 ( .A1(n7000), .A2(n6982), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6991), .ZN(n6983) );
  XNOR2_X1 U3855 ( .A(n4102), .B(n4103), .ZN(n5087) );
  NOR2_X2 U3856 ( .A1(n5208), .A2(n5360), .ZN(n5361) );
  OAI21_X2 U3857 ( .B1(n5088), .B2(STATE2_REG_0__SCAN_IN), .A(n4005), .ZN(
        n4059) );
  NOR2_X4 U3858 ( .A1(n5710), .A2(n3783), .ZN(n6240) );
  OAI21_X2 U3859 ( .B1(n6272), .B2(n6273), .A(n4653), .ZN(n6302) );
  NAND2_X2 U3860 ( .A1(n4577), .A2(n4576), .ZN(n5710) );
  AND2_X1 U3861 ( .A1(n3820), .A2(n5274), .ZN(n3670) );
  AND2_X2 U3862 ( .A1(n3820), .A2(n5274), .ZN(n4025) );
  NAND2_X1 U3863 ( .A1(n5249), .A2(n3965), .ZN(n3671) );
  INV_X4 U3864 ( .A(n4301), .ZN(n3933) );
  AND2_X4 U3865 ( .A1(n5271), .A2(n5144), .ZN(n3672) );
  AND2_X2 U3866 ( .A1(n3820), .A2(n5274), .ZN(n3674) );
  AND2_X4 U3867 ( .A1(n3731), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5271)
         );
  NOR2_X1 U3868 ( .A1(n3965), .A2(n3669), .ZN(n3987) );
  AND2_X4 U3869 ( .A1(n3819), .A2(n5144), .ZN(n4909) );
  AOI21_X1 U3870 ( .B1(n3986), .B2(n5249), .A(n3965), .ZN(n3958) );
  NAND2_X1 U3871 ( .A1(n5851), .A2(n5019), .ZN(n6275) );
  NOR2_X1 U3872 ( .A1(n4312), .A2(n3662), .ZN(n3951) );
  OR2_X1 U3873 ( .A1(n4085), .A2(n4084), .ZN(n4091) );
  NAND2_X1 U3874 ( .A1(n3788), .A2(n6160), .ZN(n3787) );
  INV_X1 U3875 ( .A(n6045), .ZN(n3788) );
  OR2_X1 U3876 ( .A1(n4035), .A2(n4034), .ZN(n4053) );
  NAND2_X1 U3877 ( .A1(n4064), .A2(n3772), .ZN(n4065) );
  NAND2_X1 U3878 ( .A1(n3774), .A2(n3773), .ZN(n3772) );
  OR2_X1 U3879 ( .A1(n3976), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3773)
         );
  NAND2_X1 U3880 ( .A1(n4250), .A2(n7632), .ZN(n4316) );
  OR2_X1 U3881 ( .A1(n7683), .A2(n5015), .ZN(n5016) );
  AND3_X1 U3882 ( .A1(n3935), .A2(n3989), .A3(n3969), .ZN(n3966) );
  INV_X1 U3883 ( .A(n4721), .ZN(n4995) );
  NOR2_X2 U3884 ( .A1(n6962), .A2(n5046), .ZN(n6953) );
  AND2_X1 U3885 ( .A1(n7030), .A2(n6963), .ZN(n5046) );
  NOR2_X1 U3886 ( .A1(n4211), .A2(n4210), .ZN(n4212) );
  NAND2_X1 U3887 ( .A1(n6246), .A2(n6247), .ZN(n4223) );
  NAND2_X1 U3888 ( .A1(n4329), .A2(n4328), .ZN(n4472) );
  NAND2_X1 U3889 ( .A1(n4023), .A2(n3705), .ZN(n3704) );
  INV_X1 U3890 ( .A(n4022), .ZN(n3705) );
  OR2_X1 U3891 ( .A1(n6420), .A2(n5027), .ZN(n6388) );
  NAND2_X1 U3892 ( .A1(n3745), .A2(n3744), .ZN(n3743) );
  AND2_X1 U3893 ( .A1(n3662), .A2(n3952), .ZN(n3880) );
  NAND2_X1 U3894 ( .A1(n4186), .A2(n4185), .ZN(n4196) );
  AND2_X1 U3895 ( .A1(n3974), .A2(n3973), .ZN(n3975) );
  NAND2_X1 U3896 ( .A1(n3776), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U3897 ( .A1(n3662), .A2(n3954), .ZN(n3953) );
  INV_X1 U3898 ( .A(n5249), .ZN(n3989) );
  OR2_X1 U3899 ( .A1(n4864), .A2(n4863), .ZN(n4881) );
  NOR2_X1 U3900 ( .A1(n7006), .A2(n3791), .ZN(n3790) );
  INV_X1 U3901 ( .A(n6535), .ZN(n3791) );
  NOR2_X1 U3902 ( .A1(n4689), .A2(n7691), .ZN(n4991) );
  NOR2_X1 U3903 ( .A1(n3787), .A2(n3786), .ZN(n3785) );
  INV_X1 U3904 ( .A(n6196), .ZN(n3786) );
  INV_X1 U3905 ( .A(n4543), .ZN(n4967) );
  NOR2_X1 U3906 ( .A1(n7143), .A2(n3717), .ZN(n3716) );
  INV_X1 U3907 ( .A(n6537), .ZN(n3717) );
  NOR2_X1 U3908 ( .A1(n6276), .A2(n6277), .ZN(n4392) );
  INV_X1 U3909 ( .A(n6215), .ZN(n3755) );
  INV_X1 U3910 ( .A(n6265), .ZN(n3758) );
  INV_X1 U3911 ( .A(n4220), .ZN(n3757) );
  AND2_X1 U3912 ( .A1(n4105), .A2(n4070), .ZN(n5592) );
  NAND2_X1 U3913 ( .A1(n4061), .A2(n4060), .ZN(n4062) );
  INV_X1 U3914 ( .A(n4086), .ZN(n4087) );
  OR2_X1 U3915 ( .A1(n4304), .A2(n3935), .ZN(n4689) );
  AOI21_X1 U3916 ( .B1(n3935), .B2(n3964), .A(n3981), .ZN(n3948) );
  INV_X1 U3917 ( .A(n3984), .ZN(n3703) );
  NAND2_X1 U3918 ( .A1(n5090), .A2(n7691), .ZN(n4123) );
  AND2_X1 U3919 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n7632), .ZN(n4283)
         );
  NAND2_X1 U3920 ( .A1(n4294), .A2(n4315), .ZN(n3735) );
  NAND2_X1 U3921 ( .A1(n3738), .A2(n3737), .ZN(n3736) );
  NAND2_X1 U3922 ( .A1(n3741), .A2(n3740), .ZN(n3739) );
  INV_X1 U3923 ( .A(n4282), .ZN(n3733) );
  OR2_X1 U3924 ( .A1(n3671), .A2(EBX_REG_1__SCAN_IN), .ZN(n4342) );
  AND2_X1 U3925 ( .A1(n4467), .A2(n4466), .ZN(n5183) );
  INV_X1 U3926 ( .A(n7286), .ZN(n5169) );
  NOR2_X1 U3927 ( .A1(n5167), .A2(n5071), .ZN(n5160) );
  INV_X1 U3928 ( .A(n6403), .ZN(n3792) );
  NAND2_X1 U3929 ( .A1(n4858), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4900)
         );
  AND2_X1 U3930 ( .A1(n4594), .A2(n4593), .ZN(n6045) );
  NAND2_X1 U3931 ( .A1(n6962), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U3932 ( .A1(n4241), .A2(n4240), .ZN(n4500) );
  NAND2_X1 U3933 ( .A1(n6428), .A2(n5060), .ZN(n6406) );
  NAND2_X1 U3934 ( .A1(n7031), .A2(n6963), .ZN(n6952) );
  NAND2_X1 U3935 ( .A1(n4223), .A2(n3777), .ZN(n6295) );
  AND2_X1 U3936 ( .A1(n4224), .A2(n4222), .ZN(n3777) );
  OR2_X1 U3937 ( .A1(n5363), .A2(n3724), .ZN(n6047) );
  OR2_X1 U3938 ( .A1(n3726), .A2(n3725), .ZN(n3724) );
  INV_X1 U3939 ( .A(n5712), .ZN(n3725) );
  NOR2_X1 U3940 ( .A1(n5363), .A2(n3726), .ZN(n5713) );
  NOR2_X1 U3941 ( .A1(n5363), .A2(n5364), .ZN(n5449) );
  AND2_X1 U3942 ( .A1(n4464), .A2(n6323), .ZN(n6175) );
  NAND2_X1 U3943 ( .A1(n4472), .A2(n5183), .ZN(n7462) );
  CLKBUF_X1 U3944 ( .A(n4306), .Z(n4307) );
  NAND2_X1 U3945 ( .A1(n5627), .A2(n5626), .ZN(n5638) );
  NAND2_X1 U3946 ( .A1(n7691), .A2(n5101), .ZN(n5591) );
  INV_X1 U3947 ( .A(n5553), .ZN(n5548) );
  NAND2_X1 U3948 ( .A1(n4048), .A2(n4037), .ZN(n4052) );
  NAND2_X1 U3949 ( .A1(n4047), .A2(n4049), .ZN(n4048) );
  AND2_X1 U3950 ( .A1(n7422), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4321) );
  AND2_X1 U3951 ( .A1(n7668), .A2(n7667), .ZN(n7673) );
  INV_X1 U3952 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7696) );
  INV_X1 U3953 ( .A(n5038), .ZN(n3729) );
  NOR2_X1 U3954 ( .A1(n6385), .A2(n6384), .ZN(n6386) );
  NAND2_X1 U3955 ( .A1(n6487), .A2(n3681), .ZN(n6420) );
  NOR2_X1 U3956 ( .A1(n5849), .A2(n5033), .ZN(n7520) );
  INV_X1 U3957 ( .A(n7376), .ZN(n6541) );
  AND2_X1 U3958 ( .A1(n7376), .A2(n6391), .ZN(n7369) );
  AND2_X1 U3959 ( .A1(n6392), .A2(n5077), .ZN(n7733) );
  XNOR2_X1 U3960 ( .A(n5049), .B(n3797), .ZN(n5059) );
  INV_X1 U3961 ( .A(n7495), .ZN(n7479) );
  AND2_X1 U3962 ( .A1(n4472), .A2(n4455), .ZN(n7495) );
  CLKBUF_X1 U3963 ( .A(n5083), .Z(n5626) );
  NAND2_X1 U3964 ( .A1(n4288), .A2(n4255), .ZN(n3744) );
  INV_X1 U3965 ( .A(n4042), .ZN(n4018) );
  NAND2_X1 U3966 ( .A1(n4271), .A2(n4270), .ZN(n3742) );
  OR2_X1 U3967 ( .A1(n4314), .A2(n7691), .ZN(n4268) );
  AND2_X1 U3968 ( .A1(n5629), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4261)
         );
  OR2_X1 U3969 ( .A1(n4138), .A2(n4137), .ZN(n4163) );
  AND2_X1 U3970 ( .A1(n4303), .A2(n4302), .ZN(n4457) );
  NAND2_X1 U3971 ( .A1(n3983), .A2(n3982), .ZN(n4462) );
  NAND2_X1 U3972 ( .A1(n5249), .A2(n3969), .ZN(n3981) );
  AOI21_X1 U3973 ( .B1(n4273), .B2(n4272), .A(n4246), .ZN(n4252) );
  NAND2_X1 U3974 ( .A1(n3742), .A2(n4278), .ZN(n3741) );
  NOR2_X1 U3975 ( .A1(n4277), .A2(n4313), .ZN(n3740) );
  INV_X1 U3976 ( .A(n3742), .ZN(n3738) );
  INV_X1 U3977 ( .A(n4276), .ZN(n3737) );
  NOR2_X1 U3978 ( .A1(n6453), .A2(n3721), .ZN(n3720) );
  INV_X1 U3979 ( .A(n6465), .ZN(n3721) );
  AND2_X1 U3980 ( .A1(n4775), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4776)
         );
  INV_X1 U3981 ( .A(n6505), .ZN(n4724) );
  XNOR2_X1 U3982 ( .A(n4173), .B(n4171), .ZN(n4548) );
  NAND2_X1 U3983 ( .A1(n6463), .A2(n3718), .ZN(n3723) );
  NOR2_X1 U3984 ( .A1(n3719), .A2(n6441), .ZN(n3718) );
  INV_X1 U3985 ( .A(n3720), .ZN(n3719) );
  NAND2_X1 U3986 ( .A1(n3770), .A2(n3689), .ZN(n3768) );
  NOR2_X1 U3987 ( .A1(n4038), .A2(n7691), .ZN(n4209) );
  NAND2_X1 U3988 ( .A1(n4392), .A2(n3713), .ZN(n3712) );
  INV_X1 U3989 ( .A(n6309), .ZN(n3713) );
  NAND2_X1 U3990 ( .A1(n4370), .A2(n3727), .ZN(n3726) );
  INV_X1 U3991 ( .A(n5364), .ZN(n3727) );
  INV_X1 U3992 ( .A(n4196), .ZN(n4187) );
  INV_X1 U3993 ( .A(n3953), .ZN(n3932) );
  CLKBUF_X1 U3994 ( .A(n4323), .Z(n4324) );
  NOR2_X1 U3995 ( .A1(n3707), .A2(n3969), .ZN(n3970) );
  NAND2_X1 U3996 ( .A1(n3989), .A2(n3922), .ZN(n3707) );
  AND2_X1 U3997 ( .A1(n3936), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3833) );
  OAI21_X1 U3998 ( .B1(n7432), .B2(n7674), .A(n7229), .ZN(n5101) );
  AND2_X1 U3999 ( .A1(n4069), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5545)
         );
  INV_X1 U4000 ( .A(n5084), .ZN(n5543) );
  INV_X1 U4001 ( .A(n3675), .ZN(n7430) );
  CLKBUF_X1 U4002 ( .A(n5011), .Z(n7618) );
  NAND2_X1 U4003 ( .A1(REIP_REG_20__SCAN_IN), .A2(n7598), .ZN(n6490) );
  NOR2_X1 U4004 ( .A1(n4671), .A2(n6307), .ZN(n4688) );
  NAND2_X1 U4005 ( .A1(n6143), .A2(REIP_REG_4__SCAN_IN), .ZN(n5776) );
  INV_X1 U4006 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U4007 ( .A1(n6463), .A2(n3720), .ZN(n6451) );
  AOI21_X1 U4008 ( .B1(n5852), .B2(n5191), .A(n4349), .ZN(n5204) );
  AOI22_X1 U4009 ( .A1(n6415), .A2(n5013), .B1(n4942), .B2(n4941), .ZN(n5052)
         );
  OR2_X1 U4010 ( .A1(n6958), .A2(n4967), .ZN(n4925) );
  AOI21_X1 U4011 ( .B1(n6382), .B2(n5013), .A(n4993), .ZN(n5069) );
  OR2_X1 U4012 ( .A1(n4946), .A2(n4945), .ZN(n5000) );
  NAND2_X1 U4013 ( .A1(n4902), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4943)
         );
  NOR2_X1 U4014 ( .A1(n4857), .A2(n4856), .ZN(n4858) );
  OR2_X1 U4015 ( .A1(n6976), .A2(n4967), .ZN(n4880) );
  AND2_X1 U4016 ( .A1(n4837), .A2(n3691), .ZN(n3789) );
  OR2_X1 U4017 ( .A1(n7605), .A2(n4967), .ZN(n4792) );
  OR2_X1 U4018 ( .A1(n4741), .A2(n7034), .ZN(n4742) );
  INV_X1 U4019 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4754) );
  NOR2_X1 U4020 ( .A1(n4742), .A2(n4754), .ZN(n4775) );
  NAND2_X1 U4021 ( .A1(n4706), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4741)
         );
  NAND2_X1 U4022 ( .A1(n4688), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4705)
         );
  INV_X1 U4023 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U4024 ( .A1(n4666), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4671)
         );
  NOR2_X1 U4025 ( .A1(n4651), .A2(n7555), .ZN(n4666) );
  NAND2_X1 U4026 ( .A1(n3785), .A2(n3784), .ZN(n3783) );
  INV_X1 U4027 ( .A(n6241), .ZN(n3784) );
  NAND2_X1 U4028 ( .A1(n4623), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4651)
         );
  NOR2_X1 U4029 ( .A1(n4619), .A2(n6189), .ZN(n4623) );
  INV_X1 U4030 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U4031 ( .A1(n4578), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4595)
         );
  INV_X1 U4032 ( .A(n4562), .ZN(n4578) );
  NOR2_X1 U4033 ( .A1(n4555), .A2(n5932), .ZN(n4556) );
  NOR2_X1 U4034 ( .A1(n4534), .A2(n6147), .ZN(n4544) );
  NAND2_X1 U4035 ( .A1(n4531), .A2(n4530), .ZN(n5195) );
  NAND3_X1 U4036 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A3(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n4534) );
  INV_X1 U4037 ( .A(n5191), .ZN(n5030) );
  NAND2_X1 U4038 ( .A1(n6404), .A2(n3933), .ZN(n5028) );
  OR2_X1 U4039 ( .A1(n6406), .A2(n6407), .ZN(n6404) );
  NOR2_X1 U4040 ( .A1(n3723), .A2(n3722), .ZN(n6428) );
  INV_X1 U4041 ( .A(n6426), .ZN(n3722) );
  NAND2_X1 U4042 ( .A1(n6463), .A2(n6465), .ZN(n6464) );
  AND2_X1 U4043 ( .A1(n3716), .A2(n3715), .ZN(n3714) );
  INV_X1 U4044 ( .A(n6488), .ZN(n3715) );
  NAND2_X1 U4045 ( .A1(n7161), .A2(n3716), .ZN(n7145) );
  NOR2_X1 U4046 ( .A1(n7163), .A2(n7162), .ZN(n7161) );
  OR2_X1 U4047 ( .A1(n6506), .A2(n6499), .ZN(n7163) );
  OR2_X1 U4048 ( .A1(n6508), .A2(n6509), .ZN(n6506) );
  NOR2_X1 U4049 ( .A1(n6278), .A2(n3710), .ZN(n6355) );
  OR2_X1 U4050 ( .A1(n3712), .A2(n6341), .ZN(n3710) );
  OR2_X1 U4051 ( .A1(n7030), .A2(n6318), .ZN(n4226) );
  NAND2_X1 U4052 ( .A1(n3711), .A2(n4392), .ZN(n6308) );
  INV_X1 U4053 ( .A(n6278), .ZN(n3711) );
  NOR2_X1 U4054 ( .A1(n6278), .A2(n3712), .ZN(n6339) );
  AND2_X1 U4055 ( .A1(n4391), .A2(n4390), .ZN(n6277) );
  AOI21_X1 U4056 ( .B1(n3757), .B2(n6265), .A(n3687), .ZN(n3756) );
  OR2_X1 U4057 ( .A1(n7462), .A2(n4489), .ZN(n6322) );
  AND2_X1 U4058 ( .A1(n4385), .A2(n4384), .ZN(n6197) );
  INV_X1 U4059 ( .A(n6047), .ZN(n4378) );
  NAND2_X1 U4060 ( .A1(n4362), .A2(n4361), .ZN(n5363) );
  INV_X1 U4061 ( .A(n5212), .ZN(n4362) );
  NAND2_X1 U4062 ( .A1(n5205), .A2(n3708), .ZN(n5212) );
  NOR2_X1 U4063 ( .A1(n3709), .A2(n5197), .ZN(n3708) );
  INV_X1 U4064 ( .A(n6366), .ZN(n3709) );
  NAND2_X1 U4065 ( .A1(n5205), .A2(n6366), .ZN(n6368) );
  AOI21_X1 U4066 ( .B1(n5413), .B2(n4294), .A(n4097), .ZN(n7383) );
  AND2_X1 U4067 ( .A1(n4474), .A2(n4473), .ZN(n5861) );
  INV_X1 U4068 ( .A(n5130), .ZN(n4453) );
  OR2_X1 U4069 ( .A1(n4324), .A2(n7430), .ZN(n5164) );
  XNOR2_X1 U4070 ( .A(n4065), .B(n4066), .ZN(n5088) );
  NAND2_X1 U4071 ( .A1(n4064), .A2(n4067), .ZN(n4102) );
  OR2_X1 U4072 ( .A1(n4068), .A2(n3731), .ZN(n4072) );
  OR2_X1 U4073 ( .A1(n4068), .A2(n3804), .ZN(n4110) );
  NOR2_X1 U4074 ( .A1(n5334), .A2(n5084), .ZN(n5311) );
  OR2_X1 U4075 ( .A1(n5085), .A2(n5297), .ZN(n5334) );
  OR2_X1 U4076 ( .A1(n5626), .A2(n5625), .ZN(n5427) );
  NOR2_X1 U4077 ( .A1(n5544), .A2(n5084), .ZN(n5505) );
  AND2_X1 U4078 ( .A1(n3667), .A2(n5871), .ZN(n5800) );
  AND3_X1 U4079 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n7691), .A3(n5101), .ZN(
        n5260) );
  INV_X1 U4080 ( .A(n5871), .ZN(n5679) );
  OR2_X1 U4081 ( .A1(n5544), .A2(n5543), .ZN(n5553) );
  OR2_X1 U4082 ( .A1(n4284), .A2(n4283), .ZN(n4287) );
  AND2_X1 U4083 ( .A1(n4288), .A2(n4318), .ZN(n4289) );
  NAND2_X1 U4084 ( .A1(n3732), .A2(n4281), .ZN(n4291) );
  NAND2_X1 U4085 ( .A1(n3734), .A2(n3733), .ZN(n3732) );
  CLKBUF_X1 U4086 ( .A(n4543), .Z(n5013) );
  NAND2_X1 U4087 ( .A1(n3646), .A2(n3750), .ZN(n5108) );
  NAND2_X1 U4088 ( .A1(n7406), .A2(n7688), .ZN(n5107) );
  NAND2_X1 U4089 ( .A1(n6487), .A2(n5022), .ZN(n6482) );
  INV_X1 U4090 ( .A(n6487), .ZN(n7603) );
  NAND2_X1 U4091 ( .A1(n6512), .A2(REIP_REG_19__SCAN_IN), .ZN(n7586) );
  NOR2_X1 U4092 ( .A1(n7567), .A2(n3751), .ZN(n6512) );
  INV_X1 U4093 ( .A(n3752), .ZN(n3751) );
  OAI21_X1 U4094 ( .B1(n6356), .B2(n7313), .A(n6230), .ZN(n3752) );
  NOR2_X1 U4095 ( .A1(n5039), .A2(n6142), .ZN(n7567) );
  INV_X1 U4096 ( .A(n7520), .ZN(n7593) );
  INV_X1 U4097 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n7549) );
  INV_X1 U4098 ( .A(n7554), .ZN(n7582) );
  INV_X1 U4099 ( .A(n6143), .ZN(n6149) );
  INV_X1 U4100 ( .A(n7606), .ZN(n7579) );
  AND2_X1 U4101 ( .A1(n5785), .A2(n5784), .ZN(n7606) );
  NAND2_X1 U4102 ( .A1(n6275), .A2(n5853), .ZN(n6230) );
  INV_X1 U4103 ( .A(n6543), .ZN(n7374) );
  AND2_X1 U4104 ( .A1(n5190), .A2(n7688), .ZN(n7376) );
  INV_X1 U4105 ( .A(n7369), .ZN(n7372) );
  INV_X1 U4106 ( .A(n7374), .ZN(n6539) );
  OAI21_X1 U4107 ( .B1(n5050), .B2(n5052), .A(n5051), .ZN(n6550) );
  NOR2_X1 U4108 ( .A1(n7735), .A2(n5225), .ZN(n6569) );
  NAND2_X1 U4109 ( .A1(n5375), .A2(n5076), .ZN(n6392) );
  OAI21_X1 U4110 ( .B1(n5128), .B2(n5075), .A(n7688), .ZN(n5076) );
  INV_X1 U4111 ( .A(n6569), .ZN(n6335) );
  OR2_X1 U4112 ( .A1(n5167), .A2(n5166), .ZN(n7286) );
  CLKBUF_X1 U4113 ( .A(n5409), .Z(n5402) );
  INV_X1 U4114 ( .A(n5375), .ZN(n5410) );
  INV_X1 U4115 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n7034) );
  NAND2_X1 U4116 ( .A1(n6214), .A2(n6215), .ZN(n3759) );
  OR2_X1 U4117 ( .A1(n5167), .A2(n7654), .ZN(n7626) );
  INV_X2 U4118 ( .A(n7035), .ZN(n7396) );
  INV_X1 U4119 ( .A(n7626), .ZN(n7402) );
  NAND2_X1 U4120 ( .A1(n4498), .A2(n4497), .ZN(n4499) );
  XNOR2_X1 U4121 ( .A(n6944), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3780)
         );
  XNOR2_X1 U4122 ( .A(n7030), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3779)
         );
  OR3_X1 U4123 ( .A1(n7156), .A2(n7098), .A3(n7099), .ZN(n7087) );
  NAND2_X1 U4124 ( .A1(n6955), .A2(n6954), .ZN(n6956) );
  NAND2_X1 U4125 ( .A1(n6953), .A2(n7030), .ZN(n6954) );
  OR2_X1 U4126 ( .A1(n7130), .A2(n4486), .ZN(n7115) );
  NAND2_X1 U4127 ( .A1(n6249), .A2(n6322), .ZN(n7219) );
  NOR2_X1 U4128 ( .A1(n6175), .A2(n5220), .ZN(n7471) );
  INV_X1 U4129 ( .A(n7196), .ZN(n7176) );
  AND2_X1 U4130 ( .A1(n4472), .A2(n7639), .ZN(n7492) );
  INV_X1 U4131 ( .A(n5552), .ZN(n5637) );
  CLKBUF_X1 U4132 ( .A(n5088), .Z(n5089) );
  CLKBUF_X1 U4133 ( .A(n4502), .Z(n5084) );
  INV_X1 U4134 ( .A(n5085), .ZN(n5413) );
  CLKBUF_X1 U4135 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n7231) );
  NAND2_X1 U4136 ( .A1(n5082), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7229) );
  INV_X1 U4137 ( .A(n7693), .ZN(n5082) );
  OAI21_X1 U4138 ( .B1(n5639), .B2(n5636), .A(n5675), .ZN(n5665) );
  AND2_X1 U4139 ( .A1(n5099), .A2(n5098), .ZN(n5265) );
  NAND2_X1 U4140 ( .A1(n5100), .A2(n5637), .ZN(n5839) );
  NOR2_X1 U4141 ( .A1(n5226), .A2(n5591), .ZN(n6130) );
  INV_X1 U4142 ( .A(n6025), .ZN(n6132) );
  NOR2_X1 U4143 ( .A1(n5374), .A2(n5591), .ZN(n6098) );
  INV_X1 U4144 ( .A(n6020), .ZN(n6099) );
  NOR2_X1 U4145 ( .A1(n5496), .A2(n5591), .ZN(n6082) );
  NOR2_X1 U4146 ( .A1(n5493), .A2(n5591), .ZN(n6121) );
  INV_X1 U4147 ( .A(n6010), .ZN(n6122) );
  NOR2_X1 U4148 ( .A1(n5239), .A2(n5591), .ZN(n6090) );
  INV_X1 U4149 ( .A(n6005), .ZN(n6091) );
  NOR2_X1 U4150 ( .A1(n5491), .A2(n5591), .ZN(n6113) );
  INV_X1 U4151 ( .A(n6038), .ZN(n6114) );
  NOR2_X1 U4152 ( .A1(n5494), .A2(n5591), .ZN(n6106) );
  INV_X1 U4153 ( .A(n6000), .ZN(n6107) );
  NOR2_X1 U4154 ( .A1(n5525), .A2(n5591), .ZN(n6074) );
  INV_X1 U4155 ( .A(n6030), .ZN(n6075) );
  OAI21_X1 U4156 ( .B1(n5721), .B2(n5720), .A(n5719), .ZN(n5760) );
  INV_X1 U4157 ( .A(n6130), .ZN(n6024) );
  INV_X1 U4158 ( .A(n6082), .ZN(n6014) );
  INV_X1 U4159 ( .A(n6121), .ZN(n6009) );
  INV_X1 U4160 ( .A(n6090), .ZN(n6004) );
  INV_X1 U4161 ( .A(n6113), .ZN(n6035) );
  NOR2_X1 U4162 ( .A1(n5553), .A2(n5552), .ZN(n6067) );
  INV_X1 U4163 ( .A(n6074), .ZN(n6029) );
  OR3_X1 U4164 ( .A1(n7663), .A2(n7662), .A3(n7661), .ZN(n7689) );
  INV_X1 U4165 ( .A(n7688), .ZN(n7671) );
  INV_X1 U4166 ( .A(n7673), .ZN(n7690) );
  INV_X1 U4167 ( .A(READY_N), .ZN(n7709) );
  NAND2_X1 U4168 ( .A1(n3730), .A2(n3685), .ZN(U2796) );
  NAND2_X1 U4169 ( .A1(n7073), .A2(n7610), .ZN(n3730) );
  AND2_X1 U4170 ( .A1(n5044), .A2(n3729), .ZN(n3728) );
  NAND2_X1 U4171 ( .A1(n6388), .A2(REIP_REG_30__SCAN_IN), .ZN(n3749) );
  AND2_X1 U4172 ( .A1(n6387), .A2(n6386), .ZN(n6389) );
  NOR2_X1 U4173 ( .A1(n3748), .A2(n3747), .ZN(n3746) );
  INV_X1 U4174 ( .A(n5066), .ZN(n5067) );
  AND2_X2 U4175 ( .A1(n3814), .A2(n5274), .ZN(n4006) );
  AND2_X1 U4176 ( .A1(n3814), .A2(n3819), .ZN(n3998) );
  NAND2_X1 U4177 ( .A1(n5249), .A2(n3638), .ZN(n4301) );
  NAND2_X1 U4178 ( .A1(n3782), .A2(n3785), .ZN(n6195) );
  AND2_X1 U4179 ( .A1(n6532), .A2(n3691), .ZN(n6473) );
  AND4_X1 U4180 ( .A1(n3993), .A2(n3985), .A3(n3992), .A4(n3991), .ZN(n3679)
         );
  AND2_X1 U4181 ( .A1(n5022), .A2(n3692), .ZN(n3680) );
  INV_X1 U4182 ( .A(n5073), .ZN(n4503) );
  AND2_X1 U4183 ( .A1(n3680), .A2(n3693), .ZN(n3681) );
  INV_X1 U4184 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3809) );
  AND2_X1 U4185 ( .A1(n3690), .A2(n5052), .ZN(n3682) );
  NAND2_X1 U4186 ( .A1(n3933), .A2(n3932), .ZN(n4456) );
  NAND2_X1 U4187 ( .A1(n6532), .A2(n6535), .ZN(n6534) );
  NAND2_X1 U4188 ( .A1(n6532), .A2(n3790), .ZN(n3683) );
  AND2_X1 U4189 ( .A1(n6487), .A2(n3680), .ZN(n3684) );
  OR2_X1 U4190 ( .A1(n5020), .A2(n6142), .ZN(n6487) );
  OAI21_X1 U4191 ( .B1(n4295), .B2(n3959), .A(n3958), .ZN(n3978) );
  AND3_X1 U4192 ( .A1(n5043), .A2(n5045), .A3(n3728), .ZN(n3685) );
  INV_X1 U4193 ( .A(n3954), .ZN(n3935) );
  AND2_X1 U4194 ( .A1(n3934), .A2(n4456), .ZN(n3985) );
  NAND2_X1 U4195 ( .A1(n6971), .A2(n4236), .ZN(n6962) );
  AND2_X1 U4196 ( .A1(n4045), .A2(n7472), .ZN(n3686) );
  NAND2_X1 U4197 ( .A1(n4072), .A2(n4071), .ZN(n4103) );
  NOR2_X1 U4198 ( .A1(n7030), .A2(n7218), .ZN(n3687) );
  AND2_X1 U4199 ( .A1(n4294), .A2(n4275), .ZN(n4280) );
  INV_X1 U4200 ( .A(n4280), .ZN(n3745) );
  NOR2_X1 U4201 ( .A1(n5710), .A2(n6045), .ZN(n6044) );
  NAND2_X1 U4202 ( .A1(n7161), .A2(n6537), .ZN(n6536) );
  AND2_X1 U4203 ( .A1(n7030), .A2(n4470), .ZN(n3689) );
  NAND2_X1 U4204 ( .A1(n3753), .A2(n3756), .ZN(n6246) );
  NAND2_X1 U4205 ( .A1(n3759), .A2(n4220), .ZN(n6264) );
  NAND2_X1 U4206 ( .A1(n4503), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4686) );
  INV_X1 U4207 ( .A(n4686), .ZN(n4665) );
  AND2_X1 U4208 ( .A1(n6424), .A2(n4899), .ZN(n3690) );
  AND2_X1 U4209 ( .A1(n4809), .A2(n3790), .ZN(n3691) );
  NAND2_X1 U4210 ( .A1(n4223), .A2(n4222), .ZN(n6292) );
  OR2_X1 U4211 ( .A1(n6275), .A2(n5024), .ZN(n3692) );
  INV_X1 U4212 ( .A(n5710), .ZN(n3782) );
  NAND2_X1 U4213 ( .A1(n7510), .A2(n5025), .ZN(n3693) );
  INV_X1 U4214 ( .A(n3771), .ZN(n3770) );
  NOR2_X1 U4215 ( .A1(n7030), .A2(n4232), .ZN(n3771) );
  AND2_X1 U4216 ( .A1(n6477), .A2(n6479), .ZN(n6463) );
  AND2_X1 U4217 ( .A1(n7161), .A2(n3714), .ZN(n6477) );
  AND2_X1 U4218 ( .A1(n3682), .A2(n3792), .ZN(n3694) );
  NOR2_X1 U4219 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4543) );
  AND2_X1 U4220 ( .A1(n5204), .A2(n5203), .ZN(n5205) );
  NAND2_X1 U4221 ( .A1(n4507), .A2(n4506), .ZN(n5179) );
  NAND2_X1 U4222 ( .A1(n4046), .A2(n3686), .ZN(n5215) );
  INV_X1 U4223 ( .A(n7618), .ZN(n3750) );
  AND2_X1 U4224 ( .A1(n4665), .A2(n4650), .ZN(n3695) );
  NOR2_X1 U4225 ( .A1(n3953), .A2(n3968), .ZN(n4333) );
  NAND2_X1 U4226 ( .A1(n3935), .A2(n5073), .ZN(n5184) );
  INV_X2 U4227 ( .A(n7059), .ZN(n7392) );
  INV_X1 U4228 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3781) );
  INV_X1 U4229 ( .A(n7604), .ZN(n7577) );
  OR2_X1 U4230 ( .A1(n7501), .A2(n7669), .ZN(n5849) );
  AND2_X2 U4231 ( .A1(n3820), .A2(n5282), .ZN(n3927) );
  NAND2_X1 U4232 ( .A1(n3696), .A2(n4218), .ZN(n6169) );
  OAI21_X2 U4233 ( .B1(n5770), .B2(n3762), .A(n3697), .ZN(n3696) );
  INV_X1 U4234 ( .A(n3761), .ZN(n3697) );
  NAND2_X1 U4235 ( .A1(n4195), .A2(n4194), .ZN(n5770) );
  OR2_X1 U4236 ( .A1(n7024), .A2(n7023), .ZN(n3701) );
  NAND2_X1 U4237 ( .A1(n3698), .A2(n3800), .ZN(n7010) );
  OR2_X1 U4238 ( .A1(n7024), .A2(n3699), .ZN(n3698) );
  OR2_X1 U4239 ( .A1(n3700), .A2(n7023), .ZN(n3699) );
  INV_X1 U4240 ( .A(n3701), .ZN(n6980) );
  NOR2_X2 U4241 ( .A1(n7010), .A2(n7009), .ZN(n7152) );
  NOR2_X1 U4242 ( .A1(n7030), .A2(n7018), .ZN(n3700) );
  NAND2_X2 U4243 ( .A1(n3796), .A2(n3798), .ZN(n5249) );
  NAND4_X1 U4244 ( .A1(n3960), .A2(n3948), .A3(n3985), .A4(n3703), .ZN(n3702)
         );
  AND2_X2 U4245 ( .A1(n4066), .A2(n3704), .ZN(n4509) );
  NAND2_X1 U4246 ( .A1(n4089), .A2(n4090), .ZN(n3706) );
  INV_X1 U4247 ( .A(n3723), .ZN(n6440) );
  NAND3_X1 U4248 ( .A1(n3739), .A2(n3736), .A3(n3735), .ZN(n3734) );
  NAND3_X1 U4249 ( .A1(n3749), .A2(n6389), .A3(n3746), .ZN(U2797) );
  NOR3_X2 U4250 ( .A1(n6411), .A2(n7338), .A3(REIP_REG_30__SCAN_IN), .ZN(n3747) );
  NOR3_X2 U4251 ( .A1(n6274), .A2(n7308), .A3(n6305), .ZN(n5039) );
  NAND2_X1 U4252 ( .A1(n6214), .A2(n3754), .ZN(n3753) );
  NAND2_X1 U4253 ( .A1(n3760), .A2(n4207), .ZN(n6050) );
  NAND2_X1 U4254 ( .A1(n5770), .A2(n5771), .ZN(n3760) );
  OAI21_X1 U4255 ( .B1(n5771), .B2(n3762), .A(n6051), .ZN(n3761) );
  INV_X1 U4256 ( .A(n4207), .ZN(n3762) );
  INV_X1 U4257 ( .A(n5233), .ZN(n4145) );
  NAND2_X1 U4258 ( .A1(n3764), .A2(n3763), .ZN(n5233) );
  NAND2_X1 U4259 ( .A1(n7390), .A2(n4468), .ZN(n3763) );
  NAND2_X1 U4260 ( .A1(n4046), .A2(n4045), .ZN(n4056) );
  NAND2_X1 U4261 ( .A1(n5215), .A2(n5218), .ZN(n3765) );
  INV_X1 U4262 ( .A(n3766), .ZN(n6970) );
  INV_X1 U4263 ( .A(n3775), .ZN(n3774) );
  OAI211_X1 U4264 ( .C1(n5011), .C2(n3972), .A(n4335), .B(n4330), .ZN(n3776)
         );
  NAND2_X1 U4265 ( .A1(n4500), .A2(n3779), .ZN(n3778) );
  NOR2_X1 U4266 ( .A1(n5710), .A2(n3787), .ZN(n6161) );
  NAND2_X1 U4267 ( .A1(n6437), .A2(n3682), .ZN(n5051) );
  AND2_X1 U4268 ( .A1(n6437), .A2(n3690), .ZN(n5050) );
  AND2_X1 U4269 ( .A1(n6437), .A2(n4899), .ZN(n6423) );
  AND2_X2 U4270 ( .A1(n6437), .A2(n3694), .ZN(n6402) );
  INV_X1 U4271 ( .A(n7382), .ZN(n4099) );
  NAND2_X1 U4273 ( .A1(n6240), .A2(n3695), .ZN(n4653) );
  INV_X1 U4274 ( .A(n4148), .ZN(n4150) );
  NAND2_X1 U4275 ( .A1(n4148), .A2(n4125), .ZN(n5083) );
  XNOR2_X1 U4276 ( .A(n4148), .B(n4149), .ZN(n4523) );
  NAND2_X1 U4277 ( .A1(n4197), .A2(n4196), .ZN(n4208) );
  INV_X1 U4278 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n7555) );
  OR3_X1 U4279 ( .A1(REIP_REG_22__SCAN_IN), .A2(n7321), .A3(n6490), .ZN(n3793)
         );
  NOR2_X1 U4280 ( .A1(n3668), .A2(n5089), .ZN(n3794) );
  NAND2_X1 U4281 ( .A1(n3986), .A2(n3949), .ZN(n3795) );
  AND4_X1 U4282 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3796)
         );
  XOR2_X1 U4283 ( .A(n7030), .B(n5062), .Z(n3797) );
  AND4_X1 U4284 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(n3798)
         );
  AND2_X1 U4285 ( .A1(n7026), .A2(n7025), .ZN(n3799) );
  NAND2_X1 U4286 ( .A1(n7031), .A2(n4242), .ZN(n6944) );
  INV_X1 U4287 ( .A(n6944), .ZN(n4243) );
  AOI21_X1 U4288 ( .B1(n4548), .B2(n4665), .A(n4547), .ZN(n5209) );
  OR2_X1 U4289 ( .A1(n7031), .A2(n7154), .ZN(n3800) );
  AND3_X1 U4290 ( .A1(n3939), .A2(n3938), .A3(n3937), .ZN(n3801) );
  INV_X1 U4291 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5417) );
  AND2_X1 U4292 ( .A1(n7736), .A2(DATAI_30_), .ZN(n3802) );
  NOR2_X1 U4293 ( .A1(n3952), .A2(n7669), .ZN(n4542) );
  AND2_X1 U4294 ( .A1(n4495), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3803)
         );
  OR2_X1 U4295 ( .A1(n4004), .A2(n4003), .ZN(n4042) );
  OR2_X1 U4296 ( .A1(n4849), .A2(n4848), .ZN(n4862) );
  OR2_X1 U4297 ( .A1(n4160), .A2(n4159), .ZN(n4200) );
  AOI21_X1 U4298 ( .B1(n4006), .B2(INSTQUEUE_REG_5__6__SCAN_IN), .A(n3833), 
        .ZN(n3837) );
  NOR2_X1 U4299 ( .A1(n3981), .A2(n3954), .ZN(n3962) );
  INV_X1 U4300 ( .A(n6439), .ZN(n4899) );
  INV_X1 U4301 ( .A(n6486), .ZN(n4809) );
  OR2_X1 U4302 ( .A1(n7030), .A2(n7207), .ZN(n4229) );
  OR2_X1 U4303 ( .A1(n4184), .A2(n4183), .ZN(n4199) );
  OR2_X1 U4304 ( .A1(n4121), .A2(n4120), .ZN(n4127) );
  NAND2_X1 U4305 ( .A1(n3669), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U4306 ( .A1(n3669), .A2(n3988), .ZN(n4331) );
  INV_X1 U4307 ( .A(n7025), .ZN(n4759) );
  AND2_X1 U4308 ( .A1(n4901), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4902)
         );
  OR2_X1 U4309 ( .A1(n4810), .A2(n7001), .ZN(n4811) );
  INV_X1 U4310 ( .A(n4991), .ZN(n4964) );
  INV_X1 U4311 ( .A(n4542), .ZN(n4721) );
  INV_X1 U4312 ( .A(n6048), .ZN(n4377) );
  AND2_X1 U4313 ( .A1(n4284), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4250)
         );
  INV_X1 U4314 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6307) );
  INV_X1 U4315 ( .A(n5849), .ZN(n5851) );
  INV_X1 U4316 ( .A(n5213), .ZN(n4361) );
  OR2_X1 U4317 ( .A1(n4811), .A2(n6476), .ZN(n4857) );
  NOR2_X1 U4318 ( .A1(n4705), .A2(n6357), .ZN(n4706) );
  INV_X1 U4319 ( .A(n4850), .ZN(n4994) );
  NAND2_X1 U4320 ( .A1(n4556), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4562)
         );
  INV_X1 U4321 ( .A(n6293), .ZN(n4224) );
  INV_X1 U4322 ( .A(n4294), .ZN(n4210) );
  INV_X1 U4323 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5630) );
  AND2_X1 U4324 ( .A1(n5464), .A2(n6061), .ZN(n5944) );
  INV_X1 U4325 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7649) );
  OR2_X1 U4326 ( .A1(n5085), .A2(n5296), .ZN(n5544) );
  AND2_X1 U4327 ( .A1(n7623), .A2(n3971), .ZN(n7406) );
  NAND2_X1 U4328 ( .A1(n4287), .A2(n4286), .ZN(n4318) );
  INV_X1 U4329 ( .A(n6275), .ZN(n7510) );
  OR2_X1 U4330 ( .A1(n4595), .A2(n7549), .ZN(n4619) );
  INV_X1 U4331 ( .A(n6230), .ZN(n6142) );
  AND2_X1 U4332 ( .A1(n4925), .A2(n4924), .ZN(n6424) );
  XNOR2_X1 U4333 ( .A(n4208), .B(n4198), .ZN(n4561) );
  INV_X1 U4334 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U4335 ( .A1(n4898), .A2(n4897), .ZN(n6439) );
  NAND2_X1 U4336 ( .A1(n4776), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4810)
         );
  INV_X1 U4337 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5932) );
  OAI22_X1 U4338 ( .A1(n6953), .A2(n5048), .B1(n7031), .B2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5049) );
  INV_X1 U4339 ( .A(n6067), .ZN(n6134) );
  INV_X1 U4340 ( .A(n5591), .ZN(n5675) );
  INV_X1 U4341 ( .A(n5875), .ZN(n6063) );
  INV_X1 U4342 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5629) );
  AOI21_X1 U4343 ( .B1(n5629), .B2(STATE2_REG_3__SCAN_IN), .A(n5591), .ZN(
        n5551) );
  NOR2_X1 U4344 ( .A1(n7425), .A2(n5016), .ZN(n7501) );
  INV_X1 U4345 ( .A(n7595), .ZN(n7611) );
  XNOR2_X1 U4346 ( .A(n5002), .B(n5037), .ZN(n5785) );
  INV_X1 U4347 ( .A(n7601), .ZN(n7608) );
  NOR2_X2 U4348 ( .A1(n7735), .A2(n3968), .ZN(n7736) );
  INV_X1 U4349 ( .A(n6392), .ZN(n7735) );
  NOR2_X1 U4350 ( .A1(n5409), .A2(n5160), .ZN(n5366) );
  NAND2_X1 U4351 ( .A1(n5160), .A2(n3965), .ZN(n5375) );
  INV_X1 U4352 ( .A(n6497), .ZN(n7026) );
  NAND2_X1 U4353 ( .A1(n4544), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4555)
         );
  NAND2_X1 U4354 ( .A1(n7626), .A2(n5004), .ZN(n7035) );
  OAI21_X1 U4355 ( .B1(n6521), .B2(n7479), .A(n5065), .ZN(n5066) );
  INV_X1 U4356 ( .A(n7477), .ZN(n7460) );
  AND2_X1 U4357 ( .A1(n5111), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5218)
         );
  INV_X1 U4358 ( .A(n7212), .ZN(n7488) );
  INV_X1 U4359 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7422) );
  NOR2_X1 U4360 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5154) );
  OAI211_X1 U4361 ( .C1(n5995), .C2(n5996), .A(n5994), .B(n6063), .ZN(n6034)
         );
  INV_X1 U4362 ( .A(n5948), .ZN(n5985) );
  INV_X1 U4363 ( .A(n5709), .ZN(n5347) );
  OAI211_X1 U4364 ( .C1(n5678), .C2(n5034), .A(n5677), .B(n5994), .ZN(n5702)
         );
  OAI21_X1 U4365 ( .B1(n5595), .B2(n5594), .A(n5593), .ZN(n5617) );
  INV_X1 U4366 ( .A(n5585), .ZN(n5621) );
  OR3_X1 U4367 ( .A1(n5797), .A2(n5946), .A3(n5796), .ZN(n5847) );
  INV_X1 U4368 ( .A(n6015), .ZN(n6083) );
  AND2_X1 U4369 ( .A1(n5505), .A2(n5552), .ZN(n5840) );
  INV_X1 U4370 ( .A(n5722), .ZN(n5764) );
  AND2_X1 U4371 ( .A1(n4321), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7688) );
  INV_X1 U4372 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7420) );
  OR2_X1 U4373 ( .A1(n7501), .A2(n5034), .ZN(n7601) );
  OR2_X1 U4374 ( .A1(n5785), .A2(n5783), .ZN(n7595) );
  NAND2_X1 U4375 ( .A1(n7376), .A2(n3952), .ZN(n6543) );
  INV_X1 U4376 ( .A(n6987), .ZN(n6562) );
  INV_X1 U4377 ( .A(n7401), .ZN(n7523) );
  INV_X1 U4378 ( .A(n5008), .ZN(n5009) );
  NAND2_X1 U4379 ( .A1(n5871), .A2(n4999), .ZN(n7059) );
  AND2_X1 U4380 ( .A1(n4493), .A2(n4492), .ZN(n4494) );
  NAND2_X1 U4381 ( .A1(n4472), .A2(n4338), .ZN(n7212) );
  AND2_X1 U4382 ( .A1(n5295), .A2(n5591), .ZN(n7254) );
  INV_X1 U4383 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7632) );
  AOI21_X1 U4384 ( .B1(n6066), .B2(n6065), .A(n6064), .ZN(n6141) );
  NAND2_X1 U4385 ( .A1(n5628), .A2(n5637), .ZN(n6043) );
  NAND3_X1 U4386 ( .A1(n5626), .A2(n5463), .A3(n5637), .ZN(n5983) );
  NAND2_X1 U4387 ( .A1(n5311), .A2(n5552), .ZN(n5948) );
  NAND2_X1 U4388 ( .A1(n5311), .A2(n5637), .ZN(n5709) );
  NAND3_X1 U4389 ( .A1(n5326), .A2(n5637), .A3(n5084), .ZN(n5912) );
  NOR2_X1 U4390 ( .A1(n5878), .A2(n5877), .ZN(n5917) );
  NAND2_X1 U4391 ( .A1(n5419), .A2(n5637), .ZN(n5619) );
  AOI22_X1 U4392 ( .A1(n5589), .A2(n5595), .B1(n6069), .B2(n5723), .ZN(n5624)
         );
  INV_X1 U4393 ( .A(n6098), .ZN(n6019) );
  INV_X1 U4394 ( .A(n6106), .ZN(n5999) );
  OR2_X1 U4395 ( .A1(n5497), .A2(n5552), .ZN(n5722) );
  NAND2_X1 U4396 ( .A1(n5548), .A2(n5552), .ZN(n5769) );
  INV_X1 U4397 ( .A(n7716), .ZN(n7706) );
  NAND2_X1 U4398 ( .A1(n3944), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3808) );
  INV_X1 U4399 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U4400 ( .A1(n4006), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3807) );
  NAND2_X1 U4401 ( .A1(n3642), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3806) );
  AND2_X2 U4402 ( .A1(n5144), .A2(n5282), .ZN(n3936) );
  NAND2_X1 U4403 ( .A1(n3936), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3805)
         );
  NAND2_X1 U4404 ( .A1(n4970), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3813)
         );
  NAND2_X1 U4405 ( .A1(n3643), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3812) );
  NAND2_X1 U4406 ( .A1(n4115), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3811) );
  NAND2_X1 U4407 ( .A1(n3927), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3810)
         );
  AND2_X2 U4408 ( .A1(n5274), .A2(n5133), .ZN(n4676) );
  NAND2_X1 U4409 ( .A1(n4676), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4410 ( .A1(n3665), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3817)
         );
  NAND2_X1 U4411 ( .A1(n3676), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3816)
         );
  NAND2_X1 U4412 ( .A1(n4909), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3815) );
  NAND2_X1 U4413 ( .A1(n3998), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3824) );
  AND2_X4 U4414 ( .A1(n5271), .A2(n5144), .ZN(n4074) );
  NAND2_X1 U4415 ( .A1(n4074), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3823)
         );
  AND2_X2 U4416 ( .A1(n5133), .A2(n3819), .ZN(n4971) );
  NAND2_X1 U4417 ( .A1(n4971), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3822) );
  NAND2_X1 U4418 ( .A1(n4025), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3821) );
  NAND4_X4 U4419 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3954)
         );
  AOI22_X1 U4420 ( .A1(n4970), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3927), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4421 ( .A1(n3998), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4422 ( .A1(n4676), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4423 ( .A1(n3678), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4424 ( .A1(n3665), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4425 ( .A1(n4971), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4426 ( .A1(n3944), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3642), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U4427 ( .A1(n3643), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3843) );
  NAND2_X1 U4428 ( .A1(n4970), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3842)
         );
  NAND2_X1 U4429 ( .A1(n4115), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U4430 ( .A1(n3927), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3840)
         );
  NAND2_X1 U4431 ( .A1(n3944), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3847) );
  NAND2_X1 U4432 ( .A1(n4006), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3846) );
  NAND2_X1 U4433 ( .A1(n3642), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3845) );
  NAND2_X1 U4434 ( .A1(n3936), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3844)
         );
  NAND2_X1 U4435 ( .A1(n3998), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3851) );
  NAND2_X1 U4436 ( .A1(n3672), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3850)
         );
  NAND2_X1 U4437 ( .A1(n4971), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3849) );
  NAND2_X1 U4438 ( .A1(n3670), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3848) );
  NAND2_X1 U4439 ( .A1(n3639), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3855)
         );
  NAND2_X1 U4440 ( .A1(n4676), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3854) );
  NAND2_X1 U4441 ( .A1(n3677), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3853)
         );
  NAND2_X1 U4442 ( .A1(n3664), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3852) );
  NAND2_X1 U4443 ( .A1(n3998), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U4444 ( .A1(n3678), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3862) );
  NAND2_X1 U4445 ( .A1(n4115), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3861) );
  NAND2_X1 U4446 ( .A1(n3640), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U4447 ( .A1(n3672), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3867)
         );
  NAND2_X1 U4448 ( .A1(n3639), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3866)
         );
  NAND2_X1 U4449 ( .A1(n4025), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3865) );
  NAND2_X1 U4450 ( .A1(n3677), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3864)
         );
  NAND2_X1 U4451 ( .A1(n4676), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4452 ( .A1(n4970), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3870)
         );
  NAND2_X1 U4453 ( .A1(n4971), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4454 ( .A1(n4909), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3868) );
  NAND2_X1 U4455 ( .A1(n3944), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U4456 ( .A1(n4006), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3874) );
  NAND2_X1 U4457 ( .A1(n3936), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3873)
         );
  NAND2_X1 U4458 ( .A1(n3927), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3872)
         );
  NAND4_X4 U4459 ( .A1(n3879), .A2(n3878), .A3(n3876), .A4(n3877), .ZN(n3952)
         );
  NAND2_X1 U4460 ( .A1(n5184), .A2(n3880), .ZN(n4297) );
  NAND2_X1 U4461 ( .A1(n3678), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3884) );
  NAND2_X1 U4462 ( .A1(n4970), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3883)
         );
  NAND2_X1 U4463 ( .A1(n4115), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3882) );
  NAND2_X1 U4464 ( .A1(n3927), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3881)
         );
  NAND2_X1 U4465 ( .A1(n4074), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3888)
         );
  NAND2_X1 U4466 ( .A1(n3998), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3887) );
  NAND2_X1 U4467 ( .A1(n4971), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3886) );
  NAND2_X1 U4468 ( .A1(n4025), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3885) );
  NAND2_X1 U4469 ( .A1(n4676), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3892) );
  NAND2_X1 U4470 ( .A1(n3665), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3891)
         );
  NAND2_X1 U4471 ( .A1(n3677), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3890)
         );
  NAND2_X1 U4472 ( .A1(n3663), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3889) );
  NAND2_X1 U4473 ( .A1(n3944), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3896) );
  NAND2_X1 U4474 ( .A1(n4006), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3895) );
  NAND2_X1 U4475 ( .A1(n3641), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3894) );
  NAND2_X1 U4476 ( .A1(n3936), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3893)
         );
  NAND4_X4 U4477 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3965)
         );
  NAND2_X1 U4478 ( .A1(n4006), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3904) );
  NAND2_X1 U4479 ( .A1(n3944), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3903) );
  NAND2_X1 U4480 ( .A1(n3642), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3902) );
  NAND2_X1 U4481 ( .A1(n3936), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3901)
         );
  NAND2_X1 U4482 ( .A1(n4676), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3908) );
  NAND2_X1 U4483 ( .A1(n3665), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3907)
         );
  NAND2_X1 U4484 ( .A1(n3676), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3906)
         );
  NAND2_X1 U4485 ( .A1(n4909), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3905) );
  NAND2_X1 U4486 ( .A1(n3678), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3913) );
  NAND2_X1 U4487 ( .A1(n4970), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3912)
         );
  NAND2_X1 U4488 ( .A1(n4115), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U4489 ( .A1(n3927), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3910)
         );
  NAND2_X1 U4490 ( .A1(n4074), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3917)
         );
  NAND2_X1 U4491 ( .A1(n3998), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3916) );
  NAND2_X1 U4492 ( .A1(n4971), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3915) );
  NAND2_X1 U4493 ( .A1(n4025), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3914) );
  NAND4_X4 U4494 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n4017)
         );
  NAND2_X1 U4495 ( .A1(n4297), .A2(n3987), .ZN(n3934) );
  AOI22_X1 U4496 ( .A1(n4676), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4971), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4497 ( .A1(n3676), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4498 ( .A1(n3643), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4499 ( .A1(n3998), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4500 ( .A1(n3944), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3642), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4501 ( .A1(n4970), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3927), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4502 ( .A1(n4006), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4503 ( .A1(n3639), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3928) );
  INV_X1 U4504 ( .A(n3965), .ZN(n3988) );
  XNOR2_X1 U4505 ( .A(STATE_REG_2__SCAN_IN), .B(STATE_REG_1__SCAN_IN), .ZN(
        n4310) );
  NAND2_X1 U4506 ( .A1(n3988), .A2(n4310), .ZN(n3964) );
  AOI22_X1 U4507 ( .A1(n3678), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4508 ( .A1(n4006), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4509 ( .A1(n4970), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3927), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4510 ( .A1(n3665), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4676), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4511 ( .A1(n3998), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4512 ( .A1(n4971), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4513 ( .A1(n3677), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4514 ( .A1(n3944), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3642), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3946) );
  OAI211_X1 U4515 ( .C1(n3986), .C2(n3949), .A(n3952), .B(n5184), .ZN(n4300)
         );
  INV_X1 U4516 ( .A(n4300), .ZN(n3950) );
  NAND2_X1 U4517 ( .A1(n3950), .A2(n3795), .ZN(n3984) );
  NAND2_X2 U4518 ( .A1(n5073), .A2(n3952), .ZN(n3968) );
  NAND2_X1 U4519 ( .A1(n4333), .A2(n4312), .ZN(n3957) );
  NOR2_X1 U4520 ( .A1(n3968), .A2(n3954), .ZN(n3955) );
  NAND2_X1 U4521 ( .A1(n3955), .A2(n3969), .ZN(n3956) );
  NAND2_X1 U4522 ( .A1(n3957), .A2(n3956), .ZN(n3959) );
  NAND2_X1 U4523 ( .A1(n3978), .A2(n3922), .ZN(n3960) );
  INV_X1 U4524 ( .A(n4297), .ZN(n3961) );
  NAND2_X1 U4525 ( .A1(n3962), .A2(n3961), .ZN(n4323) );
  INV_X1 U4526 ( .A(n4323), .ZN(n3963) );
  NAND2_X1 U4527 ( .A1(n3963), .A2(n4017), .ZN(n5011) );
  INV_X1 U4528 ( .A(n3964), .ZN(n3972) );
  INV_X1 U4529 ( .A(n4331), .ZN(n3967) );
  INV_X1 U4530 ( .A(n3968), .ZN(n4452) );
  NAND2_X1 U4531 ( .A1(n4453), .A2(n4452), .ZN(n4335) );
  NAND2_X1 U4532 ( .A1(n3970), .A2(n4333), .ZN(n4306) );
  NAND2_X1 U4533 ( .A1(n5154), .A2(n7691), .ZN(n5003) );
  INV_X1 U4534 ( .A(n5003), .ZN(n4108) );
  NAND2_X1 U4535 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U4536 ( .A1(n5630), .A2(n5629), .ZN(n6061) );
  NAND2_X1 U4537 ( .A1(n4108), .A2(n5944), .ZN(n3974) );
  INV_X1 U4538 ( .A(n4321), .ZN(n4107) );
  NAND2_X1 U4539 ( .A1(n4107), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3973) );
  INV_X1 U4540 ( .A(n3975), .ZN(n3976) );
  MUX2_X1 U4541 ( .A(n4321), .B(n5003), .S(n5629), .Z(n3977) );
  NAND2_X1 U4542 ( .A1(n4294), .A2(n3662), .ZN(n3979) );
  NAND2_X1 U4543 ( .A1(n3978), .A2(n3979), .ZN(n3980) );
  NAND2_X1 U4544 ( .A1(n3980), .A2(n3922), .ZN(n3983) );
  NOR2_X1 U4545 ( .A1(n3981), .A2(n3669), .ZN(n4334) );
  INV_X1 U4546 ( .A(n4334), .ZN(n3982) );
  NAND2_X1 U4547 ( .A1(n3984), .A2(n3965), .ZN(n3993) );
  INV_X1 U4548 ( .A(n3986), .ZN(n4298) );
  NAND2_X1 U4549 ( .A1(n5154), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7672) );
  AOI21_X1 U4550 ( .B1(n4298), .B2(n3675), .A(n7672), .ZN(n3992) );
  INV_X1 U4551 ( .A(n4295), .ZN(n4304) );
  NAND2_X1 U4552 ( .A1(n4304), .A2(n3988), .ZN(n3990) );
  NAND2_X1 U4553 ( .A1(n3990), .A2(n3989), .ZN(n3991) );
  CLKBUF_X2 U4554 ( .A(n4006), .Z(n4079) );
  AOI22_X1 U4555 ( .A1(n4079), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4556 ( .A1(n3672), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4557 ( .A1(n3644), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4558 ( .A1(n3665), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3994) );
  NAND4_X1 U4559 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n4004)
         );
  AOI22_X1 U4560 ( .A1(n4978), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4561 ( .A1(n4950), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4562 ( .A1(n4979), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4563 ( .A1(n3643), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3999) );
  NAND4_X1 U4564 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4003)
         );
  OR2_X1 U4565 ( .A1(n4256), .A2(n4018), .ZN(n4005) );
  AOI22_X1 U4566 ( .A1(n4079), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4979), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4567 ( .A1(n3644), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4568 ( .A1(n3665), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4569 ( .A1(n4950), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4007) );
  NAND4_X1 U4570 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(n4016)
         );
  AOI22_X1 U4571 ( .A1(n3678), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4572 ( .A1(n4978), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4573 ( .A1(n4025), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4574 ( .A1(n4797), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4011) );
  NAND4_X1 U4575 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4015)
         );
  OR2_X1 U4576 ( .A1(n4256), .A2(n4214), .ZN(n4024) );
  NAND2_X1 U4577 ( .A1(n4275), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4020) );
  OR2_X1 U4578 ( .A1(n4073), .A2(n4018), .ZN(n4019) );
  XNOR2_X1 U4579 ( .A(n4059), .B(n4060), .ZN(n4058) );
  INV_X1 U4580 ( .A(n4021), .ZN(n4023) );
  NAND2_X1 U4581 ( .A1(n3662), .A2(n4214), .ZN(n4038) );
  INV_X1 U4582 ( .A(n4024), .ZN(n4036) );
  AOI22_X1 U4583 ( .A1(n4079), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4979), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4584 ( .A1(n3678), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4978), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4585 ( .A1(n4074), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4586 ( .A1(n4950), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U4587 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4035)
         );
  AOI22_X1 U4588 ( .A1(n3644), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4589 ( .A1(n3639), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4590 ( .A1(n3642), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4591 ( .A1(n7224), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U4592 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4034)
         );
  MUX2_X1 U4593 ( .A(n4209), .B(n4036), .S(n4053), .Z(n4050) );
  INV_X1 U4594 ( .A(n4050), .ZN(n4037) );
  NAND2_X1 U4595 ( .A1(n4047), .A2(n4037), .ZN(n4041) );
  NAND2_X1 U4596 ( .A1(n4275), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4040) );
  AOI21_X1 U4597 ( .B1(n3922), .B2(n4053), .A(n7691), .ZN(n4039) );
  NAND3_X1 U4598 ( .A1(n4040), .A2(n4039), .A3(n4038), .ZN(n4049) );
  XNOR2_X1 U4599 ( .A(n4058), .B(n4057), .ZN(n4502) );
  NAND2_X1 U4600 ( .A1(n4502), .A2(n3965), .ZN(n4046) );
  NAND2_X1 U4601 ( .A1(n4053), .A2(n4042), .ZN(n4092) );
  OAI21_X1 U4602 ( .B1(n4042), .B2(n4053), .A(n4092), .ZN(n4043) );
  INV_X1 U4603 ( .A(n3981), .ZN(n4459) );
  OAI211_X1 U4604 ( .C1(n4043), .C2(n7430), .A(n4459), .B(n3954), .ZN(n4044)
         );
  INV_X1 U4605 ( .A(n4044), .ZN(n4045) );
  NAND2_X1 U4606 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  NAND2_X1 U4607 ( .A1(n3669), .A2(n5249), .ZN(n4095) );
  OAI21_X1 U4608 ( .B1(n7430), .B2(n4053), .A(n4095), .ZN(n4054) );
  INV_X1 U4609 ( .A(n4054), .ZN(n4055) );
  OAI21_X1 U4610 ( .B1(n5552), .B2(n4210), .A(n4055), .ZN(n5111) );
  NAND2_X1 U4611 ( .A1(n4056), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5216)
         );
  NAND2_X1 U4612 ( .A1(n7382), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4098)
         );
  NAND2_X1 U4613 ( .A1(n4058), .A2(n4057), .ZN(n4063) );
  INV_X1 U4614 ( .A(n4059), .ZN(n4061) );
  NAND2_X1 U4615 ( .A1(n4063), .A2(n4062), .ZN(n4089) );
  NAND2_X1 U4616 ( .A1(n3661), .A2(n4066), .ZN(n4067) );
  INV_X1 U4617 ( .A(n5464), .ZN(n4069) );
  INV_X1 U4618 ( .A(n5545), .ZN(n4105) );
  NAND2_X1 U4619 ( .A1(n5464), .A2(n5417), .ZN(n4070) );
  AOI22_X1 U4620 ( .A1(n5592), .A2(n4108), .B1(n4107), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4621 ( .A1(n4978), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U4622 ( .A1(n3639), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U4623 ( .A1(n4971), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U4624 ( .A1(n3666), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U4625 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4085)
         );
  AOI22_X1 U4626 ( .A1(n3643), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4627 ( .A1(n4979), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U4628 ( .A1(n3673), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U4629 ( .A1(n4079), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4080) );
  NAND4_X1 U4630 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4084)
         );
  AOI22_X1 U4631 ( .A1(n4288), .A2(n4091), .B1(INSTQUEUE_REG_0__2__SCAN_IN), 
        .B2(n4275), .ZN(n4086) );
  INV_X1 U4632 ( .A(n4091), .ZN(n4093) );
  NAND2_X1 U4633 ( .A1(n4092), .A2(n4093), .ZN(n4126) );
  OAI21_X1 U4634 ( .B1(n4093), .B2(n4092), .A(n4126), .ZN(n4094) );
  NAND2_X1 U4635 ( .A1(n4094), .A2(n3675), .ZN(n4096) );
  NAND2_X1 U4636 ( .A1(n4096), .A2(n4095), .ZN(n4097) );
  NAND2_X1 U4637 ( .A1(n4098), .A2(n7383), .ZN(n4101) );
  NAND2_X1 U4638 ( .A1(n4099), .A2(n7485), .ZN(n4100) );
  INV_X1 U4639 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4468) );
  INV_X1 U4640 ( .A(n4102), .ZN(n4104) );
  NAND2_X1 U4641 ( .A1(n5545), .A2(n7649), .ZN(n5328) );
  NAND2_X1 U4642 ( .A1(n4105), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4106) );
  NAND2_X1 U4643 ( .A1(n5328), .A2(n4106), .ZN(n6071) );
  AOI22_X1 U4644 ( .A1(n6071), .A2(n4108), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4107), .ZN(n4109) );
  AOI22_X1 U4645 ( .A1(n4978), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U4646 ( .A1(n3665), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4647 ( .A1(n4908), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U4648 ( .A1(n3666), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4111) );
  NAND4_X1 U4649 ( .A1(n4114), .A2(n4113), .A3(n4112), .A4(n4111), .ZN(n4121)
         );
  AOI22_X1 U4650 ( .A1(n3678), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U4651 ( .A1(n4979), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U4652 ( .A1(n3673), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U4653 ( .A1(n4079), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4116) );
  NAND4_X1 U4654 ( .A1(n4119), .A2(n4118), .A3(n4117), .A4(n4116), .ZN(n4120)
         );
  AOI22_X1 U4655 ( .A1(n4288), .A2(n4127), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n4275), .ZN(n4122) );
  NAND2_X2 U4656 ( .A1(n3651), .A2(n5297), .ZN(n4148) );
  INV_X1 U4657 ( .A(n5297), .ZN(n5296) );
  NAND2_X1 U4658 ( .A1(n4124), .A2(n5296), .ZN(n4125) );
  NAND2_X1 U4659 ( .A1(n4126), .A2(n4127), .ZN(n4165) );
  OAI211_X1 U4660 ( .C1(n4127), .C2(n4126), .A(n4165), .B(n3675), .ZN(n4128)
         );
  AOI22_X1 U4661 ( .A1(n4978), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U4662 ( .A1(n3665), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4676), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U4663 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3674), .B1(n4908), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U4664 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3666), .B1(n4909), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4129) );
  NAND4_X1 U4665 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4138)
         );
  AOI22_X1 U4666 ( .A1(n3678), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U4667 ( .A1(n4979), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U4668 ( .A1(n3673), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U4669 ( .A1(n4079), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4133) );
  NAND4_X1 U4670 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4137)
         );
  NAND2_X1 U4671 ( .A1(n4288), .A2(n4163), .ZN(n4140) );
  NAND2_X1 U4672 ( .A1(n4275), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4139) );
  NAND2_X1 U4673 ( .A1(n4140), .A2(n4139), .ZN(n4149) );
  NAND2_X1 U4674 ( .A1(n4523), .A2(n4294), .ZN(n4143) );
  XNOR2_X1 U4675 ( .A(n4165), .B(n4163), .ZN(n4141) );
  NAND2_X1 U4676 ( .A1(n4141), .A2(n3675), .ZN(n4142) );
  NAND2_X1 U4677 ( .A1(n4143), .A2(n4142), .ZN(n4146) );
  XNOR2_X1 U4678 ( .A(n4146), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5234)
         );
  INV_X1 U4679 ( .A(n5234), .ZN(n4144) );
  NAND2_X1 U4680 ( .A1(n4145), .A2(n4144), .ZN(n5231) );
  NAND2_X1 U4681 ( .A1(n4146), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4147)
         );
  NAND2_X1 U4682 ( .A1(n5231), .A2(n4147), .ZN(n7399) );
  AOI22_X1 U4683 ( .A1(n4978), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U4684 ( .A1(n3665), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4676), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U4685 ( .A1(n4908), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U4686 ( .A1(n3666), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4151) );
  NAND4_X1 U4687 ( .A1(n4154), .A2(n4153), .A3(n4152), .A4(n4151), .ZN(n4160)
         );
  AOI22_X1 U4688 ( .A1(n3678), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U4689 ( .A1(n4979), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U4690 ( .A1(n3673), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U4691 ( .A1(n4079), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4155) );
  NAND4_X1 U4692 ( .A1(n4158), .A2(n4157), .A3(n4156), .A4(n4155), .ZN(n4159)
         );
  NAND2_X1 U4693 ( .A1(n4288), .A2(n4200), .ZN(n4162) );
  NAND2_X1 U4694 ( .A1(n4275), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4161) );
  NAND2_X1 U4695 ( .A1(n4162), .A2(n4161), .ZN(n4171) );
  NAND2_X1 U4696 ( .A1(n4548), .A2(n4294), .ZN(n4168) );
  INV_X1 U4697 ( .A(n4163), .ZN(n4164) );
  OR2_X1 U4698 ( .A1(n4165), .A2(n4164), .ZN(n4188) );
  XNOR2_X1 U4699 ( .A(n4188), .B(n4200), .ZN(n4166) );
  NAND2_X1 U4700 ( .A1(n4166), .A2(n3675), .ZN(n4167) );
  NAND2_X1 U4701 ( .A1(n4168), .A2(n4167), .ZN(n4169) );
  INV_X1 U4702 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7466) );
  XNOR2_X1 U4703 ( .A(n4169), .B(n7466), .ZN(n7398) );
  NAND2_X1 U4704 ( .A1(n7399), .A2(n7398), .ZN(n7397) );
  NAND2_X1 U4705 ( .A1(n4169), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4170)
         );
  NAND2_X1 U4706 ( .A1(n7397), .A2(n4170), .ZN(n5453) );
  INV_X1 U4707 ( .A(n4171), .ZN(n4172) );
  NOR2_X2 U4708 ( .A1(n4173), .A2(n4172), .ZN(n4197) );
  AOI22_X1 U4709 ( .A1(n4978), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U4710 ( .A1(n3665), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U4711 ( .A1(n4908), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U4712 ( .A1(n3666), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4174) );
  NAND4_X1 U4713 ( .A1(n4177), .A2(n4176), .A3(n4175), .A4(n4174), .ZN(n4184)
         );
  AOI22_X1 U4714 ( .A1(n3637), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U4716 ( .A1(n4979), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U4717 ( .A1(n3673), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4180) );
  INV_X1 U4718 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U4719 ( .A1(n4079), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4179) );
  NAND4_X1 U4720 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4183)
         );
  NAND2_X1 U4721 ( .A1(n4288), .A2(n4199), .ZN(n4186) );
  NAND2_X1 U4722 ( .A1(n4275), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4185) );
  XNOR2_X1 U4723 ( .A(n4197), .B(n4187), .ZN(n4554) );
  INV_X1 U4724 ( .A(n4188), .ZN(n4202) );
  NAND2_X1 U4725 ( .A1(n4202), .A2(n4200), .ZN(n4189) );
  XNOR2_X1 U4726 ( .A(n4189), .B(n4199), .ZN(n4190) );
  AND2_X1 U4727 ( .A1(n4190), .A2(n3675), .ZN(n4191) );
  AOI21_X1 U4728 ( .B1(n4554), .B2(n4294), .A(n4191), .ZN(n5454) );
  INV_X1 U4729 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U4730 ( .A1(n5454), .A2(n4363), .ZN(n4192) );
  NAND2_X1 U4731 ( .A1(n5453), .A2(n4192), .ZN(n4195) );
  INV_X1 U4732 ( .A(n5454), .ZN(n4193) );
  NAND2_X1 U4733 ( .A1(n4193), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4194)
         );
  AOI22_X1 U4734 ( .A1(n4288), .A2(n4214), .B1(INSTQUEUE_REG_0__7__SCAN_IN), 
        .B2(n4275), .ZN(n4198) );
  AND2_X1 U4735 ( .A1(n4200), .A2(n4199), .ZN(n4201) );
  NAND2_X1 U4736 ( .A1(n4202), .A2(n4201), .ZN(n4213) );
  XNOR2_X1 U4737 ( .A(n4213), .B(n4214), .ZN(n4203) );
  NAND2_X1 U4738 ( .A1(n4203), .A2(n3675), .ZN(n4204) );
  NAND2_X1 U4739 ( .A1(n4206), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4207)
         );
  INV_X1 U4740 ( .A(n4209), .ZN(n4211) );
  NAND2_X2 U4741 ( .A1(n4208), .A2(n4212), .ZN(n7016) );
  INV_X1 U4742 ( .A(n4213), .ZN(n4215) );
  NAND3_X1 U4743 ( .A1(n4215), .A2(n3675), .A3(n4214), .ZN(n4216) );
  NAND2_X1 U4744 ( .A1(n7016), .A2(n4216), .ZN(n4217) );
  INV_X1 U4745 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4371) );
  XNOR2_X1 U4746 ( .A(n4217), .B(n4371), .ZN(n6051) );
  NAND2_X1 U4747 ( .A1(n4217), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4218)
         );
  XNOR2_X1 U4748 ( .A(n7030), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6170)
         );
  INV_X1 U4749 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6181) );
  OR2_X1 U4750 ( .A1(n7030), .A2(n6181), .ZN(n4219) );
  XNOR2_X1 U4751 ( .A(n7016), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6215)
         );
  INV_X1 U4752 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4379) );
  OR2_X1 U4753 ( .A1(n7030), .A2(n4379), .ZN(n4220) );
  XNOR2_X1 U4754 ( .A(n7030), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6265)
         );
  INV_X1 U4755 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n7218) );
  XNOR2_X1 U4756 ( .A(n7030), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6247)
         );
  INV_X1 U4757 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4221) );
  OR2_X1 U4758 ( .A1(n7030), .A2(n4221), .ZN(n4222) );
  INV_X1 U4759 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6320) );
  XNOR2_X1 U4760 ( .A(n7030), .B(n6320), .ZN(n6293) );
  NAND2_X1 U4761 ( .A1(n7016), .A2(n6320), .ZN(n4225) );
  INV_X1 U4762 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U4763 ( .A1(n7016), .A2(n6318), .ZN(n4227) );
  INV_X1 U4764 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7207) );
  AND2_X1 U4765 ( .A1(n7030), .A2(n7207), .ZN(n4230) );
  INV_X1 U4766 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U4767 ( .A1(n7016), .A2(n7205), .ZN(n4231) );
  INV_X1 U4768 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7179) );
  INV_X1 U4769 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n7185) );
  AND3_X1 U4770 ( .A1(n7205), .A2(n7179), .A3(n7185), .ZN(n4232) );
  NAND2_X1 U4771 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4470) );
  NOR2_X1 U4772 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7155) );
  NOR2_X1 U4773 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6981) );
  INV_X1 U4774 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n7124) );
  INV_X1 U4775 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n7118) );
  AND4_X1 U4776 ( .A1(n7155), .A2(n6981), .A3(n7124), .A4(n7118), .ZN(n4233)
         );
  NOR2_X1 U4777 ( .A1(n7030), .A2(n4233), .ZN(n4235) );
  AND2_X1 U4778 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n7154) );
  AND2_X1 U4779 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4481) );
  AND2_X1 U4780 ( .A1(n7154), .A2(n4481), .ZN(n7125) );
  AND2_X1 U4781 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U4782 ( .A1(n7125), .A2(n4484), .ZN(n7098) );
  NAND2_X1 U4783 ( .A1(n7016), .A2(n7098), .ZN(n4234) );
  XNOR2_X1 U4784 ( .A(n7030), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6973)
         );
  NAND2_X2 U4785 ( .A1(n6970), .A2(n6973), .ZN(n6971) );
  INV_X1 U4786 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U4787 ( .A1(n7016), .A2(n7107), .ZN(n4236) );
  INV_X1 U4788 ( .A(n6962), .ZN(n4237) );
  AND2_X1 U4789 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n7078) );
  AND2_X1 U4790 ( .A1(n7078), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4495)
         );
  NAND2_X1 U4791 ( .A1(n4237), .A2(n3803), .ZN(n4241) );
  OAI21_X1 U4792 ( .B1(n6971), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n7031), 
        .ZN(n4239) );
  NOR2_X1 U4793 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4238) );
  OR2_X1 U4794 ( .A1(n7030), .A2(n4238), .ZN(n5047) );
  NAND2_X1 U4795 ( .A1(n4239), .A2(n5047), .ZN(n6943) );
  INV_X1 U4796 ( .A(n6943), .ZN(n4240) );
  INV_X1 U4797 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4242) );
  XNOR2_X1 U4798 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4262) );
  NAND2_X1 U4799 ( .A1(n4261), .A2(n4262), .ZN(n4245) );
  NAND2_X1 U4800 ( .A1(n5630), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U4801 ( .A1(n4245), .A2(n4244), .ZN(n4273) );
  MUX2_X1 U4802 ( .A(n5417), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4272) );
  NOR2_X1 U4803 ( .A1(n3731), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4246)
         );
  NAND2_X1 U4804 ( .A1(n7231), .A2(n7649), .ZN(n4247) );
  NAND2_X1 U4805 ( .A1(n4252), .A2(n4247), .ZN(n4249) );
  NAND2_X1 U4806 ( .A1(n3804), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4248) );
  NAND2_X1 U4807 ( .A1(n4249), .A2(n4248), .ZN(n4284) );
  MUX2_X1 U4808 ( .A(n7649), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(n3804), 
        .Z(n4251) );
  XNOR2_X1 U4809 ( .A(n4252), .B(n4251), .ZN(n4315) );
  INV_X1 U4810 ( .A(n4315), .ZN(n4253) );
  AOI21_X1 U4811 ( .B1(n4316), .B2(n4253), .A(n4275), .ZN(n4282) );
  AND2_X1 U4812 ( .A1(n3809), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4254)
         );
  NOR2_X1 U4813 ( .A1(n4261), .A2(n4254), .ZN(n4255) );
  OAI21_X1 U4814 ( .B1(n4256), .B2(n3935), .A(n4255), .ZN(n4257) );
  NAND2_X1 U4815 ( .A1(n4257), .A2(n4017), .ZN(n4259) );
  NAND2_X1 U4816 ( .A1(n3935), .A2(n4017), .ZN(n4258) );
  NAND2_X1 U4817 ( .A1(n4258), .A2(n3988), .ZN(n4278) );
  NAND2_X1 U4818 ( .A1(n4259), .A2(n4278), .ZN(n4260) );
  XNOR2_X1 U4819 ( .A(n4262), .B(n4261), .ZN(n4314) );
  INV_X1 U4820 ( .A(n4275), .ZN(n4265) );
  INV_X1 U4821 ( .A(n4314), .ZN(n4264) );
  NAND2_X1 U4822 ( .A1(n4288), .A2(n3965), .ZN(n4263) );
  OAI211_X1 U4823 ( .C1(n4265), .C2(n4264), .A(n4263), .B(n3954), .ZN(n4266)
         );
  INV_X1 U4824 ( .A(n4266), .ZN(n4267) );
  OAI21_X1 U4825 ( .B1(n4269), .B2(n4268), .A(n4267), .ZN(n4271) );
  NAND3_X1 U4826 ( .A1(n4269), .A2(n3745), .A3(n4268), .ZN(n4270) );
  XNOR2_X1 U4827 ( .A(n4273), .B(n4272), .ZN(n4313) );
  INV_X1 U4828 ( .A(n4278), .ZN(n4274) );
  AOI21_X1 U4829 ( .B1(n4275), .B2(n4313), .A(n4274), .ZN(n4276) );
  INV_X1 U4830 ( .A(n4288), .ZN(n4277) );
  INV_X1 U4831 ( .A(n4316), .ZN(n4279) );
  AOI22_X1 U4832 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n7691), .B1(n4280), .B2(n4279), .ZN(n4281) );
  INV_X1 U4833 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4285) );
  NAND2_X1 U4834 ( .A1(n4285), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4286) );
  INV_X1 U4835 ( .A(n4318), .ZN(n4290) );
  NAND2_X1 U4836 ( .A1(n4291), .A2(n4290), .ZN(n4292) );
  NAND2_X1 U4837 ( .A1(n4295), .A2(n4294), .ZN(n4465) );
  INV_X1 U4838 ( .A(n4465), .ZN(n4296) );
  NAND2_X1 U4839 ( .A1(n7693), .A2(n4296), .ZN(n4309) );
  NAND2_X1 U4840 ( .A1(n4297), .A2(n4017), .ZN(n4299) );
  MUX2_X1 U4841 ( .A(n4299), .B(n7430), .S(n4298), .Z(n4303) );
  NAND2_X1 U4842 ( .A1(n4300), .A2(n3933), .ZN(n4302) );
  OAI21_X1 U4843 ( .B1(n4689), .B2(n3989), .A(n3982), .ZN(n4305) );
  NAND2_X1 U4844 ( .A1(n4457), .A2(n4305), .ZN(n4308) );
  NAND2_X1 U4845 ( .A1(n4308), .A2(n4307), .ZN(n4467) );
  NAND2_X1 U4846 ( .A1(n4309), .A2(n4467), .ZN(n5127) );
  INV_X1 U4847 ( .A(n4310), .ZN(n4311) );
  INV_X1 U4848 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7710) );
  NAND2_X1 U4849 ( .A1(n4311), .A2(n7710), .ZN(n7428) );
  NAND2_X1 U4850 ( .A1(n3965), .A2(n7428), .ZN(n4320) );
  NOR3_X1 U4851 ( .A1(n4315), .A2(n4314), .A3(n4313), .ZN(n4317) );
  OAI21_X1 U4852 ( .B1(n4318), .B2(n4317), .A(n4316), .ZN(n7623) );
  NAND2_X1 U4853 ( .A1(n7709), .A2(n7623), .ZN(n5072) );
  INV_X1 U4854 ( .A(n5072), .ZN(n4319) );
  AND3_X1 U4855 ( .A1(n4320), .A2(n4312), .A3(n4319), .ZN(n4322) );
  OAI21_X1 U4856 ( .B1(n5127), .B2(n4322), .A(n7688), .ZN(n4329) );
  NAND2_X1 U4857 ( .A1(n3988), .A2(n7428), .ZN(n5018) );
  NAND2_X1 U4858 ( .A1(n5018), .A2(n7709), .ZN(n4326) );
  AND2_X1 U4859 ( .A1(n3968), .A2(n4017), .ZN(n4325) );
  OAI22_X1 U4860 ( .A1(n4324), .A2(n4326), .B1(n4325), .B2(n4312), .ZN(n4327)
         );
  NAND2_X1 U4861 ( .A1(n3646), .A2(n4327), .ZN(n4328) );
  INV_X1 U4862 ( .A(n4689), .ZN(n5139) );
  NOR2_X1 U4863 ( .A1(n4331), .A2(n3989), .ZN(n4332) );
  NAND2_X1 U4864 ( .A1(n5139), .A2(n4332), .ZN(n5143) );
  NAND2_X1 U4865 ( .A1(n4334), .A2(n4333), .ZN(n7654) );
  AND2_X1 U4866 ( .A1(n5143), .A2(n7654), .ZN(n7619) );
  OR2_X1 U4867 ( .A1(n4324), .A2(n5030), .ZN(n5120) );
  INV_X1 U4868 ( .A(n4335), .ZN(n4336) );
  NAND2_X1 U4869 ( .A1(n4336), .A2(n3949), .ZN(n4337) );
  NAND4_X1 U4870 ( .A1(n4330), .A2(n7619), .A3(n5120), .A4(n4337), .ZN(n4338)
         );
  INV_X1 U4871 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n7472) );
  NAND2_X1 U4872 ( .A1(n4440), .A2(n7472), .ZN(n4341) );
  INV_X1 U4873 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4339) );
  NAND2_X1 U4874 ( .A1(n5191), .A2(n4339), .ZN(n4340) );
  NAND3_X1 U4875 ( .A1(n4341), .A2(n3671), .A3(n4340), .ZN(n4343) );
  NAND2_X1 U4876 ( .A1(n4343), .A2(n4342), .ZN(n4348) );
  NAND2_X1 U4877 ( .A1(n4440), .A2(EBX_REG_0__SCAN_IN), .ZN(n4346) );
  INV_X1 U4878 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4344) );
  NAND2_X1 U4879 ( .A1(n3671), .A2(n4344), .ZN(n4345) );
  NAND2_X1 U4880 ( .A1(n4346), .A2(n4345), .ZN(n5229) );
  XNOR2_X1 U4881 ( .A(n4348), .B(n5229), .ZN(n5852) );
  INV_X1 U4882 ( .A(n5229), .ZN(n4347) );
  NOR2_X1 U4883 ( .A1(n4348), .A2(n4347), .ZN(n4349) );
  INV_X1 U4884 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n7485) );
  NAND2_X1 U4885 ( .A1(n4440), .A2(n7485), .ZN(n4351) );
  INV_X1 U4886 ( .A(EBX_REG_2__SCAN_IN), .ZN(n7512) );
  NAND2_X1 U4887 ( .A1(n5191), .A2(n7512), .ZN(n4350) );
  NAND3_X1 U4888 ( .A1(n4351), .A2(n4448), .A3(n4350), .ZN(n4353) );
  NAND2_X1 U4889 ( .A1(n3933), .A2(n7512), .ZN(n4352) );
  NAND2_X1 U4890 ( .A1(n4353), .A2(n4352), .ZN(n5203) );
  MUX2_X1 U4891 ( .A(n4437), .B(n4448), .S(EBX_REG_3__SCAN_IN), .Z(n4355) );
  OR2_X1 U4892 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4354)
         );
  AND2_X1 U4893 ( .A1(n4355), .A2(n4354), .ZN(n6366) );
  INV_X1 U4894 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4469) );
  NAND2_X1 U4895 ( .A1(n4440), .A2(n4469), .ZN(n4357) );
  INV_X1 U4896 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U4897 ( .A1(n5191), .A2(n6144), .ZN(n4356) );
  NAND3_X1 U4898 ( .A1(n4357), .A2(n4448), .A3(n4356), .ZN(n4359) );
  NAND2_X1 U4899 ( .A1(n3933), .A2(n6144), .ZN(n4358) );
  AND2_X1 U4900 ( .A1(n4359), .A2(n4358), .ZN(n5197) );
  MUX2_X1 U4901 ( .A(n4437), .B(n4448), .S(EBX_REG_5__SCAN_IN), .Z(n4360) );
  OAI21_X1 U4902 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5228), .A(n4360), 
        .ZN(n5213) );
  NAND2_X1 U4903 ( .A1(n4440), .A2(n4363), .ZN(n4365) );
  INV_X1 U4904 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U4905 ( .A1(n5191), .A2(n5937), .ZN(n4364) );
  NAND3_X1 U4906 ( .A1(n4365), .A2(n4448), .A3(n4364), .ZN(n4367) );
  NAND2_X1 U4907 ( .A1(n3933), .A2(n5937), .ZN(n4366) );
  AND2_X1 U4908 ( .A1(n4367), .A2(n4366), .ZN(n5364) );
  MUX2_X1 U4909 ( .A(n4437), .B(n4448), .S(EBX_REG_7__SCAN_IN), .Z(n4369) );
  OR2_X1 U4910 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4368)
         );
  NAND2_X1 U4911 ( .A1(n4369), .A2(n4368), .ZN(n5451) );
  INV_X1 U4912 ( .A(n5451), .ZN(n4370) );
  NAND2_X1 U4913 ( .A1(n4440), .A2(n4371), .ZN(n4373) );
  INV_X1 U4914 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U4915 ( .A1(n5191), .A2(n5789), .ZN(n4372) );
  NAND3_X1 U4916 ( .A1(n4373), .A2(n4448), .A3(n4372), .ZN(n4375) );
  NAND2_X1 U4917 ( .A1(n3933), .A2(n5789), .ZN(n4374) );
  NAND2_X1 U4918 ( .A1(n4375), .A2(n4374), .ZN(n5712) );
  MUX2_X1 U4919 ( .A(n4437), .B(n4448), .S(EBX_REG_9__SCAN_IN), .Z(n4376) );
  OAI21_X1 U4920 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5228), .A(n4376), 
        .ZN(n6048) );
  NAND2_X1 U4921 ( .A1(n4378), .A2(n4377), .ZN(n6165) );
  NAND2_X1 U4922 ( .A1(n4440), .A2(n4379), .ZN(n4381) );
  INV_X1 U4923 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U4924 ( .A1(n5191), .A2(n6186), .ZN(n4380) );
  NAND3_X1 U4925 ( .A1(n4381), .A2(n4448), .A3(n4380), .ZN(n4383) );
  NAND2_X1 U4926 ( .A1(n3933), .A2(n6186), .ZN(n4382) );
  AND2_X1 U4927 ( .A1(n4383), .A2(n4382), .ZN(n6164) );
  MUX2_X1 U4928 ( .A(n4437), .B(n4448), .S(EBX_REG_11__SCAN_IN), .Z(n4385) );
  OR2_X1 U4929 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4384)
         );
  NAND2_X1 U4930 ( .A1(n6198), .A2(n6197), .ZN(n6278) );
  MUX2_X1 U4931 ( .A(n4437), .B(n4448), .S(EBX_REG_13__SCAN_IN), .Z(n4386) );
  OAI21_X1 U4932 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5228), .A(n4386), 
        .ZN(n6276) );
  NAND2_X1 U4933 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4387) );
  NAND2_X1 U4934 ( .A1(n4440), .A2(n4387), .ZN(n4389) );
  INV_X1 U4935 ( .A(EBX_REG_12__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U4936 ( .A1(n5191), .A2(n7559), .ZN(n4388) );
  NAND2_X1 U4937 ( .A1(n4389), .A2(n4388), .ZN(n4391) );
  NAND2_X1 U4938 ( .A1(n3933), .A2(n7559), .ZN(n4390) );
  NAND2_X1 U4939 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U4940 ( .A1(n4440), .A2(n4393), .ZN(n4396) );
  INV_X1 U4941 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U4942 ( .A1(n5191), .A2(n4394), .ZN(n4395) );
  AOI22_X1 U4943 ( .A1(n4396), .A2(n4395), .B1(n3933), .B2(n4394), .ZN(n6309)
         );
  MUX2_X1 U4944 ( .A(n4437), .B(n4448), .S(EBX_REG_15__SCAN_IN), .Z(n4398) );
  OR2_X1 U4945 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4397)
         );
  NAND2_X1 U4946 ( .A1(n4398), .A2(n4397), .ZN(n6341) );
  NAND2_X1 U4947 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4399) );
  NAND2_X1 U4948 ( .A1(n4440), .A2(n4399), .ZN(n4401) );
  INV_X1 U4949 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U4950 ( .A1(n5191), .A2(n4402), .ZN(n4400) );
  NAND2_X1 U4951 ( .A1(n4401), .A2(n4400), .ZN(n4404) );
  NAND2_X1 U4952 ( .A1(n3933), .A2(n4402), .ZN(n4403) );
  NAND2_X1 U4953 ( .A1(n4404), .A2(n4403), .ZN(n6354) );
  NAND2_X1 U4954 ( .A1(n6355), .A2(n6354), .ZN(n6508) );
  MUX2_X1 U4955 ( .A(n4437), .B(n4448), .S(EBX_REG_17__SCAN_IN), .Z(n4405) );
  OAI21_X1 U4956 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5228), .A(n4405), 
        .ZN(n6509) );
  NAND2_X1 U4957 ( .A1(n4440), .A2(n7185), .ZN(n4407) );
  INV_X1 U4958 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4408) );
  NAND2_X1 U4959 ( .A1(n5191), .A2(n4408), .ZN(n4406) );
  NAND3_X1 U4960 ( .A1(n4407), .A2(n4448), .A3(n4406), .ZN(n4410) );
  NAND2_X1 U4961 ( .A1(n3933), .A2(n4408), .ZN(n4409) );
  AND2_X1 U4962 ( .A1(n4410), .A2(n4409), .ZN(n6499) );
  NAND2_X1 U4963 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4411) );
  OAI211_X1 U4964 ( .C1(n5030), .C2(EBX_REG_19__SCAN_IN), .A(n4440), .B(n4411), 
        .ZN(n4412) );
  OAI21_X1 U4965 ( .B1(n4437), .B2(EBX_REG_19__SCAN_IN), .A(n4412), .ZN(n7162)
         );
  NAND2_X1 U4966 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4413) );
  NAND2_X1 U4967 ( .A1(n4440), .A2(n4413), .ZN(n4415) );
  INV_X1 U4968 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U4969 ( .A1(n5191), .A2(n4416), .ZN(n4414) );
  NAND2_X1 U4970 ( .A1(n4415), .A2(n4414), .ZN(n4418) );
  NAND2_X1 U4971 ( .A1(n3933), .A2(n4416), .ZN(n4417) );
  NAND2_X1 U4972 ( .A1(n4418), .A2(n4417), .ZN(n6537) );
  NAND2_X1 U4973 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4419) );
  OAI211_X1 U4974 ( .C1(n5030), .C2(EBX_REG_21__SCAN_IN), .A(n4440), .B(n4419), 
        .ZN(n4420) );
  OAI21_X1 U4975 ( .B1(n4437), .B2(EBX_REG_21__SCAN_IN), .A(n4420), .ZN(n7143)
         );
  INV_X1 U4976 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U4977 ( .A1(n4440), .A2(n6998), .ZN(n4422) );
  INV_X1 U4978 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U4979 ( .A1(n5191), .A2(n6528), .ZN(n4421) );
  NAND3_X1 U4980 ( .A1(n4422), .A2(n4448), .A3(n4421), .ZN(n4424) );
  NAND2_X1 U4981 ( .A1(n3933), .A2(n6528), .ZN(n4423) );
  AND2_X1 U4982 ( .A1(n4424), .A2(n4423), .ZN(n6488) );
  MUX2_X1 U4983 ( .A(n4437), .B(n4448), .S(EBX_REG_23__SCAN_IN), .Z(n4426) );
  OR2_X1 U4984 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4425)
         );
  AND2_X1 U4985 ( .A1(n4426), .A2(n4425), .ZN(n6479) );
  NAND2_X1 U4986 ( .A1(n4440), .A2(n7118), .ZN(n4428) );
  INV_X1 U4987 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4429) );
  NAND2_X1 U4988 ( .A1(n5191), .A2(n4429), .ZN(n4427) );
  NAND3_X1 U4989 ( .A1(n4428), .A2(n4448), .A3(n4427), .ZN(n4431) );
  NAND2_X1 U4990 ( .A1(n3933), .A2(n4429), .ZN(n4430) );
  NAND2_X1 U4991 ( .A1(n4431), .A2(n4430), .ZN(n6465) );
  MUX2_X1 U4992 ( .A(n4437), .B(n4448), .S(EBX_REG_25__SCAN_IN), .Z(n4432) );
  OAI21_X1 U4993 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5228), .A(n4432), 
        .ZN(n6453) );
  INV_X1 U4994 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U4995 ( .A1(n4440), .A2(n6963), .ZN(n4433) );
  OAI211_X1 U4996 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5030), .A(n4433), .B(n4448), 
        .ZN(n4436) );
  INV_X1 U4997 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4434) );
  NAND2_X1 U4998 ( .A1(n3933), .A2(n4434), .ZN(n4435) );
  AND2_X1 U4999 ( .A1(n4436), .A2(n4435), .ZN(n6441) );
  MUX2_X1 U5000 ( .A(n4437), .B(n3671), .S(EBX_REG_27__SCAN_IN), .Z(n4439) );
  OR2_X1 U5001 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4438)
         );
  AND2_X1 U5002 ( .A1(n4439), .A2(n4438), .ZN(n6426) );
  INV_X1 U5003 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U5004 ( .A1(n4440), .A2(n5062), .ZN(n4441) );
  OAI211_X1 U5005 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5030), .A(n4441), .B(n4448), 
        .ZN(n4443) );
  INV_X1 U5006 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U5007 ( .A1(n3933), .A2(n6522), .ZN(n4442) );
  NAND2_X1 U5008 ( .A1(n4443), .A2(n4442), .ZN(n5060) );
  OR2_X1 U5009 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4446)
         );
  INV_X1 U5010 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4444) );
  NAND2_X1 U5011 ( .A1(n5191), .A2(n4444), .ZN(n4445) );
  AND2_X1 U5012 ( .A1(n4446), .A2(n4445), .ZN(n4449) );
  INV_X1 U5013 ( .A(n4449), .ZN(n4450) );
  NOR2_X1 U5014 ( .A1(n4448), .A2(EBX_REG_29__SCAN_IN), .ZN(n4447) );
  AOI21_X1 U5015 ( .B1(n4449), .B2(n4448), .A(n4447), .ZN(n6407) );
  OAI21_X1 U5016 ( .B1(n6406), .B2(n4450), .A(n5028), .ZN(n4451) );
  OAI22_X1 U5017 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n5030), .ZN(n5029) );
  NAND3_X1 U5018 ( .A1(n4453), .A2(n3662), .A3(n4452), .ZN(n4454) );
  NAND2_X1 U5019 ( .A1(n5164), .A2(n4454), .ZN(n4455) );
  NAND2_X1 U5020 ( .A1(n6381), .A2(n7495), .ZN(n4493) );
  NOR2_X1 U5021 ( .A1(n4307), .A2(n3988), .ZN(n7639) );
  INV_X1 U5022 ( .A(n7492), .ZN(n4464) );
  AOI21_X1 U5023 ( .B1(n3969), .B2(n3965), .A(n3968), .ZN(n4458) );
  OAI21_X1 U5024 ( .B1(n4459), .B2(n4458), .A(n4457), .ZN(n4460) );
  INV_X1 U5025 ( .A(n4460), .ZN(n4461) );
  AND2_X1 U5026 ( .A1(n4462), .A2(n4461), .ZN(n5132) );
  OAI21_X1 U5027 ( .B1(n4017), .B2(n4456), .A(n5132), .ZN(n4463) );
  NAND2_X1 U5028 ( .A1(n4472), .A2(n4463), .ZN(n6323) );
  NAND2_X1 U5029 ( .A1(n3922), .A2(n3965), .ZN(n5850) );
  NOR2_X1 U5030 ( .A1(n5850), .A2(n4312), .ZN(n5123) );
  NOR2_X1 U5031 ( .A1(n4465), .A2(n5123), .ZN(n4466) );
  NAND2_X1 U5032 ( .A1(n6175), .A2(n7462), .ZN(n7196) );
  NOR2_X1 U5033 ( .A1(n7485), .A2(n7472), .ZN(n5457) );
  NOR2_X1 U5034 ( .A1(n4469), .A2(n4468), .ZN(n7451) );
  AND2_X1 U5035 ( .A1(n5457), .A2(n7451), .ZN(n7467) );
  NAND3_X1 U5036 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n7467), .ZN(n5863) );
  NAND2_X1 U5037 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4476) );
  NAND2_X1 U5038 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6250) );
  NOR3_X1 U5039 ( .A1(n5863), .A2(n4476), .A3(n6250), .ZN(n4488) );
  NAND2_X1 U5040 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6324) );
  INV_X1 U5041 ( .A(n6324), .ZN(n6321) );
  NAND2_X1 U5042 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6321), .ZN(n6327) );
  NOR2_X1 U5043 ( .A1(n6318), .A2(n6327), .ZN(n7199) );
  NAND3_X1 U5044 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n7199), .ZN(n7187) );
  NOR2_X1 U5045 ( .A1(n7187), .A2(n4470), .ZN(n4490) );
  AND2_X1 U5046 ( .A1(n4488), .A2(n4490), .ZN(n4471) );
  OR2_X1 U5047 ( .A1(n6175), .A2(n4471), .ZN(n4475) );
  OR2_X1 U5048 ( .A1(n6323), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4474)
         );
  NOR2_X2 U5049 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5871) );
  NAND2_X1 U5050 ( .A1(n5871), .A2(n7422), .ZN(n7417) );
  OR2_X2 U5051 ( .A1(n7417), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7477) );
  NOR2_X1 U5052 ( .A1(n7460), .A2(n4472), .ZN(n7491) );
  INV_X1 U5053 ( .A(n7491), .ZN(n4473) );
  NAND2_X1 U5054 ( .A1(n4475), .A2(n5861), .ZN(n4480) );
  INV_X1 U5055 ( .A(n4490), .ZN(n4477) );
  INV_X1 U5056 ( .A(n4476), .ZN(n6207) );
  INV_X1 U5057 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7489) );
  OAI21_X1 U5058 ( .B1(n7472), .B2(n7489), .A(n7485), .ZN(n7453) );
  NAND2_X1 U5059 ( .A1(n7451), .A2(n7453), .ZN(n7461) );
  NOR3_X1 U5060 ( .A1(n4363), .A2(n7466), .A3(n7461), .ZN(n6203) );
  NAND2_X1 U5061 ( .A1(n6207), .A2(n6203), .ZN(n6179) );
  OR2_X1 U5062 ( .A1(n6250), .A2(n6179), .ZN(n4489) );
  NOR2_X1 U5063 ( .A1(n4477), .A2(n4489), .ZN(n4478) );
  NOR2_X1 U5064 ( .A1(n7462), .A2(n4478), .ZN(n4479) );
  OR2_X1 U5065 ( .A1(n4480), .A2(n4479), .ZN(n7168) );
  INV_X1 U5066 ( .A(n7154), .ZN(n7137) );
  OAI22_X1 U5067 ( .A1(n7168), .A2(n7137), .B1(n7196), .B2(n4480), .ZN(n7138)
         );
  INV_X1 U5068 ( .A(n4481), .ZN(n4482) );
  NAND2_X1 U5069 ( .A1(n7196), .A2(n4482), .ZN(n4483) );
  NAND2_X1 U5070 ( .A1(n7138), .A2(n4483), .ZN(n7130) );
  NOR2_X1 U5071 ( .A1(n7492), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5220)
         );
  INV_X1 U5072 ( .A(n7471), .ZN(n4485) );
  AOI21_X1 U5073 ( .B1(n4485), .B2(n7462), .A(n4484), .ZN(n4486) );
  NAND2_X1 U5074 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n7099) );
  AND2_X1 U5075 ( .A1(n7196), .A2(n7099), .ZN(n4487) );
  NOR2_X1 U5076 ( .A1(n7115), .A2(n4487), .ZN(n7077) );
  OAI21_X1 U5077 ( .B1(n4495), .B2(n7176), .A(n7077), .ZN(n7066) );
  INV_X1 U5078 ( .A(REIP_REG_30__SCAN_IN), .ZN(n7339) );
  NOR2_X1 U5079 ( .A1(n7477), .A2(n7339), .ZN(n6936) );
  NAND2_X1 U5080 ( .A1(n7471), .A2(n4488), .ZN(n6249) );
  NAND2_X1 U5081 ( .A1(n7219), .A2(n4490), .ZN(n7156) );
  INV_X1 U5082 ( .A(n4495), .ZN(n7069) );
  NOR3_X1 U5083 ( .A1(n7087), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n7069), 
        .ZN(n4491) );
  AOI211_X1 U5084 ( .C1(n7066), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n6936), .B(n4491), .ZN(n4492) );
  OAI21_X1 U5085 ( .B1(n6942), .B2(n7212), .A(n4494), .ZN(U2988) );
  NAND3_X1 U5086 ( .A1(n4495), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U5087 ( .A1(n6944), .A2(n4496), .ZN(n4497) );
  AOI21_X1 U5088 ( .B1(n4500), .B2(n7031), .A(n4499), .ZN(n4501) );
  XNOR2_X1 U5089 ( .A(n4501), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n7076)
         );
  NAND2_X1 U5090 ( .A1(n4502), .A2(n4665), .ZN(n4507) );
  NOR2_X1 U5091 ( .A1(n3968), .A2(n7669), .ZN(n4526) );
  NAND2_X1 U5092 ( .A1(n4526), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4505) );
  AOI22_X1 U5093 ( .A1(n4542), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n7669), .ZN(n4504) );
  AND2_X1 U5094 ( .A1(n4505), .A2(n4504), .ZN(n4506) );
  NAND2_X1 U5095 ( .A1(n4509), .A2(n4665), .ZN(n4513) );
  NAND2_X1 U5096 ( .A1(n4526), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U5097 ( .A1(n4542), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n7669), .ZN(n4510) );
  AND2_X1 U5098 ( .A1(n4511), .A2(n4510), .ZN(n4512) );
  NAND2_X1 U5099 ( .A1(n4513), .A2(n4512), .ZN(n5114) );
  NAND2_X1 U5100 ( .A1(n5115), .A2(n5114), .ZN(n5113) );
  INV_X1 U5101 ( .A(n5114), .ZN(n4514) );
  NAND2_X1 U5102 ( .A1(n4514), .A2(n4543), .ZN(n4515) );
  NAND2_X1 U5103 ( .A1(n5113), .A2(n4515), .ZN(n5180) );
  NAND2_X1 U5104 ( .A1(n7669), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4850) );
  NAND2_X1 U5105 ( .A1(n4526), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4519) );
  INV_X1 U5106 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U5107 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4533) );
  OAI21_X1 U5108 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4533), .ZN(n7518) );
  NAND2_X1 U5109 ( .A1(n4543), .A2(n7518), .ZN(n4516) );
  OAI21_X1 U5110 ( .B1(n4850), .B2(n7503), .A(n4516), .ZN(n4517) );
  AOI21_X1 U5111 ( .B1(n4995), .B2(EAX_REG_2__SCAN_IN), .A(n4517), .ZN(n4518)
         );
  NAND2_X1 U5112 ( .A1(n4519), .A2(n4518), .ZN(n5200) );
  NAND2_X1 U5113 ( .A1(n5201), .A2(n5200), .ZN(n4522) );
  NAND2_X1 U5114 ( .A1(n4520), .A2(n5182), .ZN(n4521) );
  NAND2_X1 U5115 ( .A1(n4523), .A2(n4665), .ZN(n4531) );
  INV_X1 U5116 ( .A(n4534), .ZN(n4525) );
  INV_X1 U5117 ( .A(n4544), .ZN(n4524) );
  OAI21_X1 U5118 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n4525), .A(n4524), 
        .ZN(n6152) );
  INV_X1 U5119 ( .A(n4526), .ZN(n4538) );
  AOI21_X1 U5120 ( .B1(n6147), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4527) );
  AOI21_X1 U5121 ( .B1(n4995), .B2(EAX_REG_4__SCAN_IN), .A(n4527), .ZN(n4528)
         );
  OAI21_X1 U5122 ( .B1(n4538), .B2(n7632), .A(n4528), .ZN(n4529) );
  OAI21_X1 U5123 ( .B1(n4967), .B2(n6152), .A(n4529), .ZN(n4530) );
  INV_X1 U5124 ( .A(n5083), .ZN(n4532) );
  NAND2_X1 U5125 ( .A1(n4532), .A2(n4665), .ZN(n4541) );
  INV_X1 U5126 ( .A(n4533), .ZN(n4535) );
  OAI21_X1 U5127 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4535), .A(n4534), 
        .ZN(n7395) );
  AOI22_X1 U5128 ( .A1(n5013), .A2(n7395), .B1(n4994), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4537) );
  NAND2_X1 U5129 ( .A1(n4995), .A2(EAX_REG_3__SCAN_IN), .ZN(n4536) );
  OAI211_X1 U5130 ( .C1(n4538), .C2(n3804), .A(n4537), .B(n4536), .ZN(n4539)
         );
  INV_X1 U5131 ( .A(n4539), .ZN(n4540) );
  NAND3_X1 U5132 ( .A1(n5194), .A2(n5195), .A3(n5492), .ZN(n5193) );
  INV_X1 U5133 ( .A(n5193), .ZN(n4550) );
  INV_X1 U5134 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4546) );
  OAI21_X1 U5135 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n4544), .A(n4555), 
        .ZN(n7530) );
  AOI22_X1 U5136 ( .A1(n5013), .A2(n7530), .B1(n4994), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4545) );
  OAI21_X1 U5137 ( .B1(n4721), .B2(n4546), .A(n4545), .ZN(n4547) );
  INV_X1 U5138 ( .A(n5209), .ZN(n4549) );
  NAND2_X1 U5139 ( .A1(n4550), .A2(n4549), .ZN(n5208) );
  NAND2_X1 U5140 ( .A1(n4995), .A2(EAX_REG_6__SCAN_IN), .ZN(n4552) );
  OAI21_X1 U5141 ( .B1(n7696), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n7669), 
        .ZN(n4551) );
  XNOR2_X1 U5142 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n4555), .ZN(n5931) );
  AOI22_X1 U5143 ( .A1(n4552), .A2(n4551), .B1(n5013), .B2(n5931), .ZN(n4553)
         );
  AOI21_X1 U5144 ( .B1(n4554), .B2(n4665), .A(n4553), .ZN(n5360) );
  INV_X1 U5145 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4558) );
  OAI21_X1 U5146 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n4556), .A(n4562), 
        .ZN(n7533) );
  NAND2_X1 U5147 ( .A1(n5013), .A2(n7533), .ZN(n4557) );
  OAI21_X1 U5148 ( .B1(n4558), .B2(n4850), .A(n4557), .ZN(n4559) );
  AOI21_X1 U5149 ( .B1(n4995), .B2(EAX_REG_7__SCAN_IN), .A(n4559), .ZN(n4560)
         );
  NAND2_X1 U5150 ( .A1(n5361), .A2(n5448), .ZN(n5447) );
  INV_X1 U5151 ( .A(n5447), .ZN(n4577) );
  XOR2_X1 U5152 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4578), .Z(n6054) );
  AOI22_X1 U5153 ( .A1(n4074), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4566) );
  AOI22_X1 U5154 ( .A1(n4977), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5155 ( .A1(n4979), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4564) );
  AOI22_X1 U5156 ( .A1(n4978), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4563) );
  NAND4_X1 U5157 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .ZN(n4572)
         );
  AOI22_X1 U5158 ( .A1(n4079), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5159 ( .A1(n3673), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5160 ( .A1(n3637), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5161 ( .A1(n4950), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4567) );
  NAND4_X1 U5162 ( .A1(n4570), .A2(n4569), .A3(n4568), .A4(n4567), .ZN(n4571)
         );
  OR2_X1 U5163 ( .A1(n4572), .A2(n4571), .ZN(n4573) );
  AOI22_X1 U5164 ( .A1(n4665), .A2(n4573), .B1(n4994), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U5165 ( .A1(n4995), .A2(EAX_REG_8__SCAN_IN), .ZN(n4574) );
  OAI211_X1 U5166 ( .C1(n6054), .C2(n4967), .A(n4575), .B(n4574), .ZN(n4576)
         );
  INV_X1 U5167 ( .A(n4576), .ZN(n5711) );
  XNOR2_X1 U5168 ( .A(n4595), .B(n7549), .ZN(n7543) );
  NAND2_X1 U5169 ( .A1(n7543), .A2(n5013), .ZN(n4594) );
  AOI22_X1 U5170 ( .A1(n4079), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4979), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4582) );
  AOI22_X1 U5171 ( .A1(n3673), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4581) );
  AOI22_X1 U5172 ( .A1(n4977), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4580) );
  AOI22_X1 U5173 ( .A1(n3637), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4579) );
  NAND4_X1 U5174 ( .A1(n4582), .A2(n4581), .A3(n4580), .A4(n4579), .ZN(n4588)
         );
  AOI22_X1 U5175 ( .A1(n4978), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4586) );
  AOI22_X1 U5176 ( .A1(n3672), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5177 ( .A1(n4797), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4584) );
  AOI22_X1 U5178 ( .A1(n4950), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4583) );
  NAND4_X1 U5179 ( .A1(n4586), .A2(n4585), .A3(n4584), .A4(n4583), .ZN(n4587)
         );
  NOR2_X1 U5180 ( .A1(n4588), .A2(n4587), .ZN(n4591) );
  NAND2_X1 U5181 ( .A1(n4995), .A2(EAX_REG_9__SCAN_IN), .ZN(n4590) );
  NAND2_X1 U5182 ( .A1(n4994), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4589)
         );
  OAI211_X1 U5183 ( .C1(n4686), .C2(n4591), .A(n4590), .B(n4589), .ZN(n4592)
         );
  INV_X1 U5184 ( .A(n4592), .ZN(n4593) );
  XOR2_X1 U5185 ( .A(n6189), .B(n4619), .Z(n6216) );
  AOI22_X1 U5186 ( .A1(n3637), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4599) );
  AOI22_X1 U5187 ( .A1(n4978), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4598) );
  AOI22_X1 U5188 ( .A1(n4908), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4597) );
  AOI22_X1 U5189 ( .A1(n7224), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4596) );
  NAND4_X1 U5190 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4605)
         );
  AOI22_X1 U5191 ( .A1(n4977), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5192 ( .A1(n4979), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4602) );
  AOI22_X1 U5193 ( .A1(n4079), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4601) );
  AOI22_X1 U5194 ( .A1(n4950), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4600) );
  NAND4_X1 U5195 ( .A1(n4603), .A2(n4602), .A3(n4601), .A4(n4600), .ZN(n4604)
         );
  OR2_X1 U5196 ( .A1(n4605), .A2(n4604), .ZN(n4606) );
  AOI22_X1 U5197 ( .A1(n4665), .A2(n4606), .B1(n4994), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U5198 ( .A1(n4995), .A2(EAX_REG_10__SCAN_IN), .ZN(n4607) );
  OAI211_X1 U5199 ( .C1(n6216), .C2(n4967), .A(n4608), .B(n4607), .ZN(n6160)
         );
  AOI22_X1 U5200 ( .A1(n4978), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4612) );
  AOI22_X1 U5201 ( .A1(n3672), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4611) );
  AOI22_X1 U5202 ( .A1(n4977), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4610) );
  AOI22_X1 U5203 ( .A1(n4979), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4609) );
  NAND4_X1 U5204 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n4609), .ZN(n4618)
         );
  AOI22_X1 U5205 ( .A1(n4079), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5206 ( .A1(n3637), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4615) );
  AOI22_X1 U5207 ( .A1(n4797), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4614) );
  AOI22_X1 U5208 ( .A1(n4950), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4613) );
  NAND4_X1 U5209 ( .A1(n4616), .A2(n4615), .A3(n4614), .A4(n4613), .ZN(n4617)
         );
  NOR2_X1 U5210 ( .A1(n4618), .A2(n4617), .ZN(n4622) );
  XNOR2_X1 U5211 ( .A(n4623), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6267)
         );
  NAND2_X1 U5212 ( .A1(n6267), .A2(n5013), .ZN(n4621) );
  AOI22_X1 U5213 ( .A1(n4995), .A2(EAX_REG_11__SCAN_IN), .B1(n4994), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4620) );
  OAI211_X1 U5214 ( .C1(n4622), .C2(n4686), .A(n4621), .B(n4620), .ZN(n6196)
         );
  XOR2_X1 U5215 ( .A(n7555), .B(n4651), .Z(n7564) );
  NAND2_X1 U5216 ( .A1(n7564), .A2(n4543), .ZN(n4639) );
  INV_X1 U5217 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4625) );
  OAI21_X1 U5218 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n7696), .A(n7669), 
        .ZN(n4624) );
  OAI21_X1 U5219 ( .B1(n4721), .B2(n4625), .A(n4624), .ZN(n4638) );
  AOI22_X1 U5220 ( .A1(n4978), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U5221 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4977), .B1(n4950), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5222 ( .A1(n4908), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4627) );
  AOI22_X1 U5223 ( .A1(n4979), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4626) );
  NAND4_X1 U5224 ( .A1(n4629), .A2(n4628), .A3(n4627), .A4(n4626), .ZN(n4635)
         );
  AOI22_X1 U5225 ( .A1(n3673), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5226 ( .A1(n4079), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4632) );
  AOI22_X1 U5227 ( .A1(n3637), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4631) );
  AOI22_X1 U5228 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3666), .B1(n3663), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4630) );
  NAND4_X1 U5229 ( .A1(n4633), .A2(n4632), .A3(n4631), .A4(n4630), .ZN(n4634)
         );
  NOR2_X1 U5230 ( .A1(n4635), .A2(n4634), .ZN(n4636) );
  NOR2_X1 U5231 ( .A1(n4686), .A2(n4636), .ZN(n4637) );
  AOI21_X1 U5232 ( .B1(n4639), .B2(n4638), .A(n4637), .ZN(n6241) );
  AOI22_X1 U5233 ( .A1(n4978), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4643) );
  AOI22_X1 U5234 ( .A1(n4977), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4642) );
  AOI22_X1 U5235 ( .A1(n4908), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4641) );
  AOI22_X1 U5236 ( .A1(n3666), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4640) );
  NAND4_X1 U5237 ( .A1(n4643), .A2(n4642), .A3(n4641), .A4(n4640), .ZN(n4649)
         );
  AOI22_X1 U5238 ( .A1(n3637), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4647) );
  AOI22_X1 U5239 ( .A1(n4979), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4646) );
  AOI22_X1 U5240 ( .A1(n3673), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4645) );
  AOI22_X1 U5241 ( .A1(n4079), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4644) );
  NAND4_X1 U5242 ( .A1(n4647), .A2(n4646), .A3(n4645), .A4(n4644), .ZN(n4648)
         );
  OR2_X1 U5243 ( .A1(n4649), .A2(n4648), .ZN(n4650) );
  XNOR2_X1 U5244 ( .A(n6240), .B(n3695), .ZN(n6272) );
  XNOR2_X1 U5245 ( .A(n4666), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6297)
         );
  INV_X1 U5246 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7283) );
  INV_X1 U5247 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6281) );
  OAI22_X1 U5248 ( .A1(n4721), .A2(n7283), .B1(n4850), .B2(n6281), .ZN(n4652)
         );
  AOI21_X1 U5249 ( .B1(n6297), .B2(n5013), .A(n4652), .ZN(n6273) );
  INV_X1 U5250 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4670) );
  AOI22_X1 U5251 ( .A1(n4977), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5252 ( .A1(n3672), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4656) );
  AOI22_X1 U5253 ( .A1(n3673), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5254 ( .A1(n3666), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4654) );
  NAND4_X1 U5255 ( .A1(n4657), .A2(n4656), .A3(n4655), .A4(n4654), .ZN(n4663)
         );
  AOI22_X1 U5256 ( .A1(n3637), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5257 ( .A1(n4978), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4660) );
  AOI22_X1 U5258 ( .A1(n4979), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5259 ( .A1(n4079), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4658) );
  NAND4_X1 U5260 ( .A1(n4661), .A2(n4660), .A3(n4659), .A4(n4658), .ZN(n4662)
         );
  OR2_X1 U5261 ( .A1(n4663), .A2(n4662), .ZN(n4664) );
  NAND2_X1 U5262 ( .A1(n4665), .A2(n4664), .ZN(n4669) );
  INV_X1 U5263 ( .A(n4671), .ZN(n4667) );
  XNOR2_X1 U5264 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4667), .ZN(n6346)
         );
  AOI22_X1 U5265 ( .A1(n4543), .A2(n6346), .B1(n4994), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4668) );
  OAI211_X1 U5266 ( .C1(n4721), .C2(n4670), .A(n4669), .B(n4668), .ZN(n6304)
         );
  NAND2_X1 U5267 ( .A1(n6302), .A2(n6304), .ZN(n6303) );
  XOR2_X1 U5268 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4688), .Z(n7568) );
  INV_X1 U5269 ( .A(n7568), .ZN(n7063) );
  AOI22_X1 U5270 ( .A1(n4074), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4675) );
  AOI22_X1 U5271 ( .A1(n4977), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5272 ( .A1(n4979), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5273 ( .A1(n3673), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4672) );
  NAND4_X1 U5274 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4682)
         );
  AOI22_X1 U5275 ( .A1(n4079), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U5276 ( .A1(n4978), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4679) );
  AOI22_X1 U5277 ( .A1(n3637), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5278 ( .A1(n4950), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4677) );
  NAND4_X1 U5279 ( .A1(n4680), .A2(n4679), .A3(n4678), .A4(n4677), .ZN(n4681)
         );
  NOR2_X1 U5280 ( .A1(n4682), .A2(n4681), .ZN(n4685) );
  NAND2_X1 U5281 ( .A1(n4995), .A2(EAX_REG_15__SCAN_IN), .ZN(n4684) );
  NAND2_X1 U5282 ( .A1(n4994), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4683)
         );
  OAI211_X1 U5283 ( .C1(n4686), .C2(n4685), .A(n4684), .B(n4683), .ZN(n4687)
         );
  AOI21_X1 U5284 ( .B1(n7063), .B2(n5013), .A(n4687), .ZN(n6337) );
  XNOR2_X1 U5285 ( .A(n4705), .B(n6357), .ZN(n7054) );
  NAND2_X1 U5286 ( .A1(n7054), .A2(n5013), .ZN(n4704) );
  AOI22_X1 U5287 ( .A1(n4079), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4979), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4693) );
  AOI22_X1 U5288 ( .A1(n3637), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4692) );
  AOI22_X1 U5289 ( .A1(n4977), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4691) );
  AOI22_X1 U5290 ( .A1(n3673), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4690) );
  NAND4_X1 U5291 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4699)
         );
  AOI22_X1 U5292 ( .A1(n4978), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U5293 ( .A1(n4950), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4696) );
  AOI22_X1 U5294 ( .A1(n4797), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4695) );
  AOI22_X1 U5295 ( .A1(n3666), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4694) );
  NAND4_X1 U5296 ( .A1(n4697), .A2(n4696), .A3(n4695), .A4(n4694), .ZN(n4698)
         );
  OR2_X1 U5297 ( .A1(n4699), .A2(n4698), .ZN(n4702) );
  INV_X1 U5298 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4700) );
  OAI22_X1 U5299 ( .A1(n4721), .A2(n4700), .B1(n6357), .B2(n4850), .ZN(n4701)
         );
  AOI21_X1 U5300 ( .B1(n4991), .B2(n4702), .A(n4701), .ZN(n4703) );
  NAND2_X1 U5301 ( .A1(n4704), .A2(n4703), .ZN(n6352) );
  NAND2_X1 U5302 ( .A1(n6336), .A2(n6352), .ZN(n6351) );
  INV_X1 U5303 ( .A(n6351), .ZN(n4725) );
  OR2_X1 U5304 ( .A1(n4706), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4707)
         );
  NAND2_X1 U5305 ( .A1(n4741), .A2(n4707), .ZN(n7049) );
  AOI22_X1 U5306 ( .A1(n4978), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U5307 ( .A1(n4977), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4710) );
  AOI22_X1 U5308 ( .A1(n4950), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4709) );
  AOI22_X1 U5309 ( .A1(n3637), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4708) );
  NAND4_X1 U5310 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n4717)
         );
  AOI22_X1 U5311 ( .A1(n3673), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4715) );
  AOI22_X1 U5312 ( .A1(n4979), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4714) );
  AOI22_X1 U5313 ( .A1(n3674), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5314 ( .A1(n4079), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4712) );
  NAND4_X1 U5315 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4716)
         );
  NOR2_X1 U5316 ( .A1(n4717), .A2(n4716), .ZN(n4718) );
  NOR2_X1 U5317 ( .A1(n4964), .A2(n4718), .ZN(n4723) );
  INV_X1 U5318 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U5319 ( .A1(n7669), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4719)
         );
  OAI211_X1 U5320 ( .C1(n4721), .C2(n4720), .A(n4967), .B(n4719), .ZN(n4722)
         );
  OAI22_X1 U5321 ( .A1(n7049), .A2(n4967), .B1(n4723), .B2(n4722), .ZN(n6505)
         );
  XNOR2_X1 U5322 ( .A(n4741), .B(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n7037)
         );
  NAND2_X1 U5323 ( .A1(n7037), .A2(n4543), .ZN(n4740) );
  AOI22_X1 U5324 ( .A1(n4079), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4729) );
  AOI22_X1 U5325 ( .A1(n3673), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4728) );
  AOI22_X1 U5326 ( .A1(n3674), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4727) );
  AOI22_X1 U5327 ( .A1(n4979), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4726) );
  NAND4_X1 U5328 ( .A1(n4729), .A2(n4728), .A3(n4727), .A4(n4726), .ZN(n4735)
         );
  AOI22_X1 U5329 ( .A1(n4977), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5330 ( .A1(n4978), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5331 ( .A1(n4950), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4731) );
  AOI22_X1 U5332 ( .A1(n3637), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4730) );
  NAND4_X1 U5333 ( .A1(n4733), .A2(n4732), .A3(n4731), .A4(n4730), .ZN(n4734)
         );
  NOR2_X1 U5334 ( .A1(n4735), .A2(n4734), .ZN(n4738) );
  OAI21_X1 U5335 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7034), .A(n4967), .ZN(
        n4736) );
  AOI21_X1 U5336 ( .B1(n4995), .B2(EAX_REG_18__SCAN_IN), .A(n4736), .ZN(n4737)
         );
  OAI21_X1 U5337 ( .B1(n4964), .B2(n4738), .A(n4737), .ZN(n4739) );
  AND2_X1 U5338 ( .A1(n4742), .A2(n4754), .ZN(n4743) );
  OR2_X1 U5339 ( .A1(n4743), .A2(n4775), .ZN(n7580) );
  AOI22_X1 U5340 ( .A1(n4079), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4747) );
  AOI22_X1 U5341 ( .A1(n4977), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4746) );
  AOI22_X1 U5342 ( .A1(n4074), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4745) );
  AOI22_X1 U5343 ( .A1(n3673), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4744) );
  NAND4_X1 U5344 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n4753)
         );
  AOI22_X1 U5345 ( .A1(n4978), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4751) );
  AOI22_X1 U5346 ( .A1(n4979), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4750) );
  AOI22_X1 U5347 ( .A1(n3666), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4749) );
  AOI22_X1 U5348 ( .A1(n7224), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4748) );
  NAND4_X1 U5349 ( .A1(n4751), .A2(n4750), .A3(n4749), .A4(n4748), .ZN(n4752)
         );
  NOR2_X1 U5350 ( .A1(n4753), .A2(n4752), .ZN(n4757) );
  OAI21_X1 U5351 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4754), .A(n4967), .ZN(
        n4755) );
  AOI21_X1 U5352 ( .B1(n4995), .B2(EAX_REG_19__SCAN_IN), .A(n4755), .ZN(n4756)
         );
  OAI21_X1 U5353 ( .B1(n4964), .B2(n4757), .A(n4756), .ZN(n4758) );
  OAI21_X1 U5354 ( .B1(n7580), .B2(n4967), .A(n4758), .ZN(n7025) );
  AND2_X2 U5355 ( .A1(n6497), .A2(n4759), .ZN(n6532) );
  INV_X1 U5356 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n7602) );
  XNOR2_X1 U5357 ( .A(n4775), .B(n7602), .ZN(n7592) );
  AOI22_X1 U5358 ( .A1(n4978), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4763) );
  AOI22_X1 U5359 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4977), .B1(n4950), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4762) );
  AOI22_X1 U5360 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4908), .B1(n3674), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4761) );
  AOI22_X1 U5361 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3666), .B1(n3664), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4760) );
  NAND4_X1 U5362 ( .A1(n4763), .A2(n4762), .A3(n4761), .A4(n4760), .ZN(n4769)
         );
  AOI22_X1 U5363 ( .A1(n3637), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4767) );
  AOI22_X1 U5364 ( .A1(n4979), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4766) );
  AOI22_X1 U5365 ( .A1(n3673), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5366 ( .A1(n4079), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4764) );
  NAND4_X1 U5367 ( .A1(n4767), .A2(n4766), .A3(n4765), .A4(n4764), .ZN(n4768)
         );
  OR2_X1 U5368 ( .A1(n4769), .A2(n4768), .ZN(n4773) );
  INV_X1 U5369 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4771) );
  OAI21_X1 U5370 ( .B1(n7696), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n7669), 
        .ZN(n4770) );
  OAI21_X1 U5371 ( .B1(n4721), .B2(n4771), .A(n4770), .ZN(n4772) );
  AOI21_X1 U5372 ( .B1(n4991), .B2(n4773), .A(n4772), .ZN(n4774) );
  AOI21_X1 U5373 ( .B1(n7592), .B2(n5013), .A(n4774), .ZN(n6535) );
  OR2_X1 U5374 ( .A1(n4776), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4777)
         );
  NAND2_X1 U5375 ( .A1(n4810), .A2(n4777), .ZN(n7605) );
  AOI22_X1 U5376 ( .A1(n4079), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5377 ( .A1(n4978), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4780) );
  AOI22_X1 U5378 ( .A1(n4977), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4779) );
  AOI22_X1 U5379 ( .A1(n4979), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4778) );
  NAND4_X1 U5380 ( .A1(n4781), .A2(n4780), .A3(n4779), .A4(n4778), .ZN(n4787)
         );
  AOI22_X1 U5381 ( .A1(n3672), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5382 ( .A1(n7224), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4784) );
  AOI22_X1 U5383 ( .A1(n3673), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4783) );
  AOI22_X1 U5384 ( .A1(n4950), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4782) );
  NAND4_X1 U5385 ( .A1(n4785), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(n4786)
         );
  NOR2_X1 U5386 ( .A1(n4787), .A2(n4786), .ZN(n4790) );
  OAI21_X1 U5387 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n7696), .A(n7669), 
        .ZN(n4789) );
  NAND2_X1 U5388 ( .A1(n4995), .A2(EAX_REG_21__SCAN_IN), .ZN(n4788) );
  OAI211_X1 U5389 ( .C1(n4964), .C2(n4790), .A(n4789), .B(n4788), .ZN(n4791)
         );
  NAND2_X1 U5390 ( .A1(n4792), .A2(n4791), .ZN(n7006) );
  XNOR2_X1 U5391 ( .A(n4810), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n7003)
         );
  NAND2_X1 U5392 ( .A1(n7003), .A2(n5013), .ZN(n4808) );
  AOI22_X1 U5393 ( .A1(n4978), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4796) );
  AOI22_X1 U5394 ( .A1(n4977), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U5395 ( .A1(n4908), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4794) );
  AOI22_X1 U5396 ( .A1(n3666), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4793) );
  NAND4_X1 U5397 ( .A1(n4796), .A2(n4795), .A3(n4794), .A4(n4793), .ZN(n4803)
         );
  AOI22_X1 U5398 ( .A1(n3637), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4801) );
  AOI22_X1 U5399 ( .A1(n4979), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4800) );
  AOI22_X1 U5400 ( .A1(n3673), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4799) );
  AOI22_X1 U5401 ( .A1(n4079), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4798) );
  NAND4_X1 U5402 ( .A1(n4801), .A2(n4800), .A3(n4799), .A4(n4798), .ZN(n4802)
         );
  NOR2_X1 U5403 ( .A1(n4803), .A2(n4802), .ZN(n4806) );
  INV_X1 U5404 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n7001) );
  AOI21_X1 U5405 ( .B1(n7001), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4804) );
  AOI21_X1 U5406 ( .B1(n4995), .B2(EAX_REG_22__SCAN_IN), .A(n4804), .ZN(n4805)
         );
  OAI21_X1 U5407 ( .B1(n4964), .B2(n4806), .A(n4805), .ZN(n4807) );
  NAND2_X1 U5408 ( .A1(n4808), .A2(n4807), .ZN(n6486) );
  INV_X1 U5409 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U5410 ( .A1(n4811), .A2(n6476), .ZN(n4812) );
  NAND2_X1 U5411 ( .A1(n4857), .A2(n4812), .ZN(n6994) );
  AOI22_X1 U5412 ( .A1(n3637), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4816) );
  AOI22_X1 U5413 ( .A1(n4977), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4815) );
  AOI22_X1 U5414 ( .A1(n4079), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4814) );
  AOI22_X1 U5415 ( .A1(n4950), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4813) );
  NAND4_X1 U5416 ( .A1(n4816), .A2(n4815), .A3(n4814), .A4(n4813), .ZN(n4822)
         );
  AOI22_X1 U5417 ( .A1(n4978), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4820) );
  AOI22_X1 U5418 ( .A1(n4908), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4819) );
  AOI22_X1 U5419 ( .A1(n4979), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3642), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4818) );
  AOI22_X1 U5420 ( .A1(n7224), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4817) );
  NAND4_X1 U5421 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .ZN(n4821)
         );
  NOR2_X1 U5422 ( .A1(n4822), .A2(n4821), .ZN(n4839) );
  AOI22_X1 U5423 ( .A1(n4978), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4826) );
  AOI22_X1 U5424 ( .A1(n4977), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4825) );
  AOI22_X1 U5425 ( .A1(n3637), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4824) );
  AOI22_X1 U5426 ( .A1(n3673), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4823) );
  NAND4_X1 U5427 ( .A1(n4826), .A2(n4825), .A3(n4824), .A4(n4823), .ZN(n4832)
         );
  AOI22_X1 U5428 ( .A1(n4079), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4830) );
  AOI22_X1 U5429 ( .A1(n3672), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U5430 ( .A1(n4979), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4828) );
  AOI22_X1 U5431 ( .A1(n4950), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4827) );
  NAND4_X1 U5432 ( .A1(n4830), .A2(n4829), .A3(n4828), .A4(n4827), .ZN(n4831)
         );
  NOR2_X1 U5433 ( .A1(n4832), .A2(n4831), .ZN(n4838) );
  XNOR2_X1 U5434 ( .A(n4839), .B(n4838), .ZN(n4835) );
  AOI21_X1 U5435 ( .B1(n6476), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4833) );
  AOI21_X1 U5436 ( .B1(n4995), .B2(EAX_REG_23__SCAN_IN), .A(n4833), .ZN(n4834)
         );
  OAI21_X1 U5437 ( .B1(n4964), .B2(n4835), .A(n4834), .ZN(n4836) );
  OAI21_X1 U5438 ( .B1(n6994), .B2(n4967), .A(n4836), .ZN(n6475) );
  INV_X1 U5439 ( .A(n6475), .ZN(n4837) );
  INV_X1 U5440 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4856) );
  XNOR2_X1 U5441 ( .A(n4857), .B(n4856), .ZN(n6985) );
  NAND2_X1 U5442 ( .A1(n6985), .A2(n5013), .ZN(n4855) );
  OR2_X1 U5443 ( .A1(n4839), .A2(n4838), .ZN(n4864) );
  AOI22_X1 U5444 ( .A1(n3637), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4978), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4843) );
  AOI22_X1 U5445 ( .A1(n7224), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4842) );
  AOI22_X1 U5446 ( .A1(n3673), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4841) );
  AOI22_X1 U5447 ( .A1(n4979), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4840) );
  NAND4_X1 U5448 ( .A1(n4843), .A2(n4842), .A3(n4841), .A4(n4840), .ZN(n4849)
         );
  AOI22_X1 U5449 ( .A1(n4977), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4847) );
  AOI22_X1 U5450 ( .A1(n4950), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4846) );
  AOI22_X1 U5451 ( .A1(n4079), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4845) );
  AOI22_X1 U5452 ( .A1(n4074), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4844) );
  NAND4_X1 U5453 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n4848)
         );
  XNOR2_X1 U5454 ( .A(n4864), .B(n4862), .ZN(n4853) );
  INV_X1 U5455 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4851) );
  OAI22_X1 U5456 ( .A1(n4721), .A2(n4851), .B1(n4856), .B2(n4850), .ZN(n4852)
         );
  AOI21_X1 U5457 ( .B1(n4991), .B2(n4853), .A(n4852), .ZN(n4854) );
  NAND2_X1 U5458 ( .A1(n4855), .A2(n4854), .ZN(n6461) );
  INV_X1 U5459 ( .A(n4858), .ZN(n4860) );
  INV_X1 U5460 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4859) );
  NAND2_X1 U5461 ( .A1(n4860), .A2(n4859), .ZN(n4861) );
  NAND2_X1 U5462 ( .A1(n4900), .A2(n4861), .ZN(n6976) );
  INV_X1 U5463 ( .A(n4862), .ZN(n4863) );
  AOI22_X1 U5464 ( .A1(n4079), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4868) );
  AOI22_X1 U5465 ( .A1(n4978), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4867) );
  AOI22_X1 U5466 ( .A1(n4977), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4866) );
  AOI22_X1 U5467 ( .A1(n4950), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4865) );
  NAND4_X1 U5468 ( .A1(n4868), .A2(n4867), .A3(n4866), .A4(n4865), .ZN(n4874)
         );
  AOI22_X1 U5469 ( .A1(n3674), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4872) );
  AOI22_X1 U5470 ( .A1(n4979), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3642), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4871) );
  AOI22_X1 U5471 ( .A1(n3672), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4870) );
  AOI22_X1 U5472 ( .A1(n7224), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4869) );
  NAND4_X1 U5473 ( .A1(n4872), .A2(n4871), .A3(n4870), .A4(n4869), .ZN(n4873)
         );
  NOR2_X1 U5474 ( .A1(n4874), .A2(n4873), .ZN(n4882) );
  XNOR2_X1 U5475 ( .A(n4881), .B(n4882), .ZN(n4878) );
  NAND2_X1 U5476 ( .A1(n7669), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4875)
         );
  NAND2_X1 U5477 ( .A1(n4967), .A2(n4875), .ZN(n4876) );
  AOI21_X1 U5478 ( .B1(n4995), .B2(EAX_REG_25__SCAN_IN), .A(n4876), .ZN(n4877)
         );
  OAI21_X1 U5479 ( .B1(n4878), .B2(n4964), .A(n4877), .ZN(n4879) );
  NAND2_X1 U5480 ( .A1(n4880), .A2(n4879), .ZN(n6450) );
  XNOR2_X1 U5481 ( .A(n4900), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6442)
         );
  NAND2_X1 U5482 ( .A1(n6442), .A2(n4543), .ZN(n4898) );
  NOR2_X1 U5483 ( .A1(n4882), .A2(n4881), .ZN(n4907) );
  AOI22_X1 U5484 ( .A1(n4978), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4886) );
  AOI22_X1 U5485 ( .A1(n4977), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4885) );
  AOI22_X1 U5486 ( .A1(n4908), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4884) );
  AOI22_X1 U5487 ( .A1(n3666), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4909), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4883) );
  NAND4_X1 U5488 ( .A1(n4886), .A2(n4885), .A3(n4884), .A4(n4883), .ZN(n4892)
         );
  AOI22_X1 U5489 ( .A1(n3637), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4890) );
  AOI22_X1 U5490 ( .A1(n4979), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4889) );
  AOI22_X1 U5491 ( .A1(n3673), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4888) );
  AOI22_X1 U5492 ( .A1(n4079), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4887) );
  NAND4_X1 U5493 ( .A1(n4890), .A2(n4889), .A3(n4888), .A4(n4887), .ZN(n4891)
         );
  OR2_X1 U5494 ( .A1(n4892), .A2(n4891), .ZN(n4906) );
  XNOR2_X1 U5495 ( .A(n4907), .B(n4906), .ZN(n4896) );
  INV_X1 U5496 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4893) );
  AOI21_X1 U5497 ( .B1(n4893), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4894) );
  AOI21_X1 U5498 ( .B1(n4995), .B2(EAX_REG_26__SCAN_IN), .A(n4894), .ZN(n4895)
         );
  OAI21_X1 U5499 ( .B1(n4896), .B2(n4964), .A(n4895), .ZN(n4897) );
  INV_X1 U5500 ( .A(n4900), .ZN(n4901) );
  INV_X1 U5501 ( .A(n4902), .ZN(n4904) );
  INV_X1 U5502 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4903) );
  NAND2_X1 U5503 ( .A1(n4904), .A2(n4903), .ZN(n4905) );
  NAND2_X1 U5504 ( .A1(n4943), .A2(n4905), .ZN(n6958) );
  NAND2_X1 U5505 ( .A1(n4907), .A2(n4906), .ZN(n4938) );
  AOI22_X1 U5506 ( .A1(n3637), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4913) );
  AOI22_X1 U5507 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4978), .B1(n3674), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4912) );
  AOI22_X1 U5508 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4977), .B1(n4908), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4911) );
  AOI22_X1 U5509 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4950), .B1(n3664), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4910) );
  NAND4_X1 U5510 ( .A1(n4913), .A2(n4912), .A3(n4911), .A4(n4910), .ZN(n4919)
         );
  AOI22_X1 U5511 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4074), .B1(n3666), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4917) );
  AOI22_X1 U5512 ( .A1(n4979), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4797), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4916) );
  AOI22_X1 U5513 ( .A1(n7224), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4915) );
  AOI22_X1 U5514 ( .A1(n4079), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4914) );
  NAND4_X1 U5515 ( .A1(n4917), .A2(n4916), .A3(n4915), .A4(n4914), .ZN(n4918)
         );
  NOR2_X1 U5516 ( .A1(n4919), .A2(n4918), .ZN(n4939) );
  XNOR2_X1 U5517 ( .A(n4938), .B(n4939), .ZN(n4923) );
  NAND2_X1 U5518 ( .A1(n7669), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4920)
         );
  NAND2_X1 U5519 ( .A1(n4967), .A2(n4920), .ZN(n4921) );
  AOI21_X1 U5520 ( .B1(n4995), .B2(EAX_REG_27__SCAN_IN), .A(n4921), .ZN(n4922)
         );
  OAI21_X1 U5521 ( .B1(n4923), .B2(n4964), .A(n4922), .ZN(n4924) );
  XNOR2_X1 U5522 ( .A(n4943), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6415)
         );
  INV_X1 U5523 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4926) );
  AOI21_X1 U5524 ( .B1(n4926), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4927) );
  AOI21_X1 U5525 ( .B1(n4995), .B2(EAX_REG_28__SCAN_IN), .A(n4927), .ZN(n4942)
         );
  AOI22_X1 U5526 ( .A1(n4978), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4931) );
  AOI22_X1 U5527 ( .A1(n4977), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4930) );
  AOI22_X1 U5528 ( .A1(n4971), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4929) );
  AOI22_X1 U5529 ( .A1(n3666), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4928) );
  NAND4_X1 U5530 ( .A1(n4931), .A2(n4930), .A3(n4929), .A4(n4928), .ZN(n4937)
         );
  AOI22_X1 U5531 ( .A1(n3637), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4935) );
  AOI22_X1 U5532 ( .A1(n4979), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4934) );
  AOI22_X1 U5533 ( .A1(n3673), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4933) );
  AOI22_X1 U5534 ( .A1(n4079), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4932) );
  NAND4_X1 U5535 ( .A1(n4935), .A2(n4934), .A3(n4933), .A4(n4932), .ZN(n4936)
         );
  OR2_X1 U5536 ( .A1(n4937), .A2(n4936), .ZN(n4948) );
  NOR2_X1 U5537 ( .A1(n4939), .A2(n4938), .ZN(n4949) );
  XOR2_X1 U5538 ( .A(n4948), .B(n4949), .Z(n4940) );
  NAND2_X1 U5539 ( .A1(n4940), .A2(n4991), .ZN(n4941) );
  INV_X1 U5540 ( .A(n4943), .ZN(n4944) );
  NAND2_X1 U5541 ( .A1(n4944), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4946)
         );
  INV_X1 U5542 ( .A(n4946), .ZN(n4947) );
  INV_X1 U5543 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4945) );
  OAI21_X1 U5544 ( .B1(n4947), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5000), 
        .ZN(n6948) );
  NAND2_X1 U5545 ( .A1(n4949), .A2(n4948), .ZN(n4968) );
  AOI22_X1 U5546 ( .A1(n3637), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4954) );
  AOI22_X1 U5547 ( .A1(n4977), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4908), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U5548 ( .A1(n4950), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4952) );
  AOI22_X1 U5549 ( .A1(n4079), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3642), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4951) );
  NAND4_X1 U5550 ( .A1(n4954), .A2(n4953), .A3(n4952), .A4(n4951), .ZN(n4961)
         );
  AOI22_X1 U5551 ( .A1(n4978), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4959) );
  AOI22_X1 U5552 ( .A1(n7224), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4958) );
  AOI22_X1 U5553 ( .A1(n3674), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U5554 ( .A1(n4979), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4956) );
  NAND4_X1 U5555 ( .A1(n4959), .A2(n4958), .A3(n4957), .A4(n4956), .ZN(n4960)
         );
  NOR2_X1 U5556 ( .A1(n4961), .A2(n4960), .ZN(n4969) );
  XNOR2_X1 U5557 ( .A(n4968), .B(n4969), .ZN(n4965) );
  AOI21_X1 U5558 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n7669), .A(n5013), 
        .ZN(n4963) );
  NAND2_X1 U5559 ( .A1(n4995), .A2(EAX_REG_29__SCAN_IN), .ZN(n4962) );
  OAI211_X1 U5560 ( .C1(n4965), .C2(n4964), .A(n4963), .B(n4962), .ZN(n4966)
         );
  OAI21_X1 U5561 ( .B1(n6948), .B2(n4967), .A(n4966), .ZN(n6403) );
  XNOR2_X1 U5562 ( .A(n5000), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6382)
         );
  NOR2_X1 U5563 ( .A1(n4969), .A2(n4968), .ZN(n4987) );
  AOI22_X1 U5564 ( .A1(n3673), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4976) );
  AOI22_X1 U5565 ( .A1(n4971), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4975) );
  AOI22_X1 U5566 ( .A1(n4079), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4974) );
  AOI22_X1 U5567 ( .A1(n3637), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4972), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4973) );
  NAND4_X1 U5568 ( .A1(n4976), .A2(n4975), .A3(n4974), .A4(n4973), .ZN(n4985)
         );
  AOI22_X1 U5569 ( .A1(n4977), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4950), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4983) );
  AOI22_X1 U5570 ( .A1(n4978), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n7224), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4982) );
  AOI22_X1 U5571 ( .A1(n4979), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4955), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4981) );
  AOI22_X1 U5572 ( .A1(n3666), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4980) );
  NAND4_X1 U5573 ( .A1(n4983), .A2(n4982), .A3(n4981), .A4(n4980), .ZN(n4984)
         );
  NOR2_X1 U5574 ( .A1(n4985), .A2(n4984), .ZN(n4986) );
  XNOR2_X1 U5575 ( .A(n4987), .B(n4986), .ZN(n4992) );
  INV_X1 U5576 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4989) );
  OAI21_X1 U5577 ( .B1(n7696), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n7669), 
        .ZN(n4988) );
  OAI21_X1 U5578 ( .B1(n4721), .B2(n4989), .A(n4988), .ZN(n4990) );
  AOI21_X1 U5579 ( .B1(n4992), .B2(n4991), .A(n4990), .ZN(n4993) );
  NAND2_X1 U5580 ( .A1(n6402), .A2(n5069), .ZN(n4998) );
  AOI22_X1 U5581 ( .A1(n4995), .A2(EAX_REG_31__SCAN_IN), .B1(n4994), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4996) );
  INV_X1 U5582 ( .A(n4996), .ZN(n4997) );
  XNOR2_X2 U5583 ( .A(n4998), .B(n4997), .ZN(n6394) );
  NAND2_X1 U5584 ( .A1(n7691), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5168) );
  INV_X1 U5585 ( .A(n5168), .ZN(n5012) );
  NAND2_X1 U5586 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5012), .ZN(n7423) );
  INV_X1 U5587 ( .A(n7423), .ZN(n4999) );
  NAND2_X1 U5588 ( .A1(n6394), .A2(n7392), .ZN(n5010) );
  INV_X1 U5589 ( .A(n5000), .ZN(n5001) );
  NAND2_X1 U5590 ( .A1(n5001), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5002)
         );
  INV_X1 U5591 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U5592 ( .A1(n5679), .A2(n5003), .ZN(n7426) );
  NAND2_X1 U5593 ( .A1(n7426), .A2(n7691), .ZN(n5004) );
  NAND2_X1 U5594 ( .A1(n7691), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U5595 ( .A1(n7696), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U5596 ( .A1(n5006), .A2(n5005), .ZN(n5110) );
  NAND2_X2 U5597 ( .A1(n7035), .A2(n5110), .ZN(n7405) );
  INV_X1 U5598 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7341) );
  NOR2_X1 U5599 ( .A1(n7477), .A2(n7341), .ZN(n7071) );
  AOI21_X1 U5600 ( .B1(n7396), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n7071), 
        .ZN(n5007) );
  OAI21_X1 U5601 ( .B1(n5785), .B2(n7405), .A(n5007), .ZN(n5008) );
  OAI211_X1 U5602 ( .C1(n7076), .C2(n7626), .A(n5010), .B(n5009), .ZN(U2955)
         );
  NOR2_X1 U5603 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n7432) );
  NAND2_X1 U5604 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n7432), .ZN(n7692) );
  NOR2_X1 U5605 ( .A1(n7691), .A2(n7692), .ZN(n7683) );
  AND2_X1 U5606 ( .A1(n5013), .A2(n5012), .ZN(n7676) );
  INV_X1 U5607 ( .A(n7676), .ZN(n5014) );
  NAND2_X1 U5608 ( .A1(n7477), .A2(n5014), .ZN(n5015) );
  OR2_X1 U5609 ( .A1(n7501), .A2(n7422), .ZN(n5783) );
  NAND2_X1 U5610 ( .A1(n6394), .A2(n7611), .ZN(n5045) );
  NAND2_X1 U5611 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n6356) );
  NAND2_X1 U5612 ( .A1(n7696), .A2(n7709), .ZN(n5779) );
  INV_X1 U5613 ( .A(n5779), .ZN(n5017) );
  AND3_X1 U5614 ( .A1(n5018), .A2(n4017), .A3(n5017), .ZN(n5019) );
  INV_X1 U5615 ( .A(n7501), .ZN(n5853) );
  INV_X1 U5616 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7313) );
  INV_X1 U5617 ( .A(REIP_REG_1__SCAN_IN), .ZN(n7506) );
  INV_X1 U5618 ( .A(REIP_REG_2__SCAN_IN), .ZN(n7507) );
  INV_X1 U5619 ( .A(REIP_REG_5__SCAN_IN), .ZN(n7293) );
  NAND4_X1 U5620 ( .A1(n5930), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .A4(REIP_REG_8__SCAN_IN), .ZN(n5778) );
  INV_X1 U5621 ( .A(REIP_REG_9__SCAN_IN), .ZN(n7300) );
  INV_X1 U5622 ( .A(REIP_REG_10__SCAN_IN), .ZN(n7302) );
  NOR3_X2 U5623 ( .A1(n5778), .A2(n7300), .A3(n7302), .ZN(n6231) );
  NAND2_X1 U5624 ( .A1(n6231), .A2(REIP_REG_11__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U5625 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n6305) );
  INV_X1 U5626 ( .A(REIP_REG_14__SCAN_IN), .ZN(n7308) );
  INV_X1 U5627 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7314) );
  INV_X1 U5628 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7319) );
  NOR3_X1 U5629 ( .A1(n7586), .A2(n7314), .A3(n7319), .ZN(n5020) );
  NAND2_X1 U5630 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5021) );
  INV_X1 U5631 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7325) );
  OAI21_X1 U5632 ( .B1(n5021), .B2(n7325), .A(n6230), .ZN(n5022) );
  AND2_X1 U5633 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5041) );
  INV_X1 U5634 ( .A(n5041), .ZN(n5023) );
  INV_X1 U5635 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7331) );
  NOR2_X1 U5636 ( .A1(n5023), .A2(n7331), .ZN(n5024) );
  NAND2_X1 U5637 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5025) );
  INV_X1 U5638 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7338) );
  NOR2_X1 U5639 ( .A1(n7339), .A2(n7338), .ZN(n5026) );
  NOR2_X1 U5640 ( .A1(n6275), .A2(n5026), .ZN(n5027) );
  NAND2_X1 U5641 ( .A1(n6388), .A2(REIP_REG_31__SCAN_IN), .ZN(n5044) );
  OAI21_X1 U5642 ( .B1(n6404), .B2(n5029), .A(n5028), .ZN(n5032) );
  AOI22_X1 U5643 ( .A1(n5228), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5030), .ZN(n5031) );
  XNOR2_X1 U5644 ( .A(n5032), .B(n5031), .ZN(n7073) );
  NAND3_X1 U5645 ( .A1(n5191), .A2(EBX_REG_31__SCAN_IN), .A3(n5779), .ZN(n5033) );
  INV_X1 U5646 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5034) );
  NOR2_X1 U5647 ( .A1(n7428), .A2(n5779), .ZN(n7665) );
  INV_X1 U5648 ( .A(n7665), .ZN(n5035) );
  NAND2_X1 U5649 ( .A1(n3675), .A2(n5035), .ZN(n5781) );
  INV_X1 U5650 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6518) );
  OR2_X1 U5651 ( .A1(n5781), .A2(n6518), .ZN(n5036) );
  OAI22_X1 U5652 ( .A1(n5037), .A2(n7601), .B1(n5849), .B2(n5036), .ZN(n5038)
         );
  INV_X1 U5653 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7317) );
  NAND3_X1 U5654 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        n7570), .ZN(n6513) );
  NAND2_X1 U5655 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6500), .ZN(n7585) );
  NAND3_X1 U5656 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_23__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5040) );
  NOR2_X2 U5657 ( .A1(n6490), .A2(n5040), .ZN(n6470) );
  NAND2_X1 U5658 ( .A1(n6470), .A2(n5041), .ZN(n6444) );
  NAND2_X1 U5659 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .ZN(
        n5042) );
  OR2_X2 U5660 ( .A1(n6444), .A2(n5042), .ZN(n6414) );
  INV_X1 U5661 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7335) );
  NOR2_X1 U5662 ( .A1(n6414), .A2(n7335), .ZN(n6380) );
  NAND4_X1 U5663 ( .A1(n6380), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n7341), .ZN(n5043) );
  INV_X1 U5664 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U5665 ( .A1(n5059), .A2(n7402), .ZN(n5058) );
  NOR2_X1 U5666 ( .A1(n7477), .A2(n7335), .ZN(n5064) );
  INV_X1 U5667 ( .A(n6415), .ZN(n5053) );
  NOR2_X1 U5668 ( .A1(n5053), .A2(n7405), .ZN(n5054) );
  AOI211_X1 U5669 ( .C1(n7396), .C2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5064), 
        .B(n5054), .ZN(n5055) );
  NAND2_X1 U5670 ( .A1(n5058), .A2(n5057), .ZN(U2958) );
  NAND2_X1 U5671 ( .A1(n5059), .A2(n7488), .ZN(n5068) );
  OR2_X1 U5672 ( .A1(n6428), .A2(n5060), .ZN(n5061) );
  NAND2_X1 U5673 ( .A1(n6406), .A2(n5061), .ZN(n6521) );
  INV_X1 U5674 ( .A(n7077), .ZN(n7094) );
  INV_X1 U5675 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n7089) );
  AOI211_X1 U5676 ( .C1(n7089), .C2(n5062), .A(n7078), .B(n7087), .ZN(n5063)
         );
  AOI211_X1 U5677 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n7094), .A(n5064), .B(n5063), .ZN(n5065) );
  NAND2_X1 U5678 ( .A1(n5068), .A2(n5067), .ZN(U2990) );
  XNOR2_X1 U5679 ( .A(n6402), .B(n5070), .ZN(n6940) );
  NAND2_X1 U5680 ( .A1(n3750), .A2(n7709), .ZN(n5071) );
  OAI22_X1 U5681 ( .A1(n7693), .A2(n5143), .B1(n5072), .B2(n4330), .ZN(n5128)
         );
  INV_X1 U5682 ( .A(n3952), .ZN(n6391) );
  NAND3_X1 U5683 ( .A1(n3662), .A2(n6391), .A3(n5073), .ZN(n5074) );
  NOR2_X1 U5684 ( .A1(n5130), .A2(n5074), .ZN(n5075) );
  NAND2_X1 U5685 ( .A1(n3986), .A2(n3952), .ZN(n5225) );
  NAND2_X2 U5686 ( .A1(n6392), .A2(n5225), .ZN(n6568) );
  NAND2_X1 U5687 ( .A1(n6940), .A2(n3645), .ZN(n5081) );
  AND2_X1 U5688 ( .A1(n3935), .A2(n3952), .ZN(n5077) );
  AOI22_X1 U5689 ( .A1(n7733), .A2(DATAI_14_), .B1(n7735), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5078) );
  INV_X1 U5690 ( .A(n5078), .ZN(n5079) );
  NOR2_X1 U5691 ( .A1(n5079), .A2(n3802), .ZN(n5080) );
  NAND2_X1 U5692 ( .A1(n5081), .A2(n5080), .ZN(U2861) );
  NAND2_X1 U5693 ( .A1(n5417), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5874) );
  OR2_X1 U5694 ( .A1(n5630), .A2(n5874), .ZN(n5590) );
  INV_X1 U5695 ( .A(n5590), .ZN(n5097) );
  NOR2_X1 U5696 ( .A1(n7422), .A2(n7669), .ZN(n7674) );
  NAND2_X1 U5697 ( .A1(n5084), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6397) );
  INV_X1 U5698 ( .A(n6397), .ZN(n5086) );
  AND2_X1 U5699 ( .A1(n5086), .A2(n5085), .ZN(n5465) );
  AOI21_X1 U5700 ( .B1(n4532), .B2(n5465), .A(n5679), .ZN(n5094) );
  AND2_X1 U5701 ( .A1(n3794), .A2(n3667), .ZN(n5595) );
  NOR2_X1 U5702 ( .A1(n5464), .A2(n5874), .ZN(n5102) );
  AOI21_X1 U5703 ( .B1(n5595), .B2(n4509), .A(n5102), .ZN(n5095) );
  NAND2_X1 U5704 ( .A1(n5094), .A2(n5095), .ZN(n5091) );
  OAI211_X1 U5705 ( .C1(n5871), .C2(n5097), .A(n5551), .B(n5091), .ZN(n5259)
         );
  INV_X1 U5706 ( .A(n5259), .ZN(n5093) );
  INV_X1 U5707 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n5092) );
  NOR2_X1 U5708 ( .A1(n5093), .A2(n5092), .ZN(n5106) );
  INV_X1 U5709 ( .A(n5094), .ZN(n5096) );
  OR2_X1 U5710 ( .A1(n5096), .A2(n5095), .ZN(n5099) );
  NAND2_X1 U5711 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5097), .ZN(n5098) );
  INV_X1 U5712 ( .A(DATAI_0_), .ZN(n5226) );
  NOR2_X1 U5713 ( .A1(n5265), .A2(n6024), .ZN(n5105) );
  NAND2_X1 U5714 ( .A1(n5085), .A2(n5084), .ZN(n5471) );
  NOR2_X1 U5715 ( .A1(n5626), .A2(n5471), .ZN(n5100) );
  NAND2_X1 U5716 ( .A1(n5100), .A2(n5552), .ZN(n5585) );
  NAND2_X1 U5717 ( .A1(n7392), .A2(DATAI_24_), .ZN(n6135) );
  NOR2_X1 U5718 ( .A1(n5585), .A2(n6135), .ZN(n5104) );
  AND2_X1 U5719 ( .A1(n7392), .A2(DATAI_16_), .ZN(n6138) );
  INV_X1 U5720 ( .A(n6138), .ZN(n5768) );
  NAND2_X1 U5721 ( .A1(n5260), .A2(n4017), .ZN(n6025) );
  INV_X1 U5722 ( .A(n5102), .ZN(n5261) );
  OAI22_X1 U5723 ( .A1(n5768), .A2(n5839), .B1(n6025), .B2(n5261), .ZN(n5103)
         );
  OR4_X1 U5724 ( .A1(n5106), .A2(n5105), .A3(n5104), .A4(n5103), .ZN(U3108) );
  INV_X1 U5725 ( .A(n5107), .ZN(n5109) );
  INV_X1 U5726 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7718) );
  OAI211_X1 U5727 ( .C1(n5109), .C2(n7718), .A(n5108), .B(n7417), .ZN(U2788)
         );
  OAI21_X1 U5728 ( .B1(n7396), .B2(n5110), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5119) );
  NOR2_X1 U5729 ( .A1(n5111), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5112)
         );
  NOR2_X1 U5730 ( .A1(n5112), .A2(n5218), .ZN(n7487) );
  OAI21_X1 U5731 ( .B1(n5115), .B2(n5114), .A(n5113), .ZN(n5923) );
  INV_X1 U5732 ( .A(REIP_REG_0__SCAN_IN), .ZN(n5116) );
  OR2_X1 U5733 ( .A1(n7477), .A2(n5116), .ZN(n7498) );
  OAI21_X1 U5734 ( .B1(n5923), .B2(n7059), .A(n7498), .ZN(n5117) );
  AOI21_X1 U5735 ( .B1(n7402), .B2(n7487), .A(n5117), .ZN(n5118) );
  NAND2_X1 U5736 ( .A1(n5119), .A2(n5118), .ZN(U2986) );
  INV_X1 U5737 ( .A(n7428), .ZN(n5165) );
  OAI21_X1 U5738 ( .B1(n7639), .B2(n3963), .A(n5165), .ZN(n5121) );
  NAND2_X1 U5739 ( .A1(n5121), .A2(n5120), .ZN(n5122) );
  NAND2_X1 U5740 ( .A1(n5122), .A2(n7709), .ZN(n5125) );
  INV_X1 U5741 ( .A(n5123), .ZN(n5124) );
  OAI21_X1 U5742 ( .B1(n7693), .B2(n5125), .A(n5124), .ZN(n5126) );
  OR3_X1 U5743 ( .A1(n5128), .A2(n5127), .A3(n5126), .ZN(n7636) );
  NAND2_X1 U5744 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7674), .ZN(n7680) );
  INV_X1 U5745 ( .A(n7680), .ZN(n7681) );
  AOI22_X1 U5746 ( .A1(n7688), .A2(n7636), .B1(FLUSH_REG_SCAN_IN), .B2(n7681), 
        .ZN(n7634) );
  OAI21_X1 U5747 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n5034), .A(n7634), .ZN(
        n7631) );
  OAI21_X1 U5748 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7229), .A(n7631), 
        .ZN(n5156) );
  INV_X1 U5749 ( .A(n5156), .ZN(n5138) );
  INV_X1 U5750 ( .A(n7639), .ZN(n5277) );
  INV_X1 U5751 ( .A(n5089), .ZN(n5420) );
  AND4_X1 U5752 ( .A1(n4456), .A2(n4330), .A3(n4324), .A4(n5130), .ZN(n5131)
         );
  NAND2_X1 U5753 ( .A1(n5132), .A2(n5131), .ZN(n5270) );
  NAND2_X1 U5754 ( .A1(n5420), .A2(n5270), .ZN(n5135) );
  OAI21_X1 U5755 ( .B1(n3814), .B2(n5133), .A(n5139), .ZN(n5134) );
  OAI211_X1 U5756 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n5277), .A(n5135), .B(n5134), .ZN(n7635) );
  INV_X1 U5757 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5136) );
  AOI22_X1 U5758 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5136), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n7472), .ZN(n5150) );
  NOR2_X1 U5759 ( .A1(n7422), .A2(n7489), .ZN(n5149) );
  NOR2_X1 U5760 ( .A1(n7229), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5155)
         );
  AOI222_X1 U5761 ( .A1(n7635), .A2(n5154), .B1(n5150), .B2(n5149), .C1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n5155), .ZN(n5137) );
  INV_X1 U5762 ( .A(n7631), .ZN(n5158) );
  OAI22_X1 U5763 ( .A1(n5138), .A2(n3781), .B1(n5137), .B2(n5158), .ZN(U3460)
         );
  AOI22_X1 U5764 ( .A1(n4509), .A2(n5270), .B1(n5139), .B2(n3809), .ZN(n7637)
         );
  INV_X1 U5765 ( .A(n5154), .ZN(n7629) );
  OAI22_X1 U5766 ( .A1(n7637), .A2(n7629), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n7422), .ZN(n5140) );
  OAI22_X1 U5767 ( .A1(n5156), .A2(n5140), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7631), .ZN(n5142) );
  NAND3_X1 U5768 ( .A1(n7639), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n5154), .ZN(n5141) );
  NAND2_X1 U5769 ( .A1(n5142), .A2(n5141), .ZN(U3461) );
  NAND2_X1 U5770 ( .A1(n3668), .A2(n5270), .ZN(n5148) );
  INV_X1 U5771 ( .A(n5183), .ZN(n7617) );
  NAND2_X1 U5772 ( .A1(n7617), .A2(n5143), .ZN(n5272) );
  INV_X1 U5773 ( .A(n5144), .ZN(n7225) );
  XNOR2_X1 U5774 ( .A(n5144), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5146)
         );
  XNOR2_X1 U5775 ( .A(n3731), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5145)
         );
  AOI22_X1 U5776 ( .A1(n5272), .A2(n5146), .B1(n7639), .B2(n5145), .ZN(n5147)
         );
  NAND2_X1 U5777 ( .A1(n5148), .A2(n5147), .ZN(n5279) );
  INV_X1 U5778 ( .A(n5149), .ZN(n5151) );
  NOR2_X1 U5779 ( .A1(n5151), .A2(n5150), .ZN(n5153) );
  NOR3_X1 U5780 ( .A1(n7229), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n7225), 
        .ZN(n5152) );
  AOI211_X1 U5781 ( .C1(n5154), .C2(n5279), .A(n5153), .B(n5152), .ZN(n5159)
         );
  OAI21_X1 U5782 ( .B1(n5156), .B2(n5155), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n5157) );
  OAI21_X1 U5783 ( .B1(n5159), .B2(n5158), .A(n5157), .ZN(U3459) );
  NOR2_X2 U5784 ( .A1(n5167), .A2(n5164), .ZN(n5409) );
  AOI22_X1 U5785 ( .A1(n5366), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n5409), .ZN(n5161) );
  NAND2_X1 U5786 ( .A1(n5410), .A2(DATAI_5_), .ZN(n5407) );
  NAND2_X1 U5787 ( .A1(n5161), .A2(n5407), .ZN(U2929) );
  AOI22_X1 U5788 ( .A1(n5366), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n5409), .ZN(n5162) );
  NAND2_X1 U5789 ( .A1(n5410), .A2(DATAI_3_), .ZN(n5378) );
  NAND2_X1 U5790 ( .A1(n5162), .A2(n5378), .ZN(U2927) );
  AOI22_X1 U5791 ( .A1(n5366), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n5409), .ZN(n5163) );
  NAND2_X1 U5792 ( .A1(n5410), .A2(DATAI_4_), .ZN(n5380) );
  NAND2_X1 U5793 ( .A1(n5163), .A2(n5380), .ZN(U2928) );
  INV_X1 U5794 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5171) );
  INV_X1 U5795 ( .A(n5164), .ZN(n7666) );
  OAI21_X1 U5796 ( .B1(n7639), .B2(n7666), .A(n5165), .ZN(n5166) );
  NAND2_X1 U5797 ( .A1(n5169), .A2(n4017), .ZN(n5541) );
  OR2_X1 U5798 ( .A1(n7669), .A2(n5168), .ZN(n7664) );
  INV_X2 U5799 ( .A(n7664), .ZN(n7427) );
  NOR2_X4 U5800 ( .A1(n7427), .A2(n5169), .ZN(n7268) );
  AOI22_X1 U5801 ( .A1(n7427), .A2(UWORD_REG_5__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5170) );
  OAI21_X1 U5802 ( .B1(n5171), .B2(n5541), .A(n5170), .ZN(U2902) );
  INV_X1 U5803 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5173) );
  AOI22_X1 U5804 ( .A1(n7427), .A2(UWORD_REG_9__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5172) );
  OAI21_X1 U5805 ( .B1(n5173), .B2(n5541), .A(n5172), .ZN(U2898) );
  INV_X1 U5806 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5175) );
  AOI22_X1 U5807 ( .A1(n7427), .A2(UWORD_REG_6__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5174) );
  OAI21_X1 U5808 ( .B1(n5175), .B2(n5541), .A(n5174), .ZN(U2901) );
  INV_X1 U5809 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5177) );
  AOI22_X1 U5810 ( .A1(n7427), .A2(UWORD_REG_7__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5176) );
  OAI21_X1 U5811 ( .B1(n5177), .B2(n5541), .A(n5176), .ZN(U2900) );
  AOI22_X1 U5812 ( .A1(n7427), .A2(UWORD_REG_8__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5178) );
  OAI21_X1 U5813 ( .B1(n4851), .B2(n5541), .A(n5178), .ZN(U2899) );
  NOR2_X1 U5814 ( .A1(n5179), .A2(n5180), .ZN(n5181) );
  NOR2_X1 U5815 ( .A1(n5182), .A2(n5181), .ZN(n7378) );
  INV_X1 U5816 ( .A(n7378), .ZN(n5860) );
  NAND2_X1 U5817 ( .A1(n7693), .A2(n5183), .ZN(n5189) );
  INV_X1 U5818 ( .A(n5184), .ZN(n5187) );
  NOR2_X1 U5819 ( .A1(n5249), .A2(n3949), .ZN(n5186) );
  NOR2_X1 U5820 ( .A1(n4312), .A2(n3952), .ZN(n5185) );
  NAND4_X1 U5821 ( .A1(n5187), .A2(n5191), .A3(n5186), .A4(n5185), .ZN(n5188)
         );
  NAND2_X1 U5822 ( .A1(n5189), .A2(n5188), .ZN(n5190) );
  XNOR2_X1 U5823 ( .A(n5852), .B(n5191), .ZN(n5223) );
  AOI22_X1 U5824 ( .A1(n7369), .A2(n5223), .B1(n6541), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5192) );
  OAI21_X1 U5825 ( .B1(n5860), .B2(n6539), .A(n5192), .ZN(U2858) );
  AOI21_X1 U5826 ( .B1(n5194), .B2(n5492), .A(n5195), .ZN(n5196) );
  NOR2_X1 U5827 ( .A1(n4550), .A2(n5196), .ZN(n6154) );
  INV_X1 U5828 ( .A(n6154), .ZN(n5227) );
  NAND2_X1 U5829 ( .A1(n6368), .A2(n5197), .ZN(n5198) );
  AND2_X1 U5830 ( .A1(n5212), .A2(n5198), .ZN(n7444) );
  AOI22_X1 U5831 ( .A1(n7369), .A2(n7444), .B1(n6541), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n5199) );
  OAI21_X1 U5832 ( .B1(n5227), .B2(n6539), .A(n5199), .ZN(U2855) );
  NOR2_X1 U5833 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  NOR2_X1 U5834 ( .A1(n5194), .A2(n5202), .ZN(n7514) );
  INV_X1 U5835 ( .A(n7514), .ZN(n5495) );
  NOR2_X1 U5836 ( .A1(n5204), .A2(n5203), .ZN(n5206) );
  NOR2_X1 U5837 ( .A1(n5206), .A2(n5205), .ZN(n7508) );
  AOI22_X1 U5838 ( .A1(n7369), .A2(n7508), .B1(n6541), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5207) );
  OAI21_X1 U5839 ( .B1(n5495), .B2(n6539), .A(n5207), .ZN(U2857) );
  NAND2_X1 U5840 ( .A1(n5193), .A2(n5209), .ZN(n5210) );
  AND2_X1 U5841 ( .A1(n5208), .A2(n5210), .ZN(n7401) );
  INV_X1 U5842 ( .A(n5363), .ZN(n5211) );
  AOI21_X1 U5843 ( .B1(n5213), .B2(n5212), .A(n5211), .ZN(n7519) );
  AOI22_X1 U5844 ( .A1(n7369), .A2(n7519), .B1(n6541), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n5214) );
  OAI21_X1 U5845 ( .B1(n7523), .B2(n6539), .A(n5214), .ZN(U2854) );
  NAND2_X1 U5846 ( .A1(n5215), .A2(n5216), .ZN(n5217) );
  XOR2_X1 U5847 ( .A(n5218), .B(n5217), .Z(n7377) );
  NAND2_X1 U5848 ( .A1(n7462), .A2(n6323), .ZN(n7490) );
  AOI21_X1 U5849 ( .B1(n7489), .B2(n7490), .A(n7491), .ZN(n5219) );
  OAI22_X1 U5850 ( .A1(n7477), .A2(n7506), .B1(n5219), .B2(n7472), .ZN(n5222)
         );
  NOR3_X1 U5851 ( .A1(n7176), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n5220), 
        .ZN(n5221) );
  AOI211_X1 U5852 ( .C1(n7495), .C2(n5223), .A(n5222), .B(n5221), .ZN(n5224)
         );
  OAI21_X1 U5853 ( .B1(n7212), .B2(n7377), .A(n5224), .ZN(U3017) );
  INV_X1 U5854 ( .A(EAX_REG_0__SCAN_IN), .ZN(n7258) );
  OAI222_X1 U5855 ( .A1(n6335), .A2(n5226), .B1(n6392), .B2(n7258), .C1(n6568), 
        .C2(n5923), .ZN(U2891) );
  INV_X1 U5856 ( .A(DATAI_4_), .ZN(n5239) );
  INV_X1 U5857 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7266) );
  OAI222_X1 U5858 ( .A1(n6335), .A2(n5239), .B1(n6392), .B2(n7266), .C1(n6568), 
        .C2(n5227), .ZN(U2887) );
  OR2_X1 U5859 ( .A1(n5228), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5230)
         );
  NAND2_X1 U5860 ( .A1(n5230), .A2(n5229), .ZN(n7493) );
  OAI222_X1 U5861 ( .A1(n7493), .A2(n7372), .B1(n4344), .B2(n7376), .C1(n5923), 
        .C2(n6539), .ZN(U2859) );
  INV_X1 U5862 ( .A(n5231), .ZN(n5232) );
  AOI21_X1 U5863 ( .B1(n5234), .B2(n5233), .A(n5232), .ZN(n7447) );
  INV_X1 U5864 ( .A(n7447), .ZN(n5238) );
  AOI22_X1 U5865 ( .A1(n7396), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n7460), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n5235) );
  OAI21_X1 U5866 ( .B1(n6152), .B2(n7405), .A(n5235), .ZN(n5236) );
  AOI21_X1 U5867 ( .B1(n6154), .B2(n7392), .A(n5236), .ZN(n5237) );
  OAI21_X1 U5868 ( .B1(n5238), .B2(n7626), .A(n5237), .ZN(U2982) );
  NAND2_X1 U5869 ( .A1(n5259), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n5242)
         );
  NAND2_X1 U5870 ( .A1(n7392), .A2(DATAI_28_), .ZN(n6093) );
  INV_X1 U5871 ( .A(n6093), .ZN(n5736) );
  AND2_X1 U5872 ( .A1(n7392), .A2(DATAI_20_), .ZN(n6095) );
  INV_X1 U5873 ( .A(n6095), .ZN(n5739) );
  NAND2_X1 U5874 ( .A1(n5260), .A2(n3949), .ZN(n6005) );
  OAI22_X1 U5875 ( .A1(n5739), .A2(n5839), .B1(n6005), .B2(n5261), .ZN(n5240)
         );
  AOI21_X1 U5876 ( .B1(n5736), .B2(n5621), .A(n5240), .ZN(n5241) );
  OAI211_X1 U5877 ( .C1(n5265), .C2(n6004), .A(n5242), .B(n5241), .ZN(U3112)
         );
  INV_X1 U5878 ( .A(DATAI_6_), .ZN(n5494) );
  NAND2_X1 U5879 ( .A1(n5259), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5245)
         );
  NAND2_X1 U5880 ( .A1(n7392), .A2(DATAI_30_), .ZN(n6109) );
  INV_X1 U5881 ( .A(n6109), .ZN(n5746) );
  AND2_X1 U5882 ( .A1(n7392), .A2(DATAI_22_), .ZN(n6111) );
  INV_X1 U5883 ( .A(n6111), .ZN(n5749) );
  NAND2_X1 U5884 ( .A1(n5260), .A2(n5073), .ZN(n6000) );
  OAI22_X1 U5885 ( .A1(n5749), .A2(n5839), .B1(n6000), .B2(n5261), .ZN(n5243)
         );
  AOI21_X1 U5886 ( .B1(n5746), .B2(n5621), .A(n5243), .ZN(n5244) );
  OAI211_X1 U5887 ( .C1(n5265), .C2(n5999), .A(n5245), .B(n5244), .ZN(U3114)
         );
  INV_X1 U5888 ( .A(DATAI_1_), .ZN(n5374) );
  NAND2_X1 U5889 ( .A1(n5259), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n5248)
         );
  NAND2_X1 U5890 ( .A1(n7392), .A2(DATAI_25_), .ZN(n6101) );
  INV_X1 U5891 ( .A(n6101), .ZN(n5741) );
  AND2_X1 U5892 ( .A1(n7392), .A2(DATAI_17_), .ZN(n6103) );
  INV_X1 U5893 ( .A(n6103), .ZN(n5744) );
  NAND2_X1 U5894 ( .A1(n5260), .A2(n3965), .ZN(n6020) );
  OAI22_X1 U5895 ( .A1(n5744), .A2(n5839), .B1(n6020), .B2(n5261), .ZN(n5246)
         );
  AOI21_X1 U5896 ( .B1(n5741), .B2(n5621), .A(n5246), .ZN(n5247) );
  OAI211_X1 U5897 ( .C1(n5265), .C2(n6019), .A(n5248), .B(n5247), .ZN(U3109)
         );
  INV_X1 U5898 ( .A(DATAI_3_), .ZN(n5493) );
  NAND2_X1 U5899 ( .A1(n5259), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5252)
         );
  NAND2_X1 U5900 ( .A1(n7392), .A2(DATAI_27_), .ZN(n6124) );
  INV_X1 U5901 ( .A(n6124), .ZN(n5756) );
  AND2_X1 U5902 ( .A1(n7392), .A2(DATAI_19_), .ZN(n6126) );
  INV_X1 U5903 ( .A(n6126), .ZN(n5759) );
  NAND2_X1 U5904 ( .A1(n5260), .A2(n5249), .ZN(n6010) );
  OAI22_X1 U5905 ( .A1(n5759), .A2(n5839), .B1(n6010), .B2(n5261), .ZN(n5250)
         );
  AOI21_X1 U5906 ( .B1(n5756), .B2(n5621), .A(n5250), .ZN(n5251) );
  OAI211_X1 U5907 ( .C1(n5265), .C2(n6009), .A(n5252), .B(n5251), .ZN(U3111)
         );
  INV_X1 U5908 ( .A(DATAI_2_), .ZN(n5496) );
  NAND2_X1 U5909 ( .A1(n5259), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5255)
         );
  NAND2_X1 U5910 ( .A1(n7392), .A2(DATAI_26_), .ZN(n6085) );
  INV_X1 U5911 ( .A(n6085), .ZN(n5726) );
  AND2_X1 U5912 ( .A1(n7392), .A2(DATAI_18_), .ZN(n6087) );
  INV_X1 U5913 ( .A(n6087), .ZN(n5729) );
  NAND2_X1 U5914 ( .A1(n5260), .A2(n4312), .ZN(n6015) );
  OAI22_X1 U5915 ( .A1(n5729), .A2(n5839), .B1(n6015), .B2(n5261), .ZN(n5253)
         );
  AOI21_X1 U5916 ( .B1(n5726), .B2(n5621), .A(n5253), .ZN(n5254) );
  OAI211_X1 U5917 ( .C1(n5265), .C2(n6014), .A(n5255), .B(n5254), .ZN(U3110)
         );
  INV_X1 U5918 ( .A(DATAI_5_), .ZN(n5491) );
  NAND2_X1 U5919 ( .A1(n5259), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5258)
         );
  NAND2_X1 U5920 ( .A1(n7392), .A2(DATAI_29_), .ZN(n6116) );
  INV_X1 U5921 ( .A(n6116), .ZN(n5751) );
  AND2_X1 U5922 ( .A1(n7392), .A2(DATAI_21_), .ZN(n6118) );
  INV_X1 U5923 ( .A(n6118), .ZN(n5754) );
  NAND2_X1 U5924 ( .A1(n5260), .A2(n3954), .ZN(n6038) );
  OAI22_X1 U5925 ( .A1(n5754), .A2(n5839), .B1(n6038), .B2(n5261), .ZN(n5256)
         );
  AOI21_X1 U5926 ( .B1(n5751), .B2(n5621), .A(n5256), .ZN(n5257) );
  OAI211_X1 U5927 ( .C1(n5265), .C2(n6035), .A(n5258), .B(n5257), .ZN(U3113)
         );
  INV_X1 U5928 ( .A(DATAI_7_), .ZN(n5525) );
  NAND2_X1 U5929 ( .A1(n5259), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5264)
         );
  NAND2_X1 U5930 ( .A1(n7392), .A2(DATAI_31_), .ZN(n6077) );
  INV_X1 U5931 ( .A(n6077), .ZN(n5731) );
  AND2_X1 U5932 ( .A1(n7392), .A2(DATAI_23_), .ZN(n6079) );
  INV_X1 U5933 ( .A(n6079), .ZN(n5734) );
  NAND2_X1 U5934 ( .A1(n5260), .A2(n3952), .ZN(n6030) );
  OAI22_X1 U5935 ( .A1(n5734), .A2(n5839), .B1(n6030), .B2(n5261), .ZN(n5262)
         );
  AOI21_X1 U5936 ( .B1(n5731), .B2(n5621), .A(n5262), .ZN(n5263) );
  OAI211_X1 U5937 ( .C1(n5265), .C2(n6029), .A(n5264), .B(n5263), .ZN(U3115)
         );
  AOI22_X1 U5938 ( .A1(n5366), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n5402), .ZN(n5266) );
  NAND2_X1 U5939 ( .A1(n5410), .A2(DATAI_6_), .ZN(n5383) );
  NAND2_X1 U5940 ( .A1(n5266), .A2(n5383), .ZN(U2930) );
  AOI22_X1 U5941 ( .A1(n5366), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n5402), .ZN(n5267) );
  NAND2_X1 U5942 ( .A1(n5410), .A2(DATAI_8_), .ZN(n5371) );
  NAND2_X1 U5943 ( .A1(n5267), .A2(n5371), .ZN(U2932) );
  AOI22_X1 U5944 ( .A1(n5366), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n5402), .ZN(n5268) );
  NAND2_X1 U5945 ( .A1(n5410), .A2(DATAI_7_), .ZN(n5385) );
  NAND2_X1 U5946 ( .A1(n5268), .A2(n5385), .ZN(U2931) );
  INV_X1 U5947 ( .A(n3667), .ZN(n6374) );
  NAND2_X1 U5948 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5269) );
  AOI22_X1 U5949 ( .A1(n5274), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n7231), .B2(n5269), .ZN(n5278) );
  NAND2_X1 U5950 ( .A1(n3667), .A2(n5270), .ZN(n5276) );
  MUX2_X1 U5951 ( .A(n5271), .B(n3804), .S(n5144), .Z(n5273) );
  OAI21_X1 U5952 ( .B1(n5274), .B2(n5273), .A(n5272), .ZN(n5275) );
  OAI211_X1 U5953 ( .C1(n5278), .C2(n5277), .A(n5276), .B(n5275), .ZN(n7226)
         );
  MUX2_X1 U5954 ( .A(n7231), .B(n7226), .S(n7636), .Z(n7650) );
  NAND2_X1 U5955 ( .A1(n7636), .A2(n5279), .ZN(n5280) );
  OAI21_X1 U5956 ( .B1(n7636), .B2(n3731), .A(n5280), .ZN(n7644) );
  NAND3_X1 U5957 ( .A1(n7650), .A2(n7422), .A3(n7644), .ZN(n5284) );
  NOR2_X1 U5958 ( .A1(FLUSH_REG_SCAN_IN), .A2(n7422), .ZN(n5281) );
  NAND2_X1 U5959 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  NAND2_X1 U5960 ( .A1(n5284), .A2(n5283), .ZN(n7662) );
  INV_X1 U5961 ( .A(n3820), .ZN(n5285) );
  NAND2_X1 U5962 ( .A1(n7662), .A2(n5285), .ZN(n5294) );
  MUX2_X1 U5963 ( .A(n7636), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n5286) );
  INV_X1 U5964 ( .A(n5286), .ZN(n5293) );
  INV_X1 U5965 ( .A(n5287), .ZN(n5288) );
  OR2_X1 U5966 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  XNOR2_X1 U5967 ( .A(n5290), .B(n7632), .ZN(n7630) );
  OR2_X1 U5968 ( .A1(n4330), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5291) );
  NOR2_X1 U5969 ( .A1(n7630), .A2(n5291), .ZN(n5292) );
  AOI21_X1 U5970 ( .B1(n5293), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n5292), 
        .ZN(n7660) );
  NAND2_X1 U5971 ( .A1(n5294), .A2(n7660), .ZN(n5301) );
  OAI21_X1 U5972 ( .B1(n5301), .B2(FLUSH_REG_SCAN_IN), .A(n7681), .ZN(n5295)
         );
  INV_X1 U5973 ( .A(n7254), .ZN(n5418) );
  OAI21_X1 U5974 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7422), .A(n5418), .ZN(
        n6401) );
  NOR2_X1 U5975 ( .A1(n7254), .A2(n5679), .ZN(n6398) );
  INV_X1 U5976 ( .A(n5505), .ZN(n5497) );
  NOR2_X1 U5977 ( .A1(n5497), .A2(n7696), .ZN(n5498) );
  NOR2_X1 U5978 ( .A1(n5334), .A2(n6397), .ZN(n5327) );
  AOI21_X1 U5979 ( .B1(n5413), .B2(STATEBS16_REG_SCAN_IN), .A(n5626), .ZN(
        n5298) );
  OR3_X1 U5980 ( .A1(n5498), .A2(n5327), .A3(n5298), .ZN(n5299) );
  AOI22_X1 U5981 ( .A1(n6398), .A2(n5299), .B1(n7254), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5300) );
  OAI21_X1 U5982 ( .B1(n6374), .B2(n6401), .A(n5300), .ZN(U3462) );
  INV_X1 U5983 ( .A(n4509), .ZN(n5918) );
  INV_X1 U5984 ( .A(n5301), .ZN(n7682) );
  NAND2_X1 U5985 ( .A1(n7682), .A2(n7674), .ZN(n5303) );
  NAND2_X1 U5986 ( .A1(n7254), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5302) );
  OAI21_X1 U5987 ( .B1(n7254), .B2(n5303), .A(n5302), .ZN(n5304) );
  AOI21_X1 U5988 ( .B1(n6398), .B2(n5637), .A(n5304), .ZN(n5305) );
  OAI21_X1 U5989 ( .B1(n5918), .B2(n6401), .A(n5305), .ZN(U3465) );
  INV_X1 U5990 ( .A(n5334), .ZN(n5326) );
  NOR2_X1 U5991 ( .A1(n5084), .A2(n7696), .ZN(n5306) );
  AOI21_X1 U5992 ( .B1(n5326), .B2(n5306), .A(n5679), .ZN(n5308) );
  NOR2_X1 U5993 ( .A1(n3667), .A2(n5918), .ZN(n5633) );
  NAND2_X1 U5994 ( .A1(n3668), .A2(n5089), .ZN(n5951) );
  INV_X1 U5995 ( .A(n5951), .ZN(n5799) );
  NAND3_X1 U5996 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7649), .A3(n5630), .ZN(n5943) );
  NOR2_X1 U5997 ( .A1(n5629), .A2(n5943), .ZN(n5348) );
  AOI21_X1 U5998 ( .B1(n5633), .B2(n5799), .A(n5348), .ZN(n5310) );
  AOI22_X1 U5999 ( .A1(n5308), .A2(n5310), .B1(n5679), .B2(n5943), .ZN(n5307)
         );
  NAND2_X1 U6000 ( .A1(n5551), .A2(n5307), .ZN(n5346) );
  INV_X1 U6001 ( .A(n5308), .ZN(n5309) );
  OAI22_X1 U6002 ( .A1(n5310), .A2(n5309), .B1(n7669), .B2(n5943), .ZN(n5345)
         );
  AOI22_X1 U6003 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5346), .B1(n6082), 
        .B2(n5345), .ZN(n5313) );
  AOI22_X1 U6004 ( .A1(n6083), .A2(n5348), .B1(n5347), .B2(n6087), .ZN(n5312)
         );
  OAI211_X1 U6005 ( .C1(n6085), .C2(n5948), .A(n5313), .B(n5312), .ZN(U3062)
         );
  AOI22_X1 U6006 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5346), .B1(n6121), 
        .B2(n5345), .ZN(n5315) );
  AOI22_X1 U6007 ( .A1(n6122), .A2(n5348), .B1(n5347), .B2(n6126), .ZN(n5314)
         );
  OAI211_X1 U6008 ( .C1(n6124), .C2(n5948), .A(n5315), .B(n5314), .ZN(U3063)
         );
  AOI22_X1 U6009 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5346), .B1(n6113), 
        .B2(n5345), .ZN(n5317) );
  AOI22_X1 U6010 ( .A1(n6114), .A2(n5348), .B1(n5347), .B2(n6118), .ZN(n5316)
         );
  OAI211_X1 U6011 ( .C1(n6116), .C2(n5948), .A(n5317), .B(n5316), .ZN(U3065)
         );
  AOI22_X1 U6012 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5346), .B1(n6106), 
        .B2(n5345), .ZN(n5319) );
  AOI22_X1 U6013 ( .A1(n6107), .A2(n5348), .B1(n5347), .B2(n6111), .ZN(n5318)
         );
  OAI211_X1 U6014 ( .C1(n6109), .C2(n5948), .A(n5319), .B(n5318), .ZN(U3066)
         );
  AOI22_X1 U6015 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5346), .B1(n6090), 
        .B2(n5345), .ZN(n5321) );
  AOI22_X1 U6016 ( .A1(n6091), .A2(n5348), .B1(n5347), .B2(n6095), .ZN(n5320)
         );
  OAI211_X1 U6017 ( .C1(n6093), .C2(n5948), .A(n5321), .B(n5320), .ZN(U3064)
         );
  AOI22_X1 U6018 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5346), .B1(n6130), 
        .B2(n5345), .ZN(n5323) );
  AOI22_X1 U6019 ( .A1(n6132), .A2(n5348), .B1(n5347), .B2(n6138), .ZN(n5322)
         );
  OAI211_X1 U6020 ( .C1(n6135), .C2(n5948), .A(n5323), .B(n5322), .ZN(U3060)
         );
  AOI22_X1 U6021 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5346), .B1(n6098), 
        .B2(n5345), .ZN(n5325) );
  AOI22_X1 U6022 ( .A1(n6099), .A2(n5348), .B1(n5347), .B2(n6103), .ZN(n5324)
         );
  OAI211_X1 U6023 ( .C1(n6101), .C2(n5948), .A(n5325), .B(n5324), .ZN(U3061)
         );
  NOR2_X1 U6024 ( .A1(n5327), .A2(n5679), .ZN(n5330) );
  AND2_X1 U6025 ( .A1(n3668), .A2(n5420), .ZN(n5724) );
  INV_X1 U6026 ( .A(n5328), .ZN(n5357) );
  AOI21_X1 U6027 ( .B1(n5633), .B2(n5724), .A(n5357), .ZN(n5332) );
  NAND3_X1 U6028 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7649), .ZN(n5671) );
  AOI22_X1 U6029 ( .A1(n5330), .A2(n5332), .B1(n5679), .B2(n5671), .ZN(n5329)
         );
  NAND2_X1 U6030 ( .A1(n5551), .A2(n5329), .ZN(n5356) );
  INV_X1 U6031 ( .A(n5330), .ZN(n5331) );
  OAI22_X1 U6032 ( .A1(n5332), .A2(n5331), .B1(n7669), .B2(n5671), .ZN(n5355)
         );
  AOI22_X1 U6033 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5356), .B1(n6082), 
        .B2(n5355), .ZN(n5336) );
  NAND2_X1 U6034 ( .A1(n5084), .A2(n5552), .ZN(n5333) );
  NOR2_X2 U6035 ( .A1(n5334), .A2(n5333), .ZN(n5706) );
  AOI22_X1 U6036 ( .A1(n6083), .A2(n5357), .B1(n5726), .B2(n5706), .ZN(n5335)
         );
  OAI211_X1 U6037 ( .C1(n5729), .C2(n5912), .A(n5336), .B(n5335), .ZN(U3078)
         );
  AOI22_X1 U6038 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5356), .B1(n6121), 
        .B2(n5355), .ZN(n5338) );
  AOI22_X1 U6039 ( .A1(n6122), .A2(n5357), .B1(n5756), .B2(n5706), .ZN(n5337)
         );
  OAI211_X1 U6040 ( .C1(n5759), .C2(n5912), .A(n5338), .B(n5337), .ZN(U3079)
         );
  AOI22_X1 U6041 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5356), .B1(n6090), 
        .B2(n5355), .ZN(n5340) );
  AOI22_X1 U6042 ( .A1(n6091), .A2(n5357), .B1(n5736), .B2(n5706), .ZN(n5339)
         );
  OAI211_X1 U6043 ( .C1(n5739), .C2(n5912), .A(n5340), .B(n5339), .ZN(U3080)
         );
  AOI22_X1 U6044 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5356), .B1(n6113), 
        .B2(n5355), .ZN(n5342) );
  AOI22_X1 U6045 ( .A1(n6114), .A2(n5357), .B1(n5751), .B2(n5706), .ZN(n5341)
         );
  OAI211_X1 U6046 ( .C1(n5754), .C2(n5912), .A(n5342), .B(n5341), .ZN(U3081)
         );
  AOI22_X1 U6047 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5356), .B1(n6074), 
        .B2(n5355), .ZN(n5344) );
  AOI22_X1 U6048 ( .A1(n6075), .A2(n5357), .B1(n5731), .B2(n5706), .ZN(n5343)
         );
  OAI211_X1 U6049 ( .C1(n5734), .C2(n5912), .A(n5344), .B(n5343), .ZN(U3083)
         );
  AOI22_X1 U6050 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5346), .B1(n6074), 
        .B2(n5345), .ZN(n5350) );
  AOI22_X1 U6051 ( .A1(n6075), .A2(n5348), .B1(n5347), .B2(n6079), .ZN(n5349)
         );
  OAI211_X1 U6052 ( .C1(n6077), .C2(n5948), .A(n5350), .B(n5349), .ZN(U3067)
         );
  AOI22_X1 U6053 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5356), .B1(n6130), 
        .B2(n5355), .ZN(n5352) );
  INV_X1 U6054 ( .A(n6135), .ZN(n5765) );
  AOI22_X1 U6055 ( .A1(n6132), .A2(n5357), .B1(n5765), .B2(n5706), .ZN(n5351)
         );
  OAI211_X1 U6056 ( .C1(n5768), .C2(n5912), .A(n5352), .B(n5351), .ZN(U3076)
         );
  AOI22_X1 U6057 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5356), .B1(n6098), 
        .B2(n5355), .ZN(n5354) );
  AOI22_X1 U6058 ( .A1(n6099), .A2(n5357), .B1(n5741), .B2(n5706), .ZN(n5353)
         );
  OAI211_X1 U6059 ( .C1(n5744), .C2(n5912), .A(n5354), .B(n5353), .ZN(U3077)
         );
  AOI22_X1 U6060 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5356), .B1(n6106), 
        .B2(n5355), .ZN(n5359) );
  AOI22_X1 U6061 ( .A1(n6107), .A2(n5357), .B1(n5746), .B2(n5706), .ZN(n5358)
         );
  OAI211_X1 U6062 ( .C1(n5749), .C2(n5912), .A(n5359), .B(n5358), .ZN(U3082)
         );
  AND2_X1 U6063 ( .A1(n5360), .A2(n5208), .ZN(n5362) );
  OR2_X1 U6064 ( .A1(n5362), .A2(n5361), .ZN(n5940) );
  AOI21_X1 U6065 ( .B1(n5364), .B2(n5363), .A(n5449), .ZN(n5934) );
  AOI22_X1 U6066 ( .A1(n7369), .A2(n5934), .B1(n6541), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n5365) );
  OAI21_X1 U6067 ( .B1(n5940), .B2(n6543), .A(n5365), .ZN(U2853) );
  AOI22_X1 U6068 ( .A1(n5411), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n5402), .ZN(n5367) );
  NAND2_X1 U6069 ( .A1(n5410), .A2(DATAI_9_), .ZN(n5389) );
  NAND2_X1 U6070 ( .A1(n5367), .A2(n5389), .ZN(U2933) );
  AOI22_X1 U6071 ( .A1(n5411), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n5402), .ZN(n5368) );
  NAND2_X1 U6072 ( .A1(n5410), .A2(DATAI_11_), .ZN(n5392) );
  NAND2_X1 U6073 ( .A1(n5368), .A2(n5392), .ZN(U2935) );
  AOI22_X1 U6074 ( .A1(n5411), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n5402), .ZN(n5369) );
  INV_X1 U6075 ( .A(DATAI_12_), .ZN(n6242) );
  OR2_X1 U6076 ( .A1(n5375), .A2(n6242), .ZN(n5394) );
  NAND2_X1 U6077 ( .A1(n5369), .A2(n5394), .ZN(U2936) );
  AOI22_X1 U6078 ( .A1(n5411), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n5402), .ZN(n5370) );
  NAND2_X1 U6079 ( .A1(n5410), .A2(DATAI_13_), .ZN(n5396) );
  NAND2_X1 U6080 ( .A1(n5370), .A2(n5396), .ZN(U2937) );
  AOI22_X1 U6081 ( .A1(n5411), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n5402), .ZN(n5372) );
  NAND2_X1 U6082 ( .A1(n5372), .A2(n5371), .ZN(U2947) );
  AOI22_X1 U6083 ( .A1(n5411), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n5402), .ZN(n5373) );
  NAND2_X1 U6084 ( .A1(n5410), .A2(DATAI_0_), .ZN(n5403) );
  NAND2_X1 U6085 ( .A1(n5373), .A2(n5403), .ZN(U2939) );
  AOI22_X1 U6086 ( .A1(n5411), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n5402), .ZN(n5376) );
  OR2_X1 U6087 ( .A1(n5375), .A2(n5374), .ZN(n5405) );
  NAND2_X1 U6088 ( .A1(n5376), .A2(n5405), .ZN(U2940) );
  AOI22_X1 U6089 ( .A1(n5411), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n5409), .ZN(n5377) );
  NAND2_X1 U6090 ( .A1(n5410), .A2(DATAI_2_), .ZN(n5387) );
  NAND2_X1 U6091 ( .A1(n5377), .A2(n5387), .ZN(U2941) );
  AOI22_X1 U6092 ( .A1(n5411), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n5409), .ZN(n5379) );
  NAND2_X1 U6093 ( .A1(n5379), .A2(n5378), .ZN(U2942) );
  AOI22_X1 U6094 ( .A1(n5411), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n5409), .ZN(n5381) );
  NAND2_X1 U6095 ( .A1(n5381), .A2(n5380), .ZN(U2943) );
  AOI22_X1 U6096 ( .A1(n5411), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n5402), .ZN(n5382) );
  NAND2_X1 U6097 ( .A1(n5410), .A2(DATAI_14_), .ZN(n5398) );
  NAND2_X1 U6098 ( .A1(n5382), .A2(n5398), .ZN(U2938) );
  AOI22_X1 U6099 ( .A1(n5411), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n5409), .ZN(n5384) );
  NAND2_X1 U6100 ( .A1(n5384), .A2(n5383), .ZN(U2945) );
  AOI22_X1 U6101 ( .A1(n5411), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n5402), .ZN(n5386) );
  NAND2_X1 U6102 ( .A1(n5386), .A2(n5385), .ZN(U2946) );
  AOI22_X1 U6103 ( .A1(n5411), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n5409), .ZN(n5388) );
  NAND2_X1 U6104 ( .A1(n5388), .A2(n5387), .ZN(U2926) );
  AOI22_X1 U6105 ( .A1(n5411), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n5402), .ZN(n5390) );
  NAND2_X1 U6106 ( .A1(n5390), .A2(n5389), .ZN(U2948) );
  AOI22_X1 U6107 ( .A1(n5411), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n5402), .ZN(n5391) );
  NAND2_X1 U6108 ( .A1(n5410), .A2(DATAI_10_), .ZN(n5400) );
  NAND2_X1 U6109 ( .A1(n5391), .A2(n5400), .ZN(U2934) );
  AOI22_X1 U6110 ( .A1(n5411), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n5402), .ZN(n5393) );
  NAND2_X1 U6111 ( .A1(n5393), .A2(n5392), .ZN(U2950) );
  AOI22_X1 U6112 ( .A1(n5411), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n5402), .ZN(n5395) );
  NAND2_X1 U6113 ( .A1(n5395), .A2(n5394), .ZN(U2951) );
  AOI22_X1 U6114 ( .A1(n5411), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n5402), .ZN(n5397) );
  NAND2_X1 U6115 ( .A1(n5397), .A2(n5396), .ZN(U2952) );
  AOI22_X1 U6116 ( .A1(n5411), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n5402), .ZN(n5399) );
  NAND2_X1 U6117 ( .A1(n5399), .A2(n5398), .ZN(U2953) );
  AOI22_X1 U6118 ( .A1(n5411), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n5402), .ZN(n5401) );
  NAND2_X1 U6119 ( .A1(n5401), .A2(n5400), .ZN(U2949) );
  AOI22_X1 U6120 ( .A1(n5411), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n5402), .ZN(n5404) );
  NAND2_X1 U6121 ( .A1(n5404), .A2(n5403), .ZN(U2924) );
  AOI22_X1 U6122 ( .A1(n5411), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n5409), .ZN(n5406) );
  NAND2_X1 U6123 ( .A1(n5406), .A2(n5405), .ZN(U2925) );
  AOI22_X1 U6124 ( .A1(n5411), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n5409), .ZN(n5408) );
  NAND2_X1 U6125 ( .A1(n5408), .A2(n5407), .ZN(U2944) );
  AOI222_X1 U6126 ( .A1(n5411), .A2(LWORD_REG_15__SCAN_IN), .B1(n5410), .B2(
        DATAI_15_), .C1(EAX_REG_15__SCAN_IN), .C2(n5409), .ZN(n5412) );
  INV_X1 U6127 ( .A(n5412), .ZN(U2954) );
  INV_X1 U6128 ( .A(n3668), .ZN(n5416) );
  INV_X1 U6129 ( .A(n6398), .ZN(n5415) );
  AOI21_X1 U6130 ( .B1(n5413), .B2(n6397), .A(n5465), .ZN(n5414) );
  OAI222_X1 U6131 ( .A1(n5418), .A2(n5417), .B1(n6401), .B2(n5416), .C1(n5415), 
        .C2(n5414), .ZN(U3463) );
  NAND2_X1 U6132 ( .A1(n5085), .A2(n5543), .ZN(n5625) );
  INV_X1 U6133 ( .A(n5427), .ZN(n5419) );
  NOR2_X1 U6134 ( .A1(n5874), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5423)
         );
  OAI21_X1 U6135 ( .B1(n5427), .B2(n7696), .A(n5871), .ZN(n5425) );
  INV_X1 U6136 ( .A(n5425), .ZN(n5421) );
  AND2_X1 U6137 ( .A1(n3667), .A2(n4509), .ZN(n5546) );
  OR2_X1 U6138 ( .A1(n3668), .A2(n5420), .ZN(n6072) );
  INV_X1 U6139 ( .A(n6072), .ZN(n5632) );
  INV_X1 U6140 ( .A(n5423), .ZN(n5424) );
  NOR2_X1 U6141 ( .A1(n5629), .A2(n5424), .ZN(n5444) );
  AOI21_X1 U6142 ( .B1(n5546), .B2(n5632), .A(n5444), .ZN(n5426) );
  NAND2_X1 U6143 ( .A1(n5421), .A2(n5426), .ZN(n5422) );
  OAI211_X1 U6144 ( .C1(n5871), .C2(n5423), .A(n5551), .B(n5422), .ZN(n5443)
         );
  OAI22_X1 U6145 ( .A1(n5426), .A2(n5425), .B1(n7669), .B2(n5424), .ZN(n5442)
         );
  AOI22_X1 U6146 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5443), .B1(n6082), 
        .B2(n5442), .ZN(n5429) );
  NOR2_X2 U6147 ( .A1(n5427), .A2(n5637), .ZN(n5914) );
  AOI22_X1 U6148 ( .A1(n6083), .A2(n5444), .B1(n5914), .B2(n5726), .ZN(n5428)
         );
  OAI211_X1 U6149 ( .C1(n5619), .C2(n5729), .A(n5429), .B(n5428), .ZN(U3094)
         );
  AOI22_X1 U6150 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5443), .B1(n6074), 
        .B2(n5442), .ZN(n5431) );
  AOI22_X1 U6151 ( .A1(n6075), .A2(n5444), .B1(n5914), .B2(n5731), .ZN(n5430)
         );
  OAI211_X1 U6152 ( .C1(n5619), .C2(n5734), .A(n5431), .B(n5430), .ZN(U3099)
         );
  AOI22_X1 U6153 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5443), .B1(n6121), 
        .B2(n5442), .ZN(n5433) );
  AOI22_X1 U6154 ( .A1(n6122), .A2(n5444), .B1(n5914), .B2(n5756), .ZN(n5432)
         );
  OAI211_X1 U6155 ( .C1(n5619), .C2(n5759), .A(n5433), .B(n5432), .ZN(U3095)
         );
  AOI22_X1 U6156 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5443), .B1(n6130), 
        .B2(n5442), .ZN(n5435) );
  AOI22_X1 U6157 ( .A1(n6132), .A2(n5444), .B1(n5914), .B2(n5765), .ZN(n5434)
         );
  OAI211_X1 U6158 ( .C1(n5768), .C2(n5619), .A(n5435), .B(n5434), .ZN(U3092)
         );
  AOI22_X1 U6159 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5443), .B1(n6106), 
        .B2(n5442), .ZN(n5437) );
  AOI22_X1 U6160 ( .A1(n6107), .A2(n5444), .B1(n5914), .B2(n5746), .ZN(n5436)
         );
  OAI211_X1 U6161 ( .C1(n5619), .C2(n5749), .A(n5437), .B(n5436), .ZN(U3098)
         );
  AOI22_X1 U6162 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5443), .B1(n6090), 
        .B2(n5442), .ZN(n5439) );
  AOI22_X1 U6163 ( .A1(n6091), .A2(n5444), .B1(n5914), .B2(n5736), .ZN(n5438)
         );
  OAI211_X1 U6164 ( .C1(n5619), .C2(n5739), .A(n5439), .B(n5438), .ZN(U3096)
         );
  AOI22_X1 U6165 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5443), .B1(n6113), 
        .B2(n5442), .ZN(n5441) );
  AOI22_X1 U6166 ( .A1(n6114), .A2(n5444), .B1(n5914), .B2(n5751), .ZN(n5440)
         );
  OAI211_X1 U6167 ( .C1(n5619), .C2(n5754), .A(n5441), .B(n5440), .ZN(U3097)
         );
  AOI22_X1 U6168 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5443), .B1(n6098), 
        .B2(n5442), .ZN(n5446) );
  AOI22_X1 U6169 ( .A1(n6099), .A2(n5444), .B1(n5914), .B2(n5741), .ZN(n5445)
         );
  OAI211_X1 U6170 ( .C1(n5619), .C2(n5744), .A(n5446), .B(n5445), .ZN(U3093)
         );
  OAI21_X1 U6171 ( .B1(n5361), .B2(n5448), .A(n5447), .ZN(n7532) );
  INV_X1 U6172 ( .A(n5449), .ZN(n5450) );
  AOI21_X1 U6173 ( .B1(n5451), .B2(n5450), .A(n5713), .ZN(n7531) );
  AOI22_X1 U6174 ( .A1(n7369), .A2(n7531), .B1(n6541), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5452) );
  OAI21_X1 U6175 ( .B1(n7532), .B2(n6543), .A(n5452), .ZN(U2852) );
  XNOR2_X1 U6176 ( .A(n5454), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5455)
         );
  XNOR2_X1 U6177 ( .A(n5453), .B(n5455), .ZN(n5929) );
  NOR2_X1 U6178 ( .A1(n7466), .A2(n7461), .ZN(n5456) );
  OAI21_X1 U6179 ( .B1(n6175), .B2(n5457), .A(n5861), .ZN(n7473) );
  INV_X1 U6180 ( .A(n7473), .ZN(n7446) );
  OAI21_X1 U6181 ( .B1(n7176), .B2(n5456), .A(n7446), .ZN(n7464) );
  INV_X1 U6182 ( .A(n5934), .ZN(n5460) );
  INV_X1 U6183 ( .A(n7462), .ZN(n7475) );
  AOI21_X1 U6184 ( .B1(n7471), .B2(n5457), .A(n7475), .ZN(n6180) );
  NOR3_X1 U6185 ( .A1(n6180), .A2(n7461), .A3(n7466), .ZN(n5458) );
  AOI22_X1 U6186 ( .A1(n7460), .A2(REIP_REG_6__SCAN_IN), .B1(n5458), .B2(n4363), .ZN(n5459) );
  OAI21_X1 U6187 ( .B1(n7479), .B2(n5460), .A(n5459), .ZN(n5461) );
  AOI21_X1 U6188 ( .B1(n7464), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n5461), 
        .ZN(n5462) );
  OAI21_X1 U6189 ( .B1(n5929), .B2(n7212), .A(n5462), .ZN(U3012) );
  INV_X1 U6190 ( .A(n5471), .ZN(n5463) );
  NAND2_X1 U6191 ( .A1(n7649), .A2(n5417), .ZN(n6060) );
  NOR2_X1 U6192 ( .A1(n5464), .A2(n6060), .ZN(n5488) );
  AOI21_X1 U6193 ( .B1(n5633), .B2(n3794), .A(n5488), .ZN(n5470) );
  INV_X1 U6194 ( .A(n5470), .ZN(n5468) );
  INV_X1 U6195 ( .A(n5465), .ZN(n5466) );
  OAI21_X1 U6196 ( .B1(n5466), .B2(n4532), .A(n5871), .ZN(n5469) );
  INV_X1 U6197 ( .A(n6060), .ZN(n5631) );
  NAND2_X1 U6198 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5631), .ZN(n5993) );
  INV_X1 U6199 ( .A(n5551), .ZN(n5499) );
  AOI21_X1 U6200 ( .B1(n5679), .B2(n5993), .A(n5499), .ZN(n5467) );
  OAI21_X1 U6201 ( .B1(n5468), .B2(n5469), .A(n5467), .ZN(n5487) );
  OAI22_X1 U6202 ( .A1(n5470), .A2(n5469), .B1(n7669), .B2(n5993), .ZN(n5486)
         );
  AOI22_X1 U6203 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n5487), .B1(n6121), 
        .B2(n5486), .ZN(n5473) );
  NOR3_X4 U6204 ( .A1(n4532), .A2(n5637), .A3(n5471), .ZN(n6040) );
  AOI22_X1 U6205 ( .A1(n6040), .A2(n5756), .B1(n6122), .B2(n5488), .ZN(n5472)
         );
  OAI211_X1 U6206 ( .C1(n5759), .C2(n5983), .A(n5473), .B(n5472), .ZN(U3047)
         );
  AOI22_X1 U6207 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5487), .B1(n6113), 
        .B2(n5486), .ZN(n5475) );
  AOI22_X1 U6208 ( .A1(n6040), .A2(n5751), .B1(n6114), .B2(n5488), .ZN(n5474)
         );
  OAI211_X1 U6209 ( .C1(n5754), .C2(n5983), .A(n5475), .B(n5474), .ZN(U3049)
         );
  AOI22_X1 U6210 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5487), .B1(n6106), 
        .B2(n5486), .ZN(n5477) );
  AOI22_X1 U6211 ( .A1(n6040), .A2(n5746), .B1(n6107), .B2(n5488), .ZN(n5476)
         );
  OAI211_X1 U6212 ( .C1(n5749), .C2(n5983), .A(n5477), .B(n5476), .ZN(U3050)
         );
  AOI22_X1 U6213 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5487), .B1(n6098), 
        .B2(n5486), .ZN(n5479) );
  AOI22_X1 U6214 ( .A1(n6040), .A2(n5741), .B1(n6099), .B2(n5488), .ZN(n5478)
         );
  OAI211_X1 U6215 ( .C1(n5744), .C2(n5983), .A(n5479), .B(n5478), .ZN(U3045)
         );
  AOI22_X1 U6216 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5487), .B1(n6130), 
        .B2(n5486), .ZN(n5481) );
  AOI22_X1 U6217 ( .A1(n6040), .A2(n5765), .B1(n6132), .B2(n5488), .ZN(n5480)
         );
  OAI211_X1 U6218 ( .C1(n5768), .C2(n5983), .A(n5481), .B(n5480), .ZN(U3044)
         );
  AOI22_X1 U6219 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5487), .B1(n6082), 
        .B2(n5486), .ZN(n5483) );
  AOI22_X1 U6220 ( .A1(n6040), .A2(n5726), .B1(n6083), .B2(n5488), .ZN(n5482)
         );
  OAI211_X1 U6221 ( .C1(n5729), .C2(n5983), .A(n5483), .B(n5482), .ZN(U3046)
         );
  AOI22_X1 U6222 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5487), .B1(n6074), 
        .B2(n5486), .ZN(n5485) );
  AOI22_X1 U6223 ( .A1(n6040), .A2(n5731), .B1(n6075), .B2(n5488), .ZN(n5484)
         );
  OAI211_X1 U6224 ( .C1(n5734), .C2(n5983), .A(n5485), .B(n5484), .ZN(U3051)
         );
  AOI22_X1 U6225 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5487), .B1(n6090), 
        .B2(n5486), .ZN(n5490) );
  AOI22_X1 U6226 ( .A1(n6040), .A2(n5736), .B1(n6091), .B2(n5488), .ZN(n5489)
         );
  OAI211_X1 U6227 ( .C1(n5739), .C2(n5983), .A(n5490), .B(n5489), .ZN(U3048)
         );
  OAI222_X1 U6228 ( .A1(n6335), .A2(n5491), .B1(n6392), .B2(n4546), .C1(n6568), 
        .C2(n7523), .ZN(U2886) );
  INV_X1 U6229 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7264) );
  XNOR2_X1 U6230 ( .A(n5194), .B(n5492), .ZN(n7387) );
  OAI222_X1 U6231 ( .A1(n6335), .A2(n5493), .B1(n6392), .B2(n7264), .C1(n6568), 
        .C2(n7387), .ZN(U2888) );
  INV_X1 U6232 ( .A(EAX_REG_6__SCAN_IN), .ZN(n7270) );
  OAI222_X1 U6233 ( .A1(n6335), .A2(n5494), .B1(n6392), .B2(n7270), .C1(n6568), 
        .C2(n5940), .ZN(U2885) );
  INV_X1 U6234 ( .A(EAX_REG_2__SCAN_IN), .ZN(n7262) );
  OAI222_X1 U6235 ( .A1(n6335), .A2(n5496), .B1(n6392), .B2(n7262), .C1(n6568), 
        .C2(n5495), .ZN(U2889) );
  NOR3_X1 U6236 ( .A1(n5417), .A2(n7649), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5501) );
  NOR2_X1 U6237 ( .A1(n5498), .A2(n5679), .ZN(n5502) );
  INV_X1 U6238 ( .A(n5501), .ZN(n5795) );
  NOR2_X1 U6239 ( .A1(n5629), .A2(n5795), .ZN(n5522) );
  AOI21_X1 U6240 ( .B1(n5546), .B2(n5799), .A(n5522), .ZN(n5504) );
  AOI21_X1 U6241 ( .B1(n5502), .B2(n5504), .A(n5499), .ZN(n5500) );
  OAI21_X1 U6242 ( .B1(n5871), .B2(n5501), .A(n5500), .ZN(n5521) );
  INV_X1 U6243 ( .A(n5502), .ZN(n5503) );
  OAI22_X1 U6244 ( .A1(n5504), .A2(n5503), .B1(n7669), .B2(n5795), .ZN(n5520)
         );
  AOI22_X1 U6245 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5521), .B1(n6106), 
        .B2(n5520), .ZN(n5507) );
  AOI22_X1 U6246 ( .A1(n6107), .A2(n5522), .B1(n5746), .B2(n5840), .ZN(n5506)
         );
  OAI211_X1 U6247 ( .C1(n5749), .C2(n5722), .A(n5507), .B(n5506), .ZN(U3130)
         );
  AOI22_X1 U6248 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5521), .B1(n6113), 
        .B2(n5520), .ZN(n5509) );
  AOI22_X1 U6249 ( .A1(n6114), .A2(n5522), .B1(n5751), .B2(n5840), .ZN(n5508)
         );
  OAI211_X1 U6250 ( .C1(n5754), .C2(n5722), .A(n5509), .B(n5508), .ZN(U3129)
         );
  AOI22_X1 U6251 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5521), .B1(n6074), 
        .B2(n5520), .ZN(n5511) );
  AOI22_X1 U6252 ( .A1(n6075), .A2(n5522), .B1(n5731), .B2(n5840), .ZN(n5510)
         );
  OAI211_X1 U6253 ( .C1(n5734), .C2(n5722), .A(n5511), .B(n5510), .ZN(U3131)
         );
  AOI22_X1 U6254 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5521), .B1(n6090), 
        .B2(n5520), .ZN(n5513) );
  AOI22_X1 U6255 ( .A1(n6091), .A2(n5522), .B1(n5736), .B2(n5840), .ZN(n5512)
         );
  OAI211_X1 U6256 ( .C1(n5739), .C2(n5722), .A(n5513), .B(n5512), .ZN(U3128)
         );
  AOI22_X1 U6257 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5521), .B1(n6082), 
        .B2(n5520), .ZN(n5515) );
  AOI22_X1 U6258 ( .A1(n6083), .A2(n5522), .B1(n5726), .B2(n5840), .ZN(n5514)
         );
  OAI211_X1 U6259 ( .C1(n5729), .C2(n5722), .A(n5515), .B(n5514), .ZN(U3126)
         );
  AOI22_X1 U6260 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5521), .B1(n6121), 
        .B2(n5520), .ZN(n5517) );
  AOI22_X1 U6261 ( .A1(n6122), .A2(n5522), .B1(n5756), .B2(n5840), .ZN(n5516)
         );
  OAI211_X1 U6262 ( .C1(n5759), .C2(n5722), .A(n5517), .B(n5516), .ZN(U3127)
         );
  AOI22_X1 U6263 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5521), .B1(n6130), 
        .B2(n5520), .ZN(n5519) );
  AOI22_X1 U6264 ( .A1(n6132), .A2(n5522), .B1(n5765), .B2(n5840), .ZN(n5518)
         );
  OAI211_X1 U6265 ( .C1(n5768), .C2(n5722), .A(n5519), .B(n5518), .ZN(U3124)
         );
  AOI22_X1 U6266 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5521), .B1(n6098), 
        .B2(n5520), .ZN(n5524) );
  AOI22_X1 U6267 ( .A1(n6099), .A2(n5522), .B1(n5741), .B2(n5840), .ZN(n5523)
         );
  OAI211_X1 U6268 ( .C1(n5744), .C2(n5722), .A(n5524), .B(n5523), .ZN(U3125)
         );
  INV_X1 U6269 ( .A(EAX_REG_7__SCAN_IN), .ZN(n7272) );
  OAI222_X1 U6270 ( .A1(n6335), .A2(n5525), .B1(n6392), .B2(n7272), .C1(n6568), 
        .C2(n7532), .ZN(U2884) );
  AOI22_X1 U6271 ( .A1(n7427), .A2(UWORD_REG_14__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5526) );
  OAI21_X1 U6272 ( .B1(n4989), .B2(n5541), .A(n5526), .ZN(U2893) );
  INV_X1 U6273 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5528) );
  AOI22_X1 U6274 ( .A1(n7427), .A2(UWORD_REG_10__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5527) );
  OAI21_X1 U6275 ( .B1(n5528), .B2(n5541), .A(n5527), .ZN(U2897) );
  INV_X1 U6276 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5530) );
  AOI22_X1 U6277 ( .A1(n7427), .A2(UWORD_REG_3__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5529) );
  OAI21_X1 U6278 ( .B1(n5530), .B2(n5541), .A(n5529), .ZN(U2904) );
  AOI22_X1 U6279 ( .A1(n7427), .A2(UWORD_REG_1__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5531) );
  OAI21_X1 U6280 ( .B1(n4720), .B2(n5541), .A(n5531), .ZN(U2906) );
  INV_X1 U6281 ( .A(EAX_REG_29__SCAN_IN), .ZN(n5533) );
  AOI22_X1 U6282 ( .A1(n7427), .A2(UWORD_REG_13__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5532) );
  OAI21_X1 U6283 ( .B1(n5533), .B2(n5541), .A(n5532), .ZN(U2894) );
  INV_X1 U6284 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5535) );
  AOI22_X1 U6285 ( .A1(n7427), .A2(UWORD_REG_12__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5534) );
  OAI21_X1 U6286 ( .B1(n5535), .B2(n5541), .A(n5534), .ZN(U2895) );
  INV_X1 U6287 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5537) );
  AOI22_X1 U6288 ( .A1(n7427), .A2(UWORD_REG_11__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5536) );
  OAI21_X1 U6289 ( .B1(n5537), .B2(n5541), .A(n5536), .ZN(U2896) );
  AOI22_X1 U6290 ( .A1(n7427), .A2(UWORD_REG_4__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5538) );
  OAI21_X1 U6291 ( .B1(n4771), .B2(n5541), .A(n5538), .ZN(U2903) );
  AOI22_X1 U6292 ( .A1(n7427), .A2(UWORD_REG_0__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5539) );
  OAI21_X1 U6293 ( .B1(n4700), .B2(n5541), .A(n5539), .ZN(U2907) );
  INV_X1 U6294 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5542) );
  AOI22_X1 U6295 ( .A1(n7427), .A2(UWORD_REG_2__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5540) );
  OAI21_X1 U6296 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(U2905) );
  AND2_X1 U6297 ( .A1(n5545), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5554)
         );
  AOI21_X1 U6298 ( .B1(n5546), .B2(n5724), .A(n5554), .ZN(n5555) );
  NOR2_X1 U6299 ( .A1(n5679), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5989) );
  INV_X1 U6300 ( .A(n5989), .ZN(n5547) );
  OAI21_X1 U6301 ( .B1(n5548), .B2(n7059), .A(n5547), .ZN(n5549) );
  NAND3_X1 U6302 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5717) );
  AOI22_X1 U6303 ( .A1(n5555), .A2(n5549), .B1(n5679), .B2(n5717), .ZN(n5550)
         );
  NAND2_X1 U6304 ( .A1(n5551), .A2(n5550), .ZN(n5579) );
  NAND2_X1 U6305 ( .A1(n5579), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5560)
         );
  INV_X1 U6306 ( .A(n5554), .ZN(n5581) );
  INV_X1 U6307 ( .A(n5555), .ZN(n5557) );
  INV_X1 U6308 ( .A(n5717), .ZN(n5556) );
  AOI22_X1 U6309 ( .A1(n5557), .A2(n5871), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5556), .ZN(n5580) );
  OAI22_X1 U6310 ( .A1(n6015), .A2(n5581), .B1(n5580), .B2(n6014), .ZN(n5558)
         );
  AOI21_X1 U6311 ( .B1(n6087), .B2(n6067), .A(n5558), .ZN(n5559) );
  OAI211_X1 U6312 ( .C1(n5769), .C2(n6085), .A(n5560), .B(n5559), .ZN(U3142)
         );
  NAND2_X1 U6313 ( .A1(n5579), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5563)
         );
  OAI22_X1 U6314 ( .A1(n6000), .A2(n5581), .B1(n5580), .B2(n5999), .ZN(n5561)
         );
  AOI21_X1 U6315 ( .B1(n6111), .B2(n6067), .A(n5561), .ZN(n5562) );
  OAI211_X1 U6316 ( .C1(n5769), .C2(n6109), .A(n5563), .B(n5562), .ZN(U3146)
         );
  NAND2_X1 U6317 ( .A1(n5579), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5566)
         );
  OAI22_X1 U6318 ( .A1(n6020), .A2(n5581), .B1(n5580), .B2(n6019), .ZN(n5564)
         );
  AOI21_X1 U6319 ( .B1(n6103), .B2(n6067), .A(n5564), .ZN(n5565) );
  OAI211_X1 U6320 ( .C1(n5769), .C2(n6101), .A(n5566), .B(n5565), .ZN(U3141)
         );
  NAND2_X1 U6321 ( .A1(n5579), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5569)
         );
  OAI22_X1 U6322 ( .A1(n6038), .A2(n5581), .B1(n5580), .B2(n6035), .ZN(n5567)
         );
  AOI21_X1 U6323 ( .B1(n6118), .B2(n6067), .A(n5567), .ZN(n5568) );
  OAI211_X1 U6324 ( .C1(n5769), .C2(n6116), .A(n5569), .B(n5568), .ZN(U3145)
         );
  NAND2_X1 U6325 ( .A1(n5579), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5572)
         );
  OAI22_X1 U6326 ( .A1(n6025), .A2(n5581), .B1(n5580), .B2(n6024), .ZN(n5570)
         );
  AOI21_X1 U6327 ( .B1(n6138), .B2(n6067), .A(n5570), .ZN(n5571) );
  OAI211_X1 U6328 ( .C1(n6135), .C2(n5769), .A(n5572), .B(n5571), .ZN(U3140)
         );
  NAND2_X1 U6329 ( .A1(n5579), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5575)
         );
  OAI22_X1 U6330 ( .A1(n6005), .A2(n5581), .B1(n5580), .B2(n6004), .ZN(n5573)
         );
  AOI21_X1 U6331 ( .B1(n6095), .B2(n6067), .A(n5573), .ZN(n5574) );
  OAI211_X1 U6332 ( .C1(n5769), .C2(n6093), .A(n5575), .B(n5574), .ZN(U3144)
         );
  NAND2_X1 U6333 ( .A1(n5579), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5578)
         );
  OAI22_X1 U6334 ( .A1(n6010), .A2(n5581), .B1(n5580), .B2(n6009), .ZN(n5576)
         );
  AOI21_X1 U6335 ( .B1(n6126), .B2(n6067), .A(n5576), .ZN(n5577) );
  OAI211_X1 U6336 ( .C1(n5769), .C2(n6124), .A(n5578), .B(n5577), .ZN(U3143)
         );
  NAND2_X1 U6337 ( .A1(n5579), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5584)
         );
  OAI22_X1 U6338 ( .A1(n6030), .A2(n5581), .B1(n5580), .B2(n6029), .ZN(n5582)
         );
  AOI21_X1 U6339 ( .B1(n6079), .B2(n6067), .A(n5582), .ZN(n5583) );
  OAI211_X1 U6340 ( .C1(n5769), .C2(n6077), .A(n5584), .B(n5583), .ZN(U3147)
         );
  NAND2_X1 U6341 ( .A1(n5619), .A2(n5585), .ZN(n5586) );
  NAND2_X1 U6342 ( .A1(n5586), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5587) );
  NAND2_X1 U6343 ( .A1(n5587), .A2(n5871), .ZN(n5594) );
  INV_X1 U6344 ( .A(n5594), .ZN(n5589) );
  INV_X1 U6345 ( .A(n5592), .ZN(n5588) );
  NAND2_X1 U6346 ( .A1(n5588), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5880) );
  INV_X1 U6347 ( .A(n5880), .ZN(n6069) );
  INV_X1 U6348 ( .A(n5944), .ZN(n6068) );
  NOR2_X1 U6349 ( .A1(n6068), .A2(n7649), .ZN(n5723) );
  OR2_X1 U6350 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5590), .ZN(n5618)
         );
  AOI21_X1 U6351 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n5944), .A(n7669), 
        .ZN(n5718) );
  NAND2_X1 U6352 ( .A1(n5592), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U6353 ( .A1(n5675), .A2(n5801), .ZN(n5875) );
  AOI211_X1 U6354 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5618), .A(n5718), .B(
        n5875), .ZN(n5593) );
  NAND2_X1 U6355 ( .A1(n5617), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5598)
         );
  OAI22_X1 U6356 ( .A1(n5619), .A2(n6116), .B1(n6038), .B2(n5618), .ZN(n5596)
         );
  AOI21_X1 U6357 ( .B1(n6118), .B2(n5621), .A(n5596), .ZN(n5597) );
  OAI211_X1 U6358 ( .C1(n5624), .C2(n6035), .A(n5598), .B(n5597), .ZN(U3105)
         );
  NAND2_X1 U6359 ( .A1(n5617), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5601)
         );
  OAI22_X1 U6360 ( .A1(n5619), .A2(n6093), .B1(n6005), .B2(n5618), .ZN(n5599)
         );
  AOI21_X1 U6361 ( .B1(n6095), .B2(n5621), .A(n5599), .ZN(n5600) );
  OAI211_X1 U6362 ( .C1(n5624), .C2(n6004), .A(n5601), .B(n5600), .ZN(U3104)
         );
  NAND2_X1 U6363 ( .A1(n5617), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5604)
         );
  OAI22_X1 U6364 ( .A1(n5619), .A2(n6109), .B1(n6000), .B2(n5618), .ZN(n5602)
         );
  AOI21_X1 U6365 ( .B1(n6111), .B2(n5621), .A(n5602), .ZN(n5603) );
  OAI211_X1 U6366 ( .C1(n5624), .C2(n5999), .A(n5604), .B(n5603), .ZN(U3106)
         );
  NAND2_X1 U6367 ( .A1(n5617), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5607)
         );
  OAI22_X1 U6368 ( .A1(n5619), .A2(n6085), .B1(n6015), .B2(n5618), .ZN(n5605)
         );
  AOI21_X1 U6369 ( .B1(n6087), .B2(n5621), .A(n5605), .ZN(n5606) );
  OAI211_X1 U6370 ( .C1(n5624), .C2(n6014), .A(n5607), .B(n5606), .ZN(U3102)
         );
  NAND2_X1 U6371 ( .A1(n5617), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5610)
         );
  OAI22_X1 U6372 ( .A1(n5619), .A2(n6077), .B1(n6030), .B2(n5618), .ZN(n5608)
         );
  AOI21_X1 U6373 ( .B1(n6079), .B2(n5621), .A(n5608), .ZN(n5609) );
  OAI211_X1 U6374 ( .C1(n5624), .C2(n6029), .A(n5610), .B(n5609), .ZN(U3107)
         );
  NAND2_X1 U6375 ( .A1(n5617), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5613)
         );
  OAI22_X1 U6376 ( .A1(n5619), .A2(n6101), .B1(n6020), .B2(n5618), .ZN(n5611)
         );
  AOI21_X1 U6377 ( .B1(n6103), .B2(n5621), .A(n5611), .ZN(n5612) );
  OAI211_X1 U6378 ( .C1(n5624), .C2(n6019), .A(n5613), .B(n5612), .ZN(U3101)
         );
  NAND2_X1 U6379 ( .A1(n5617), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5616)
         );
  OAI22_X1 U6380 ( .A1(n5619), .A2(n6135), .B1(n6025), .B2(n5618), .ZN(n5614)
         );
  AOI21_X1 U6381 ( .B1(n6138), .B2(n5621), .A(n5614), .ZN(n5615) );
  OAI211_X1 U6382 ( .C1(n5624), .C2(n6024), .A(n5616), .B(n5615), .ZN(U3100)
         );
  NAND2_X1 U6383 ( .A1(n5617), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5623)
         );
  OAI22_X1 U6384 ( .A1(n5619), .A2(n6124), .B1(n6010), .B2(n5618), .ZN(n5620)
         );
  AOI21_X1 U6385 ( .B1(n6126), .B2(n5621), .A(n5620), .ZN(n5622) );
  OAI211_X1 U6386 ( .C1(n5624), .C2(n6009), .A(n5623), .B(n5622), .ZN(U3103)
         );
  INV_X1 U6387 ( .A(n5625), .ZN(n5627) );
  INV_X1 U6388 ( .A(n5638), .ZN(n5628) );
  NOR3_X1 U6389 ( .A1(n5629), .A2(n6060), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5639) );
  NAND3_X1 U6390 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5631), .A3(n5630), .ZN(
        n5641) );
  OR2_X1 U6391 ( .A1(n5638), .A2(n7696), .ZN(n5634) );
  NAND2_X1 U6392 ( .A1(n5633), .A2(n5632), .ZN(n5640) );
  AND2_X1 U6393 ( .A1(n5634), .A2(n5640), .ZN(n5635) );
  OAI22_X1 U6394 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5641), .B1(n5635), .B2(
        n5679), .ZN(n5636) );
  NAND2_X1 U6395 ( .A1(n5665), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5646) );
  NOR2_X2 U6396 ( .A1(n5638), .A2(n5637), .ZN(n6137) );
  INV_X1 U6397 ( .A(n5639), .ZN(n5667) );
  AOI21_X1 U6398 ( .B1(n5640), .B2(n5667), .A(n5679), .ZN(n5643) );
  INV_X1 U6399 ( .A(n5641), .ZN(n5642) );
  NOR2_X1 U6400 ( .A1(n5643), .A2(n5642), .ZN(n5666) );
  OAI22_X1 U6401 ( .A1(n6005), .A2(n5667), .B1(n5666), .B2(n6004), .ZN(n5644)
         );
  AOI21_X1 U6402 ( .B1(n5736), .B2(n6137), .A(n5644), .ZN(n5645) );
  OAI211_X1 U6403 ( .C1(n6043), .C2(n5739), .A(n5646), .B(n5645), .ZN(U3032)
         );
  NAND2_X1 U6404 ( .A1(n5665), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5649) );
  OAI22_X1 U6405 ( .A1(n6030), .A2(n5667), .B1(n5666), .B2(n6029), .ZN(n5647)
         );
  AOI21_X1 U6406 ( .B1(n5731), .B2(n6137), .A(n5647), .ZN(n5648) );
  OAI211_X1 U6407 ( .C1(n6043), .C2(n5734), .A(n5649), .B(n5648), .ZN(U3035)
         );
  NAND2_X1 U6408 ( .A1(n5665), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5652) );
  OAI22_X1 U6409 ( .A1(n6015), .A2(n5667), .B1(n5666), .B2(n6014), .ZN(n5650)
         );
  AOI21_X1 U6410 ( .B1(n5726), .B2(n6137), .A(n5650), .ZN(n5651) );
  OAI211_X1 U6411 ( .C1(n6043), .C2(n5729), .A(n5652), .B(n5651), .ZN(U3030)
         );
  NAND2_X1 U6412 ( .A1(n5665), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5655) );
  OAI22_X1 U6413 ( .A1(n6038), .A2(n5667), .B1(n5666), .B2(n6035), .ZN(n5653)
         );
  AOI21_X1 U6414 ( .B1(n5751), .B2(n6137), .A(n5653), .ZN(n5654) );
  OAI211_X1 U6415 ( .C1(n6043), .C2(n5754), .A(n5655), .B(n5654), .ZN(U3033)
         );
  NAND2_X1 U6416 ( .A1(n5665), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5658) );
  OAI22_X1 U6417 ( .A1(n6000), .A2(n5667), .B1(n5666), .B2(n5999), .ZN(n5656)
         );
  AOI21_X1 U6418 ( .B1(n5746), .B2(n6137), .A(n5656), .ZN(n5657) );
  OAI211_X1 U6419 ( .C1(n6043), .C2(n5749), .A(n5658), .B(n5657), .ZN(U3034)
         );
  NAND2_X1 U6420 ( .A1(n5665), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5661) );
  OAI22_X1 U6421 ( .A1(n6020), .A2(n5667), .B1(n5666), .B2(n6019), .ZN(n5659)
         );
  AOI21_X1 U6422 ( .B1(n5741), .B2(n6137), .A(n5659), .ZN(n5660) );
  OAI211_X1 U6423 ( .C1(n6043), .C2(n5744), .A(n5661), .B(n5660), .ZN(U3029)
         );
  NAND2_X1 U6424 ( .A1(n5665), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5664) );
  OAI22_X1 U6425 ( .A1(n6010), .A2(n5667), .B1(n5666), .B2(n6009), .ZN(n5662)
         );
  AOI21_X1 U6426 ( .B1(n5756), .B2(n6137), .A(n5662), .ZN(n5663) );
  OAI211_X1 U6427 ( .C1(n6043), .C2(n5759), .A(n5664), .B(n5663), .ZN(U3031)
         );
  NAND2_X1 U6428 ( .A1(n5665), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5670) );
  OAI22_X1 U6429 ( .A1(n6025), .A2(n5667), .B1(n5666), .B2(n6024), .ZN(n5668)
         );
  AOI21_X1 U6430 ( .B1(n5765), .B2(n6137), .A(n5668), .ZN(n5669) );
  OAI211_X1 U6431 ( .C1(n5768), .C2(n6043), .A(n5670), .B(n5669), .ZN(U3028)
         );
  NOR2_X1 U6432 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5671), .ZN(n5678)
         );
  INV_X1 U6433 ( .A(n5800), .ZN(n6059) );
  NOR2_X1 U6434 ( .A1(n5724), .A2(n5679), .ZN(n5716) );
  INV_X1 U6435 ( .A(n5716), .ZN(n5674) );
  INV_X1 U6436 ( .A(n5706), .ZN(n5672) );
  AOI21_X1 U6437 ( .B1(n5672), .B2(n5709), .A(n7696), .ZN(n5673) );
  AOI21_X1 U6438 ( .B1(n6059), .B2(n5674), .A(n5673), .ZN(n5676) );
  NAND2_X1 U6439 ( .A1(n5675), .A2(n5880), .ZN(n5946) );
  NOR2_X1 U6440 ( .A1(n5676), .A2(n5946), .ZN(n5677) );
  NAND2_X1 U6441 ( .A1(n5944), .A2(n7649), .ZN(n5680) );
  NAND2_X1 U6442 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5680), .ZN(n5994) );
  NAND2_X1 U6443 ( .A1(n5702), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5683) );
  INV_X1 U6444 ( .A(n5678), .ZN(n5704) );
  NOR2_X1 U6445 ( .A1(n3667), .A2(n5679), .ZN(n5998) );
  INV_X1 U6446 ( .A(n5801), .ZN(n5949) );
  INV_X1 U6447 ( .A(n5680), .ZN(n5997) );
  AOI22_X1 U6448 ( .A1(n5998), .A2(n5724), .B1(n5949), .B2(n5997), .ZN(n5703)
         );
  OAI22_X1 U6449 ( .A1(n6038), .A2(n5704), .B1(n5703), .B2(n6035), .ZN(n5681)
         );
  AOI21_X1 U6450 ( .B1(n6118), .B2(n5706), .A(n5681), .ZN(n5682) );
  OAI211_X1 U6451 ( .C1(n5709), .C2(n6116), .A(n5683), .B(n5682), .ZN(U3073)
         );
  NAND2_X1 U6452 ( .A1(n5702), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5686) );
  OAI22_X1 U6453 ( .A1(n6000), .A2(n5704), .B1(n5703), .B2(n5999), .ZN(n5684)
         );
  AOI21_X1 U6454 ( .B1(n6111), .B2(n5706), .A(n5684), .ZN(n5685) );
  OAI211_X1 U6455 ( .C1(n5709), .C2(n6109), .A(n5686), .B(n5685), .ZN(U3074)
         );
  NAND2_X1 U6456 ( .A1(n5702), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5689) );
  OAI22_X1 U6457 ( .A1(n6025), .A2(n5704), .B1(n5703), .B2(n6024), .ZN(n5687)
         );
  AOI21_X1 U6458 ( .B1(n6138), .B2(n5706), .A(n5687), .ZN(n5688) );
  OAI211_X1 U6459 ( .C1(n6135), .C2(n5709), .A(n5689), .B(n5688), .ZN(U3068)
         );
  NAND2_X1 U6460 ( .A1(n5702), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5692) );
  OAI22_X1 U6461 ( .A1(n6005), .A2(n5704), .B1(n5703), .B2(n6004), .ZN(n5690)
         );
  AOI21_X1 U6462 ( .B1(n6095), .B2(n5706), .A(n5690), .ZN(n5691) );
  OAI211_X1 U6463 ( .C1(n5709), .C2(n6093), .A(n5692), .B(n5691), .ZN(U3072)
         );
  NAND2_X1 U6464 ( .A1(n5702), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5695) );
  OAI22_X1 U6465 ( .A1(n6030), .A2(n5704), .B1(n5703), .B2(n6029), .ZN(n5693)
         );
  AOI21_X1 U6466 ( .B1(n6079), .B2(n5706), .A(n5693), .ZN(n5694) );
  OAI211_X1 U6467 ( .C1(n5709), .C2(n6077), .A(n5695), .B(n5694), .ZN(U3075)
         );
  NAND2_X1 U6468 ( .A1(n5702), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5698) );
  OAI22_X1 U6469 ( .A1(n6010), .A2(n5704), .B1(n5703), .B2(n6009), .ZN(n5696)
         );
  AOI21_X1 U6470 ( .B1(n6126), .B2(n5706), .A(n5696), .ZN(n5697) );
  OAI211_X1 U6471 ( .C1(n5709), .C2(n6124), .A(n5698), .B(n5697), .ZN(U3071)
         );
  NAND2_X1 U6472 ( .A1(n5702), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5701) );
  OAI22_X1 U6473 ( .A1(n6020), .A2(n5704), .B1(n5703), .B2(n6019), .ZN(n5699)
         );
  AOI21_X1 U6474 ( .B1(n6103), .B2(n5706), .A(n5699), .ZN(n5700) );
  OAI211_X1 U6475 ( .C1(n5709), .C2(n6101), .A(n5701), .B(n5700), .ZN(U3069)
         );
  NAND2_X1 U6476 ( .A1(n5702), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5708) );
  OAI22_X1 U6477 ( .A1(n6015), .A2(n5704), .B1(n5703), .B2(n6014), .ZN(n5705)
         );
  AOI21_X1 U6478 ( .B1(n6087), .B2(n5706), .A(n5705), .ZN(n5707) );
  OAI211_X1 U6479 ( .C1(n5709), .C2(n6085), .A(n5708), .B(n5707), .ZN(U3070)
         );
  AOI21_X1 U6480 ( .B1(n5711), .B2(n5447), .A(n3782), .ZN(n6055) );
  INV_X1 U6481 ( .A(n6055), .ZN(n5924) );
  OR2_X1 U6482 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  AND2_X1 U6483 ( .A1(n6047), .A2(n5714), .ZN(n6205) );
  AOI22_X1 U6484 ( .A1(n7369), .A2(n6205), .B1(n6541), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5715) );
  OAI21_X1 U6485 ( .B1(n5924), .B2(n6539), .A(n5715), .ZN(U2851) );
  AOI21_X1 U6486 ( .B1(n5769), .B2(n5722), .A(n7696), .ZN(n5721) );
  NOR2_X1 U6487 ( .A1(n5716), .A2(n5998), .ZN(n5720) );
  OR2_X1 U6488 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5717), .ZN(n5762)
         );
  AOI211_X1 U6489 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5762), .A(n5718), .B(
        n5946), .ZN(n5719) );
  NAND2_X1 U6490 ( .A1(n5760), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5728)
         );
  AOI22_X1 U6491 ( .A1(n5800), .A2(n5724), .B1(n5949), .B2(n5723), .ZN(n5761)
         );
  OAI22_X1 U6492 ( .A1(n6015), .A2(n5762), .B1(n5761), .B2(n6014), .ZN(n5725)
         );
  AOI21_X1 U6493 ( .B1(n5726), .B2(n5764), .A(n5725), .ZN(n5727) );
  OAI211_X1 U6494 ( .C1(n5769), .C2(n5729), .A(n5728), .B(n5727), .ZN(U3134)
         );
  NAND2_X1 U6495 ( .A1(n5760), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5733)
         );
  OAI22_X1 U6496 ( .A1(n6030), .A2(n5762), .B1(n5761), .B2(n6029), .ZN(n5730)
         );
  AOI21_X1 U6497 ( .B1(n5731), .B2(n5764), .A(n5730), .ZN(n5732) );
  OAI211_X1 U6498 ( .C1(n5769), .C2(n5734), .A(n5733), .B(n5732), .ZN(U3139)
         );
  NAND2_X1 U6499 ( .A1(n5760), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5738)
         );
  OAI22_X1 U6500 ( .A1(n6005), .A2(n5762), .B1(n5761), .B2(n6004), .ZN(n5735)
         );
  AOI21_X1 U6501 ( .B1(n5736), .B2(n5764), .A(n5735), .ZN(n5737) );
  OAI211_X1 U6502 ( .C1(n5769), .C2(n5739), .A(n5738), .B(n5737), .ZN(U3136)
         );
  NAND2_X1 U6503 ( .A1(n5760), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5743)
         );
  OAI22_X1 U6504 ( .A1(n6020), .A2(n5762), .B1(n5761), .B2(n6019), .ZN(n5740)
         );
  AOI21_X1 U6505 ( .B1(n5741), .B2(n5764), .A(n5740), .ZN(n5742) );
  OAI211_X1 U6506 ( .C1(n5769), .C2(n5744), .A(n5743), .B(n5742), .ZN(U3133)
         );
  NAND2_X1 U6507 ( .A1(n5760), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5748)
         );
  OAI22_X1 U6508 ( .A1(n6000), .A2(n5762), .B1(n5761), .B2(n5999), .ZN(n5745)
         );
  AOI21_X1 U6509 ( .B1(n5746), .B2(n5764), .A(n5745), .ZN(n5747) );
  OAI211_X1 U6510 ( .C1(n5769), .C2(n5749), .A(n5748), .B(n5747), .ZN(U3138)
         );
  NAND2_X1 U6511 ( .A1(n5760), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5753)
         );
  OAI22_X1 U6512 ( .A1(n6038), .A2(n5762), .B1(n5761), .B2(n6035), .ZN(n5750)
         );
  AOI21_X1 U6513 ( .B1(n5751), .B2(n5764), .A(n5750), .ZN(n5752) );
  OAI211_X1 U6514 ( .C1(n5769), .C2(n5754), .A(n5753), .B(n5752), .ZN(U3137)
         );
  NAND2_X1 U6515 ( .A1(n5760), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5758)
         );
  OAI22_X1 U6516 ( .A1(n6010), .A2(n5762), .B1(n5761), .B2(n6009), .ZN(n5755)
         );
  AOI21_X1 U6517 ( .B1(n5756), .B2(n5764), .A(n5755), .ZN(n5757) );
  OAI211_X1 U6518 ( .C1(n5769), .C2(n5759), .A(n5758), .B(n5757), .ZN(U3135)
         );
  NAND2_X1 U6519 ( .A1(n5760), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5767)
         );
  OAI22_X1 U6520 ( .A1(n6025), .A2(n5762), .B1(n5761), .B2(n6024), .ZN(n5763)
         );
  AOI21_X1 U6521 ( .B1(n5765), .B2(n5764), .A(n5763), .ZN(n5766) );
  OAI211_X1 U6522 ( .C1(n5769), .C2(n5768), .A(n5767), .B(n5766), .ZN(U3132)
         );
  XNOR2_X1 U6523 ( .A(n5770), .B(n5771), .ZN(n5870) );
  INV_X1 U6524 ( .A(n7532), .ZN(n5774) );
  INV_X1 U6525 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7537) );
  NOR2_X1 U6526 ( .A1(n7477), .A2(n7537), .ZN(n5867) );
  AOI21_X1 U6527 ( .B1(n7396), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5867), 
        .ZN(n5772) );
  OAI21_X1 U6528 ( .B1(n7533), .B2(n7405), .A(n5772), .ZN(n5773) );
  AOI21_X1 U6529 ( .B1(n5774), .B2(n7392), .A(n5773), .ZN(n5775) );
  OAI21_X1 U6530 ( .B1(n5870), .B2(n7626), .A(n5775), .ZN(U2979) );
  INV_X1 U6531 ( .A(REIP_REG_8__SCAN_IN), .ZN(n7298) );
  NOR2_X1 U6532 ( .A1(n5776), .A2(n6275), .ZN(n7527) );
  INV_X1 U6533 ( .A(n7527), .ZN(n5777) );
  NOR2_X1 U6534 ( .A1(n5777), .A2(n7293), .ZN(n7538) );
  NAND3_X1 U6535 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n7538), .ZN(n6187) );
  NAND2_X1 U6536 ( .A1(n7298), .A2(n6187), .ZN(n5791) );
  AND2_X1 U6537 ( .A1(n5778), .A2(n6230), .ZN(n7547) );
  NAND3_X1 U6538 ( .A1(n4017), .A2(n5779), .A3(n6518), .ZN(n5780) );
  AND2_X1 U6539 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  NOR2_X2 U6540 ( .A1(n5849), .A2(n5782), .ZN(n7604) );
  INV_X1 U6541 ( .A(n5783), .ZN(n5784) );
  NAND2_X1 U6542 ( .A1(n7606), .A2(n6054), .ZN(n5788) );
  INV_X1 U6543 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6052) );
  OR2_X1 U6544 ( .A1(n7501), .A2(n7417), .ZN(n7554) );
  OAI21_X1 U6545 ( .B1(n7601), .B2(n6052), .A(n7554), .ZN(n5786) );
  AOI21_X1 U6546 ( .B1(n7520), .B2(n6205), .A(n5786), .ZN(n5787) );
  OAI211_X1 U6547 ( .C1(n5789), .C2(n7577), .A(n5788), .B(n5787), .ZN(n5790)
         );
  AOI21_X1 U6548 ( .B1(n5791), .B2(n7547), .A(n5790), .ZN(n5792) );
  OAI21_X1 U6549 ( .B1(n5924), .B2(n7595), .A(n5792), .ZN(U2819) );
  INV_X1 U6550 ( .A(n5998), .ZN(n6073) );
  NAND2_X1 U6551 ( .A1(n5951), .A2(n5871), .ZN(n5942) );
  INV_X1 U6552 ( .A(n5840), .ZN(n5793) );
  AOI21_X1 U6553 ( .B1(n5793), .B2(n5839), .A(n7696), .ZN(n5794) );
  AOI21_X1 U6554 ( .B1(n6073), .B2(n5942), .A(n5794), .ZN(n5797) );
  NOR2_X1 U6555 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5795), .ZN(n5798)
         );
  NAND2_X1 U6556 ( .A1(n6071), .A2(n6068), .ZN(n5879) );
  NAND2_X1 U6557 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5879), .ZN(n5876) );
  OAI21_X1 U6558 ( .B1(n5798), .B2(n5034), .A(n5876), .ZN(n5796) );
  NOR2_X1 U6559 ( .A1(n5839), .A2(n6124), .ZN(n5807) );
  INV_X1 U6560 ( .A(n5798), .ZN(n5844) );
  NAND2_X1 U6561 ( .A1(n5840), .A2(n6126), .ZN(n5805) );
  NAND2_X1 U6562 ( .A1(n5800), .A2(n5799), .ZN(n5803) );
  OR2_X1 U6563 ( .A1(n5879), .A2(n5801), .ZN(n5802) );
  NAND2_X1 U6564 ( .A1(n5803), .A2(n5802), .ZN(n5841) );
  NAND2_X1 U6565 ( .A1(n5841), .A2(n6121), .ZN(n5804) );
  OAI211_X1 U6566 ( .C1(n6010), .C2(n5844), .A(n5805), .B(n5804), .ZN(n5806)
         );
  AOI211_X1 U6567 ( .C1(n5847), .C2(INSTQUEUE_REG_12__3__SCAN_IN), .A(n5807), 
        .B(n5806), .ZN(n5808) );
  INV_X1 U6568 ( .A(n5808), .ZN(U3119) );
  NOR2_X1 U6569 ( .A1(n5839), .A2(n6135), .ZN(n5812) );
  NAND2_X1 U6570 ( .A1(n5840), .A2(n6138), .ZN(n5810) );
  NAND2_X1 U6571 ( .A1(n5841), .A2(n6130), .ZN(n5809) );
  OAI211_X1 U6572 ( .C1(n6025), .C2(n5844), .A(n5810), .B(n5809), .ZN(n5811)
         );
  AOI211_X1 U6573 ( .C1(n5847), .C2(INSTQUEUE_REG_12__0__SCAN_IN), .A(n5812), 
        .B(n5811), .ZN(n5813) );
  INV_X1 U6574 ( .A(n5813), .ZN(U3116) );
  NOR2_X1 U6575 ( .A1(n5839), .A2(n6077), .ZN(n5817) );
  NAND2_X1 U6576 ( .A1(n5840), .A2(n6079), .ZN(n5815) );
  NAND2_X1 U6577 ( .A1(n5841), .A2(n6074), .ZN(n5814) );
  OAI211_X1 U6578 ( .C1(n6030), .C2(n5844), .A(n5815), .B(n5814), .ZN(n5816)
         );
  AOI211_X1 U6579 ( .C1(n5847), .C2(INSTQUEUE_REG_12__7__SCAN_IN), .A(n5817), 
        .B(n5816), .ZN(n5818) );
  INV_X1 U6580 ( .A(n5818), .ZN(U3123) );
  NOR2_X1 U6581 ( .A1(n5839), .A2(n6116), .ZN(n5822) );
  NAND2_X1 U6582 ( .A1(n5840), .A2(n6118), .ZN(n5820) );
  NAND2_X1 U6583 ( .A1(n5841), .A2(n6113), .ZN(n5819) );
  OAI211_X1 U6584 ( .C1(n6038), .C2(n5844), .A(n5820), .B(n5819), .ZN(n5821)
         );
  AOI211_X1 U6585 ( .C1(n5847), .C2(INSTQUEUE_REG_12__5__SCAN_IN), .A(n5822), 
        .B(n5821), .ZN(n5823) );
  INV_X1 U6586 ( .A(n5823), .ZN(U3121) );
  NOR2_X1 U6587 ( .A1(n5839), .A2(n6093), .ZN(n5827) );
  NAND2_X1 U6588 ( .A1(n5840), .A2(n6095), .ZN(n5825) );
  NAND2_X1 U6589 ( .A1(n5841), .A2(n6090), .ZN(n5824) );
  OAI211_X1 U6590 ( .C1(n6005), .C2(n5844), .A(n5825), .B(n5824), .ZN(n5826)
         );
  AOI211_X1 U6591 ( .C1(n5847), .C2(INSTQUEUE_REG_12__4__SCAN_IN), .A(n5827), 
        .B(n5826), .ZN(n5828) );
  INV_X1 U6592 ( .A(n5828), .ZN(U3120) );
  NOR2_X1 U6593 ( .A1(n5839), .A2(n6085), .ZN(n5832) );
  NAND2_X1 U6594 ( .A1(n5840), .A2(n6087), .ZN(n5830) );
  NAND2_X1 U6595 ( .A1(n5841), .A2(n6082), .ZN(n5829) );
  OAI211_X1 U6596 ( .C1(n6015), .C2(n5844), .A(n5830), .B(n5829), .ZN(n5831)
         );
  AOI211_X1 U6597 ( .C1(n5847), .C2(INSTQUEUE_REG_12__2__SCAN_IN), .A(n5832), 
        .B(n5831), .ZN(n5833) );
  INV_X1 U6598 ( .A(n5833), .ZN(U3118) );
  NOR2_X1 U6599 ( .A1(n5839), .A2(n6109), .ZN(n5837) );
  NAND2_X1 U6600 ( .A1(n5840), .A2(n6111), .ZN(n5835) );
  NAND2_X1 U6601 ( .A1(n5841), .A2(n6106), .ZN(n5834) );
  OAI211_X1 U6602 ( .C1(n6000), .C2(n5844), .A(n5835), .B(n5834), .ZN(n5836)
         );
  AOI211_X1 U6603 ( .C1(n5847), .C2(INSTQUEUE_REG_12__6__SCAN_IN), .A(n5837), 
        .B(n5836), .ZN(n5838) );
  INV_X1 U6604 ( .A(n5838), .ZN(U3122) );
  NOR2_X1 U6605 ( .A1(n5839), .A2(n6101), .ZN(n5846) );
  NAND2_X1 U6606 ( .A1(n5840), .A2(n6103), .ZN(n5843) );
  NAND2_X1 U6607 ( .A1(n5841), .A2(n6098), .ZN(n5842) );
  OAI211_X1 U6608 ( .C1(n6020), .C2(n5844), .A(n5843), .B(n5842), .ZN(n5845)
         );
  AOI211_X1 U6609 ( .C1(n5847), .C2(INSTQUEUE_REG_12__1__SCAN_IN), .A(n5846), 
        .B(n5845), .ZN(n5848) );
  INV_X1 U6610 ( .A(n5848), .ZN(U3117) );
  OAI21_X1 U6611 ( .B1(n4331), .B2(n5849), .A(n7595), .ZN(n7515) );
  INV_X1 U6612 ( .A(n7515), .ZN(n7524) );
  INV_X1 U6613 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5858) );
  INV_X1 U6614 ( .A(n5850), .ZN(n7414) );
  NAND2_X1 U6615 ( .A1(n5851), .A2(n7414), .ZN(n7500) );
  AOI22_X1 U6616 ( .A1(EBX_REG_1__SCAN_IN), .A2(n7604), .B1(n7520), .B2(n5852), 
        .ZN(n5856) );
  OAI22_X1 U6617 ( .A1(n5858), .A2(n7601), .B1(n5853), .B2(n7506), .ZN(n5854)
         );
  AOI21_X1 U6618 ( .B1(n7510), .B2(n7506), .A(n5854), .ZN(n5855) );
  OAI211_X1 U6619 ( .C1(n5089), .C2(n7500), .A(n5856), .B(n5855), .ZN(n5857)
         );
  AOI21_X1 U6620 ( .B1(n7606), .B2(n5858), .A(n5857), .ZN(n5859) );
  OAI21_X1 U6621 ( .B1(n7524), .B2(n5860), .A(n5859), .ZN(U2826) );
  INV_X1 U6622 ( .A(n6175), .ZN(n5864) );
  INV_X1 U6623 ( .A(n5861), .ZN(n5862) );
  AOI21_X1 U6624 ( .B1(n5864), .B2(n5863), .A(n5862), .ZN(n6174) );
  OAI21_X1 U6625 ( .B1(n6203), .B2(n7462), .A(n6174), .ZN(n6212) );
  INV_X1 U6626 ( .A(n6180), .ZN(n7452) );
  AND2_X1 U6627 ( .A1(n7452), .A2(n6203), .ZN(n5866) );
  INV_X1 U6628 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5865) );
  AOI22_X1 U6629 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n6212), .B1(n5866), 
        .B2(n5865), .ZN(n5869) );
  AOI21_X1 U6630 ( .B1(n7495), .B2(n7531), .A(n5867), .ZN(n5868) );
  OAI211_X1 U6631 ( .C1(n5870), .C2(n7212), .A(n5869), .B(n5868), .ZN(U3011)
         );
  NAND2_X1 U6632 ( .A1(n6072), .A2(n5871), .ZN(n6058) );
  INV_X1 U6633 ( .A(n5914), .ZN(n5872) );
  AOI21_X1 U6634 ( .B1(n5872), .B2(n5912), .A(n7696), .ZN(n5873) );
  AOI21_X1 U6635 ( .B1(n6073), .B2(n6058), .A(n5873), .ZN(n5878) );
  NOR2_X1 U6636 ( .A1(n6061), .A2(n5874), .ZN(n5910) );
  OAI211_X1 U6637 ( .C1(n5034), .C2(n5910), .A(n6063), .B(n5876), .ZN(n5877)
         );
  INV_X1 U6638 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5884) );
  OAI22_X1 U6639 ( .A1(n6059), .A2(n6072), .B1(n5880), .B2(n5879), .ZN(n5909)
         );
  AOI22_X1 U6640 ( .A1(n6114), .A2(n5910), .B1(n6113), .B2(n5909), .ZN(n5881)
         );
  OAI21_X1 U6641 ( .B1(n6116), .B2(n5912), .A(n5881), .ZN(n5882) );
  AOI21_X1 U6642 ( .B1(n5914), .B2(n6118), .A(n5882), .ZN(n5883) );
  OAI21_X1 U6643 ( .B1(n5917), .B2(n5884), .A(n5883), .ZN(U3089) );
  INV_X1 U6644 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5888) );
  AOI22_X1 U6645 ( .A1(n6107), .A2(n5910), .B1(n6106), .B2(n5909), .ZN(n5885)
         );
  OAI21_X1 U6646 ( .B1(n6109), .B2(n5912), .A(n5885), .ZN(n5886) );
  AOI21_X1 U6647 ( .B1(n5914), .B2(n6111), .A(n5886), .ZN(n5887) );
  OAI21_X1 U6648 ( .B1(n5917), .B2(n5888), .A(n5887), .ZN(U3090) );
  INV_X1 U6649 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5892) );
  AOI22_X1 U6650 ( .A1(n6075), .A2(n5910), .B1(n6074), .B2(n5909), .ZN(n5889)
         );
  OAI21_X1 U6651 ( .B1(n6077), .B2(n5912), .A(n5889), .ZN(n5890) );
  AOI21_X1 U6652 ( .B1(n5914), .B2(n6079), .A(n5890), .ZN(n5891) );
  OAI21_X1 U6653 ( .B1(n5917), .B2(n5892), .A(n5891), .ZN(U3091) );
  INV_X1 U6654 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5896) );
  AOI22_X1 U6655 ( .A1(n6091), .A2(n5910), .B1(n6090), .B2(n5909), .ZN(n5893)
         );
  OAI21_X1 U6656 ( .B1(n6093), .B2(n5912), .A(n5893), .ZN(n5894) );
  AOI21_X1 U6657 ( .B1(n5914), .B2(n6095), .A(n5894), .ZN(n5895) );
  OAI21_X1 U6658 ( .B1(n5917), .B2(n5896), .A(n5895), .ZN(U3088) );
  INV_X1 U6659 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5900) );
  AOI22_X1 U6660 ( .A1(n6122), .A2(n5910), .B1(n6121), .B2(n5909), .ZN(n5897)
         );
  OAI21_X1 U6661 ( .B1(n6124), .B2(n5912), .A(n5897), .ZN(n5898) );
  AOI21_X1 U6662 ( .B1(n5914), .B2(n6126), .A(n5898), .ZN(n5899) );
  OAI21_X1 U6663 ( .B1(n5917), .B2(n5900), .A(n5899), .ZN(U3087) );
  INV_X1 U6664 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5904) );
  AOI22_X1 U6665 ( .A1(n6083), .A2(n5910), .B1(n6082), .B2(n5909), .ZN(n5901)
         );
  OAI21_X1 U6666 ( .B1(n6085), .B2(n5912), .A(n5901), .ZN(n5902) );
  AOI21_X1 U6667 ( .B1(n5914), .B2(n6087), .A(n5902), .ZN(n5903) );
  OAI21_X1 U6668 ( .B1(n5917), .B2(n5904), .A(n5903), .ZN(U3086) );
  INV_X1 U6669 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5908) );
  AOI22_X1 U6670 ( .A1(n6099), .A2(n5910), .B1(n6098), .B2(n5909), .ZN(n5905)
         );
  OAI21_X1 U6671 ( .B1(n6101), .B2(n5912), .A(n5905), .ZN(n5906) );
  AOI21_X1 U6672 ( .B1(n5914), .B2(n6103), .A(n5906), .ZN(n5907) );
  OAI21_X1 U6673 ( .B1(n5917), .B2(n5908), .A(n5907), .ZN(U3085) );
  INV_X1 U6674 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5916) );
  AOI22_X1 U6675 ( .A1(n6132), .A2(n5910), .B1(n6130), .B2(n5909), .ZN(n5911)
         );
  OAI21_X1 U6676 ( .B1(n6135), .B2(n5912), .A(n5911), .ZN(n5913) );
  AOI21_X1 U6677 ( .B1(n6138), .B2(n5914), .A(n5913), .ZN(n5915) );
  OAI21_X1 U6678 ( .B1(n5917), .B2(n5916), .A(n5915), .ZN(U3084) );
  NOR2_X1 U6679 ( .A1(n7500), .A2(n5918), .ZN(n5920) );
  OAI22_X1 U6680 ( .A1(n7577), .A2(n4344), .B1(n7593), .B2(n7493), .ZN(n5919)
         );
  AOI211_X1 U6681 ( .C1(REIP_REG_0__SCAN_IN), .C2(n6230), .A(n5920), .B(n5919), 
        .ZN(n5922) );
  OAI21_X1 U6682 ( .B1(n7606), .B2(n7608), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5921) );
  OAI211_X1 U6683 ( .C1(n7524), .C2(n5923), .A(n5922), .B(n5921), .ZN(U2827)
         );
  INV_X1 U6684 ( .A(DATAI_8_), .ZN(n5925) );
  INV_X1 U6685 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7274) );
  OAI222_X1 U6686 ( .A1(n6335), .A2(n5925), .B1(n6392), .B2(n7274), .C1(n6568), 
        .C2(n5924), .ZN(U2883) );
  INV_X1 U6687 ( .A(n7405), .ZN(n7038) );
  OAI22_X1 U6688 ( .A1(n7035), .A2(n5932), .B1(n7477), .B2(n7295), .ZN(n5927)
         );
  NOR2_X1 U6689 ( .A1(n5940), .A2(n7059), .ZN(n5926) );
  AOI211_X1 U6690 ( .C1(n7038), .C2(n5931), .A(n5927), .B(n5926), .ZN(n5928)
         );
  OAI21_X1 U6691 ( .B1(n7626), .B2(n5929), .A(n5928), .ZN(U2980) );
  NOR2_X1 U6692 ( .A1(n5930), .A2(n6142), .ZN(n7536) );
  NAND2_X1 U6693 ( .A1(n7606), .A2(n5931), .ZN(n5936) );
  INV_X1 U6694 ( .A(REIP_REG_6__SCAN_IN), .ZN(n7295) );
  AND2_X1 U6695 ( .A1(n7295), .A2(n7538), .ZN(n7535) );
  OAI21_X1 U6696 ( .B1(n7601), .B2(n5932), .A(n7554), .ZN(n5933) );
  AOI211_X1 U6697 ( .C1(n7520), .C2(n5934), .A(n7535), .B(n5933), .ZN(n5935)
         );
  OAI211_X1 U6698 ( .C1(n5937), .C2(n7577), .A(n5936), .B(n5935), .ZN(n5938)
         );
  AOI21_X1 U6699 ( .B1(n7536), .B2(REIP_REG_6__SCAN_IN), .A(n5938), .ZN(n5939)
         );
  OAI21_X1 U6700 ( .B1(n7595), .B2(n5940), .A(n5939), .ZN(U2821) );
  AOI21_X1 U6701 ( .B1(n5948), .B2(n5983), .A(n7696), .ZN(n5941) );
  AOI21_X1 U6702 ( .B1(n5942), .B2(n6059), .A(n5941), .ZN(n5947) );
  NOR2_X1 U6703 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5943), .ZN(n5981)
         );
  OAI21_X1 U6704 ( .B1(n5944), .B2(n6071), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6062) );
  OAI21_X1 U6705 ( .B1(n5981), .B2(n5034), .A(n6062), .ZN(n5945) );
  NOR3_X2 U6706 ( .A1(n5947), .A2(n5946), .A3(n5945), .ZN(n5988) );
  INV_X1 U6707 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U6708 ( .A1(n5949), .A2(n6068), .ZN(n5950) );
  OAI22_X1 U6709 ( .A1(n6073), .A2(n5951), .B1(n6071), .B2(n5950), .ZN(n5980)
         );
  AOI22_X1 U6710 ( .A1(n6099), .A2(n5981), .B1(n6098), .B2(n5980), .ZN(n5952)
         );
  OAI21_X1 U6711 ( .B1(n6101), .B2(n5983), .A(n5952), .ZN(n5953) );
  AOI21_X1 U6712 ( .B1(n6103), .B2(n5985), .A(n5953), .ZN(n5954) );
  OAI21_X1 U6713 ( .B1(n5988), .B2(n5955), .A(n5954), .ZN(U3053) );
  INV_X1 U6714 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5959) );
  AOI22_X1 U6715 ( .A1(n6075), .A2(n5981), .B1(n6074), .B2(n5980), .ZN(n5956)
         );
  OAI21_X1 U6716 ( .B1(n6077), .B2(n5983), .A(n5956), .ZN(n5957) );
  AOI21_X1 U6717 ( .B1(n6079), .B2(n5985), .A(n5957), .ZN(n5958) );
  OAI21_X1 U6718 ( .B1(n5988), .B2(n5959), .A(n5958), .ZN(U3059) );
  INV_X1 U6719 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5963) );
  AOI22_X1 U6720 ( .A1(n6107), .A2(n5981), .B1(n6106), .B2(n5980), .ZN(n5960)
         );
  OAI21_X1 U6721 ( .B1(n6109), .B2(n5983), .A(n5960), .ZN(n5961) );
  AOI21_X1 U6722 ( .B1(n6111), .B2(n5985), .A(n5961), .ZN(n5962) );
  OAI21_X1 U6723 ( .B1(n5988), .B2(n5963), .A(n5962), .ZN(U3058) );
  INV_X1 U6724 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5967) );
  AOI22_X1 U6725 ( .A1(n6114), .A2(n5981), .B1(n6113), .B2(n5980), .ZN(n5964)
         );
  OAI21_X1 U6726 ( .B1(n6116), .B2(n5983), .A(n5964), .ZN(n5965) );
  AOI21_X1 U6727 ( .B1(n6118), .B2(n5985), .A(n5965), .ZN(n5966) );
  OAI21_X1 U6728 ( .B1(n5988), .B2(n5967), .A(n5966), .ZN(U3057) );
  INV_X1 U6729 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5971) );
  AOI22_X1 U6730 ( .A1(n6091), .A2(n5981), .B1(n6090), .B2(n5980), .ZN(n5968)
         );
  OAI21_X1 U6731 ( .B1(n6093), .B2(n5983), .A(n5968), .ZN(n5969) );
  AOI21_X1 U6732 ( .B1(n6095), .B2(n5985), .A(n5969), .ZN(n5970) );
  OAI21_X1 U6733 ( .B1(n5988), .B2(n5971), .A(n5970), .ZN(U3056) );
  INV_X1 U6734 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5975) );
  AOI22_X1 U6735 ( .A1(n6122), .A2(n5981), .B1(n6121), .B2(n5980), .ZN(n5972)
         );
  OAI21_X1 U6736 ( .B1(n6124), .B2(n5983), .A(n5972), .ZN(n5973) );
  AOI21_X1 U6737 ( .B1(n6126), .B2(n5985), .A(n5973), .ZN(n5974) );
  OAI21_X1 U6738 ( .B1(n5988), .B2(n5975), .A(n5974), .ZN(U3055) );
  INV_X1 U6739 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5979) );
  AOI22_X1 U6740 ( .A1(n6083), .A2(n5981), .B1(n6082), .B2(n5980), .ZN(n5976)
         );
  OAI21_X1 U6741 ( .B1(n6085), .B2(n5983), .A(n5976), .ZN(n5977) );
  AOI21_X1 U6742 ( .B1(n6087), .B2(n5985), .A(n5977), .ZN(n5978) );
  OAI21_X1 U6743 ( .B1(n5988), .B2(n5979), .A(n5978), .ZN(U3054) );
  INV_X1 U6744 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5987) );
  AOI22_X1 U6745 ( .A1(n6132), .A2(n5981), .B1(n6130), .B2(n5980), .ZN(n5982)
         );
  OAI21_X1 U6746 ( .B1(n6135), .B2(n5983), .A(n5982), .ZN(n5984) );
  AOI21_X1 U6747 ( .B1(n6138), .B2(n5985), .A(n5984), .ZN(n5986) );
  OAI21_X1 U6748 ( .B1(n5988), .B2(n5987), .A(n5986), .ZN(U3052) );
  INV_X1 U6749 ( .A(n6040), .ZN(n5990) );
  AOI21_X1 U6750 ( .B1(n5990), .B2(n6043), .A(n5989), .ZN(n5991) );
  AOI21_X1 U6751 ( .B1(n3794), .B2(n6374), .A(n5991), .ZN(n5992) );
  NOR2_X1 U6752 ( .A1(n5992), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5995) );
  NOR2_X1 U6753 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5993), .ZN(n5996)
         );
  NAND2_X1 U6754 ( .A1(n6034), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6003) );
  INV_X1 U6755 ( .A(n5996), .ZN(n6037) );
  AOI22_X1 U6756 ( .A1(n5998), .A2(n3794), .B1(n5997), .B2(n6069), .ZN(n6036)
         );
  OAI22_X1 U6757 ( .A1(n6000), .A2(n6037), .B1(n6036), .B2(n5999), .ZN(n6001)
         );
  AOI21_X1 U6758 ( .B1(n6111), .B2(n6040), .A(n6001), .ZN(n6002) );
  OAI211_X1 U6759 ( .C1(n6043), .C2(n6109), .A(n6003), .B(n6002), .ZN(U3042)
         );
  NAND2_X1 U6760 ( .A1(n6034), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6008) );
  OAI22_X1 U6761 ( .A1(n6005), .A2(n6037), .B1(n6036), .B2(n6004), .ZN(n6006)
         );
  AOI21_X1 U6762 ( .B1(n6095), .B2(n6040), .A(n6006), .ZN(n6007) );
  OAI211_X1 U6763 ( .C1(n6043), .C2(n6093), .A(n6008), .B(n6007), .ZN(U3040)
         );
  NAND2_X1 U6764 ( .A1(n6034), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6013) );
  OAI22_X1 U6765 ( .A1(n6010), .A2(n6037), .B1(n6036), .B2(n6009), .ZN(n6011)
         );
  AOI21_X1 U6766 ( .B1(n6126), .B2(n6040), .A(n6011), .ZN(n6012) );
  OAI211_X1 U6767 ( .C1(n6043), .C2(n6124), .A(n6013), .B(n6012), .ZN(U3039)
         );
  NAND2_X1 U6768 ( .A1(n6034), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6018) );
  OAI22_X1 U6769 ( .A1(n6015), .A2(n6037), .B1(n6036), .B2(n6014), .ZN(n6016)
         );
  AOI21_X1 U6770 ( .B1(n6087), .B2(n6040), .A(n6016), .ZN(n6017) );
  OAI211_X1 U6771 ( .C1(n6043), .C2(n6085), .A(n6018), .B(n6017), .ZN(U3038)
         );
  NAND2_X1 U6772 ( .A1(n6034), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6023) );
  OAI22_X1 U6773 ( .A1(n6020), .A2(n6037), .B1(n6036), .B2(n6019), .ZN(n6021)
         );
  AOI21_X1 U6774 ( .B1(n6103), .B2(n6040), .A(n6021), .ZN(n6022) );
  OAI211_X1 U6775 ( .C1(n6043), .C2(n6101), .A(n6023), .B(n6022), .ZN(U3037)
         );
  NAND2_X1 U6776 ( .A1(n6034), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6028) );
  OAI22_X1 U6777 ( .A1(n6025), .A2(n6037), .B1(n6036), .B2(n6024), .ZN(n6026)
         );
  AOI21_X1 U6778 ( .B1(n6138), .B2(n6040), .A(n6026), .ZN(n6027) );
  OAI211_X1 U6779 ( .C1(n6043), .C2(n6135), .A(n6028), .B(n6027), .ZN(U3036)
         );
  NAND2_X1 U6780 ( .A1(n6034), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6033) );
  OAI22_X1 U6781 ( .A1(n6030), .A2(n6037), .B1(n6036), .B2(n6029), .ZN(n6031)
         );
  AOI21_X1 U6782 ( .B1(n6079), .B2(n6040), .A(n6031), .ZN(n6032) );
  OAI211_X1 U6783 ( .C1(n6043), .C2(n6077), .A(n6033), .B(n6032), .ZN(U3043)
         );
  NAND2_X1 U6784 ( .A1(n6034), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6042) );
  OAI22_X1 U6785 ( .A1(n6038), .A2(n6037), .B1(n6036), .B2(n6035), .ZN(n6039)
         );
  AOI21_X1 U6786 ( .B1(n6118), .B2(n6040), .A(n6039), .ZN(n6041) );
  OAI211_X1 U6787 ( .C1(n6043), .C2(n6116), .A(n6042), .B(n6041), .ZN(U3041)
         );
  AOI21_X1 U6788 ( .B1(n6045), .B2(n5710), .A(n6044), .ZN(n7545) );
  INV_X1 U6789 ( .A(n7545), .ZN(n6158) );
  INV_X1 U6790 ( .A(n6165), .ZN(n6046) );
  AOI21_X1 U6791 ( .B1(n6048), .B2(n6047), .A(n6046), .ZN(n7546) );
  AOI22_X1 U6792 ( .A1(n7369), .A2(n7546), .B1(n6541), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n6049) );
  OAI21_X1 U6793 ( .B1(n6158), .B2(n6539), .A(n6049), .ZN(U2850) );
  XNOR2_X1 U6794 ( .A(n6051), .B(n6050), .ZN(n6209) );
  NOR2_X1 U6795 ( .A1(n7477), .A2(n7298), .ZN(n6204) );
  NOR2_X1 U6796 ( .A1(n7035), .A2(n6052), .ZN(n6053) );
  AOI211_X1 U6797 ( .C1(n6054), .C2(n7038), .A(n6204), .B(n6053), .ZN(n6057)
         );
  NAND2_X1 U6798 ( .A1(n6055), .A2(n7392), .ZN(n6056) );
  OAI211_X1 U6799 ( .C1(n6209), .C2(n7626), .A(n6057), .B(n6056), .ZN(U2978)
         );
  OAI21_X1 U6800 ( .B1(n6137), .B2(n6067), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6066) );
  NAND2_X1 U6801 ( .A1(n6059), .A2(n6058), .ZN(n6065) );
  NOR2_X1 U6802 ( .A1(n6061), .A2(n6060), .ZN(n6131) );
  OAI211_X1 U6803 ( .C1(n5034), .C2(n6131), .A(n6063), .B(n6062), .ZN(n6064)
         );
  INV_X1 U6804 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U6805 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  OAI22_X1 U6806 ( .A1(n6073), .A2(n6072), .B1(n6071), .B2(n6070), .ZN(n6129)
         );
  AOI22_X1 U6807 ( .A1(n6075), .A2(n6131), .B1(n6074), .B2(n6129), .ZN(n6076)
         );
  OAI21_X1 U6808 ( .B1(n6077), .B2(n6134), .A(n6076), .ZN(n6078) );
  AOI21_X1 U6809 ( .B1(n6079), .B2(n6137), .A(n6078), .ZN(n6080) );
  OAI21_X1 U6810 ( .B1(n6141), .B2(n6081), .A(n6080), .ZN(U3027) );
  INV_X1 U6811 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6089) );
  AOI22_X1 U6812 ( .A1(n6083), .A2(n6131), .B1(n6082), .B2(n6129), .ZN(n6084)
         );
  OAI21_X1 U6813 ( .B1(n6085), .B2(n6134), .A(n6084), .ZN(n6086) );
  AOI21_X1 U6814 ( .B1(n6087), .B2(n6137), .A(n6086), .ZN(n6088) );
  OAI21_X1 U6815 ( .B1(n6141), .B2(n6089), .A(n6088), .ZN(U3022) );
  INV_X1 U6816 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6097) );
  AOI22_X1 U6817 ( .A1(n6091), .A2(n6131), .B1(n6090), .B2(n6129), .ZN(n6092)
         );
  OAI21_X1 U6818 ( .B1(n6093), .B2(n6134), .A(n6092), .ZN(n6094) );
  AOI21_X1 U6819 ( .B1(n6095), .B2(n6137), .A(n6094), .ZN(n6096) );
  OAI21_X1 U6820 ( .B1(n6141), .B2(n6097), .A(n6096), .ZN(U3024) );
  INV_X1 U6821 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6105) );
  AOI22_X1 U6822 ( .A1(n6099), .A2(n6131), .B1(n6098), .B2(n6129), .ZN(n6100)
         );
  OAI21_X1 U6823 ( .B1(n6101), .B2(n6134), .A(n6100), .ZN(n6102) );
  AOI21_X1 U6824 ( .B1(n6103), .B2(n6137), .A(n6102), .ZN(n6104) );
  OAI21_X1 U6825 ( .B1(n6141), .B2(n6105), .A(n6104), .ZN(U3021) );
  AOI22_X1 U6826 ( .A1(n6107), .A2(n6131), .B1(n6106), .B2(n6129), .ZN(n6108)
         );
  OAI21_X1 U6827 ( .B1(n6109), .B2(n6134), .A(n6108), .ZN(n6110) );
  AOI21_X1 U6828 ( .B1(n6111), .B2(n6137), .A(n6110), .ZN(n6112) );
  OAI21_X1 U6829 ( .B1(n6141), .B2(n4178), .A(n6112), .ZN(U3026) );
  INV_X1 U6830 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6120) );
  AOI22_X1 U6831 ( .A1(n6114), .A2(n6131), .B1(n6113), .B2(n6129), .ZN(n6115)
         );
  OAI21_X1 U6832 ( .B1(n6116), .B2(n6134), .A(n6115), .ZN(n6117) );
  AOI21_X1 U6833 ( .B1(n6118), .B2(n6137), .A(n6117), .ZN(n6119) );
  OAI21_X1 U6834 ( .B1(n6141), .B2(n6120), .A(n6119), .ZN(U3025) );
  INV_X1 U6835 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6128) );
  AOI22_X1 U6836 ( .A1(n6122), .A2(n6131), .B1(n6121), .B2(n6129), .ZN(n6123)
         );
  OAI21_X1 U6837 ( .B1(n6124), .B2(n6134), .A(n6123), .ZN(n6125) );
  AOI21_X1 U6838 ( .B1(n6126), .B2(n6137), .A(n6125), .ZN(n6127) );
  OAI21_X1 U6839 ( .B1(n6141), .B2(n6128), .A(n6127), .ZN(U3023) );
  INV_X1 U6840 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6140) );
  AOI22_X1 U6841 ( .A1(n6132), .A2(n6131), .B1(n6130), .B2(n6129), .ZN(n6133)
         );
  OAI21_X1 U6842 ( .B1(n6135), .B2(n6134), .A(n6133), .ZN(n6136) );
  AOI21_X1 U6843 ( .B1(n6138), .B2(n6137), .A(n6136), .ZN(n6139) );
  OAI21_X1 U6844 ( .B1(n6141), .B2(n6140), .A(n6139), .ZN(U3020) );
  NOR2_X1 U6845 ( .A1(n6143), .A2(n6142), .ZN(n6370) );
  INV_X1 U6846 ( .A(n6370), .ZN(n6157) );
  INV_X1 U6847 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6156) );
  OAI22_X1 U6848 ( .A1(n6144), .A2(n7577), .B1(n7630), .B2(n7500), .ZN(n6145)
         );
  INV_X1 U6849 ( .A(n6145), .ZN(n6146) );
  OAI211_X1 U6850 ( .C1(n7601), .C2(n6147), .A(n7554), .B(n6146), .ZN(n6148)
         );
  AOI21_X1 U6851 ( .B1(n7610), .B2(n7444), .A(n6148), .ZN(n6151) );
  OR3_X1 U6852 ( .A1(n6149), .A2(REIP_REG_4__SCAN_IN), .A3(n6275), .ZN(n6150)
         );
  OAI211_X1 U6853 ( .C1(n7579), .C2(n6152), .A(n6151), .B(n6150), .ZN(n6153)
         );
  AOI21_X1 U6854 ( .B1(n6154), .B2(n7515), .A(n6153), .ZN(n6155) );
  OAI21_X1 U6855 ( .B1(n6157), .B2(n6156), .A(n6155), .ZN(U2823) );
  INV_X1 U6856 ( .A(DATAI_9_), .ZN(n6159) );
  INV_X1 U6857 ( .A(EAX_REG_9__SCAN_IN), .ZN(n7276) );
  OAI222_X1 U6858 ( .A1(n6335), .A2(n6159), .B1(n6392), .B2(n7276), .C1(n6568), 
        .C2(n6158), .ZN(U2882) );
  INV_X1 U6859 ( .A(n6160), .ZN(n6163) );
  INV_X1 U6860 ( .A(n6044), .ZN(n6162) );
  AOI21_X1 U6861 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(n6220) );
  INV_X1 U6862 ( .A(n6220), .ZN(n6201) );
  AND2_X1 U6863 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  OR2_X1 U6864 ( .A1(n6198), .A2(n6166), .ZN(n6222) );
  INV_X1 U6865 ( .A(n6222), .ZN(n6167) );
  AOI22_X1 U6866 ( .A1(n7369), .A2(n6167), .B1(n6541), .B2(EBX_REG_10__SCAN_IN), .ZN(n6168) );
  OAI21_X1 U6867 ( .B1(n6201), .B2(n6543), .A(n6168), .ZN(U2849) );
  XNOR2_X1 U6868 ( .A(n6169), .B(n6170), .ZN(n6185) );
  AND2_X1 U6869 ( .A1(n7460), .A2(REIP_REG_9__SCAN_IN), .ZN(n6182) );
  AOI21_X1 U6870 ( .B1(n7396), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6182), 
        .ZN(n6171) );
  OAI21_X1 U6871 ( .B1(n7543), .B2(n7405), .A(n6171), .ZN(n6172) );
  AOI21_X1 U6872 ( .B1(n7545), .B2(n7392), .A(n6172), .ZN(n6173) );
  OAI21_X1 U6873 ( .B1(n6185), .B2(n7626), .A(n6173), .ZN(U2977) );
  OAI21_X1 U6874 ( .B1(n6175), .B2(n6207), .A(n6174), .ZN(n6176) );
  INV_X1 U6875 ( .A(n6176), .ZN(n6252) );
  INV_X1 U6876 ( .A(n6179), .ZN(n6177) );
  OR2_X1 U6877 ( .A1(n7462), .A2(n6177), .ZN(n6178) );
  NAND2_X1 U6878 ( .A1(n6252), .A2(n6178), .ZN(n6251) );
  NOR2_X1 U6879 ( .A1(n6180), .A2(n6179), .ZN(n6223) );
  AOI22_X1 U6880 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n6251), .B1(n6223), 
        .B2(n6181), .ZN(n6184) );
  AOI21_X1 U6881 ( .B1(n7495), .B2(n7546), .A(n6182), .ZN(n6183) );
  OAI211_X1 U6882 ( .C1(n6185), .C2(n7212), .A(n6184), .B(n6183), .ZN(U3009)
         );
  OAI22_X1 U6883 ( .A1(n7577), .A2(n6186), .B1(n7593), .B2(n6222), .ZN(n6191)
         );
  NOR2_X1 U6884 ( .A1(n7298), .A2(n6187), .ZN(n6192) );
  NAND3_X1 U6885 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6192), .A3(n7302), .ZN(n6188) );
  OAI211_X1 U6886 ( .C1(n7601), .C2(n6189), .A(n7554), .B(n6188), .ZN(n6190)
         );
  AOI211_X1 U6887 ( .C1(n6216), .C2(n7606), .A(n6191), .B(n6190), .ZN(n6194)
         );
  AND2_X1 U6888 ( .A1(n7300), .A2(n6192), .ZN(n7551) );
  OAI21_X1 U6889 ( .B1(n7551), .B2(n7547), .A(REIP_REG_10__SCAN_IN), .ZN(n6193) );
  OAI211_X1 U6890 ( .C1(n7595), .C2(n6201), .A(n6194), .B(n6193), .ZN(U2817)
         );
  OAI21_X1 U6891 ( .B1(n6161), .B2(n6196), .A(n6195), .ZN(n6271) );
  OR2_X1 U6892 ( .A1(n6198), .A2(n6197), .ZN(n6199) );
  AND2_X1 U6893 ( .A1(n6278), .A2(n6199), .ZN(n7216) );
  AOI22_X1 U6894 ( .A1(n7369), .A2(n7216), .B1(n6541), .B2(EBX_REG_11__SCAN_IN), .ZN(n6200) );
  OAI21_X1 U6895 ( .B1(n6271), .B2(n6543), .A(n6200), .ZN(U2848) );
  INV_X1 U6896 ( .A(DATAI_10_), .ZN(n6202) );
  INV_X1 U6897 ( .A(EAX_REG_10__SCAN_IN), .ZN(n7278) );
  OAI222_X1 U6898 ( .A1(n6335), .A2(n6202), .B1(n6392), .B2(n7278), .C1(n6568), 
        .C2(n6201), .ZN(U2881) );
  OAI211_X1 U6899 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6203), .B(n7452), .ZN(n6208) );
  AOI21_X1 U6900 ( .B1(n7495), .B2(n6205), .A(n6204), .ZN(n6206) );
  OAI21_X1 U6901 ( .B1(n6208), .B2(n6207), .A(n6206), .ZN(n6211) );
  NOR2_X1 U6902 ( .A1(n6209), .A2(n7212), .ZN(n6210) );
  AOI211_X1 U6903 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n6212), .A(n6211), 
        .B(n6210), .ZN(n6213) );
  INV_X1 U6904 ( .A(n6213), .ZN(U3010) );
  XNOR2_X1 U6905 ( .A(n6214), .B(n6215), .ZN(n6228) );
  INV_X1 U6906 ( .A(n6216), .ZN(n6218) );
  AOI22_X1 U6907 ( .A1(n7396), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n7460), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n6217) );
  OAI21_X1 U6908 ( .B1(n7405), .B2(n6218), .A(n6217), .ZN(n6219) );
  AOI21_X1 U6909 ( .B1(n6220), .B2(n7392), .A(n6219), .ZN(n6221) );
  OAI21_X1 U6910 ( .B1(n6228), .B2(n7626), .A(n6221), .ZN(U2976) );
  OAI22_X1 U6911 ( .A1(n7479), .A2(n6222), .B1(n7302), .B2(n7477), .ZN(n6226)
         );
  OAI211_X1 U6912 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6223), .B(n6250), .ZN(n6224) );
  INV_X1 U6913 ( .A(n6224), .ZN(n6225) );
  AOI211_X1 U6914 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6251), .A(n6226), .B(n6225), .ZN(n6227) );
  OAI21_X1 U6915 ( .B1(n6228), .B2(n7212), .A(n6227), .ZN(U3008) );
  INV_X1 U6916 ( .A(DATAI_11_), .ZN(n6229) );
  INV_X1 U6917 ( .A(EAX_REG_11__SCAN_IN), .ZN(n7280) );
  OAI222_X1 U6918 ( .A1(n6335), .A2(n6229), .B1(n6392), .B2(n7280), .C1(n6568), 
        .C2(n6271), .ZN(U2880) );
  INV_X1 U6919 ( .A(n6267), .ZN(n6238) );
  INV_X1 U6920 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6236) );
  AND2_X1 U6921 ( .A1(n6274), .A2(n6230), .ZN(n7563) );
  NAND2_X1 U6922 ( .A1(n7510), .A2(n6231), .ZN(n6233) );
  AOI22_X1 U6923 ( .A1(n7610), .A2(n7216), .B1(n7604), .B2(EBX_REG_11__SCAN_IN), .ZN(n6232) );
  OAI21_X1 U6924 ( .B1(REIP_REG_11__SCAN_IN), .B2(n6233), .A(n6232), .ZN(n6234) );
  AOI211_X1 U6925 ( .C1(REIP_REG_11__SCAN_IN), .C2(n7563), .A(n6234), .B(n7582), .ZN(n6235) );
  OAI21_X1 U6926 ( .B1(n6236), .B2(n7601), .A(n6235), .ZN(n6237) );
  AOI21_X1 U6927 ( .B1(n6238), .B2(n7606), .A(n6237), .ZN(n6239) );
  OAI21_X1 U6928 ( .B1(n6271), .B2(n7595), .A(n6239), .ZN(U2816) );
  AOI21_X1 U6929 ( .B1(n6241), .B2(n6195), .A(n6240), .ZN(n7562) );
  INV_X1 U6930 ( .A(n7562), .ZN(n6245) );
  OAI222_X1 U6931 ( .A1(n6245), .A2(n6568), .B1(n6335), .B2(n6242), .C1(n6392), 
        .C2(n4625), .ZN(U2879) );
  INV_X1 U6932 ( .A(n6277), .ZN(n6243) );
  XNOR2_X1 U6933 ( .A(n6278), .B(n6243), .ZN(n7557) );
  INV_X1 U6934 ( .A(n7557), .ZN(n6244) );
  OAI222_X1 U6935 ( .A1(n6245), .A2(n6543), .B1(n7559), .B2(n7376), .C1(n7372), 
        .C2(n6244), .ZN(U2847) );
  XNOR2_X1 U6936 ( .A(n6246), .B(n6247), .ZN(n6263) );
  INV_X1 U6937 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6248) );
  NOR2_X1 U6938 ( .A1(n7477), .A2(n6248), .ZN(n6260) );
  NAND2_X1 U6939 ( .A1(n6249), .A2(n7462), .ZN(n7177) );
  OR2_X1 U6940 ( .A1(n6251), .A2(n6250), .ZN(n6254) );
  NAND2_X1 U6941 ( .A1(n6252), .A2(n7176), .ZN(n6253) );
  NAND2_X1 U6942 ( .A1(n6254), .A2(n6253), .ZN(n7174) );
  INV_X1 U6943 ( .A(n7174), .ZN(n7217) );
  AOI21_X1 U6944 ( .B1(n7177), .B2(n6324), .A(n7217), .ZN(n6256) );
  AOI21_X1 U6945 ( .B1(n7219), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6255) );
  NOR2_X1 U6946 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  AOI211_X1 U6947 ( .C1(n7495), .C2(n7557), .A(n6260), .B(n6257), .ZN(n6258)
         );
  OAI21_X1 U6948 ( .B1(n6263), .B2(n7212), .A(n6258), .ZN(U3006) );
  NOR2_X1 U6949 ( .A1(n7035), .A2(n7555), .ZN(n6259) );
  AOI211_X1 U6950 ( .C1(n7038), .C2(n7564), .A(n6260), .B(n6259), .ZN(n6262)
         );
  NAND2_X1 U6951 ( .A1(n7562), .A2(n7392), .ZN(n6261) );
  OAI211_X1 U6952 ( .C1(n6263), .C2(n7626), .A(n6262), .B(n6261), .ZN(U2974)
         );
  XOR2_X1 U6953 ( .A(n6264), .B(n6265), .Z(n7214) );
  NAND2_X1 U6954 ( .A1(n7214), .A2(n7402), .ZN(n6270) );
  INV_X1 U6955 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6266) );
  NOR2_X1 U6956 ( .A1(n7477), .A2(n6266), .ZN(n7215) );
  NOR2_X1 U6957 ( .A1(n7405), .A2(n6267), .ZN(n6268) );
  AOI211_X1 U6958 ( .C1(n7396), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n7215), 
        .B(n6268), .ZN(n6269) );
  OAI211_X1 U6959 ( .C1(n7059), .C2(n6271), .A(n6270), .B(n6269), .ZN(U2975)
         );
  XNOR2_X1 U6960 ( .A(n6272), .B(n6273), .ZN(n6301) );
  INV_X1 U6961 ( .A(n6297), .ZN(n6286) );
  OR2_X1 U6962 ( .A1(n6275), .A2(n6274), .ZN(n6306) );
  INV_X1 U6963 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U6964 ( .A1(n6296), .A2(REIP_REG_12__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U6965 ( .B1(n6278), .B2(n6277), .A(n6276), .ZN(n6279) );
  NAND2_X1 U6966 ( .A1(n6279), .A2(n6308), .ZN(n6290) );
  INV_X1 U6967 ( .A(n6290), .ZN(n7437) );
  AOI22_X1 U6968 ( .A1(n7610), .A2(n7437), .B1(n7604), .B2(EBX_REG_13__SCAN_IN), .ZN(n6280) );
  OAI211_X1 U6969 ( .C1(n7601), .C2(n6281), .A(n6280), .B(n7554), .ZN(n6282)
         );
  INV_X1 U6970 ( .A(n6282), .ZN(n6283) );
  OAI21_X1 U6971 ( .B1(n6306), .B2(n6284), .A(n6283), .ZN(n6285) );
  AOI21_X1 U6972 ( .B1(n7606), .B2(n6286), .A(n6285), .ZN(n6288) );
  NOR2_X1 U6973 ( .A1(n6306), .A2(REIP_REG_12__SCAN_IN), .ZN(n7561) );
  OAI21_X1 U6974 ( .B1(n7561), .B2(n7563), .A(REIP_REG_13__SCAN_IN), .ZN(n6287) );
  OAI211_X1 U6975 ( .C1(n6301), .C2(n7595), .A(n6288), .B(n6287), .ZN(U2814)
         );
  INV_X1 U6976 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6289) );
  OAI222_X1 U6977 ( .A1(n6290), .A2(n7372), .B1(n6289), .B2(n7376), .C1(n6539), 
        .C2(n6301), .ZN(U2846) );
  INV_X1 U6978 ( .A(DATAI_13_), .ZN(n6291) );
  OAI222_X1 U6979 ( .A1(n6335), .A2(n6291), .B1(n6568), .B2(n6301), .C1(n7283), 
        .C2(n6392), .ZN(U2878) );
  NAND2_X1 U6980 ( .A1(n6292), .A2(n6293), .ZN(n6294) );
  NAND2_X1 U6981 ( .A1(n6295), .A2(n6294), .ZN(n7439) );
  NAND2_X1 U6982 ( .A1(n7439), .A2(n7402), .ZN(n6300) );
  NOR2_X1 U6983 ( .A1(n7477), .A2(n6296), .ZN(n7436) );
  NOR2_X1 U6984 ( .A1(n7405), .A2(n6297), .ZN(n6298) );
  AOI211_X1 U6985 ( .C1(n7396), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n7436), 
        .B(n6298), .ZN(n6299) );
  OAI211_X1 U6986 ( .C1(n6301), .C2(n7059), .A(n6300), .B(n6299), .ZN(U2973)
         );
  OAI21_X1 U6987 ( .B1(n6302), .B2(n6304), .A(n6303), .ZN(n6344) );
  INV_X1 U6988 ( .A(n6346), .ZN(n6315) );
  NOR3_X1 U6989 ( .A1(n6306), .A2(REIP_REG_14__SCAN_IN), .A3(n6305), .ZN(n6314) );
  OAI21_X1 U6990 ( .B1(n7601), .B2(n6307), .A(n7554), .ZN(n6311) );
  AOI21_X1 U6991 ( .B1(n6309), .B2(n6308), .A(n6339), .ZN(n6330) );
  INV_X1 U6992 ( .A(n6330), .ZN(n6333) );
  NOR2_X1 U6993 ( .A1(n7593), .A2(n6333), .ZN(n6310) );
  AOI211_X1 U6994 ( .C1(n7567), .C2(REIP_REG_14__SCAN_IN), .A(n6311), .B(n6310), .ZN(n6312) );
  OAI21_X1 U6995 ( .B1(n4394), .B2(n7577), .A(n6312), .ZN(n6313) );
  AOI211_X1 U6996 ( .C1(n7606), .C2(n6315), .A(n6314), .B(n6313), .ZN(n6316)
         );
  OAI21_X1 U6997 ( .B1(n6344), .B2(n7595), .A(n6316), .ZN(U2813) );
  XNOR2_X1 U6998 ( .A(n7030), .B(n6318), .ZN(n6319) );
  XNOR2_X1 U6999 ( .A(n6317), .B(n6319), .ZN(n6350) );
  NAND2_X1 U7000 ( .A1(n6321), .A2(n6320), .ZN(n7442) );
  AOI21_X1 U7001 ( .B1(n6323), .B2(n6322), .A(n7442), .ZN(n6326) );
  AOI22_X1 U7002 ( .A1(n7492), .A2(n6327), .B1(n7490), .B2(n6324), .ZN(n6325)
         );
  NAND2_X1 U7003 ( .A1(n7174), .A2(n6325), .ZN(n7438) );
  OAI21_X1 U7004 ( .B1(n6326), .B2(n7438), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n6332) );
  NOR2_X1 U7005 ( .A1(n7477), .A2(n7308), .ZN(n6329) );
  INV_X1 U7006 ( .A(n7219), .ZN(n7443) );
  NOR3_X1 U7007 ( .A1(n7443), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n6327), 
        .ZN(n6328) );
  AOI211_X1 U7008 ( .C1(n7495), .C2(n6330), .A(n6329), .B(n6328), .ZN(n6331)
         );
  OAI211_X1 U7009 ( .C1(n6350), .C2(n7212), .A(n6332), .B(n6331), .ZN(U3004)
         );
  OAI222_X1 U7010 ( .A1(n6344), .A2(n6543), .B1(n7376), .B2(n4394), .C1(n6333), 
        .C2(n7372), .ZN(U2845) );
  INV_X1 U7011 ( .A(DATAI_14_), .ZN(n6334) );
  OAI222_X1 U7012 ( .A1(n6335), .A2(n6334), .B1(n6392), .B2(n4670), .C1(n6568), 
        .C2(n6344), .ZN(U2877) );
  AOI21_X1 U7013 ( .B1(n6337), .B2(n6303), .A(n6336), .ZN(n7572) );
  INV_X1 U7014 ( .A(n7572), .ZN(n6343) );
  AOI22_X1 U7015 ( .A1(n6569), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n7735), .ZN(n6338) );
  OAI21_X1 U7016 ( .B1(n6343), .B2(n6568), .A(n6338), .ZN(U2876) );
  INV_X1 U7017 ( .A(n6339), .ZN(n6340) );
  AOI21_X1 U7018 ( .B1(n6341), .B2(n6340), .A(n6355), .ZN(n7569) );
  AOI22_X1 U7019 ( .A1(n7569), .A2(n7369), .B1(EBX_REG_15__SCAN_IN), .B2(n6541), .ZN(n6342) );
  OAI21_X1 U7020 ( .B1(n6343), .B2(n6543), .A(n6342), .ZN(U2844) );
  INV_X1 U7021 ( .A(n6344), .ZN(n6348) );
  AOI22_X1 U7022 ( .A1(n7396), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n7460), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n6345) );
  OAI21_X1 U7023 ( .B1(n6346), .B2(n7405), .A(n6345), .ZN(n6347) );
  AOI21_X1 U7024 ( .B1(n6348), .B2(n7392), .A(n6347), .ZN(n6349) );
  OAI21_X1 U7025 ( .B1(n6350), .B2(n7626), .A(n6349), .ZN(U2972) );
  OR2_X1 U7026 ( .A1(n6336), .A2(n6352), .ZN(n6353) );
  NAND2_X1 U7027 ( .A1(n6351), .A2(n6353), .ZN(n7058) );
  INV_X1 U7028 ( .A(n7054), .ZN(n6362) );
  OAI21_X1 U7029 ( .B1(n6355), .B2(n6354), .A(n6508), .ZN(n7198) );
  OAI211_X1 U7030 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n7570), .B(n6356), .ZN(n6360) );
  OAI22_X1 U7031 ( .A1(n6357), .A2(n7601), .B1(n4402), .B2(n7577), .ZN(n6358)
         );
  AOI211_X1 U7032 ( .C1(REIP_REG_16__SCAN_IN), .C2(n7567), .A(n6358), .B(n7582), .ZN(n6359) );
  OAI211_X1 U7033 ( .C1(n7198), .C2(n7593), .A(n6360), .B(n6359), .ZN(n6361)
         );
  AOI21_X1 U7034 ( .B1(n7606), .B2(n6362), .A(n6361), .ZN(n6363) );
  OAI21_X1 U7035 ( .B1(n7058), .B2(n7595), .A(n6363), .ZN(U2811) );
  AOI22_X1 U7036 ( .A1(n7733), .A2(DATAI_0_), .B1(n7735), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U7037 ( .A1(n7736), .A2(DATAI_16_), .ZN(n6364) );
  OAI211_X1 U7038 ( .C1(n7058), .C2(n6568), .A(n6365), .B(n6364), .ZN(U2875)
         );
  OAI222_X1 U7039 ( .A1(n7198), .A2(n7372), .B1(n7376), .B2(n4402), .C1(n7058), 
        .C2(n6539), .ZN(U2843) );
  OR2_X1 U7040 ( .A1(n5205), .A2(n6366), .ZN(n6367) );
  AND2_X1 U7041 ( .A1(n6368), .A2(n6367), .ZN(n7454) );
  AOI22_X1 U7042 ( .A1(n7369), .A2(n7454), .B1(n6541), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n6369) );
  OAI21_X1 U7043 ( .B1(n7387), .B2(n6543), .A(n6369), .ZN(U2856) );
  OAI21_X1 U7044 ( .B1(n6371), .B2(REIP_REG_3__SCAN_IN), .A(n6370), .ZN(n6378)
         );
  INV_X1 U7045 ( .A(n7395), .ZN(n6376) );
  AOI22_X1 U7046 ( .A1(n7520), .A2(n7454), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n7608), .ZN(n6373) );
  NAND2_X1 U7047 ( .A1(n7604), .A2(EBX_REG_3__SCAN_IN), .ZN(n6372) );
  OAI211_X1 U7048 ( .C1(n6374), .C2(n7500), .A(n6373), .B(n6372), .ZN(n6375)
         );
  AOI21_X1 U7049 ( .B1(n6376), .B2(n7606), .A(n6375), .ZN(n6377) );
  OAI211_X1 U7050 ( .C1(n7524), .C2(n7387), .A(n6378), .B(n6377), .ZN(U2824)
         );
  INV_X1 U7051 ( .A(n6940), .ZN(n6390) );
  AOI22_X1 U7052 ( .A1(n6381), .A2(n7369), .B1(EBX_REG_30__SCAN_IN), .B2(n6541), .ZN(n6379) );
  OAI21_X1 U7053 ( .B1(n6390), .B2(n6543), .A(n6379), .ZN(U2829) );
  INV_X1 U7054 ( .A(n6380), .ZN(n6411) );
  NAND2_X1 U7055 ( .A1(n6381), .A2(n7520), .ZN(n6387) );
  INV_X1 U7056 ( .A(n6382), .ZN(n6938) );
  NOR2_X1 U7057 ( .A1(n7579), .A2(n6938), .ZN(n6385) );
  AOI22_X1 U7058 ( .A1(n7604), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n7608), .ZN(n6383) );
  INV_X1 U7059 ( .A(n6383), .ZN(n6384) );
  AND2_X1 U7060 ( .A1(n6392), .A2(n6391), .ZN(n6393) );
  NAND2_X1 U7061 ( .A1(n6394), .A2(n6393), .ZN(n6396) );
  AOI22_X1 U7062 ( .A1(n7736), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7735), .ZN(n6395) );
  NAND2_X1 U7063 ( .A1(n6396), .A2(n6395), .ZN(U2860) );
  OAI211_X1 U7064 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5084), .A(n6398), .B(
        n6397), .ZN(n6400) );
  NAND2_X1 U7065 ( .A1(n7254), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6399) );
  OAI211_X1 U7066 ( .C1(n6401), .C2(n5089), .A(n6400), .B(n6399), .ZN(U3464)
         );
  AOI21_X1 U7067 ( .B1(n6403), .B2(n5051), .A(n6402), .ZN(n6950) );
  INV_X1 U7068 ( .A(n6950), .ZN(n6547) );
  INV_X1 U7069 ( .A(n6404), .ZN(n6405) );
  AOI21_X1 U7070 ( .B1(n6407), .B2(n6406), .A(n6405), .ZN(n7083) );
  AOI22_X1 U7071 ( .A1(n7604), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n7608), .ZN(n6408) );
  OAI21_X1 U7072 ( .B1(n7579), .B2(n6948), .A(n6408), .ZN(n6409) );
  AOI21_X1 U7073 ( .B1(n7083), .B2(n7520), .A(n6409), .ZN(n6410) );
  OAI21_X1 U7074 ( .B1(n6411), .B2(REIP_REG_29__SCAN_IN), .A(n6410), .ZN(n6412) );
  AOI21_X1 U7075 ( .B1(REIP_REG_29__SCAN_IN), .B2(n6420), .A(n6412), .ZN(n6413) );
  OAI21_X1 U7076 ( .B1(n6547), .B2(n7595), .A(n6413), .ZN(U2798) );
  INV_X1 U7077 ( .A(n6414), .ZN(n6419) );
  AOI22_X1 U7078 ( .A1(n7604), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n7608), .ZN(n6417) );
  NAND2_X1 U7079 ( .A1(n7606), .A2(n6415), .ZN(n6416) );
  OAI211_X1 U7080 ( .C1(n6521), .C2(n7593), .A(n6417), .B(n6416), .ZN(n6418)
         );
  AOI21_X1 U7081 ( .B1(n6419), .B2(n7335), .A(n6418), .ZN(n6422) );
  NAND2_X1 U7082 ( .A1(n6420), .A2(REIP_REG_28__SCAN_IN), .ZN(n6421) );
  OAI211_X1 U7083 ( .C1(n6550), .C2(n7595), .A(n6422), .B(n6421), .ZN(U2799)
         );
  INV_X1 U7084 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7333) );
  NOR2_X1 U7085 ( .A1(n6423), .A2(n6424), .ZN(n6425) );
  OR2_X2 U7086 ( .A1(n5050), .A2(n6425), .ZN(n6553) );
  INV_X1 U7087 ( .A(n6553), .ZN(n6960) );
  NAND2_X1 U7088 ( .A1(n6960), .A2(n7611), .ZN(n6436) );
  INV_X1 U7089 ( .A(n6444), .ZN(n6434) );
  NOR2_X1 U7090 ( .A1(n7331), .A2(REIP_REG_27__SCAN_IN), .ZN(n6433) );
  NOR2_X1 U7091 ( .A1(n6440), .A2(n6426), .ZN(n6427) );
  OR2_X1 U7092 ( .A1(n6428), .A2(n6427), .ZN(n7092) );
  AOI22_X1 U7093 ( .A1(n7604), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n7608), .ZN(n6431) );
  INV_X1 U7094 ( .A(n6958), .ZN(n6429) );
  NAND2_X1 U7095 ( .A1(n7606), .A2(n6429), .ZN(n6430) );
  OAI211_X1 U7096 ( .C1(n7092), .C2(n7593), .A(n6431), .B(n6430), .ZN(n6432)
         );
  AOI21_X1 U7097 ( .B1(n6434), .B2(n6433), .A(n6432), .ZN(n6435) );
  OAI211_X1 U7098 ( .C1(n3684), .C2(n7333), .A(n6436), .B(n6435), .ZN(U2800)
         );
  INV_X1 U7099 ( .A(n6438), .ZN(n6449) );
  AOI21_X1 U7100 ( .B1(n6439), .B2(n6449), .A(n6423), .ZN(n6968) );
  INV_X1 U7101 ( .A(n6968), .ZN(n6556) );
  AOI21_X1 U7102 ( .B1(n6441), .B2(n6451), .A(n6440), .ZN(n7097) );
  INV_X1 U7103 ( .A(n6442), .ZN(n6966) );
  AOI22_X1 U7104 ( .A1(n7604), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n7608), .ZN(n6443) );
  OAI21_X1 U7105 ( .B1(n7579), .B2(n6966), .A(n6443), .ZN(n6446) );
  AOI21_X1 U7106 ( .B1(n7331), .B2(n6444), .A(n3684), .ZN(n6445) );
  AOI211_X1 U7107 ( .C1(n7610), .C2(n7097), .A(n6446), .B(n6445), .ZN(n6447)
         );
  OAI21_X1 U7108 ( .B1(n6556), .B2(n7595), .A(n6447), .ZN(U2801) );
  AOI21_X1 U7109 ( .B1(n6450), .B2(n6448), .A(n6438), .ZN(n6978) );
  INV_X1 U7110 ( .A(n6978), .ZN(n6559) );
  XOR2_X1 U7111 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .Z(n6457) );
  INV_X1 U7112 ( .A(n6451), .ZN(n6452) );
  AOI21_X1 U7113 ( .B1(n6453), .B2(n6464), .A(n6452), .ZN(n7106) );
  NAND2_X1 U7114 ( .A1(n7106), .A2(n7610), .ZN(n6455) );
  AOI22_X1 U7115 ( .A1(n7604), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n7608), .ZN(n6454) );
  OAI211_X1 U7116 ( .C1(n7579), .C2(n6976), .A(n6455), .B(n6454), .ZN(n6456)
         );
  AOI21_X1 U7117 ( .B1(n6470), .B2(n6457), .A(n6456), .ZN(n6459) );
  NAND2_X1 U7118 ( .A1(n6482), .A2(REIP_REG_25__SCAN_IN), .ZN(n6458) );
  OAI211_X1 U7119 ( .C1(n6559), .C2(n7595), .A(n6459), .B(n6458), .ZN(U2802)
         );
  OR2_X1 U7120 ( .A1(n6460), .A2(n6461), .ZN(n6462) );
  AND2_X1 U7121 ( .A1(n6448), .A2(n6462), .ZN(n6987) );
  INV_X1 U7122 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7326) );
  OAI21_X1 U7123 ( .B1(n6463), .B2(n6465), .A(n6464), .ZN(n6466) );
  INV_X1 U7124 ( .A(n6466), .ZN(n7121) );
  NAND2_X1 U7125 ( .A1(n7121), .A2(n7520), .ZN(n6468) );
  AOI22_X1 U7126 ( .A1(n7604), .A2(EBX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n7608), .ZN(n6467) );
  OAI211_X1 U7127 ( .C1(n7579), .C2(n6985), .A(n6468), .B(n6467), .ZN(n6469)
         );
  AOI21_X1 U7128 ( .B1(n6470), .B2(n7326), .A(n6469), .ZN(n6472) );
  NAND2_X1 U7129 ( .A1(n6482), .A2(REIP_REG_24__SCAN_IN), .ZN(n6471) );
  OAI211_X1 U7130 ( .C1(n6562), .C2(n7595), .A(n6472), .B(n6471), .ZN(U2803)
         );
  INV_X1 U7131 ( .A(n6473), .ZN(n6474) );
  AOI21_X1 U7132 ( .B1(n6475), .B2(n6474), .A(n6460), .ZN(n6996) );
  INV_X1 U7133 ( .A(n6996), .ZN(n6565) );
  OAI22_X1 U7134 ( .A1(n6476), .A2(n7601), .B1(n6994), .B2(n7579), .ZN(n6481)
         );
  INV_X1 U7135 ( .A(n6463), .ZN(n6478) );
  OAI21_X1 U7136 ( .B1(n6479), .B2(n6477), .A(n6478), .ZN(n7128) );
  NOR2_X1 U7137 ( .A1(n7128), .A2(n7593), .ZN(n6480) );
  AOI211_X1 U7138 ( .C1(n7604), .C2(EBX_REG_23__SCAN_IN), .A(n6481), .B(n6480), 
        .ZN(n6485) );
  INV_X1 U7139 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7322) );
  INV_X1 U7140 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7321) );
  NOR3_X1 U7141 ( .A1(n6490), .A2(n7322), .A3(n7321), .ZN(n6483) );
  OAI21_X1 U7142 ( .B1(n6483), .B2(REIP_REG_23__SCAN_IN), .A(n6482), .ZN(n6484) );
  OAI211_X1 U7143 ( .C1(n6565), .C2(n7595), .A(n6485), .B(n6484), .ZN(U2804)
         );
  AOI21_X1 U7144 ( .B1(n6486), .B2(n3683), .A(n6473), .ZN(n7734) );
  INV_X1 U7145 ( .A(n7734), .ZN(n6531) );
  NOR2_X1 U7146 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6490), .ZN(n7612) );
  OAI21_X1 U7147 ( .B1(n7603), .B2(n7612), .A(REIP_REG_22__SCAN_IN), .ZN(n6494) );
  AND2_X1 U7148 ( .A1(n7145), .A2(n6488), .ZN(n6489) );
  NOR2_X1 U7149 ( .A1(n6477), .A2(n6489), .ZN(n7136) );
  AOI22_X1 U7150 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n7608), .B1(n7003), 
        .B2(n7606), .ZN(n6491) );
  OAI211_X1 U7151 ( .C1(n7577), .C2(n6528), .A(n6491), .B(n3793), .ZN(n6492)
         );
  AOI21_X1 U7152 ( .B1(n7136), .B2(n7610), .A(n6492), .ZN(n6493) );
  OAI211_X1 U7153 ( .C1(n6531), .C2(n7595), .A(n6494), .B(n6493), .ZN(U2805)
         );
  OAI21_X1 U7154 ( .B1(n6495), .B2(n6496), .A(n7026), .ZN(n7723) );
  INV_X1 U7155 ( .A(n7163), .ZN(n6498) );
  AOI21_X1 U7156 ( .B1(n6499), .B2(n6506), .A(n6498), .ZN(n7182) );
  AND2_X1 U7157 ( .A1(n6500), .A2(n7314), .ZN(n7587) );
  AOI21_X1 U7158 ( .B1(n7608), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n7582), 
        .ZN(n6502) );
  AOI22_X1 U7159 ( .A1(n7037), .A2(n7606), .B1(EBX_REG_18__SCAN_IN), .B2(n7604), .ZN(n6501) );
  OAI211_X1 U7160 ( .C1(n6512), .C2(n7314), .A(n6502), .B(n6501), .ZN(n6503)
         );
  AOI211_X1 U7161 ( .C1(n7182), .C2(n7610), .A(n7587), .B(n6503), .ZN(n6504)
         );
  OAI21_X1 U7162 ( .B1(n7723), .B2(n7595), .A(n6504), .ZN(U2809) );
  AOI21_X1 U7163 ( .B1(n6505), .B2(n6351), .A(n6495), .ZN(n7720) );
  INV_X1 U7164 ( .A(n7720), .ZN(n6544) );
  INV_X1 U7165 ( .A(n7049), .ZN(n6516) );
  INV_X1 U7166 ( .A(n6506), .ZN(n6507) );
  AOI21_X1 U7167 ( .B1(n6509), .B2(n6508), .A(n6507), .ZN(n7190) );
  INV_X1 U7168 ( .A(n7190), .ZN(n6511) );
  AOI22_X1 U7169 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n7608), .B1(
        EBX_REG_17__SCAN_IN), .B2(n7604), .ZN(n6510) );
  OAI211_X1 U7170 ( .C1(n6511), .C2(n7593), .A(n6510), .B(n7554), .ZN(n6515)
         );
  AOI21_X1 U7171 ( .B1(n7313), .B2(n6513), .A(n6512), .ZN(n6514) );
  AOI211_X1 U7172 ( .C1(n7606), .C2(n6516), .A(n6515), .B(n6514), .ZN(n6517)
         );
  OAI21_X1 U7173 ( .B1(n6544), .B2(n7595), .A(n6517), .ZN(U2810) );
  INV_X1 U7174 ( .A(n7073), .ZN(n6519) );
  OAI22_X1 U7175 ( .A1(n6519), .A2(n7372), .B1(n7376), .B2(n6518), .ZN(U2828)
         );
  AOI22_X1 U7176 ( .A1(n7083), .A2(n7369), .B1(EBX_REG_29__SCAN_IN), .B2(n6541), .ZN(n6520) );
  OAI21_X1 U7177 ( .B1(n6547), .B2(n6543), .A(n6520), .ZN(U2830) );
  OAI222_X1 U7178 ( .A1(n6539), .A2(n6550), .B1(n6522), .B2(n7376), .C1(n6521), 
        .C2(n7372), .ZN(U2831) );
  INV_X1 U7179 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6523) );
  OAI222_X1 U7180 ( .A1(n6539), .A2(n6553), .B1(n6523), .B2(n7376), .C1(n7092), 
        .C2(n7372), .ZN(U2832) );
  AOI22_X1 U7181 ( .A1(n7097), .A2(n7369), .B1(EBX_REG_26__SCAN_IN), .B2(n6541), .ZN(n6524) );
  OAI21_X1 U7182 ( .B1(n6556), .B2(n6543), .A(n6524), .ZN(U2833) );
  AOI22_X1 U7183 ( .A1(n7106), .A2(n7369), .B1(EBX_REG_25__SCAN_IN), .B2(n6541), .ZN(n6525) );
  OAI21_X1 U7184 ( .B1(n6559), .B2(n6539), .A(n6525), .ZN(U2834) );
  AOI22_X1 U7185 ( .A1(n7121), .A2(n7369), .B1(EBX_REG_24__SCAN_IN), .B2(n6541), .ZN(n6526) );
  OAI21_X1 U7186 ( .B1(n6562), .B2(n6539), .A(n6526), .ZN(U2835) );
  INV_X1 U7187 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6527) );
  OAI222_X1 U7188 ( .A1(n6539), .A2(n6565), .B1(n6527), .B2(n7376), .C1(n7128), 
        .C2(n7372), .ZN(U2836) );
  NOR2_X1 U7189 ( .A1(n7376), .A2(n6528), .ZN(n6529) );
  AOI21_X1 U7190 ( .B1(n7136), .B2(n7369), .A(n6529), .ZN(n6530) );
  OAI21_X1 U7191 ( .B1(n6531), .B2(n6543), .A(n6530), .ZN(U2837) );
  OAI21_X1 U7192 ( .B1(n6533), .B2(n6535), .A(n6534), .ZN(n7596) );
  OR2_X1 U7193 ( .A1(n7161), .A2(n6537), .ZN(n6538) );
  NAND2_X1 U7194 ( .A1(n6536), .A2(n6538), .ZN(n7594) );
  OAI222_X1 U7195 ( .A1(n6539), .A2(n7596), .B1(n7376), .B2(n4416), .C1(n7594), 
        .C2(n7372), .ZN(U2839) );
  AOI22_X1 U7196 ( .A1(n7182), .A2(n7369), .B1(EBX_REG_18__SCAN_IN), .B2(n6541), .ZN(n6540) );
  OAI21_X1 U7197 ( .B1(n7723), .B2(n6543), .A(n6540), .ZN(U2841) );
  AOI22_X1 U7198 ( .A1(n7190), .A2(n7369), .B1(EBX_REG_17__SCAN_IN), .B2(n6541), .ZN(n6542) );
  OAI21_X1 U7199 ( .B1(n6544), .B2(n6543), .A(n6542), .ZN(U2842) );
  AOI22_X1 U7200 ( .A1(n7733), .A2(DATAI_13_), .B1(n7735), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U7201 ( .A1(n7736), .A2(DATAI_29_), .ZN(n6545) );
  OAI211_X1 U7202 ( .C1(n6547), .C2(n6568), .A(n6546), .B(n6545), .ZN(U2862)
         );
  AOI22_X1 U7203 ( .A1(n7733), .A2(DATAI_12_), .B1(n7735), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U7204 ( .A1(n7736), .A2(DATAI_28_), .ZN(n6548) );
  OAI211_X1 U7205 ( .C1(n6550), .C2(n6568), .A(n6549), .B(n6548), .ZN(U2863)
         );
  AOI22_X1 U7206 ( .A1(n7733), .A2(DATAI_11_), .B1(n7735), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U7207 ( .A1(n7736), .A2(DATAI_27_), .ZN(n6551) );
  OAI211_X1 U7208 ( .C1(n6553), .C2(n6568), .A(n6552), .B(n6551), .ZN(U2864)
         );
  AOI22_X1 U7209 ( .A1(n7733), .A2(DATAI_10_), .B1(n7735), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7210 ( .A1(n7736), .A2(DATAI_26_), .ZN(n6554) );
  OAI211_X1 U7211 ( .C1(n6556), .C2(n6568), .A(n6555), .B(n6554), .ZN(U2865)
         );
  AOI22_X1 U7212 ( .A1(n7733), .A2(DATAI_9_), .B1(n7735), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U7213 ( .A1(n7736), .A2(DATAI_25_), .ZN(n6557) );
  OAI211_X1 U7214 ( .C1(n6559), .C2(n6568), .A(n6558), .B(n6557), .ZN(U2866)
         );
  AOI22_X1 U7215 ( .A1(n7733), .A2(DATAI_8_), .B1(n7735), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U7216 ( .A1(n7736), .A2(DATAI_24_), .ZN(n6560) );
  OAI211_X1 U7217 ( .C1(n6562), .C2(n6568), .A(n6561), .B(n6560), .ZN(U2867)
         );
  AOI22_X1 U7218 ( .A1(n7733), .A2(DATAI_7_), .B1(n7735), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U7219 ( .A1(n7736), .A2(DATAI_23_), .ZN(n6563) );
  OAI211_X1 U7220 ( .C1(n6565), .C2(n6568), .A(n6564), .B(n6563), .ZN(U2868)
         );
  AOI22_X1 U7221 ( .A1(n7733), .A2(DATAI_4_), .B1(n7735), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U7222 ( .A1(n7736), .A2(DATAI_20_), .ZN(n6566) );
  OAI211_X1 U7223 ( .C1(n7596), .C2(n6568), .A(n6567), .B(n6566), .ZN(U2871)
         );
  AOI222_X1 U7224 ( .A1(n6569), .A2(DATAI_1_), .B1(n3645), .B2(n7378), .C1(
        n7735), .C2(EAX_REG_1__SCAN_IN), .ZN(n6935) );
  XOR2_X1 U7225 ( .A(DATAI_28_), .B(keyinput_131), .Z(n6572) );
  XNOR2_X1 U7226 ( .A(DATAI_27_), .B(keyinput_132), .ZN(n6571) );
  XNOR2_X1 U7227 ( .A(DATAI_31_), .B(keyinput_128), .ZN(n6570) );
  NOR3_X1 U7228 ( .A1(n6572), .A2(n6571), .A3(n6570), .ZN(n6575) );
  XOR2_X1 U7229 ( .A(DATAI_29_), .B(keyinput_130), .Z(n6574) );
  XOR2_X1 U7230 ( .A(DATAI_30_), .B(keyinput_129), .Z(n6573) );
  NAND3_X1 U7231 ( .A1(n6575), .A2(n6574), .A3(n6573), .ZN(n6579) );
  XOR2_X1 U7232 ( .A(DATAI_26_), .B(keyinput_133), .Z(n6578) );
  XOR2_X1 U7233 ( .A(DATAI_24_), .B(keyinput_135), .Z(n6577) );
  XNOR2_X1 U7234 ( .A(DATAI_25_), .B(keyinput_134), .ZN(n6576) );
  NAND4_X1 U7235 ( .A1(n6579), .A2(n6578), .A3(n6577), .A4(n6576), .ZN(n6583)
         );
  XOR2_X1 U7236 ( .A(DATAI_23_), .B(keyinput_136), .Z(n6582) );
  XNOR2_X1 U7237 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n6581) );
  XNOR2_X1 U7238 ( .A(DATAI_21_), .B(keyinput_138), .ZN(n6580) );
  AOI211_X1 U7239 ( .C1(n6583), .C2(n6582), .A(n6581), .B(n6580), .ZN(n6586)
         );
  XOR2_X1 U7240 ( .A(DATAI_19_), .B(keyinput_140), .Z(n6585) );
  XNOR2_X1 U7241 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n6584) );
  NOR3_X1 U7242 ( .A1(n6586), .A2(n6585), .A3(n6584), .ZN(n6590) );
  XOR2_X1 U7243 ( .A(DATAI_18_), .B(keyinput_141), .Z(n6589) );
  XOR2_X1 U7244 ( .A(DATAI_17_), .B(keyinput_142), .Z(n6588) );
  XNOR2_X1 U7245 ( .A(DATAI_16_), .B(keyinput_143), .ZN(n6587) );
  OAI211_X1 U7246 ( .C1(n6590), .C2(n6589), .A(n6588), .B(n6587), .ZN(n6594)
         );
  XNOR2_X1 U7247 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n6593) );
  XNOR2_X1 U7248 ( .A(DATAI_14_), .B(keyinput_145), .ZN(n6592) );
  XNOR2_X1 U7249 ( .A(DATAI_15_), .B(keyinput_144), .ZN(n6591) );
  NAND4_X1 U7250 ( .A1(n6594), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(n6597)
         );
  XOR2_X1 U7251 ( .A(DATAI_12_), .B(keyinput_147), .Z(n6596) );
  XOR2_X1 U7252 ( .A(DATAI_11_), .B(keyinput_148), .Z(n6595) );
  NAND3_X1 U7253 ( .A1(n6597), .A2(n6596), .A3(n6595), .ZN(n6601) );
  XNOR2_X1 U7254 ( .A(DATAI_8_), .B(keyinput_151), .ZN(n6600) );
  XNOR2_X1 U7255 ( .A(DATAI_10_), .B(keyinput_149), .ZN(n6599) );
  XNOR2_X1 U7256 ( .A(DATAI_9_), .B(keyinput_150), .ZN(n6598) );
  NAND4_X1 U7257 ( .A1(n6601), .A2(n6600), .A3(n6599), .A4(n6598), .ZN(n6605)
         );
  XOR2_X1 U7258 ( .A(DATAI_7_), .B(keyinput_152), .Z(n6604) );
  XNOR2_X1 U7259 ( .A(DATAI_5_), .B(keyinput_154), .ZN(n6603) );
  XNOR2_X1 U7260 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n6602) );
  NAND4_X1 U7261 ( .A1(n6605), .A2(n6604), .A3(n6603), .A4(n6602), .ZN(n6609)
         );
  XNOR2_X1 U7262 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n6608) );
  XOR2_X1 U7263 ( .A(DATAI_2_), .B(keyinput_157), .Z(n6607) );
  XOR2_X1 U7264 ( .A(DATAI_3_), .B(keyinput_156), .Z(n6606) );
  AOI211_X1 U7265 ( .C1(n6609), .C2(n6608), .A(n6607), .B(n6606), .ZN(n6612)
         );
  XNOR2_X1 U7266 ( .A(DATAI_1_), .B(keyinput_158), .ZN(n6611) );
  XNOR2_X1 U7267 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n6610) );
  OAI21_X1 U7268 ( .B1(n6612), .B2(n6611), .A(n6610), .ZN(n6615) );
  XNOR2_X1 U7269 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_160), .ZN(n6614)
         );
  XNOR2_X1 U7270 ( .A(NA_N), .B(keyinput_161), .ZN(n6613) );
  NAND3_X1 U7271 ( .A1(n6615), .A2(n6614), .A3(n6613), .ZN(n6618) );
  XOR2_X1 U7272 ( .A(BS16_N), .B(keyinput_162), .Z(n6617) );
  XNOR2_X1 U7273 ( .A(n7709), .B(keyinput_163), .ZN(n6616) );
  AOI21_X1 U7274 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(n6624) );
  XOR2_X1 U7275 ( .A(HOLD), .B(keyinput_164), .Z(n6623) );
  XOR2_X1 U7276 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_165), .Z(n6621) );
  XNOR2_X1 U7277 ( .A(CODEFETCH_REG_SCAN_IN), .B(keyinput_167), .ZN(n6620) );
  XNOR2_X1 U7278 ( .A(ADS_N_REG_SCAN_IN), .B(keyinput_166), .ZN(n6619) );
  NOR3_X1 U7279 ( .A1(n6621), .A2(n6620), .A3(n6619), .ZN(n6622) );
  OAI21_X1 U7280 ( .B1(n6624), .B2(n6623), .A(n6622), .ZN(n6631) );
  XOR2_X1 U7281 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_169), .Z(n6628) );
  INV_X1 U7282 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7717) );
  XNOR2_X1 U7283 ( .A(n7717), .B(keyinput_168), .ZN(n6627) );
  XNOR2_X1 U7284 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_170), .ZN(n6626) );
  XNOR2_X1 U7285 ( .A(STATEBS16_REG_SCAN_IN), .B(keyinput_171), .ZN(n6625) );
  NOR4_X1 U7286 ( .A1(n6628), .A2(n6627), .A3(n6626), .A4(n6625), .ZN(n6630)
         );
  XOR2_X1 U7287 ( .A(MORE_REG_SCAN_IN), .B(keyinput_172), .Z(n6629) );
  AOI21_X1 U7288 ( .B1(n6631), .B2(n6630), .A(n6629), .ZN(n6635) );
  INV_X1 U7289 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7365) );
  XNOR2_X1 U7290 ( .A(n7365), .B(keyinput_175), .ZN(n6634) );
  XNOR2_X1 U7291 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_173), .ZN(n6633) );
  XNOR2_X1 U7292 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_174), .ZN(n6632) );
  NOR4_X1 U7293 ( .A1(n6635), .A2(n6634), .A3(n6633), .A4(n6632), .ZN(n6639)
         );
  XNOR2_X1 U7294 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_176), .ZN(n6638)
         );
  XNOR2_X1 U7295 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_177), .ZN(n6637)
         );
  XNOR2_X1 U7296 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_178), .ZN(n6636)
         );
  OAI211_X1 U7297 ( .C1(n6639), .C2(n6638), .A(n6637), .B(n6636), .ZN(n6645)
         );
  XNOR2_X1 U7298 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_179), .ZN(n6644) );
  XOR2_X1 U7299 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_180), .Z(n6642) );
  XNOR2_X1 U7300 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_182), .ZN(n6641) );
  XNOR2_X1 U7301 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_181), .ZN(n6640) );
  NAND3_X1 U7302 ( .A1(n6642), .A2(n6641), .A3(n6640), .ZN(n6643) );
  AOI21_X1 U7303 ( .B1(n6645), .B2(n6644), .A(n6643), .ZN(n6649) );
  XNOR2_X1 U7304 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_183), .ZN(n6648) );
  XOR2_X1 U7305 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_185), .Z(n6647) );
  XNOR2_X1 U7306 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_184), .ZN(n6646) );
  OAI211_X1 U7307 ( .C1(n6649), .C2(n6648), .A(n6647), .B(n6646), .ZN(n6655)
         );
  XNOR2_X1 U7308 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_186), .ZN(n6654) );
  XOR2_X1 U7309 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_189), .Z(n6652) );
  XNOR2_X1 U7310 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_188), .ZN(n6651) );
  XNOR2_X1 U7311 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_187), .ZN(n6650) );
  NAND3_X1 U7312 ( .A1(n6652), .A2(n6651), .A3(n6650), .ZN(n6653) );
  AOI21_X1 U7313 ( .B1(n6655), .B2(n6654), .A(n6653), .ZN(n6658) );
  XOR2_X1 U7314 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_190), .Z(n6657) );
  XOR2_X1 U7315 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_191), .Z(n6656) );
  OAI21_X1 U7316 ( .B1(n6658), .B2(n6657), .A(n6656), .ZN(n6661) );
  XOR2_X1 U7317 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_193), .Z(n6660) );
  XNOR2_X1 U7318 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_192), .ZN(n6659) );
  NAND3_X1 U7319 ( .A1(n6661), .A2(n6660), .A3(n6659), .ZN(n6665) );
  INV_X1 U7320 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n7355) );
  XNOR2_X1 U7321 ( .A(n7355), .B(keyinput_196), .ZN(n6664) );
  XOR2_X1 U7322 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_194), .Z(n6663) );
  XNOR2_X1 U7323 ( .A(BE_N_REG_3__SCAN_IN), .B(keyinput_195), .ZN(n6662) );
  NAND4_X1 U7324 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6672)
         );
  INV_X1 U7325 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n7359) );
  XNOR2_X1 U7326 ( .A(n7359), .B(keyinput_197), .ZN(n6671) );
  INV_X1 U7327 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7336) );
  XNOR2_X1 U7328 ( .A(n7336), .B(keyinput_201), .ZN(n6668) );
  INV_X1 U7329 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7340) );
  XNOR2_X1 U7330 ( .A(n7340), .B(keyinput_199), .ZN(n6667) );
  XNOR2_X1 U7331 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_198), .ZN(n6666) );
  NOR3_X1 U7332 ( .A1(n6668), .A2(n6667), .A3(n6666), .ZN(n6670) );
  XNOR2_X1 U7333 ( .A(ADDRESS_REG_28__SCAN_IN), .B(keyinput_200), .ZN(n6669)
         );
  NAND4_X1 U7334 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6679)
         );
  XNOR2_X1 U7335 ( .A(ADDRESS_REG_26__SCAN_IN), .B(keyinput_202), .ZN(n6678)
         );
  XOR2_X1 U7336 ( .A(ADDRESS_REG_23__SCAN_IN), .B(keyinput_205), .Z(n6676) );
  INV_X1 U7337 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7324) );
  XNOR2_X1 U7338 ( .A(n7324), .B(keyinput_206), .ZN(n6675) );
  XNOR2_X1 U7339 ( .A(ADDRESS_REG_24__SCAN_IN), .B(keyinput_204), .ZN(n6674)
         );
  XNOR2_X1 U7340 ( .A(ADDRESS_REG_25__SCAN_IN), .B(keyinput_203), .ZN(n6673)
         );
  NAND4_X1 U7341 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6677)
         );
  AOI21_X1 U7342 ( .B1(n6679), .B2(n6678), .A(n6677), .ZN(n6685) );
  XNOR2_X1 U7343 ( .A(ADDRESS_REG_21__SCAN_IN), .B(keyinput_207), .ZN(n6684)
         );
  INV_X1 U7344 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7318) );
  XNOR2_X1 U7345 ( .A(n7318), .B(keyinput_209), .ZN(n6682) );
  INV_X1 U7346 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7320) );
  XNOR2_X1 U7347 ( .A(n7320), .B(keyinput_208), .ZN(n6681) );
  XNOR2_X1 U7348 ( .A(ADDRESS_REG_18__SCAN_IN), .B(keyinput_210), .ZN(n6680)
         );
  NOR3_X1 U7349 ( .A1(n6682), .A2(n6681), .A3(n6680), .ZN(n6683) );
  OAI21_X1 U7350 ( .B1(n6685), .B2(n6684), .A(n6683), .ZN(n6690) );
  INV_X1 U7351 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n7312) );
  OAI22_X1 U7352 ( .A1(n7312), .A2(keyinput_212), .B1(keyinput_213), .B2(
        ADDRESS_REG_15__SCAN_IN), .ZN(n6686) );
  AOI21_X1 U7353 ( .B1(n7312), .B2(keyinput_212), .A(n6686), .ZN(n6689) );
  XNOR2_X1 U7354 ( .A(ADDRESS_REG_17__SCAN_IN), .B(keyinput_211), .ZN(n6688)
         );
  NAND2_X1 U7355 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(keyinput_213), .ZN(n6687)
         );
  NAND4_X1 U7356 ( .A1(n6690), .A2(n6689), .A3(n6688), .A4(n6687), .ZN(n6693)
         );
  INV_X1 U7357 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7309) );
  XNOR2_X1 U7358 ( .A(n7309), .B(keyinput_214), .ZN(n6692) );
  XNOR2_X1 U7359 ( .A(ADDRESS_REG_13__SCAN_IN), .B(keyinput_215), .ZN(n6691)
         );
  AOI21_X1 U7360 ( .B1(n6693), .B2(n6692), .A(n6691), .ZN(n6697) );
  INV_X1 U7361 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n7304) );
  XNOR2_X1 U7362 ( .A(n7304), .B(keyinput_218), .ZN(n6696) );
  XNOR2_X1 U7363 ( .A(ADDRESS_REG_11__SCAN_IN), .B(keyinput_217), .ZN(n6695)
         );
  XNOR2_X1 U7364 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_216), .ZN(n6694)
         );
  NOR4_X1 U7365 ( .A1(n6697), .A2(n6696), .A3(n6695), .A4(n6694), .ZN(n6700)
         );
  XNOR2_X1 U7366 ( .A(ADDRESS_REG_8__SCAN_IN), .B(keyinput_220), .ZN(n6699) );
  XNOR2_X1 U7367 ( .A(ADDRESS_REG_9__SCAN_IN), .B(keyinput_219), .ZN(n6698) );
  NOR3_X1 U7368 ( .A1(n6700), .A2(n6699), .A3(n6698), .ZN(n6706) );
  INV_X1 U7369 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7299) );
  XNOR2_X1 U7370 ( .A(n7299), .B(keyinput_221), .ZN(n6705) );
  INV_X1 U7371 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7296) );
  XNOR2_X1 U7372 ( .A(n7296), .B(keyinput_223), .ZN(n6703) );
  XNOR2_X1 U7373 ( .A(ADDRESS_REG_4__SCAN_IN), .B(keyinput_224), .ZN(n6702) );
  XNOR2_X1 U7374 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_222), .ZN(n6701) );
  NOR3_X1 U7375 ( .A1(n6703), .A2(n6702), .A3(n6701), .ZN(n6704) );
  OAI21_X1 U7376 ( .B1(n6706), .B2(n6705), .A(n6704), .ZN(n6713) );
  INV_X1 U7377 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7288) );
  XNOR2_X1 U7378 ( .A(n7288), .B(keyinput_228), .ZN(n6710) );
  INV_X1 U7379 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7291) );
  XNOR2_X1 U7380 ( .A(n7291), .B(keyinput_226), .ZN(n6709) );
  INV_X1 U7381 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7292) );
  XNOR2_X1 U7382 ( .A(n7292), .B(keyinput_225), .ZN(n6708) );
  XNOR2_X1 U7383 ( .A(ADDRESS_REG_1__SCAN_IN), .B(keyinput_227), .ZN(n6707) );
  NOR4_X1 U7384 ( .A1(n6710), .A2(n6709), .A3(n6708), .A4(n6707), .ZN(n6712)
         );
  XOR2_X1 U7385 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_229), .Z(n6711) );
  AOI21_X1 U7386 ( .B1(n6713), .B2(n6712), .A(n6711), .ZN(n6719) );
  INV_X1 U7387 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n7234) );
  AOI22_X1 U7388 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput_231), .B1(n7234), 
        .B2(keyinput_234), .ZN(n6714) );
  OAI221_X1 U7389 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput_231), .C1(n7234), 
        .C2(keyinput_234), .A(n6714), .ZN(n6718) );
  AOI22_X1 U7390 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(keyinput_233), .B1(n7420), .B2(keyinput_230), .ZN(n6715) );
  OAI221_X1 U7391 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput_233), .C1(
        n7420), .C2(keyinput_230), .A(n6715), .ZN(n6717) );
  XNOR2_X1 U7392 ( .A(DATAWIDTH_REG_0__SCAN_IN), .B(keyinput_232), .ZN(n6716)
         );
  NOR4_X1 U7393 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6722)
         );
  XNOR2_X1 U7394 ( .A(DATAWIDTH_REG_3__SCAN_IN), .B(keyinput_235), .ZN(n6721)
         );
  XNOR2_X1 U7395 ( .A(DATAWIDTH_REG_4__SCAN_IN), .B(keyinput_236), .ZN(n6720)
         );
  OAI21_X1 U7396 ( .B1(n6722), .B2(n6721), .A(n6720), .ZN(n6726) );
  INV_X1 U7397 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7239) );
  XNOR2_X1 U7398 ( .A(n7239), .B(keyinput_239), .ZN(n6725) );
  XNOR2_X1 U7399 ( .A(DATAWIDTH_REG_5__SCAN_IN), .B(keyinput_237), .ZN(n6724)
         );
  XNOR2_X1 U7400 ( .A(DATAWIDTH_REG_6__SCAN_IN), .B(keyinput_238), .ZN(n6723)
         );
  NAND4_X1 U7401 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6729)
         );
  INV_X1 U7402 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n7240) );
  XNOR2_X1 U7403 ( .A(n7240), .B(keyinput_240), .ZN(n6728) );
  XNOR2_X1 U7404 ( .A(DATAWIDTH_REG_9__SCAN_IN), .B(keyinput_241), .ZN(n6727)
         );
  NAND3_X1 U7405 ( .A1(n6729), .A2(n6728), .A3(n6727), .ZN(n6732) );
  INV_X1 U7406 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n7242) );
  XNOR2_X1 U7407 ( .A(n7242), .B(keyinput_242), .ZN(n6731) );
  XNOR2_X1 U7408 ( .A(DATAWIDTH_REG_11__SCAN_IN), .B(keyinput_243), .ZN(n6730)
         );
  NAND3_X1 U7409 ( .A1(n6732), .A2(n6731), .A3(n6730), .ZN(n6735) );
  XOR2_X1 U7410 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(keyinput_245), .Z(n6734)
         );
  INV_X1 U7411 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7244) );
  XNOR2_X1 U7412 ( .A(n7244), .B(keyinput_244), .ZN(n6733) );
  NAND3_X1 U7413 ( .A1(n6735), .A2(n6734), .A3(n6733), .ZN(n6737) );
  XNOR2_X1 U7414 ( .A(DATAWIDTH_REG_14__SCAN_IN), .B(keyinput_246), .ZN(n6736)
         );
  NAND2_X1 U7415 ( .A1(n6737), .A2(n6736), .ZN(n6743) );
  INV_X1 U7416 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7249) );
  OAI22_X1 U7417 ( .A1(n7249), .A2(keyinput_251), .B1(
        DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput_247), .ZN(n6738) );
  AOI221_X1 U7418 ( .B1(n7249), .B2(keyinput_251), .C1(keyinput_247), .C2(
        DATAWIDTH_REG_15__SCAN_IN), .A(n6738), .ZN(n6742) );
  XOR2_X1 U7419 ( .A(DATAWIDTH_REG_16__SCAN_IN), .B(keyinput_248), .Z(n6741)
         );
  INV_X1 U7420 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n7247) );
  OAI22_X1 U7421 ( .A1(n7247), .A2(keyinput_249), .B1(keyinput_250), .B2(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6739) );
  AOI221_X1 U7422 ( .B1(n7247), .B2(keyinput_249), .C1(
        DATAWIDTH_REG_18__SCAN_IN), .C2(keyinput_250), .A(n6739), .ZN(n6740)
         );
  NAND4_X1 U7423 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6746)
         );
  XNOR2_X1 U7424 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_252), .ZN(n6745)
         );
  XNOR2_X1 U7425 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_253), .ZN(n6744)
         );
  AOI21_X1 U7426 ( .B1(n6746), .B2(n6745), .A(n6744), .ZN(n6933) );
  INV_X1 U7427 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n7252) );
  XNOR2_X1 U7428 ( .A(n7252), .B(keyinput_254), .ZN(n6932) );
  XOR2_X1 U7429 ( .A(DATAI_27_), .B(keyinput_4), .Z(n6749) );
  XNOR2_X1 U7430 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n6748) );
  XNOR2_X1 U7431 ( .A(DATAI_30_), .B(keyinput_1), .ZN(n6747) );
  NOR3_X1 U7432 ( .A1(n6749), .A2(n6748), .A3(n6747), .ZN(n6752) );
  XOR2_X1 U7433 ( .A(DATAI_28_), .B(keyinput_3), .Z(n6751) );
  XOR2_X1 U7434 ( .A(DATAI_31_), .B(keyinput_0), .Z(n6750) );
  NAND3_X1 U7435 ( .A1(n6752), .A2(n6751), .A3(n6750), .ZN(n6756) );
  XOR2_X1 U7436 ( .A(DATAI_24_), .B(keyinput_7), .Z(n6755) );
  XOR2_X1 U7437 ( .A(DATAI_25_), .B(keyinput_6), .Z(n6754) );
  XNOR2_X1 U7438 ( .A(DATAI_26_), .B(keyinput_5), .ZN(n6753) );
  NAND4_X1 U7439 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(n6760)
         );
  XOR2_X1 U7440 ( .A(DATAI_23_), .B(keyinput_8), .Z(n6759) );
  XOR2_X1 U7441 ( .A(keyinput_10), .B(DATAI_21_), .Z(n6758) );
  XNOR2_X1 U7442 ( .A(keyinput_9), .B(DATAI_22_), .ZN(n6757) );
  AOI211_X1 U7443 ( .C1(n6760), .C2(n6759), .A(n6758), .B(n6757), .ZN(n6763)
         );
  XNOR2_X1 U7444 ( .A(DATAI_20_), .B(keyinput_11), .ZN(n6762) );
  XNOR2_X1 U7445 ( .A(keyinput_12), .B(DATAI_19_), .ZN(n6761) );
  NOR3_X1 U7446 ( .A1(n6763), .A2(n6762), .A3(n6761), .ZN(n6767) );
  XNOR2_X1 U7447 ( .A(keyinput_13), .B(DATAI_18_), .ZN(n6766) );
  XOR2_X1 U7448 ( .A(keyinput_14), .B(DATAI_17_), .Z(n6765) );
  XOR2_X1 U7449 ( .A(DATAI_16_), .B(keyinput_15), .Z(n6764) );
  OAI211_X1 U7450 ( .C1(n6767), .C2(n6766), .A(n6765), .B(n6764), .ZN(n6771)
         );
  XNOR2_X1 U7451 ( .A(DATAI_13_), .B(keyinput_18), .ZN(n6770) );
  XNOR2_X1 U7452 ( .A(DATAI_14_), .B(keyinput_17), .ZN(n6769) );
  XNOR2_X1 U7453 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n6768) );
  NAND4_X1 U7454 ( .A1(n6771), .A2(n6770), .A3(n6769), .A4(n6768), .ZN(n6774)
         );
  XOR2_X1 U7455 ( .A(DATAI_12_), .B(keyinput_19), .Z(n6773) );
  XNOR2_X1 U7456 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n6772) );
  NAND3_X1 U7457 ( .A1(n6774), .A2(n6773), .A3(n6772), .ZN(n6778) );
  XOR2_X1 U7458 ( .A(DATAI_9_), .B(keyinput_22), .Z(n6777) );
  XOR2_X1 U7459 ( .A(DATAI_10_), .B(keyinput_21), .Z(n6776) );
  XNOR2_X1 U7460 ( .A(DATAI_8_), .B(keyinput_23), .ZN(n6775) );
  NAND4_X1 U7461 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6782)
         );
  XOR2_X1 U7462 ( .A(DATAI_6_), .B(keyinput_25), .Z(n6781) );
  XOR2_X1 U7463 ( .A(DATAI_5_), .B(keyinput_26), .Z(n6780) );
  XNOR2_X1 U7464 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n6779) );
  NAND4_X1 U7465 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6779), .ZN(n6786)
         );
  XNOR2_X1 U7466 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n6785) );
  XOR2_X1 U7467 ( .A(DATAI_2_), .B(keyinput_29), .Z(n6784) );
  XNOR2_X1 U7468 ( .A(DATAI_3_), .B(keyinput_28), .ZN(n6783) );
  AOI211_X1 U7469 ( .C1(n6786), .C2(n6785), .A(n6784), .B(n6783), .ZN(n6789)
         );
  XNOR2_X1 U7470 ( .A(DATAI_1_), .B(keyinput_30), .ZN(n6788) );
  XNOR2_X1 U7471 ( .A(DATAI_0_), .B(keyinput_31), .ZN(n6787) );
  OAI21_X1 U7472 ( .B1(n6789), .B2(n6788), .A(n6787), .ZN(n6792) );
  XOR2_X1 U7473 ( .A(keyinput_33), .B(NA_N), .Z(n6791) );
  XOR2_X1 U7474 ( .A(keyinput_32), .B(MEMORYFETCH_REG_SCAN_IN), .Z(n6790) );
  NAND3_X1 U7475 ( .A1(n6792), .A2(n6791), .A3(n6790), .ZN(n6795) );
  XOR2_X1 U7476 ( .A(BS16_N), .B(keyinput_34), .Z(n6794) );
  XNOR2_X1 U7477 ( .A(n7709), .B(keyinput_35), .ZN(n6793) );
  AOI21_X1 U7478 ( .B1(n6795), .B2(n6794), .A(n6793), .ZN(n6801) );
  XNOR2_X1 U7479 ( .A(HOLD), .B(keyinput_36), .ZN(n6800) );
  XOR2_X1 U7480 ( .A(keyinput_37), .B(READREQUEST_REG_SCAN_IN), .Z(n6798) );
  INV_X1 U7481 ( .A(ADS_N_REG_SCAN_IN), .ZN(n7256) );
  XNOR2_X1 U7482 ( .A(n7256), .B(keyinput_38), .ZN(n6797) );
  XNOR2_X1 U7483 ( .A(keyinput_39), .B(CODEFETCH_REG_SCAN_IN), .ZN(n6796) );
  NOR3_X1 U7484 ( .A1(n6798), .A2(n6797), .A3(n6796), .ZN(n6799) );
  OAI21_X1 U7485 ( .B1(n6801), .B2(n6800), .A(n6799), .ZN(n6807) );
  XNOR2_X1 U7486 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_41), .ZN(n6803) );
  XNOR2_X1 U7487 ( .A(STATEBS16_REG_SCAN_IN), .B(keyinput_43), .ZN(n6802) );
  NOR2_X1 U7488 ( .A1(n6803), .A2(n6802), .ZN(n6806) );
  XNOR2_X1 U7489 ( .A(keyinput_42), .B(REQUESTPENDING_REG_SCAN_IN), .ZN(n6805)
         );
  XNOR2_X1 U7490 ( .A(keyinput_40), .B(M_IO_N_REG_SCAN_IN), .ZN(n6804) );
  NAND4_X1 U7491 ( .A1(n6807), .A2(n6806), .A3(n6805), .A4(n6804), .ZN(n6813)
         );
  XOR2_X1 U7492 ( .A(keyinput_44), .B(MORE_REG_SCAN_IN), .Z(n6812) );
  XOR2_X1 U7493 ( .A(keyinput_45), .B(FLUSH_REG_SCAN_IN), .Z(n6810) );
  XNOR2_X1 U7494 ( .A(n7365), .B(keyinput_47), .ZN(n6809) );
  XNOR2_X1 U7495 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_46), .ZN(n6808) );
  NAND3_X1 U7496 ( .A1(n6810), .A2(n6809), .A3(n6808), .ZN(n6811) );
  AOI21_X1 U7497 ( .B1(n6813), .B2(n6812), .A(n6811), .ZN(n6817) );
  XOR2_X1 U7498 ( .A(keyinput_48), .B(BYTEENABLE_REG_1__SCAN_IN), .Z(n6816) );
  XOR2_X1 U7499 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_50), .Z(n6815) );
  XNOR2_X1 U7500 ( .A(keyinput_49), .B(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6814)
         );
  OAI211_X1 U7501 ( .C1(n6817), .C2(n6816), .A(n6815), .B(n6814), .ZN(n6823)
         );
  XNOR2_X1 U7502 ( .A(n7341), .B(keyinput_51), .ZN(n6822) );
  XNOR2_X1 U7503 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_54), .ZN(n6820) );
  XNOR2_X1 U7504 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_52), .ZN(n6819) );
  XNOR2_X1 U7505 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_53), .ZN(n6818) );
  NAND3_X1 U7506 ( .A1(n6820), .A2(n6819), .A3(n6818), .ZN(n6821) );
  AOI21_X1 U7507 ( .B1(n6823), .B2(n6822), .A(n6821), .ZN(n6827) );
  XNOR2_X1 U7508 ( .A(n7333), .B(keyinput_55), .ZN(n6826) );
  XNOR2_X1 U7509 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_57), .ZN(n6825) );
  XNOR2_X1 U7510 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_56), .ZN(n6824) );
  OAI211_X1 U7511 ( .C1(n6827), .C2(n6826), .A(n6825), .B(n6824), .ZN(n6833)
         );
  XNOR2_X1 U7512 ( .A(n7326), .B(keyinput_58), .ZN(n6832) );
  XNOR2_X1 U7513 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_60), .ZN(n6830) );
  XNOR2_X1 U7514 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_61), .ZN(n6829) );
  XNOR2_X1 U7515 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_59), .ZN(n6828) );
  NAND3_X1 U7516 ( .A1(n6830), .A2(n6829), .A3(n6828), .ZN(n6831) );
  AOI21_X1 U7517 ( .B1(n6833), .B2(n6832), .A(n6831), .ZN(n6836) );
  XNOR2_X1 U7518 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_62), .ZN(n6835) );
  XNOR2_X1 U7519 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_63), .ZN(n6834) );
  OAI21_X1 U7520 ( .B1(n6836), .B2(n6835), .A(n6834), .ZN(n6839) );
  XNOR2_X1 U7521 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_64), .ZN(n6838) );
  XNOR2_X1 U7522 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_65), .ZN(n6837) );
  NAND3_X1 U7523 ( .A1(n6839), .A2(n6838), .A3(n6837), .ZN(n6843) );
  XNOR2_X1 U7524 ( .A(keyinput_68), .B(BE_N_REG_2__SCAN_IN), .ZN(n6842) );
  XNOR2_X1 U7525 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_66), .ZN(n6841) );
  XNOR2_X1 U7526 ( .A(BE_N_REG_3__SCAN_IN), .B(keyinput_67), .ZN(n6840) );
  NAND4_X1 U7527 ( .A1(n6843), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n6852)
         );
  XNOR2_X1 U7528 ( .A(n7340), .B(keyinput_71), .ZN(n6849) );
  XNOR2_X1 U7529 ( .A(n7336), .B(keyinput_73), .ZN(n6848) );
  XNOR2_X1 U7530 ( .A(keyinput_69), .B(BE_N_REG_1__SCAN_IN), .ZN(n6845) );
  XNOR2_X1 U7531 ( .A(keyinput_72), .B(ADDRESS_REG_28__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U7532 ( .A1(n6845), .A2(n6844), .ZN(n6847) );
  XNOR2_X1 U7533 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_70), .ZN(n6846) );
  NOR4_X1 U7534 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n6851)
         );
  INV_X1 U7535 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7332) );
  XNOR2_X1 U7536 ( .A(n7332), .B(keyinput_74), .ZN(n6850) );
  AOI21_X1 U7537 ( .B1(n6852), .B2(n6851), .A(n6850), .ZN(n6859) );
  XOR2_X1 U7538 ( .A(ADDRESS_REG_23__SCAN_IN), .B(keyinput_77), .Z(n6856) );
  INV_X1 U7539 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7328) );
  XNOR2_X1 U7540 ( .A(n7328), .B(keyinput_76), .ZN(n6855) );
  XNOR2_X1 U7541 ( .A(keyinput_75), .B(ADDRESS_REG_25__SCAN_IN), .ZN(n6854) );
  XNOR2_X1 U7542 ( .A(keyinput_78), .B(ADDRESS_REG_22__SCAN_IN), .ZN(n6853) );
  NAND4_X1 U7543 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6858)
         );
  XNOR2_X1 U7544 ( .A(keyinput_79), .B(ADDRESS_REG_21__SCAN_IN), .ZN(n6857) );
  OAI21_X1 U7545 ( .B1(n6859), .B2(n6858), .A(n6857), .ZN(n6863) );
  XNOR2_X1 U7546 ( .A(n7318), .B(keyinput_81), .ZN(n6862) );
  XNOR2_X1 U7547 ( .A(keyinput_80), .B(ADDRESS_REG_20__SCAN_IN), .ZN(n6861) );
  XNOR2_X1 U7548 ( .A(keyinput_82), .B(ADDRESS_REG_18__SCAN_IN), .ZN(n6860) );
  NAND4_X1 U7549 ( .A1(n6863), .A2(n6862), .A3(n6861), .A4(n6860), .ZN(n6867)
         );
  XOR2_X1 U7550 ( .A(keyinput_84), .B(ADDRESS_REG_16__SCAN_IN), .Z(n6866) );
  INV_X1 U7551 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7315) );
  XNOR2_X1 U7552 ( .A(n7315), .B(keyinput_83), .ZN(n6865) );
  XNOR2_X1 U7553 ( .A(keyinput_85), .B(ADDRESS_REG_15__SCAN_IN), .ZN(n6864) );
  NAND4_X1 U7554 ( .A1(n6867), .A2(n6866), .A3(n6865), .A4(n6864), .ZN(n6870)
         );
  XNOR2_X1 U7555 ( .A(n7309), .B(keyinput_86), .ZN(n6869) );
  XNOR2_X1 U7556 ( .A(keyinput_87), .B(ADDRESS_REG_13__SCAN_IN), .ZN(n6868) );
  AOI21_X1 U7557 ( .B1(n6870), .B2(n6869), .A(n6868), .ZN(n6874) );
  INV_X1 U7558 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n7306) );
  XNOR2_X1 U7559 ( .A(n7306), .B(keyinput_88), .ZN(n6873) );
  XNOR2_X1 U7560 ( .A(keyinput_90), .B(ADDRESS_REG_10__SCAN_IN), .ZN(n6872) );
  XNOR2_X1 U7561 ( .A(ADDRESS_REG_11__SCAN_IN), .B(keyinput_89), .ZN(n6871) );
  NOR4_X1 U7562 ( .A1(n6874), .A2(n6873), .A3(n6872), .A4(n6871), .ZN(n6877)
         );
  INV_X1 U7563 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7301) );
  XNOR2_X1 U7564 ( .A(n7301), .B(keyinput_92), .ZN(n6876) );
  INV_X1 U7565 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7303) );
  XNOR2_X1 U7566 ( .A(n7303), .B(keyinput_91), .ZN(n6875) );
  NOR3_X1 U7567 ( .A1(n6877), .A2(n6876), .A3(n6875), .ZN(n6883) );
  XNOR2_X1 U7568 ( .A(keyinput_93), .B(ADDRESS_REG_7__SCAN_IN), .ZN(n6882) );
  INV_X1 U7569 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7297) );
  XNOR2_X1 U7570 ( .A(n7297), .B(keyinput_94), .ZN(n6880) );
  XNOR2_X1 U7571 ( .A(ADDRESS_REG_4__SCAN_IN), .B(keyinput_96), .ZN(n6879) );
  XNOR2_X1 U7572 ( .A(keyinput_95), .B(ADDRESS_REG_5__SCAN_IN), .ZN(n6878) );
  NOR3_X1 U7573 ( .A1(n6880), .A2(n6879), .A3(n6878), .ZN(n6881) );
  OAI21_X1 U7574 ( .B1(n6883), .B2(n6882), .A(n6881), .ZN(n6890) );
  XNOR2_X1 U7575 ( .A(n7288), .B(keyinput_100), .ZN(n6887) );
  INV_X1 U7576 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7289) );
  XNOR2_X1 U7577 ( .A(n7289), .B(keyinput_99), .ZN(n6886) );
  XNOR2_X1 U7578 ( .A(keyinput_97), .B(ADDRESS_REG_3__SCAN_IN), .ZN(n6885) );
  XNOR2_X1 U7579 ( .A(keyinput_98), .B(ADDRESS_REG_2__SCAN_IN), .ZN(n6884) );
  NOR4_X1 U7580 ( .A1(n6887), .A2(n6886), .A3(n6885), .A4(n6884), .ZN(n6889)
         );
  XOR2_X1 U7581 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_101), .Z(n6888) );
  AOI21_X1 U7582 ( .B1(n6890), .B2(n6889), .A(n6888), .ZN(n6899) );
  XNOR2_X1 U7583 ( .A(DATAWIDTH_REG_2__SCAN_IN), .B(keyinput_106), .ZN(n6898)
         );
  XNOR2_X1 U7584 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_105), .ZN(n6897)
         );
  INV_X1 U7585 ( .A(keyinput_102), .ZN(n6891) );
  XNOR2_X1 U7586 ( .A(n6891), .B(STATE_REG_1__SCAN_IN), .ZN(n6895) );
  INV_X1 U7587 ( .A(keyinput_104), .ZN(n6892) );
  XNOR2_X1 U7588 ( .A(n6892), .B(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6894) );
  XNOR2_X1 U7589 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_103), .ZN(n6893) );
  NAND3_X1 U7590 ( .A1(n6895), .A2(n6894), .A3(n6893), .ZN(n6896) );
  NOR4_X1 U7591 ( .A1(n6899), .A2(n6898), .A3(n6897), .A4(n6896), .ZN(n6902)
         );
  INV_X1 U7592 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n7235) );
  XNOR2_X1 U7593 ( .A(n7235), .B(keyinput_107), .ZN(n6901) );
  INV_X1 U7594 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7236) );
  XNOR2_X1 U7595 ( .A(n7236), .B(keyinput_108), .ZN(n6900) );
  OAI21_X1 U7596 ( .B1(n6902), .B2(n6901), .A(n6900), .ZN(n6906) );
  INV_X1 U7597 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7237) );
  XNOR2_X1 U7598 ( .A(n7237), .B(keyinput_109), .ZN(n6905) );
  XNOR2_X1 U7599 ( .A(keyinput_111), .B(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6904)
         );
  XNOR2_X1 U7600 ( .A(keyinput_110), .B(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6903)
         );
  NAND4_X1 U7601 ( .A1(n6906), .A2(n6905), .A3(n6904), .A4(n6903), .ZN(n6909)
         );
  XNOR2_X1 U7602 ( .A(keyinput_113), .B(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6908)
         );
  XNOR2_X1 U7603 ( .A(keyinput_112), .B(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6907)
         );
  NAND3_X1 U7604 ( .A1(n6909), .A2(n6908), .A3(n6907), .ZN(n6912) );
  INV_X1 U7605 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7243) );
  XNOR2_X1 U7606 ( .A(n7243), .B(keyinput_115), .ZN(n6911) );
  XNOR2_X1 U7607 ( .A(keyinput_114), .B(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6910)
         );
  NAND3_X1 U7608 ( .A1(n6912), .A2(n6911), .A3(n6910), .ZN(n6915) );
  XOR2_X1 U7609 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(keyinput_117), .Z(n6914)
         );
  XNOR2_X1 U7610 ( .A(keyinput_116), .B(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6913)
         );
  NAND3_X1 U7611 ( .A1(n6915), .A2(n6914), .A3(n6913), .ZN(n6917) );
  XNOR2_X1 U7612 ( .A(keyinput_118), .B(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6916)
         );
  NAND2_X1 U7613 ( .A1(n6917), .A2(n6916), .ZN(n6923) );
  INV_X1 U7614 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n7248) );
  OAI22_X1 U7615 ( .A1(n7248), .A2(keyinput_122), .B1(
        DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput_121), .ZN(n6918) );
  AOI221_X1 U7616 ( .B1(n7248), .B2(keyinput_122), .C1(keyinput_121), .C2(
        DATAWIDTH_REG_17__SCAN_IN), .A(n6918), .ZN(n6922) );
  XOR2_X1 U7617 ( .A(DATAWIDTH_REG_15__SCAN_IN), .B(keyinput_119), .Z(n6921)
         );
  INV_X1 U7618 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n7246) );
  OAI22_X1 U7619 ( .A1(n7246), .A2(keyinput_120), .B1(
        DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput_123), .ZN(n6919) );
  AOI221_X1 U7620 ( .B1(n7246), .B2(keyinput_120), .C1(keyinput_123), .C2(
        DATAWIDTH_REG_19__SCAN_IN), .A(n6919), .ZN(n6920) );
  NAND4_X1 U7621 ( .A1(n6923), .A2(n6922), .A3(n6921), .A4(n6920), .ZN(n6926)
         );
  INV_X1 U7622 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n7250) );
  XNOR2_X1 U7623 ( .A(n7250), .B(keyinput_124), .ZN(n6925) );
  XNOR2_X1 U7624 ( .A(keyinput_125), .B(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6924)
         );
  AOI21_X1 U7625 ( .B1(n6926), .B2(n6925), .A(n6924), .ZN(n6929) );
  XNOR2_X1 U7626 ( .A(n7252), .B(keyinput_126), .ZN(n6928) );
  XNOR2_X1 U7627 ( .A(DATAWIDTH_REG_23__SCAN_IN), .B(keyinput_127), .ZN(n6927)
         );
  OAI21_X1 U7628 ( .B1(n6929), .B2(n6928), .A(n6927), .ZN(n6931) );
  XNOR2_X1 U7629 ( .A(DATAWIDTH_REG_23__SCAN_IN), .B(keyinput_255), .ZN(n6930)
         );
  OAI211_X1 U7630 ( .C1(n6933), .C2(n6932), .A(n6931), .B(n6930), .ZN(n6934)
         );
  XOR2_X1 U7631 ( .A(n6935), .B(n6934), .Z(U2890) );
  AOI21_X1 U7632 ( .B1(n7396), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6936), 
        .ZN(n6937) );
  OAI21_X1 U7633 ( .B1(n6938), .B2(n7405), .A(n6937), .ZN(n6939) );
  AOI21_X1 U7634 ( .B1(n6940), .B2(n7392), .A(n6939), .ZN(n6941) );
  OAI21_X1 U7635 ( .B1(n6942), .B2(n7626), .A(n6941), .ZN(U2956) );
  AOI21_X1 U7636 ( .B1(n6953), .B2(n7078), .A(n6943), .ZN(n6946) );
  AOI21_X1 U7637 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n7030), .A(n4243), 
        .ZN(n6945) );
  XNOR2_X1 U7638 ( .A(n6946), .B(n6945), .ZN(n7086) );
  NOR2_X1 U7639 ( .A1(n7477), .A2(n7338), .ZN(n7081) );
  AOI21_X1 U7640 ( .B1(n7396), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n7081), 
        .ZN(n6947) );
  OAI21_X1 U7641 ( .B1(n6948), .B2(n7405), .A(n6947), .ZN(n6949) );
  AOI21_X1 U7642 ( .B1(n6950), .B2(n7392), .A(n6949), .ZN(n6951) );
  OAI21_X1 U7643 ( .B1(n7626), .B2(n7086), .A(n6951), .ZN(U2957) );
  XNOR2_X1 U7644 ( .A(n6956), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n7096)
         );
  NOR2_X1 U7645 ( .A1(n7477), .A2(n7333), .ZN(n7088) );
  AOI21_X1 U7646 ( .B1(n7396), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n7088), 
        .ZN(n6957) );
  OAI21_X1 U7647 ( .B1(n6958), .B2(n7405), .A(n6957), .ZN(n6959) );
  AOI21_X1 U7648 ( .B1(n6960), .B2(n7392), .A(n6959), .ZN(n6961) );
  OAI21_X1 U7649 ( .B1(n7096), .B2(n7626), .A(n6961), .ZN(U2959) );
  XNOR2_X1 U7650 ( .A(n7030), .B(n6963), .ZN(n6964) );
  XNOR2_X1 U7651 ( .A(n6962), .B(n6964), .ZN(n7105) );
  OR2_X1 U7652 ( .A1(n7477), .A2(n7331), .ZN(n7101) );
  NAND2_X1 U7653 ( .A1(n7396), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6965)
         );
  OAI211_X1 U7654 ( .C1(n6966), .C2(n7405), .A(n7101), .B(n6965), .ZN(n6967)
         );
  AOI21_X1 U7655 ( .B1(n6968), .B2(n7392), .A(n6967), .ZN(n6969) );
  OAI21_X1 U7656 ( .B1(n7626), .B2(n7105), .A(n6969), .ZN(U2960) );
  OAI21_X1 U7657 ( .B1(n6970), .B2(n6973), .A(n6971), .ZN(n6974) );
  INV_X1 U7658 ( .A(n6974), .ZN(n7114) );
  INV_X1 U7659 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7329) );
  OR2_X1 U7660 ( .A1(n7477), .A2(n7329), .ZN(n7110) );
  NAND2_X1 U7661 ( .A1(n7396), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6975)
         );
  OAI211_X1 U7662 ( .C1(n7405), .C2(n6976), .A(n7110), .B(n6975), .ZN(n6977)
         );
  AOI21_X1 U7663 ( .B1(n6978), .B2(n7392), .A(n6977), .ZN(n6979) );
  OAI21_X1 U7664 ( .B1(n7114), .B2(n7626), .A(n6979), .ZN(U2961) );
  INV_X1 U7665 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n7018) );
  XNOR2_X1 U7666 ( .A(n7031), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7023)
         );
  XNOR2_X1 U7667 ( .A(n7031), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n7009)
         );
  AOI21_X1 U7668 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n7031), .A(n7152), 
        .ZN(n7000) );
  NAND3_X1 U7669 ( .A1(n7030), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6982) );
  NAND4_X1 U7670 ( .A1(n6980), .A2(n6981), .A3(n7031), .A4(n7018), .ZN(n6991)
         );
  XNOR2_X1 U7671 ( .A(n6983), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n7123)
         );
  NOR2_X1 U7672 ( .A1(n7477), .A2(n7326), .ZN(n7120) );
  AOI21_X1 U7673 ( .B1(n7396), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n7120), 
        .ZN(n6984) );
  OAI21_X1 U7674 ( .B1(n6985), .B2(n7405), .A(n6984), .ZN(n6986) );
  AOI21_X1 U7675 ( .B1(n6987), .B2(n7392), .A(n6986), .ZN(n6988) );
  OAI21_X1 U7676 ( .B1(n7123), .B2(n7626), .A(n6988), .ZN(U2962) );
  NAND2_X1 U7677 ( .A1(n7016), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7041) );
  NOR2_X1 U7678 ( .A1(n6989), .A2(n7041), .ZN(n7032) );
  NAND3_X1 U7679 ( .A1(n7032), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n7125), .ZN(n6990) );
  NAND2_X1 U7680 ( .A1(n6991), .A2(n6990), .ZN(n6992) );
  XNOR2_X1 U7681 ( .A(n6992), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n7132)
         );
  NAND2_X1 U7682 ( .A1(n7460), .A2(REIP_REG_23__SCAN_IN), .ZN(n7127) );
  NAND2_X1 U7683 ( .A1(n7396), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6993)
         );
  OAI211_X1 U7684 ( .C1(n7405), .C2(n6994), .A(n7127), .B(n6993), .ZN(n6995)
         );
  AOI21_X1 U7685 ( .B1(n6996), .B2(n7392), .A(n6995), .ZN(n6997) );
  OAI21_X1 U7686 ( .B1(n7132), .B2(n7626), .A(n6997), .ZN(U2963) );
  XNOR2_X1 U7687 ( .A(n7030), .B(n6998), .ZN(n6999) );
  XNOR2_X1 U7688 ( .A(n7000), .B(n6999), .ZN(n7141) );
  NOR2_X1 U7689 ( .A1(n7477), .A2(n7322), .ZN(n7135) );
  NOR2_X1 U7690 ( .A1(n7035), .A2(n7001), .ZN(n7002) );
  AOI211_X1 U7691 ( .C1(n7038), .C2(n7003), .A(n7135), .B(n7002), .ZN(n7005)
         );
  NAND2_X1 U7692 ( .A1(n7734), .A2(n7392), .ZN(n7004) );
  OAI211_X1 U7693 ( .C1(n7141), .C2(n7626), .A(n7005), .B(n7004), .ZN(U2964)
         );
  INV_X1 U7694 ( .A(n6534), .ZN(n7008) );
  INV_X1 U7695 ( .A(n7006), .ZN(n7007) );
  OAI21_X1 U7696 ( .B1(n7008), .B2(n7007), .A(n3683), .ZN(n7367) );
  INV_X1 U7697 ( .A(n7152), .ZN(n7011) );
  NAND2_X1 U7698 ( .A1(n7010), .A2(n7009), .ZN(n7142) );
  NAND3_X1 U7699 ( .A1(n7011), .A2(n7402), .A3(n7142), .ZN(n7015) );
  NAND2_X1 U7700 ( .A1(n7460), .A2(REIP_REG_21__SCAN_IN), .ZN(n7146) );
  INV_X1 U7701 ( .A(n7146), .ZN(n7013) );
  NOR2_X1 U7702 ( .A1(n7405), .A2(n7605), .ZN(n7012) );
  AOI211_X1 U7703 ( .C1(n7396), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n7013), 
        .B(n7012), .ZN(n7014) );
  OAI211_X1 U7704 ( .C1(n7059), .C2(n7367), .A(n7015), .B(n7014), .ZN(U2965)
         );
  NAND2_X1 U7705 ( .A1(n7016), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7017) );
  MUX2_X1 U7706 ( .A(n7017), .B(n7030), .S(n6980), .Z(n7019) );
  XNOR2_X1 U7707 ( .A(n7019), .B(n7018), .ZN(n7160) );
  OR2_X1 U7708 ( .A1(n7477), .A2(n7319), .ZN(n7153) );
  OAI21_X1 U7709 ( .B1(n7035), .B2(n7602), .A(n7153), .ZN(n7021) );
  NOR2_X1 U7710 ( .A1(n7596), .A2(n7059), .ZN(n7020) );
  AOI211_X1 U7711 ( .C1(n7038), .C2(n7592), .A(n7021), .B(n7020), .ZN(n7022)
         );
  OAI21_X1 U7712 ( .B1(n7160), .B2(n7626), .A(n7022), .ZN(U2966) );
  AOI21_X1 U7713 ( .B1(n7024), .B2(n7023), .A(n6980), .ZN(n7173) );
  NOR2_X1 U7714 ( .A1(n6533), .A2(n3799), .ZN(n7727) );
  NOR2_X1 U7715 ( .A1(n7477), .A2(n7317), .ZN(n7167) );
  AOI21_X1 U7716 ( .B1(n7396), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n7167), 
        .ZN(n7027) );
  OAI21_X1 U7717 ( .B1(n7580), .B2(n7405), .A(n7027), .ZN(n7028) );
  AOI21_X1 U7718 ( .B1(n7727), .B2(n7392), .A(n7028), .ZN(n7029) );
  OAI21_X1 U7719 ( .B1(n7173), .B2(n7626), .A(n7029), .ZN(U2967) );
  OAI21_X1 U7720 ( .B1(n7030), .B2(n7205), .A(n6989), .ZN(n7043) );
  NAND2_X1 U7721 ( .A1(n7031), .A2(n7179), .ZN(n7042) );
  NOR2_X1 U7722 ( .A1(n7043), .A2(n7042), .ZN(n7046) );
  NOR2_X1 U7723 ( .A1(n7046), .A2(n7032), .ZN(n7033) );
  XNOR2_X1 U7724 ( .A(n7033), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n7178)
         );
  NAND2_X1 U7725 ( .A1(n7178), .A2(n7402), .ZN(n7040) );
  NOR2_X1 U7726 ( .A1(n7477), .A2(n7314), .ZN(n7181) );
  NOR2_X1 U7727 ( .A1(n7035), .A2(n7034), .ZN(n7036) );
  AOI211_X1 U7728 ( .C1(n7038), .C2(n7037), .A(n7181), .B(n7036), .ZN(n7039)
         );
  OAI211_X1 U7729 ( .C1(n7059), .C2(n7723), .A(n7040), .B(n7039), .ZN(U2968)
         );
  INV_X1 U7730 ( .A(n7041), .ZN(n7045) );
  AND2_X1 U7731 ( .A1(n7042), .A2(n7041), .ZN(n7044) );
  MUX2_X1 U7732 ( .A(n7045), .B(n7044), .S(n7043), .Z(n7047) );
  NOR2_X1 U7733 ( .A1(n7047), .A2(n7046), .ZN(n7194) );
  NOR2_X1 U7734 ( .A1(n7477), .A2(n7313), .ZN(n7189) );
  AOI21_X1 U7735 ( .B1(n7396), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n7189), 
        .ZN(n7048) );
  OAI21_X1 U7736 ( .B1(n7049), .B2(n7405), .A(n7048), .ZN(n7050) );
  AOI21_X1 U7737 ( .B1(n7720), .B2(n7392), .A(n7050), .ZN(n7051) );
  OAI21_X1 U7738 ( .B1(n7194), .B2(n7626), .A(n7051), .ZN(U2969) );
  XNOR2_X1 U7739 ( .A(n7016), .B(n7205), .ZN(n7053) );
  XNOR2_X1 U7740 ( .A(n7052), .B(n7053), .ZN(n7197) );
  NAND2_X1 U7741 ( .A1(n7197), .A2(n7402), .ZN(n7057) );
  INV_X1 U7742 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7310) );
  NOR2_X1 U7743 ( .A1(n7477), .A2(n7310), .ZN(n7201) );
  NOR2_X1 U7744 ( .A1(n7405), .A2(n7054), .ZN(n7055) );
  AOI211_X1 U7745 ( .C1(n7396), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n7201), 
        .B(n7055), .ZN(n7056) );
  OAI211_X1 U7746 ( .C1(n7059), .C2(n7058), .A(n7057), .B(n7056), .ZN(U2970)
         );
  XNOR2_X1 U7747 ( .A(n7016), .B(n7207), .ZN(n7061) );
  XNOR2_X1 U7748 ( .A(n7060), .B(n7061), .ZN(n7213) );
  AOI22_X1 U7749 ( .A1(n7396), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n7460), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n7062) );
  OAI21_X1 U7750 ( .B1(n7063), .B2(n7405), .A(n7062), .ZN(n7064) );
  AOI21_X1 U7751 ( .B1(n7572), .B2(n7392), .A(n7064), .ZN(n7065) );
  OAI21_X1 U7752 ( .B1(n7213), .B2(n7626), .A(n7065), .ZN(U2971) );
  INV_X1 U7753 ( .A(n7066), .ZN(n7067) );
  OAI21_X1 U7754 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n7176), .A(n7067), 
        .ZN(n7072) );
  INV_X1 U7755 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n7068) );
  NOR4_X1 U7756 ( .A1(n7087), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n7069), 
        .A4(n7068), .ZN(n7070) );
  AOI211_X1 U7757 ( .C1(n7072), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n7071), .B(n7070), .ZN(n7075) );
  NAND2_X1 U7758 ( .A1(n7073), .A2(n7495), .ZN(n7074) );
  OAI211_X1 U7759 ( .C1(n7076), .C2(n7212), .A(n7075), .B(n7074), .ZN(U2987)
         );
  OAI21_X1 U7760 ( .B1(n7078), .B2(n7176), .A(n7077), .ZN(n7082) );
  INV_X1 U7761 ( .A(n7078), .ZN(n7079) );
  NOR3_X1 U7762 ( .A1(n7087), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n7079), 
        .ZN(n7080) );
  AOI211_X1 U7763 ( .C1(n7082), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n7081), .B(n7080), .ZN(n7085) );
  NAND2_X1 U7764 ( .A1(n7083), .A2(n7495), .ZN(n7084) );
  OAI211_X1 U7765 ( .C1(n7086), .C2(n7212), .A(n7085), .B(n7084), .ZN(U2989)
         );
  INV_X1 U7766 ( .A(n7087), .ZN(n7090) );
  AOI21_X1 U7767 ( .B1(n7090), .B2(n7089), .A(n7088), .ZN(n7091) );
  OAI21_X1 U7768 ( .B1(n7092), .B2(n7479), .A(n7091), .ZN(n7093) );
  AOI21_X1 U7769 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n7094), .A(n7093), 
        .ZN(n7095) );
  OAI21_X1 U7770 ( .B1(n7096), .B2(n7212), .A(n7095), .ZN(U2991) );
  INV_X1 U7771 ( .A(n7097), .ZN(n7102) );
  NOR2_X1 U7772 ( .A1(n7156), .A2(n7098), .ZN(n7108) );
  OAI211_X1 U7773 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n7108), .B(n7099), .ZN(n7100) );
  OAI211_X1 U7774 ( .C1(n7102), .C2(n7479), .A(n7101), .B(n7100), .ZN(n7103)
         );
  AOI21_X1 U7775 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n7115), .A(n7103), 
        .ZN(n7104) );
  OAI21_X1 U7776 ( .B1(n7105), .B2(n7212), .A(n7104), .ZN(U2992) );
  INV_X1 U7777 ( .A(n7106), .ZN(n7111) );
  NAND2_X1 U7778 ( .A1(n7108), .A2(n7107), .ZN(n7109) );
  OAI211_X1 U7779 ( .C1(n7111), .C2(n7479), .A(n7110), .B(n7109), .ZN(n7112)
         );
  AOI21_X1 U7780 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n7115), .A(n7112), 
        .ZN(n7113) );
  OAI21_X1 U7781 ( .B1(n7114), .B2(n7212), .A(n7113), .ZN(U2993) );
  INV_X1 U7782 ( .A(n7156), .ZN(n7170) );
  NAND3_X1 U7783 ( .A1(n7170), .A2(n7125), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n7117) );
  INV_X1 U7784 ( .A(n7115), .ZN(n7116) );
  AOI21_X1 U7785 ( .B1(n7118), .B2(n7117), .A(n7116), .ZN(n7119) );
  AOI211_X1 U7786 ( .C1(n7495), .C2(n7121), .A(n7120), .B(n7119), .ZN(n7122)
         );
  OAI21_X1 U7787 ( .B1(n7123), .B2(n7212), .A(n7122), .ZN(U2994) );
  NAND3_X1 U7788 ( .A1(n7170), .A2(n7125), .A3(n7124), .ZN(n7126) );
  OAI211_X1 U7789 ( .C1(n7128), .C2(n7479), .A(n7127), .B(n7126), .ZN(n7129)
         );
  AOI21_X1 U7790 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n7130), .A(n7129), 
        .ZN(n7131) );
  OAI21_X1 U7791 ( .B1(n7132), .B2(n7212), .A(n7131), .ZN(U2995) );
  INV_X1 U7792 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n7133) );
  NOR4_X1 U7793 ( .A1(n7156), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n7137), 
        .A4(n7133), .ZN(n7134) );
  AOI211_X1 U7794 ( .C1(n7495), .C2(n7136), .A(n7135), .B(n7134), .ZN(n7140)
         );
  NOR3_X1 U7795 ( .A1(n7156), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n7137), 
        .ZN(n7147) );
  INV_X1 U7796 ( .A(n7138), .ZN(n7149) );
  OAI21_X1 U7797 ( .B1(n7147), .B2(n7149), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n7139) );
  OAI211_X1 U7798 ( .C1(n7141), .C2(n7212), .A(n7140), .B(n7139), .ZN(U2996)
         );
  NAND2_X1 U7799 ( .A1(n7142), .A2(n7488), .ZN(n7151) );
  NAND2_X1 U7800 ( .A1(n6536), .A2(n7143), .ZN(n7144) );
  NAND2_X1 U7801 ( .A1(n7145), .A2(n7144), .ZN(n7368) );
  OAI21_X1 U7802 ( .B1(n7368), .B2(n7479), .A(n7146), .ZN(n7148) );
  AOI211_X1 U7803 ( .C1(n7149), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n7148), .B(n7147), .ZN(n7150) );
  OAI21_X1 U7804 ( .B1(n7152), .B2(n7151), .A(n7150), .ZN(U2997) );
  OAI21_X1 U7805 ( .B1(n7594), .B2(n7479), .A(n7153), .ZN(n7158) );
  NOR3_X1 U7806 ( .A1(n7156), .A2(n7155), .A3(n7154), .ZN(n7157) );
  AOI211_X1 U7807 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n7168), .A(n7158), .B(n7157), .ZN(n7159) );
  OAI21_X1 U7808 ( .B1(n7160), .B2(n7212), .A(n7159), .ZN(U2998) );
  INV_X1 U7809 ( .A(n7161), .ZN(n7165) );
  NAND2_X1 U7810 ( .A1(n7163), .A2(n7162), .ZN(n7164) );
  NAND2_X1 U7811 ( .A1(n7165), .A2(n7164), .ZN(n7583) );
  NOR2_X1 U7812 ( .A1(n7583), .A2(n7479), .ZN(n7166) );
  AOI211_X1 U7813 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n7168), .A(n7167), .B(n7166), .ZN(n7172) );
  INV_X1 U7814 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7169) );
  NAND2_X1 U7815 ( .A1(n7170), .A2(n7169), .ZN(n7171) );
  OAI211_X1 U7816 ( .C1(n7173), .C2(n7212), .A(n7172), .B(n7171), .ZN(U2999)
         );
  INV_X1 U7817 ( .A(n7187), .ZN(n7175) );
  OAI21_X1 U7818 ( .B1(n7176), .B2(n7175), .A(n7174), .ZN(n7191) );
  AOI21_X1 U7819 ( .B1(n7179), .B2(n7177), .A(n7191), .ZN(n7186) );
  NAND2_X1 U7820 ( .A1(n7178), .A2(n7488), .ZN(n7184) );
  NOR4_X1 U7821 ( .A1(n7443), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n7179), 
        .A4(n7187), .ZN(n7180) );
  AOI211_X1 U7822 ( .C1(n7495), .C2(n7182), .A(n7181), .B(n7180), .ZN(n7183)
         );
  OAI211_X1 U7823 ( .C1(n7186), .C2(n7185), .A(n7184), .B(n7183), .ZN(U3000)
         );
  NOR3_X1 U7824 ( .A1(n7443), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n7187), 
        .ZN(n7188) );
  AOI211_X1 U7825 ( .C1(n7495), .C2(n7190), .A(n7189), .B(n7188), .ZN(n7193)
         );
  NAND2_X1 U7826 ( .A1(n7191), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7192) );
  OAI211_X1 U7827 ( .C1(n7194), .C2(n7212), .A(n7193), .B(n7192), .ZN(U3001)
         );
  INV_X1 U7828 ( .A(n7199), .ZN(n7195) );
  AOI21_X1 U7829 ( .B1(n7196), .B2(n7195), .A(n7217), .ZN(n7208) );
  NAND2_X1 U7830 ( .A1(n7197), .A2(n7488), .ZN(n7204) );
  INV_X1 U7831 ( .A(n7198), .ZN(n7202) );
  NAND2_X1 U7832 ( .A1(n7199), .A2(n7219), .ZN(n7206) );
  AOI221_X1 U7833 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C1(n7205), .C2(n7207), .A(n7206), 
        .ZN(n7200) );
  AOI211_X1 U7834 ( .C1(n7202), .C2(n7495), .A(n7201), .B(n7200), .ZN(n7203)
         );
  OAI211_X1 U7835 ( .C1(n7208), .C2(n7205), .A(n7204), .B(n7203), .ZN(U3002)
         );
  INV_X1 U7836 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7571) );
  OAI22_X1 U7837 ( .A1(n7477), .A2(n7571), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n7206), .ZN(n7210) );
  NOR2_X1 U7838 ( .A1(n7208), .A2(n7207), .ZN(n7209) );
  AOI211_X1 U7839 ( .C1(n7495), .C2(n7569), .A(n7210), .B(n7209), .ZN(n7211)
         );
  OAI21_X1 U7840 ( .B1(n7213), .B2(n7212), .A(n7211), .ZN(U3003) );
  NAND2_X1 U7841 ( .A1(n7214), .A2(n7488), .ZN(n7223) );
  AOI21_X1 U7842 ( .B1(n7495), .B2(n7216), .A(n7215), .ZN(n7222) );
  NAND2_X1 U7843 ( .A1(n7217), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n7221) );
  NAND2_X1 U7844 ( .A1(n7219), .A2(n7218), .ZN(n7220) );
  NAND4_X1 U7845 ( .A1(n7223), .A2(n7222), .A3(n7221), .A4(n7220), .ZN(U3007)
         );
  AOI211_X1 U7846 ( .C1(n7231), .C2(n7225), .A(n5271), .B(n7224), .ZN(n7228)
         );
  INV_X1 U7847 ( .A(n7226), .ZN(n7227) );
  OAI22_X1 U7848 ( .A1(n7229), .A2(n7228), .B1(n7227), .B2(n7629), .ZN(n7230)
         );
  MUX2_X1 U7849 ( .A(n7231), .B(n7230), .S(n7631), .Z(U3456) );
  NOR2_X1 U7850 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7420), .ZN(n7232) );
  OR2_X1 U7851 ( .A1(n7420), .A2(STATE_REG_0__SCAN_IN), .ZN(n7716) );
  OAI21_X1 U7852 ( .B1(n7232), .B2(n7710), .A(n7716), .ZN(n7255) );
  INV_X1 U7853 ( .A(n7255), .ZN(n7699) );
  NOR2_X1 U7854 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n7411) );
  OAI21_X1 U7855 ( .B1(BS16_N), .B2(n7411), .A(n7699), .ZN(n7697) );
  OAI21_X1 U7856 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n7699), .A(n7697), .ZN(
        n7233) );
  INV_X1 U7857 ( .A(n7233), .ZN(U3451) );
  NOR2_X1 U7858 ( .A1(n7699), .A2(n7234), .ZN(U3180) );
  NOR2_X1 U7859 ( .A1(n7699), .A2(n7235), .ZN(U3179) );
  NOR2_X1 U7860 ( .A1(n7699), .A2(n7236), .ZN(U3178) );
  NOR2_X1 U7861 ( .A1(n7699), .A2(n7237), .ZN(U3177) );
  INV_X1 U7862 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7238) );
  NOR2_X1 U7863 ( .A1(n7699), .A2(n7238), .ZN(U3176) );
  NOR2_X1 U7864 ( .A1(n7699), .A2(n7239), .ZN(U3175) );
  NOR2_X1 U7865 ( .A1(n7699), .A2(n7240), .ZN(U3174) );
  INV_X1 U7866 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7241) );
  NOR2_X1 U7867 ( .A1(n7699), .A2(n7241), .ZN(U3173) );
  NOR2_X1 U7868 ( .A1(n7699), .A2(n7242), .ZN(U3172) );
  NOR2_X1 U7869 ( .A1(n7699), .A2(n7243), .ZN(U3171) );
  NOR2_X1 U7870 ( .A1(n7699), .A2(n7244), .ZN(U3170) );
  AND2_X1 U7871 ( .A1(n7255), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  INV_X1 U7872 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7245) );
  NOR2_X1 U7873 ( .A1(n7699), .A2(n7245), .ZN(U3168) );
  AND2_X1 U7874 ( .A1(n7255), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  NOR2_X1 U7875 ( .A1(n7699), .A2(n7246), .ZN(U3166) );
  NOR2_X1 U7876 ( .A1(n7699), .A2(n7247), .ZN(U3165) );
  NOR2_X1 U7877 ( .A1(n7699), .A2(n7248), .ZN(U3164) );
  NOR2_X1 U7878 ( .A1(n7699), .A2(n7249), .ZN(U3163) );
  NOR2_X1 U7879 ( .A1(n7699), .A2(n7250), .ZN(U3162) );
  INV_X1 U7880 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n7251) );
  NOR2_X1 U7881 ( .A1(n7699), .A2(n7251), .ZN(U3161) );
  NOR2_X1 U7882 ( .A1(n7699), .A2(n7252), .ZN(U3160) );
  INV_X1 U7883 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n7253) );
  NOR2_X1 U7884 ( .A1(n7699), .A2(n7253), .ZN(U3159) );
  AND2_X1 U7885 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7255), .ZN(U3158) );
  AND2_X1 U7886 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n7255), .ZN(U3157) );
  AND2_X1 U7887 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n7255), .ZN(U3156) );
  AND2_X1 U7888 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n7255), .ZN(U3155) );
  AND2_X1 U7889 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n7255), .ZN(U3154) );
  AND2_X1 U7890 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n7255), .ZN(U3153) );
  AND2_X1 U7891 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7255), .ZN(U3152) );
  AND2_X1 U7892 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7255), .ZN(U3151) );
  AND2_X1 U7893 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n7254), .ZN(U3019)
         );
  AND2_X1 U7894 ( .A1(n7268), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OAI21_X1 U7895 ( .B1(n7706), .B2(n7256), .A(n7255), .ZN(U2789) );
  AOI22_X1 U7896 ( .A1(n7427), .A2(LWORD_REG_0__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n7257) );
  OAI21_X1 U7897 ( .B1(n7258), .B2(n7286), .A(n7257), .ZN(U2923) );
  INV_X1 U7898 ( .A(EAX_REG_1__SCAN_IN), .ZN(n7260) );
  AOI22_X1 U7899 ( .A1(n7427), .A2(LWORD_REG_1__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n7259) );
  OAI21_X1 U7900 ( .B1(n7260), .B2(n7286), .A(n7259), .ZN(U2922) );
  AOI22_X1 U7901 ( .A1(n7427), .A2(LWORD_REG_2__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n7261) );
  OAI21_X1 U7902 ( .B1(n7262), .B2(n7286), .A(n7261), .ZN(U2921) );
  AOI22_X1 U7903 ( .A1(n7427), .A2(LWORD_REG_3__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n7263) );
  OAI21_X1 U7904 ( .B1(n7264), .B2(n7286), .A(n7263), .ZN(U2920) );
  AOI22_X1 U7905 ( .A1(n7427), .A2(LWORD_REG_4__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n7265) );
  OAI21_X1 U7906 ( .B1(n7266), .B2(n7286), .A(n7265), .ZN(U2919) );
  AOI22_X1 U7907 ( .A1(n7427), .A2(LWORD_REG_5__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n7267) );
  OAI21_X1 U7908 ( .B1(n4546), .B2(n7286), .A(n7267), .ZN(U2918) );
  AOI22_X1 U7909 ( .A1(n7427), .A2(LWORD_REG_6__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n7269) );
  OAI21_X1 U7910 ( .B1(n7270), .B2(n7286), .A(n7269), .ZN(U2917) );
  AOI22_X1 U7911 ( .A1(n7427), .A2(LWORD_REG_7__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n7271) );
  OAI21_X1 U7912 ( .B1(n7272), .B2(n7286), .A(n7271), .ZN(U2916) );
  AOI22_X1 U7913 ( .A1(n7427), .A2(LWORD_REG_8__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n7273) );
  OAI21_X1 U7914 ( .B1(n7274), .B2(n7286), .A(n7273), .ZN(U2915) );
  AOI22_X1 U7915 ( .A1(n7427), .A2(LWORD_REG_9__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n7275) );
  OAI21_X1 U7916 ( .B1(n7276), .B2(n7286), .A(n7275), .ZN(U2914) );
  AOI22_X1 U7917 ( .A1(n7427), .A2(LWORD_REG_10__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n7277) );
  OAI21_X1 U7918 ( .B1(n7278), .B2(n7286), .A(n7277), .ZN(U2913) );
  AOI22_X1 U7919 ( .A1(n7427), .A2(LWORD_REG_11__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n7279) );
  OAI21_X1 U7920 ( .B1(n7280), .B2(n7286), .A(n7279), .ZN(U2912) );
  AOI22_X1 U7921 ( .A1(n7427), .A2(LWORD_REG_12__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n7281) );
  OAI21_X1 U7922 ( .B1(n4625), .B2(n7286), .A(n7281), .ZN(U2911) );
  AOI22_X1 U7923 ( .A1(n7427), .A2(LWORD_REG_13__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n7282) );
  OAI21_X1 U7924 ( .B1(n7283), .B2(n7286), .A(n7282), .ZN(U2910) );
  AOI22_X1 U7925 ( .A1(n7427), .A2(LWORD_REG_14__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n7284) );
  OAI21_X1 U7926 ( .B1(n4670), .B2(n7286), .A(n7284), .ZN(U2909) );
  INV_X1 U7927 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7287) );
  AOI22_X1 U7928 ( .A1(n7427), .A2(LWORD_REG_15__SCAN_IN), .B1(n7268), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n7285) );
  OAI21_X1 U7929 ( .B1(n7287), .B2(n7286), .A(n7285), .ZN(U2908) );
  INV_X1 U7930 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7702) );
  INV_X1 U7931 ( .A(n7716), .ZN(n7719) );
  OAI222_X1 U7932 ( .A1(n7342), .A2(n7507), .B1(n7288), .B2(n7719), .C1(n7506), 
        .C2(n7334), .ZN(U3184) );
  INV_X1 U7933 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7290) );
  OAI222_X1 U7934 ( .A1(n7342), .A2(n7290), .B1(n7289), .B2(n7719), .C1(n7507), 
        .C2(n7334), .ZN(U3185) );
  OAI222_X1 U7935 ( .A1(n7342), .A2(n6156), .B1(n7291), .B2(n7719), .C1(n7290), 
        .C2(n7334), .ZN(U3186) );
  OAI222_X1 U7936 ( .A1(n7342), .A2(n7293), .B1(n7292), .B2(n7719), .C1(n6156), 
        .C2(n7334), .ZN(U3187) );
  INV_X1 U7937 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n7294) );
  OAI222_X1 U7938 ( .A1(n7342), .A2(n7295), .B1(n7294), .B2(n7719), .C1(n7293), 
        .C2(n7334), .ZN(U3188) );
  OAI222_X1 U7939 ( .A1(n7342), .A2(n7537), .B1(n7296), .B2(n7719), .C1(n7295), 
        .C2(n7334), .ZN(U3189) );
  OAI222_X1 U7940 ( .A1(n7342), .A2(n7298), .B1(n7297), .B2(n7719), .C1(n7537), 
        .C2(n7334), .ZN(U3190) );
  OAI222_X1 U7941 ( .A1(n7342), .A2(n7300), .B1(n7299), .B2(n7706), .C1(n7298), 
        .C2(n7334), .ZN(U3191) );
  OAI222_X1 U7942 ( .A1(n7342), .A2(n7302), .B1(n7301), .B2(n7719), .C1(n7300), 
        .C2(n7334), .ZN(U3192) );
  OAI222_X1 U7943 ( .A1(n7342), .A2(n6266), .B1(n7303), .B2(n7706), .C1(n7302), 
        .C2(n7334), .ZN(U3193) );
  OAI222_X1 U7944 ( .A1(n7342), .A2(n6248), .B1(n7304), .B2(n7706), .C1(n6266), 
        .C2(n7334), .ZN(U3194) );
  INV_X1 U7945 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7305) );
  OAI222_X1 U7946 ( .A1(n7334), .A2(n6248), .B1(n7305), .B2(n7706), .C1(n6296), 
        .C2(n7342), .ZN(U3195) );
  OAI222_X1 U7947 ( .A1(n7342), .A2(n7308), .B1(n7306), .B2(n7706), .C1(n6296), 
        .C2(n7334), .ZN(U3196) );
  INV_X1 U7948 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n7307) );
  OAI222_X1 U7949 ( .A1(n7334), .A2(n7308), .B1(n7307), .B2(n7706), .C1(n7571), 
        .C2(n7342), .ZN(U3197) );
  OAI222_X1 U7950 ( .A1(n7334), .A2(n7571), .B1(n7309), .B2(n7706), .C1(n7310), 
        .C2(n7342), .ZN(U3198) );
  INV_X1 U7951 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7311) );
  OAI222_X1 U7952 ( .A1(n7342), .A2(n7313), .B1(n7311), .B2(n7706), .C1(n7310), 
        .C2(n7334), .ZN(U3199) );
  OAI222_X1 U7953 ( .A1(n7334), .A2(n7313), .B1(n7312), .B2(n7706), .C1(n7314), 
        .C2(n7342), .ZN(U3200) );
  OAI222_X1 U7954 ( .A1(n7342), .A2(n7317), .B1(n7315), .B2(n7706), .C1(n7314), 
        .C2(n7334), .ZN(U3201) );
  INV_X1 U7955 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7316) );
  OAI222_X1 U7956 ( .A1(n7334), .A2(n7317), .B1(n7316), .B2(n7719), .C1(n7319), 
        .C2(n7342), .ZN(U3202) );
  OAI222_X1 U7957 ( .A1(n7334), .A2(n7319), .B1(n7318), .B2(n7719), .C1(n7321), 
        .C2(n7342), .ZN(U3203) );
  OAI222_X1 U7958 ( .A1(n7334), .A2(n7321), .B1(n7320), .B2(n7719), .C1(n7322), 
        .C2(n7342), .ZN(U3204) );
  INV_X1 U7959 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7323) );
  OAI222_X1 U7960 ( .A1(n7342), .A2(n7325), .B1(n7323), .B2(n7719), .C1(n7322), 
        .C2(n7334), .ZN(U3205) );
  OAI222_X1 U7961 ( .A1(n7334), .A2(n7325), .B1(n7324), .B2(n7706), .C1(n7326), 
        .C2(n7342), .ZN(U3206) );
  INV_X1 U7962 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7327) );
  OAI222_X1 U7963 ( .A1(n7342), .A2(n7329), .B1(n7327), .B2(n7719), .C1(n7326), 
        .C2(n7334), .ZN(U3207) );
  OAI222_X1 U7964 ( .A1(n7334), .A2(n7329), .B1(n7328), .B2(n7719), .C1(n7331), 
        .C2(n7342), .ZN(U3208) );
  INV_X1 U7965 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7330) );
  OAI222_X1 U7966 ( .A1(n7334), .A2(n7331), .B1(n7330), .B2(n7719), .C1(n7333), 
        .C2(n7342), .ZN(U3209) );
  OAI222_X1 U7967 ( .A1(n7334), .A2(n7333), .B1(n7332), .B2(n7719), .C1(n7335), 
        .C2(n7342), .ZN(U3210) );
  OAI222_X1 U7968 ( .A1(n7342), .A2(n7338), .B1(n7336), .B2(n7706), .C1(n7335), 
        .C2(n7334), .ZN(U3211) );
  INV_X1 U7969 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7337) );
  OAI222_X1 U7970 ( .A1(n7334), .A2(n7338), .B1(n7337), .B2(n7719), .C1(n7339), 
        .C2(n7342), .ZN(U3212) );
  OAI222_X1 U7971 ( .A1(n7342), .A2(n7341), .B1(n7340), .B2(n7719), .C1(n7339), 
        .C2(n7334), .ZN(U3213) );
  OAI22_X1 U7972 ( .A1(n7716), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7719), .ZN(n7343) );
  INV_X1 U7973 ( .A(n7343), .ZN(U3445) );
  AOI221_X1 U7974 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n7354) );
  NOR4_X1 U7975 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n7347) );
  NOR4_X1 U7976 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n7346) );
  NOR4_X1 U7977 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n7345) );
  NOR4_X1 U7978 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n7344) );
  NAND4_X1 U7979 ( .A1(n7347), .A2(n7346), .A3(n7345), .A4(n7344), .ZN(n7353)
         );
  NOR4_X1 U7980 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n7351) );
  AOI211_X1 U7981 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_6__SCAN_IN), .B(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n7350) );
  NOR4_X1 U7982 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(
        n7349) );
  NOR4_X1 U7983 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_17__SCAN_IN), .ZN(
        n7348) );
  NAND4_X1 U7984 ( .A1(n7351), .A2(n7350), .A3(n7349), .A4(n7348), .ZN(n7352)
         );
  NOR2_X1 U7985 ( .A1(n7353), .A2(n7352), .ZN(n7366) );
  MUX2_X1 U7986 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n7354), .S(n7366), .Z(
        U2795) );
  INV_X1 U7987 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7358) );
  AOI22_X1 U7988 ( .A1(n7719), .A2(n7358), .B1(n7355), .B2(n7716), .ZN(U3446)
         );
  AOI21_X1 U7989 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7356) );
  OAI221_X1 U7990 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7356), .C1(n7506), .C2(
        REIP_REG_0__SCAN_IN), .A(n7366), .ZN(n7357) );
  OAI21_X1 U7991 ( .B1(n7366), .B2(n7358), .A(n7357), .ZN(U3468) );
  INV_X1 U7992 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7362) );
  AOI22_X1 U7993 ( .A1(n7719), .A2(n7362), .B1(n7359), .B2(n7716), .ZN(U3447)
         );
  NOR3_X1 U7994 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n7360) );
  OAI21_X1 U7995 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7360), .A(n7366), .ZN(n7361)
         );
  OAI21_X1 U7996 ( .B1(n7366), .B2(n7362), .A(n7361), .ZN(U2794) );
  OAI22_X1 U7997 ( .A1(n7716), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        BE_N_REG_0__SCAN_IN), .B2(n7719), .ZN(n7363) );
  INV_X1 U7998 ( .A(n7363), .ZN(U3448) );
  OAI21_X1 U7999 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .A(
        n7366), .ZN(n7364) );
  OAI21_X1 U8000 ( .B1(n7366), .B2(n7365), .A(n7364), .ZN(U3469) );
  INV_X1 U8001 ( .A(EBX_REG_21__SCAN_IN), .ZN(n7371) );
  INV_X1 U8002 ( .A(n7367), .ZN(n7730) );
  INV_X1 U8003 ( .A(n7368), .ZN(n7609) );
  AOI22_X1 U8004 ( .A1(n7730), .A2(n7374), .B1(n7369), .B2(n7609), .ZN(n7370)
         );
  OAI21_X1 U8005 ( .B1(n7376), .B2(n7371), .A(n7370), .ZN(U2838) );
  INV_X1 U8006 ( .A(EBX_REG_19__SCAN_IN), .ZN(n7578) );
  NOR2_X1 U8007 ( .A1(n7583), .A2(n7372), .ZN(n7373) );
  AOI21_X1 U8008 ( .B1(n7727), .B2(n7374), .A(n7373), .ZN(n7375) );
  OAI21_X1 U8009 ( .B1(n7376), .B2(n7578), .A(n7375), .ZN(U2840) );
  AOI22_X1 U8010 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n7396), .B1(n7460), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n7381) );
  INV_X1 U8011 ( .A(n7377), .ZN(n7379) );
  AOI22_X1 U8012 ( .A1(n7379), .A2(n7402), .B1(n7392), .B2(n7378), .ZN(n7380)
         );
  OAI211_X1 U8013 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n7405), .A(n7381), 
        .B(n7380), .ZN(U2985) );
  AOI22_X1 U8014 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7396), .B1(n7460), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n7386) );
  XNOR2_X1 U8015 ( .A(n7383), .B(n7485), .ZN(n7384) );
  XNOR2_X1 U8016 ( .A(n7382), .B(n7384), .ZN(n7482) );
  AOI22_X1 U8017 ( .A1(n7392), .A2(n7514), .B1(n7482), .B2(n7402), .ZN(n7385)
         );
  OAI211_X1 U8018 ( .C1(n7405), .C2(n7518), .A(n7386), .B(n7385), .ZN(U2984)
         );
  AOI22_X1 U8019 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n7396), .B1(n7460), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n7394) );
  INV_X1 U8020 ( .A(n7387), .ZN(n7391) );
  XNOR2_X1 U8021 ( .A(n7388), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n7389)
         );
  XNOR2_X1 U8022 ( .A(n7390), .B(n7389), .ZN(n7455) );
  AOI22_X1 U8023 ( .A1(n7392), .A2(n7391), .B1(n7455), .B2(n7402), .ZN(n7393)
         );
  OAI211_X1 U8024 ( .C1(n7405), .C2(n7395), .A(n7394), .B(n7393), .ZN(U2983)
         );
  AOI22_X1 U8025 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n7396), .B1(n7460), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n7404) );
  OAI21_X1 U8026 ( .B1(n3660), .B2(n7398), .A(n7397), .ZN(n7400) );
  INV_X1 U8027 ( .A(n7400), .ZN(n7465) );
  AOI22_X1 U8028 ( .A1(n7465), .A2(n7402), .B1(n7392), .B2(n7401), .ZN(n7403)
         );
  OAI211_X1 U8029 ( .C1(n7405), .C2(n7530), .A(n7404), .B(n7403), .ZN(U2981)
         );
  NAND2_X1 U8030 ( .A1(n7693), .A2(n4331), .ZN(n7409) );
  INV_X1 U8031 ( .A(n7406), .ZN(n7407) );
  NAND2_X1 U8032 ( .A1(n7407), .A2(n7618), .ZN(n7408) );
  NAND2_X1 U8033 ( .A1(n7409), .A2(n7408), .ZN(n7625) );
  OAI21_X1 U8034 ( .B1(n7625), .B2(n7671), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n7410) );
  OAI21_X1 U8035 ( .B1(n7417), .B2(n7691), .A(n7410), .ZN(U2790) );
  INV_X1 U8036 ( .A(n7411), .ZN(n7413) );
  NOR2_X1 U8037 ( .A1(n7706), .A2(D_C_N_REG_SCAN_IN), .ZN(n7412) );
  AOI22_X1 U8038 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7706), .B1(n7413), .B2(
        n7412), .ZN(U2791) );
  INV_X1 U8039 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n7418) );
  OR2_X1 U8040 ( .A1(n3675), .A2(n7414), .ZN(n7429) );
  INV_X1 U8041 ( .A(n7429), .ZN(n7415) );
  NAND2_X1 U8042 ( .A1(n7425), .A2(n7415), .ZN(n7416) );
  OAI211_X1 U8043 ( .C1(n7425), .C2(n7418), .A(n7417), .B(n7416), .ZN(U3474)
         );
  OAI22_X1 U8044 ( .A1(n7716), .A2(n7418), .B1(W_R_N_REG_SCAN_IN), .B2(n7719), 
        .ZN(n7419) );
  INV_X1 U8045 ( .A(n7419), .ZN(U3470) );
  AND2_X1 U8046 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n7701) );
  INV_X1 U8047 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7700) );
  NOR2_X1 U8048 ( .A1(n7710), .A2(n7700), .ZN(n7708) );
  AOI21_X1 U8049 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n7708), .ZN(n7421)
         );
  NOR2_X1 U8050 ( .A1(n7420), .A2(n7709), .ZN(n7703) );
  INV_X1 U8051 ( .A(n7703), .ZN(n7714) );
  OAI211_X1 U8052 ( .C1(n7701), .C2(n7421), .A(n7428), .B(n7714), .ZN(U3182)
         );
  NOR2_X1 U8053 ( .A1(n7691), .A2(n7422), .ZN(n7670) );
  AOI21_X1 U8054 ( .B1(n7670), .B2(n7709), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n7424) );
  OAI21_X1 U8055 ( .B1(n7681), .B2(n7424), .A(n7423), .ZN(U3150) );
  AOI211_X1 U8056 ( .C1(n7427), .C2(n7709), .A(n7426), .B(n7425), .ZN(n7435)
         );
  AOI21_X1 U8057 ( .B1(n7429), .B2(n7428), .A(READY_N), .ZN(n7624) );
  OAI211_X1 U8058 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n7430), .A(n7624), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n7431) );
  NAND2_X1 U8059 ( .A1(n7431), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7434) );
  NOR2_X1 U8060 ( .A1(n7435), .A2(n7432), .ZN(n7433) );
  AOI22_X1 U8061 ( .A1(n7700), .A2(n7435), .B1(n7434), .B2(n7433), .ZN(U3472)
         );
  AOI21_X1 U8062 ( .B1(n7495), .B2(n7437), .A(n7436), .ZN(n7441) );
  AOI22_X1 U8063 ( .A1(n7439), .A2(n7488), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n7438), .ZN(n7440) );
  OAI211_X1 U8064 ( .C1(n7443), .C2(n7442), .A(n7441), .B(n7440), .ZN(U3005)
         );
  OAI211_X1 U8065 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n7452), .B(n7453), .ZN(n7450) );
  AOI22_X1 U8066 ( .A1(n7495), .A2(n7444), .B1(n7460), .B2(REIP_REG_4__SCAN_IN), .ZN(n7449) );
  INV_X1 U8067 ( .A(n7453), .ZN(n7445) );
  NAND2_X1 U8068 ( .A1(n7475), .A2(n7445), .ZN(n7476) );
  NAND2_X1 U8069 ( .A1(n7446), .A2(n7476), .ZN(n7456) );
  AOI22_X1 U8070 ( .A1(n7447), .A2(n7488), .B1(INSTADDRPOINTER_REG_4__SCAN_IN), 
        .B2(n7456), .ZN(n7448) );
  OAI211_X1 U8071 ( .C1(n7451), .C2(n7450), .A(n7449), .B(n7448), .ZN(U3014)
         );
  NAND2_X1 U8072 ( .A1(n7453), .A2(n7452), .ZN(n7459) );
  AOI22_X1 U8073 ( .A1(n7495), .A2(n7454), .B1(n7460), .B2(REIP_REG_3__SCAN_IN), .ZN(n7458) );
  AOI22_X1 U8074 ( .A1(n7456), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n7488), 
        .B2(n7455), .ZN(n7457) );
  OAI211_X1 U8075 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n7459), .A(n7458), 
        .B(n7457), .ZN(U3015) );
  AOI22_X1 U8076 ( .A1(n7495), .A2(n7519), .B1(n7460), .B2(REIP_REG_5__SCAN_IN), .ZN(n7470) );
  OAI21_X1 U8077 ( .B1(n7462), .B2(n7461), .A(n7466), .ZN(n7463) );
  AOI22_X1 U8078 ( .A1(n7465), .A2(n7488), .B1(n7464), .B2(n7463), .ZN(n7469)
         );
  NAND3_X1 U8079 ( .A1(n7471), .A2(n7467), .A3(n7466), .ZN(n7468) );
  NAND3_X1 U8080 ( .A1(n7470), .A2(n7469), .A3(n7468), .ZN(U3013) );
  NAND2_X1 U8081 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n7471), .ZN(n7486)
         );
  NOR2_X1 U8082 ( .A1(n7472), .A2(n7489), .ZN(n7474) );
  AOI21_X1 U8083 ( .B1(n7475), .B2(n7474), .A(n7473), .ZN(n7484) );
  INV_X1 U8084 ( .A(n7476), .ZN(n7481) );
  INV_X1 U8085 ( .A(n7508), .ZN(n7478) );
  OAI22_X1 U8086 ( .A1(n7479), .A2(n7478), .B1(n7507), .B2(n7477), .ZN(n7480)
         );
  AOI211_X1 U8087 ( .C1(n7488), .C2(n7482), .A(n7481), .B(n7480), .ZN(n7483)
         );
  OAI221_X1 U8088 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n7486), .C1(n7485), .C2(n7484), .A(n7483), .ZN(U3016) );
  AOI22_X1 U8089 ( .A1(n7490), .A2(n7489), .B1(n7488), .B2(n7487), .ZN(n7499)
         );
  OAI21_X1 U8090 ( .B1(n7492), .B2(n7491), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n7497) );
  INV_X1 U8091 ( .A(n7493), .ZN(n7494) );
  NAND2_X1 U8092 ( .A1(n7495), .A2(n7494), .ZN(n7496) );
  NAND4_X1 U8093 ( .A1(n7499), .A2(n7498), .A3(n7497), .A4(n7496), .ZN(U3018)
         );
  INV_X1 U8094 ( .A(n7500), .ZN(n7505) );
  NAND2_X1 U8095 ( .A1(n7501), .A2(REIP_REG_2__SCAN_IN), .ZN(n7502) );
  OAI21_X1 U8096 ( .B1(n7601), .B2(n7503), .A(n7502), .ZN(n7504) );
  AOI21_X1 U8097 ( .B1(n7505), .B2(n3668), .A(n7504), .ZN(n7517) );
  AOI22_X1 U8098 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .B1(
        n7507), .B2(n7506), .ZN(n7509) );
  AOI22_X1 U8099 ( .A1(n7510), .A2(n7509), .B1(n7520), .B2(n7508), .ZN(n7511)
         );
  OAI21_X1 U8100 ( .B1(n7512), .B2(n7577), .A(n7511), .ZN(n7513) );
  AOI21_X1 U8101 ( .B1(n7515), .B2(n7514), .A(n7513), .ZN(n7516) );
  OAI211_X1 U8102 ( .C1(n7518), .C2(n7579), .A(n7517), .B(n7516), .ZN(U2825)
         );
  INV_X1 U8103 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U8104 ( .A1(n7520), .A2(n7519), .ZN(n7521) );
  OAI211_X1 U8105 ( .C1(n7522), .C2(n7601), .A(n7521), .B(n7554), .ZN(n7526)
         );
  NOR2_X1 U8106 ( .A1(n7524), .A2(n7523), .ZN(n7525) );
  AOI211_X1 U8107 ( .C1(n7604), .C2(EBX_REG_5__SCAN_IN), .A(n7526), .B(n7525), 
        .ZN(n7529) );
  OAI21_X1 U8108 ( .B1(REIP_REG_5__SCAN_IN), .B2(n7527), .A(n7536), .ZN(n7528)
         );
  OAI211_X1 U8109 ( .C1(n7579), .C2(n7530), .A(n7529), .B(n7528), .ZN(U2822)
         );
  AOI21_X1 U8110 ( .B1(n7608), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n7582), 
        .ZN(n7542) );
  AOI22_X1 U8111 ( .A1(n7604), .A2(EBX_REG_7__SCAN_IN), .B1(n7610), .B2(n7531), 
        .ZN(n7541) );
  OAI22_X1 U8112 ( .A1(n7579), .A2(n7533), .B1(n7532), .B2(n7595), .ZN(n7534)
         );
  AOI221_X1 U8113 ( .B1(n7536), .B2(REIP_REG_7__SCAN_IN), .C1(n7535), .C2(
        REIP_REG_7__SCAN_IN), .A(n7534), .ZN(n7540) );
  NAND3_X1 U8114 ( .A1(REIP_REG_6__SCAN_IN), .A2(n7538), .A3(n7537), .ZN(n7539) );
  NAND4_X1 U8115 ( .A1(n7542), .A2(n7541), .A3(n7540), .A4(n7539), .ZN(U2820)
         );
  INV_X1 U8116 ( .A(n7543), .ZN(n7544) );
  AOI22_X1 U8117 ( .A1(n7545), .A2(n7611), .B1(n7606), .B2(n7544), .ZN(n7553)
         );
  AOI22_X1 U8118 ( .A1(n7547), .A2(REIP_REG_9__SCAN_IN), .B1(n7610), .B2(n7546), .ZN(n7548) );
  OAI211_X1 U8119 ( .C1(n7601), .C2(n7549), .A(n7548), .B(n7554), .ZN(n7550)
         );
  AOI211_X1 U8120 ( .C1(n7604), .C2(EBX_REG_9__SCAN_IN), .A(n7551), .B(n7550), 
        .ZN(n7552) );
  NAND2_X1 U8121 ( .A1(n7553), .A2(n7552), .ZN(U2818) );
  OAI21_X1 U8122 ( .B1(n7601), .B2(n7555), .A(n7554), .ZN(n7556) );
  AOI21_X1 U8123 ( .B1(n7610), .B2(n7557), .A(n7556), .ZN(n7558) );
  OAI21_X1 U8124 ( .B1(n7577), .B2(n7559), .A(n7558), .ZN(n7560) );
  AOI211_X1 U8125 ( .C1(n7562), .C2(n7611), .A(n7561), .B(n7560), .ZN(n7566)
         );
  AOI22_X1 U8126 ( .A1(n7564), .A2(n7606), .B1(REIP_REG_12__SCAN_IN), .B2(
        n7563), .ZN(n7565) );
  NAND2_X1 U8127 ( .A1(n7566), .A2(n7565), .ZN(U2815) );
  AOI22_X1 U8128 ( .A1(n7568), .A2(n7606), .B1(REIP_REG_15__SCAN_IN), .B2(
        n7567), .ZN(n7576) );
  AOI22_X1 U8129 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n7608), .B1(
        EBX_REG_15__SCAN_IN), .B2(n7604), .ZN(n7575) );
  AOI21_X1 U8130 ( .B1(n7610), .B2(n7569), .A(n7582), .ZN(n7574) );
  AOI22_X1 U8131 ( .A1(n7572), .A2(n7611), .B1(n7571), .B2(n7570), .ZN(n7573)
         );
  NAND4_X1 U8132 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(U2812)
         );
  OAI22_X1 U8133 ( .A1(n7580), .A2(n7579), .B1(n7578), .B2(n7577), .ZN(n7581)
         );
  AOI211_X1 U8134 ( .C1(n7608), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n7582), 
        .B(n7581), .ZN(n7591) );
  NOR2_X1 U8135 ( .A1(n7583), .A2(n7593), .ZN(n7584) );
  AOI21_X1 U8136 ( .B1(n7727), .B2(n7611), .A(n7584), .ZN(n7590) );
  INV_X1 U8137 ( .A(n7585), .ZN(n7588) );
  OAI22_X1 U8138 ( .A1(REIP_REG_19__SCAN_IN), .A2(n7588), .B1(n7587), .B2(
        n7586), .ZN(n7589) );
  NAND3_X1 U8139 ( .A1(n7591), .A2(n7590), .A3(n7589), .ZN(U2808) );
  AOI22_X1 U8140 ( .A1(n7592), .A2(n7606), .B1(EBX_REG_20__SCAN_IN), .B2(n7604), .ZN(n7600) );
  OAI22_X1 U8141 ( .A1(n7596), .A2(n7595), .B1(n7594), .B2(n7593), .ZN(n7597)
         );
  AOI221_X1 U8142 ( .B1(REIP_REG_20__SCAN_IN), .B2(n7603), .C1(n7598), .C2(
        n7603), .A(n7597), .ZN(n7599) );
  OAI211_X1 U8143 ( .C1(n7602), .C2(n7601), .A(n7600), .B(n7599), .ZN(U2807)
         );
  AOI22_X1 U8144 ( .A1(EBX_REG_21__SCAN_IN), .A2(n7604), .B1(
        REIP_REG_21__SCAN_IN), .B2(n7603), .ZN(n7616) );
  INV_X1 U8145 ( .A(n7605), .ZN(n7607) );
  AOI22_X1 U8146 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n7608), .B1(n7607), 
        .B2(n7606), .ZN(n7615) );
  AOI22_X1 U8147 ( .A1(n7730), .A2(n7611), .B1(n7610), .B2(n7609), .ZN(n7614)
         );
  INV_X1 U8148 ( .A(n7612), .ZN(n7613) );
  NAND4_X1 U8149 ( .A1(n7616), .A2(n7615), .A3(n7614), .A4(n7613), .ZN(U2806)
         );
  OR2_X1 U8150 ( .A1(n7693), .A2(n7617), .ZN(n7622) );
  NAND2_X1 U8151 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  NAND2_X1 U8152 ( .A1(n7693), .A2(n7620), .ZN(n7621) );
  OAI211_X1 U8153 ( .C1(n7623), .C2(n4307), .A(n7622), .B(n7621), .ZN(n7653)
         );
  OR2_X1 U8154 ( .A1(n7625), .A2(n7624), .ZN(n7657) );
  AND2_X1 U8155 ( .A1(n7688), .A2(n7657), .ZN(n7628) );
  MUX2_X1 U8156 ( .A(MORE_REG_SCAN_IN), .B(n7653), .S(n7628), .Z(U3471) );
  INV_X1 U8157 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7627) );
  OAI21_X1 U8158 ( .B1(n7628), .B2(n7627), .A(n7626), .ZN(U2793) );
  OR3_X1 U8159 ( .A1(n7630), .A2(n4330), .A3(n7629), .ZN(n7633) );
  OAI22_X1 U8160 ( .A1(n7634), .A2(n7633), .B1(n7632), .B2(n7631), .ZN(U3455)
         );
  NAND2_X1 U8161 ( .A1(n7636), .A2(n7635), .ZN(n7641) );
  INV_X1 U8162 ( .A(n7637), .ZN(n7638) );
  AOI21_X1 U8163 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7639), .A(n7638), 
        .ZN(n7640) );
  OAI211_X1 U8164 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n7641), .A(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n7640), .ZN(n7643) );
  NAND2_X1 U8165 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7641), .ZN(n7642) );
  NAND2_X1 U8166 ( .A1(n7643), .A2(n7642), .ZN(n7646) );
  INV_X1 U8167 ( .A(n7644), .ZN(n7645) );
  AOI21_X1 U8168 ( .B1(n7646), .B2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n7645), 
        .ZN(n7648) );
  NOR2_X1 U8169 ( .A1(n7646), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7647)
         );
  OAI22_X1 U8170 ( .A1(n7648), .A2(n7647), .B1(n7649), .B2(n7650), .ZN(n7652)
         );
  NAND2_X1 U8171 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  AOI21_X1 U8172 ( .B1(n7652), .B2(n7651), .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .ZN(n7663) );
  NOR2_X1 U8173 ( .A1(MORE_REG_SCAN_IN), .A2(FLUSH_REG_SCAN_IN), .ZN(n7656) );
  INV_X1 U8174 ( .A(n7653), .ZN(n7655) );
  OAI211_X1 U8175 ( .C1(n7657), .C2(n7656), .A(n7655), .B(n7654), .ZN(n7658)
         );
  INV_X1 U8176 ( .A(n7658), .ZN(n7659) );
  NAND2_X1 U8177 ( .A1(n7660), .A2(n7659), .ZN(n7661) );
  OAI22_X1 U8178 ( .A1(n7689), .A2(n7671), .B1(n7709), .B2(n7664), .ZN(n7668)
         );
  NAND2_X1 U8179 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  AOI21_X1 U8180 ( .B1(READY_N), .B2(n7669), .A(n7673), .ZN(n7686) );
  INV_X1 U8181 ( .A(n7670), .ZN(n7679) );
  OAI21_X1 U8182 ( .B1(READY_N), .B2(n7672), .A(n7671), .ZN(n7677) );
  AND2_X1 U8183 ( .A1(n7674), .A2(n7673), .ZN(n7675) );
  AOI211_X1 U8184 ( .C1(n7690), .C2(n7677), .A(n7676), .B(n7675), .ZN(n7678)
         );
  OAI21_X1 U8185 ( .B1(n7686), .B2(n7679), .A(n7678), .ZN(U3149) );
  OAI221_X1 U8186 ( .B1(n5034), .B2(STATE2_REG_0__SCAN_IN), .C1(n5034), .C2(
        n7690), .A(n7680), .ZN(U3453) );
  NAND2_X1 U8187 ( .A1(n7682), .A2(n7681), .ZN(n7685) );
  INV_X1 U8188 ( .A(n7683), .ZN(n7684) );
  OAI211_X1 U8189 ( .C1(n7686), .C2(n7691), .A(n7685), .B(n7684), .ZN(n7687)
         );
  AOI21_X1 U8190 ( .B1(n7689), .B2(n7688), .A(n7687), .ZN(n7695) );
  OAI211_X1 U8191 ( .C1(n7693), .C2(n7692), .A(n7691), .B(n7690), .ZN(n7694)
         );
  NAND2_X1 U8192 ( .A1(n7695), .A2(n7694), .ZN(U3148) );
  OAI21_X1 U8193 ( .B1(n7699), .B2(n7696), .A(n7697), .ZN(U2792) );
  INV_X1 U8194 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7698) );
  OAI21_X1 U8195 ( .B1(n7699), .B2(n7698), .A(n7697), .ZN(U3452) );
  AOI211_X1 U8196 ( .C1(HOLD), .C2(STATE_REG_1__SCAN_IN), .A(n7701), .B(n7700), 
        .ZN(n7705) );
  INV_X1 U8197 ( .A(NA_N), .ZN(n7707) );
  AOI221_X1 U8198 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7707), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7712) );
  AOI21_X1 U8199 ( .B1(n7703), .B2(n7702), .A(n7712), .ZN(n7704) );
  OAI21_X1 U8200 ( .B1(n7706), .B2(n7705), .A(n7704), .ZN(U3181) );
  AOI21_X1 U8201 ( .B1(n7708), .B2(n7707), .A(STATE_REG_2__SCAN_IN), .ZN(n7715) );
  AOI221_X1 U8202 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7709), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7711) );
  AOI221_X1 U8203 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7711), .C2(HOLD), .A(n7710), .ZN(n7713) );
  OAI22_X1 U8204 ( .A1(n7715), .A2(n7714), .B1(n7713), .B2(n7712), .ZN(U3183)
         );
  AOI22_X1 U8205 ( .A1(n7719), .A2(n7718), .B1(n7717), .B2(n7716), .ZN(U3473)
         );
  AOI22_X1 U8206 ( .A1(n7720), .A2(n3645), .B1(n7733), .B2(DATAI_1_), .ZN(
        n7722) );
  AOI22_X1 U8207 ( .A1(n7736), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n7735), .ZN(n7721) );
  NAND2_X1 U8208 ( .A1(n7722), .A2(n7721), .ZN(U2874) );
  INV_X1 U8209 ( .A(n7723), .ZN(n7724) );
  AOI22_X1 U8210 ( .A1(n7724), .A2(n3645), .B1(n7733), .B2(DATAI_2_), .ZN(
        n7726) );
  AOI22_X1 U8211 ( .A1(n7736), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n7735), .ZN(n7725) );
  NAND2_X1 U8212 ( .A1(n7726), .A2(n7725), .ZN(U2873) );
  AOI22_X1 U8213 ( .A1(n7727), .A2(n3645), .B1(n7733), .B2(DATAI_3_), .ZN(
        n7729) );
  AOI22_X1 U8214 ( .A1(n7736), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n7735), .ZN(n7728) );
  NAND2_X1 U8215 ( .A1(n7729), .A2(n7728), .ZN(U2872) );
  AOI22_X1 U8216 ( .A1(n7730), .A2(n3645), .B1(n7733), .B2(DATAI_5_), .ZN(
        n7732) );
  AOI22_X1 U8217 ( .A1(n7736), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n7735), .ZN(n7731) );
  NAND2_X1 U8218 ( .A1(n7732), .A2(n7731), .ZN(U2870) );
  AOI22_X1 U8219 ( .A1(n7734), .A2(n3645), .B1(n7733), .B2(DATAI_6_), .ZN(
        n7738) );
  AOI22_X1 U8220 ( .A1(n7736), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n7735), .ZN(n7737) );
  NAND2_X1 U8221 ( .A1(n7738), .A2(n7737), .ZN(U2869) );
  CLKBUF_X1 U3712 ( .A(n4970), .Z(n3644) );
  CLKBUF_X1 U4272 ( .A(n3641), .Z(n4797) );
endmodule

