

module b22_C_gen_AntiSAT_k_256_4 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6663, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938;

  AND2_X1 U7411 ( .A1(n14697), .A2(n9910), .ZN(n14461) );
  INV_X1 U7412 ( .A(n14646), .ZN(n14529) );
  INV_X1 U7413 ( .A(n12532), .ZN(n7140) );
  INV_X1 U7414 ( .A(n12814), .ZN(n12840) );
  NAND2_X1 U7415 ( .A1(n11639), .A2(n11638), .ZN(n15072) );
  INV_X1 U7416 ( .A(n9858), .ZN(n9660) );
  NAND2_X1 U7417 ( .A1(n7588), .A2(n12445), .ZN(n10020) );
  NAND2_X2 U7418 ( .A1(n6687), .A2(n10154), .ZN(n9997) );
  INV_X1 U7419 ( .A(n13248), .ZN(n7086) );
  NAND2_X2 U7420 ( .A1(n7296), .A2(n13248), .ZN(n9139) );
  OR2_X1 U7421 ( .A1(n8013), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8139) );
  NAND2_X2 U7422 ( .A1(n7993), .A2(n10153), .ZN(n7990) );
  INV_X1 U7423 ( .A(n10154), .ZN(n10153) );
  INV_X1 U7424 ( .A(n13249), .ZN(n6663) );
  INV_X2 U7425 ( .A(n6663), .ZN(P3_U3151) );
  INV_X1 U7426 ( .A(P3_STATE_REG_SCAN_IN), .ZN(n13249) );
  CLKBUF_X2 U7427 ( .A(n9858), .Z(n10011) );
  INV_X2 U7428 ( .A(n10011), .ZN(n10075) );
  AND2_X1 U7429 ( .A1(n8219), .A2(n7872), .ZN(n8242) );
  NAND2_X1 U7430 ( .A1(n14505), .A2(n14332), .ZN(n14306) );
  INV_X1 U7431 ( .A(n9139), .ZN(n9151) );
  INV_X4 U7432 ( .A(n13941), .ZN(n6666) );
  NAND2_X1 U7433 ( .A1(n10540), .A2(n11674), .ZN(n10725) );
  AND4_X1 U7434 ( .A1(n8722), .A2(n8724), .A3(n8723), .A4(n8725), .ZN(n11795)
         );
  XNOR2_X1 U7435 ( .A(n12960), .B(n12897), .ZN(n12958) );
  INV_X2 U7436 ( .A(n10820), .ZN(n11580) );
  OR2_X1 U7437 ( .A1(n13260), .A2(n9465), .ZN(n7545) );
  INV_X1 U7438 ( .A(n7930), .ZN(n8538) );
  INV_X1 U7439 ( .A(n13787), .ZN(n13659) );
  NAND2_X1 U7440 ( .A1(n7993), .A2(n10154), .ZN(n7938) );
  NAND2_X1 U7441 ( .A1(n7372), .A2(n7371), .ZN(n11881) );
  NAND2_X1 U7442 ( .A1(n11881), .A2(n11880), .ZN(n11886) );
  INV_X1 U7443 ( .A(n10020), .ZN(n10012) );
  XNOR2_X1 U7444 ( .A(n14646), .B(n14330), .ZN(n14520) );
  AND2_X1 U7445 ( .A1(n10725), .A2(n10724), .ZN(n13985) );
  OAI21_X1 U7446 ( .B1(n8493), .B2(n8492), .A(n8491), .ZN(n8496) );
  NAND2_X1 U7447 ( .A1(n6845), .A2(n9082), .ZN(n13125) );
  NAND2_X1 U7448 ( .A1(n9826), .A2(n9825), .ZN(n14646) );
  NOR2_X1 U7449 ( .A1(n14696), .A2(n10540), .ZN(n10732) );
  XNOR2_X1 U7450 ( .A(n8500), .B(n8499), .ZN(n12446) );
  XNOR2_X1 U7451 ( .A(n8422), .B(n8401), .ZN(n12146) );
  AND2_X1 U7452 ( .A1(n8294), .A2(n8293), .ZN(n13744) );
  INV_X1 U7453 ( .A(n10187), .ZN(n11695) );
  AND2_X1 U7454 ( .A1(n9593), .A2(n6798), .ZN(n11524) );
  XOR2_X1 U7455 ( .A(n12926), .B(n12929), .Z(n6665) );
  INV_X1 U7456 ( .A(n8666), .ZN(n8833) );
  NOR2_X2 U7457 ( .A1(n10469), .A2(n10398), .ZN(n10465) );
  NAND2_X2 U7458 ( .A1(n7905), .A2(n7807), .ZN(n7950) );
  NAND2_X2 U7459 ( .A1(n7806), .A2(n7901), .ZN(n7905) );
  NAND2_X2 U7460 ( .A1(n15925), .A2(n14771), .ZN(n14775) );
  OAI21_X2 U7461 ( .B1(n9035), .B2(n9034), .A(n9036), .ZN(n9047) );
  AOI21_X2 U7462 ( .B1(n7812), .B2(n7986), .A(n7985), .ZN(n7813) );
  NAND2_X1 U7463 ( .A1(n7809), .A2(SI_3_), .ZN(n7986) );
  AOI21_X2 U7464 ( .B1(n8192), .B2(n8191), .A(n8190), .ZN(n8211) );
  OR2_X2 U7465 ( .A1(n11728), .A2(n7250), .ZN(n7248) );
  XNOR2_X2 U7466 ( .A(n7883), .B(n7882), .ZN(n12461) );
  OR2_X2 U7467 ( .A1(n7881), .A2(n7874), .ZN(n7883) );
  AND2_X2 U7468 ( .A1(n8016), .A2(n8139), .ZN(n13399) );
  OR2_X2 U7469 ( .A1(n14411), .A2(n7503), .ZN(n7502) );
  NAND2_X2 U7470 ( .A1(n14677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9549) );
  INV_X4 U7471 ( .A(n13940), .ZN(n14045) );
  INV_X4 U7472 ( .A(n9910), .ZN(n10177) );
  AOI21_X2 U7473 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11727), .A(n11726), .ZN(
        n11950) );
  XNOR2_X2 U7474 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8676) );
  NAND2_X2 U7475 ( .A1(n8467), .A2(n8466), .ZN(n8500) );
  OR2_X4 U7476 ( .A1(n9368), .A2(n13492), .ZN(n11933) );
  XNOR2_X2 U7477 ( .A(n7876), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13492) );
  XNOR2_X2 U7478 ( .A(n8034), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13410) );
  XNOR2_X2 U7479 ( .A(n8647), .B(n8646), .ZN(n13243) );
  NOR3_X2 U7480 ( .A1(n12177), .A2(n12176), .A3(n12175), .ZN(n12720) );
  NOR3_X2 U7481 ( .A1(n11960), .A2(n11959), .A3(n11962), .ZN(n12177) );
  AOI21_X4 U7482 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n14795), .A(n15015), .ZN(
        n14829) );
  AND3_X1 U7483 ( .A1(n8447), .A2(n7614), .A3(n8446), .ZN(n7274) );
  NAND2_X1 U7484 ( .A1(n7225), .A2(n6678), .ZN(n14444) );
  OAI21_X1 U7485 ( .B1(n9064), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n9065), .ZN(
        n9078) );
  AOI211_X1 U7486 ( .C1(n9510), .C2(n12063), .A(n12062), .B(n12061), .ZN(
        n12069) );
  AOI211_X1 U7487 ( .C1(n9510), .C2(n14948), .A(n14947), .B(n14946), .ZN(
        n14951) );
  NOR2_X1 U7488 ( .A1(n12815), .A2(n7090), .ZN(n12839) );
  NOR2_X1 U7489 ( .A1(n12803), .A2(n12804), .ZN(n12815) );
  AOI211_X1 U7490 ( .C1(n9510), .C2(n15385), .A(n15384), .B(n15383), .ZN(
        n15390) );
  OAI21_X1 U7491 ( .B1(n12802), .B2(n12801), .A(n12800), .ZN(n12803) );
  NAND2_X1 U7492 ( .A1(n9711), .A2(n9710), .ZN(n11912) );
  INV_X2 U7493 ( .A(n9464), .ZN(n11089) );
  NAND2_X2 U7494 ( .A1(n14042), .A2(n15205), .ZN(n13940) );
  INV_X1 U7495 ( .A(n15424), .ZN(n11575) );
  INV_X1 U7496 ( .A(n8525), .ZN(n7173) );
  INV_X2 U7497 ( .A(n11661), .ZN(n11488) );
  CLKBUF_X2 U7498 ( .A(n7798), .Z(n14928) );
  CLKBUF_X1 U7499 ( .A(n13492), .Z(n6686) );
  CLKBUF_X2 U7500 ( .A(n9878), .Z(n6690) );
  INV_X4 U7501 ( .A(n13985), .ZN(n14043) );
  INV_X2 U7502 ( .A(n7001), .ZN(n9138) );
  NAND2_X2 U7503 ( .A1(n7086), .A2(n7296), .ZN(n9123) );
  NAND2_X1 U7506 ( .A1(n8242), .A2(n7873), .ZN(n8244) );
  OR2_X2 U7507 ( .A1(n10752), .A2(n10783), .ZN(n7257) );
  NOR2_X1 U7508 ( .A1(n6685), .A2(n9534), .ZN(n6684) );
  OAI21_X1 U7509 ( .B1(n8603), .B2(n10187), .A(n8602), .ZN(n8631) );
  OR2_X1 U7510 ( .A1(n13191), .A2(n15530), .ZN(n7118) );
  AOI21_X1 U7511 ( .B1(n9342), .B2(n6742), .A(n9346), .ZN(n7417) );
  OR2_X1 U7512 ( .A1(n13334), .A2(n13333), .ZN(n13331) );
  NAND2_X1 U7513 ( .A1(n6835), .A2(n9478), .ZN(n13334) );
  AOI21_X1 U7514 ( .B1(n8568), .B2(n6713), .A(n8567), .ZN(n7613) );
  NAND2_X1 U7515 ( .A1(n13287), .A2(n13286), .ZN(n6835) );
  NAND2_X1 U7516 ( .A1(n9137), .A2(n9136), .ZN(n13183) );
  NAND2_X1 U7517 ( .A1(n9474), .A2(n9473), .ZN(n13287) );
  NAND2_X1 U7518 ( .A1(n6675), .A2(n7606), .ZN(n14376) );
  NAND2_X1 U7519 ( .A1(n6675), .A2(n6673), .ZN(n14582) );
  NAND2_X1 U7520 ( .A1(n6676), .A2(n7607), .ZN(n6675) );
  NOR2_X1 U7521 ( .A1(n8557), .A2(n7802), .ZN(n8563) );
  INV_X1 U7522 ( .A(n14398), .ZN(n6676) );
  NAND2_X1 U7523 ( .A1(n14600), .A2(n14316), .ZN(n14398) );
  OAI22_X1 U7524 ( .A1(n13193), .A2(n13168), .B1(n15532), .B2(n13124), .ZN(
        n7117) );
  OAI21_X1 U7525 ( .B1(n12894), .B2(n7766), .A(n7764), .ZN(n12942) );
  NAND2_X1 U7526 ( .A1(n7603), .A2(n6755), .ZN(n14600) );
  NAND2_X1 U7527 ( .A1(n14444), .A2(n7601), .ZN(n7603) );
  NAND2_X1 U7528 ( .A1(n7225), .A2(n14312), .ZN(n14446) );
  NOR2_X1 U7529 ( .A1(n6674), .A2(n14375), .ZN(n6673) );
  OAI21_X1 U7530 ( .B1(n9089), .B2(n9088), .A(n9090), .ZN(n9104) );
  INV_X1 U7531 ( .A(n7606), .ZN(n6674) );
  NAND2_X1 U7532 ( .A1(n9053), .A2(n9052), .ZN(n12974) );
  NAND2_X1 U7533 ( .A1(n13527), .A2(n13526), .ZN(n13663) );
  CLKBUF_X1 U7534 ( .A(n14501), .Z(n7063) );
  NOR3_X2 U7535 ( .A1(n13694), .A2(n7233), .A3(n13858), .ZN(n13641) );
  NAND2_X1 U7536 ( .A1(n14902), .A2(n9441), .ZN(n13323) );
  NAND2_X1 U7537 ( .A1(n6834), .A2(n14897), .ZN(n14902) );
  INV_X1 U7538 ( .A(n6672), .ZN(n6671) );
  AND2_X1 U7539 ( .A1(n14442), .A2(n14312), .ZN(n6678) );
  OAI21_X1 U7540 ( .B1(n6801), .B2(n14546), .A(n14303), .ZN(n6672) );
  NAND2_X1 U7541 ( .A1(n14547), .A2(n14546), .ZN(n7599) );
  NAND2_X1 U7542 ( .A1(n9435), .A2(n9434), .ZN(n14900) );
  AND2_X1 U7543 ( .A1(n13725), .A2(n13735), .ZN(n13719) );
  NAND2_X1 U7544 ( .A1(n9928), .A2(n9927), .ZN(n14452) );
  NAND2_X1 U7545 ( .A1(n9016), .A2(n9015), .ZN(n13010) );
  NAND2_X1 U7546 ( .A1(n6729), .A2(n14301), .ZN(n6801) );
  OR2_X1 U7547 ( .A1(n14959), .A2(n14325), .ZN(n14960) );
  NAND2_X1 U7548 ( .A1(n12490), .A2(n9430), .ZN(n7567) );
  OAI21_X1 U7549 ( .B1(n14290), .B2(n14322), .A(n14293), .ZN(n14959) );
  NAND2_X1 U7550 ( .A1(n9012), .A2(n9011), .ZN(n9024) );
  NAND2_X1 U7551 ( .A1(n6677), .A2(n12245), .ZN(n14290) );
  NAND2_X1 U7552 ( .A1(n9894), .A2(n9893), .ZN(n14484) );
  NAND2_X1 U7553 ( .A1(n12237), .A2(n6836), .ZN(n12490) );
  NAND2_X1 U7554 ( .A1(n6837), .A2(n7064), .ZN(n12237) );
  NAND2_X1 U7555 ( .A1(n12053), .A2(n12052), .ZN(n12244) );
  NOR2_X1 U7556 ( .A1(n12766), .A2(n7035), .ZN(n12802) );
  OR2_X1 U7557 ( .A1(n8329), .A2(n10495), .ZN(n8305) );
  OAI21_X1 U7558 ( .B1(n8955), .B2(n7396), .A(n7393), .ZN(n8975) );
  NAND2_X1 U7559 ( .A1(n11507), .A2(n11508), .ZN(n11681) );
  NAND2_X1 U7560 ( .A1(n8942), .A2(n8941), .ZN(n8955) );
  NAND2_X1 U7561 ( .A1(n6681), .A2(n11746), .ZN(n11840) );
  OAI211_X1 U7562 ( .C1(n7227), .C2(n15072), .A(n6682), .B(n11821), .ZN(n6681)
         );
  NAND2_X1 U7563 ( .A1(n11506), .A2(n11505), .ZN(n11507) );
  OR2_X1 U7564 ( .A1(n11379), .A2(n11501), .ZN(n11506) );
  INV_X1 U7565 ( .A(n12985), .ZN(n13007) );
  OR2_X1 U7566 ( .A1(n7227), .A2(n7589), .ZN(n6682) );
  NAND2_X1 U7567 ( .A1(n8902), .A2(n8901), .ZN(n8905) );
  XNOR2_X1 U7568 ( .A(n11437), .B(n11438), .ZN(n11153) );
  NAND2_X1 U7569 ( .A1(n9723), .A2(n9722), .ZN(n11978) );
  NAND2_X1 U7570 ( .A1(n7380), .A2(n7378), .ZN(n14021) );
  NAND2_X1 U7571 ( .A1(n15929), .A2(n14779), .ZN(n14808) );
  AND2_X1 U7572 ( .A1(n11384), .A2(n11504), .ZN(n11512) );
  NAND2_X1 U7573 ( .A1(n8122), .A2(n8121), .ZN(n12064) );
  INV_X1 U7574 ( .A(n11744), .ZN(n6667) );
  NAND2_X1 U7575 ( .A1(n7833), .A2(n8118), .ZN(n10185) );
  NOR2_X1 U7576 ( .A1(n11111), .A2(n11375), .ZN(n11384) );
  NAND2_X1 U7577 ( .A1(n9697), .A2(n9696), .ZN(n11879) );
  AND2_X1 U7578 ( .A1(n8077), .A2(n8076), .ZN(n11504) );
  NAND2_X1 U7579 ( .A1(n10712), .A2(n10711), .ZN(n11272) );
  OR2_X1 U7580 ( .A1(n11110), .A2(n11211), .ZN(n11111) );
  NAND2_X1 U7581 ( .A1(n9609), .A2(n6679), .ZN(n7062) );
  AND2_X1 U7582 ( .A1(n10576), .A2(n11201), .ZN(n10905) );
  OR2_X1 U7583 ( .A1(n11004), .A2(n11005), .ZN(n7468) );
  AND2_X1 U7584 ( .A1(n11491), .A2(n9594), .ZN(n11529) );
  NAND2_X1 U7585 ( .A1(n7011), .A2(n7010), .ZN(n11491) );
  OAI21_X1 U7586 ( .B1(n11658), .B2(n11657), .A(n11473), .ZN(n6679) );
  INV_X2 U7587 ( .A(n8565), .ZN(n8545) );
  AND2_X2 U7588 ( .A1(n10865), .A2(n10864), .ZN(n12532) );
  NAND2_X1 U7589 ( .A1(n11473), .A2(n10053), .ZN(n11658) );
  AND2_X1 U7590 ( .A1(n10966), .A2(n10965), .ZN(n11003) );
  INV_X1 U7591 ( .A(n11524), .ZN(n7010) );
  BUF_X4 U7592 ( .A(n7173), .Z(n8565) );
  NAND2_X1 U7593 ( .A1(n7959), .A2(n7958), .ZN(n10580) );
  NAND2_X1 U7594 ( .A1(n7942), .A2(n7941), .ZN(n10469) );
  AND3_X1 U7595 ( .A1(n8697), .A2(n8696), .A3(n8695), .ZN(n11574) );
  CLKBUF_X1 U7596 ( .A(n8525), .Z(n7079) );
  INV_X2 U7597 ( .A(n9379), .ZN(n9464) );
  OR2_X1 U7598 ( .A1(n11661), .A2(n15142), .ZN(n11473) );
  AND3_X1 U7599 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(n12612) );
  OR2_X2 U7600 ( .A1(n10110), .A2(P2_U3088), .ZN(n13356) );
  NAND4_X1 U7601 ( .A1(n9554), .A2(n9553), .A3(n9552), .A4(n9551), .ZN(n14182)
         );
  AND4_X1 U7602 ( .A1(n9624), .A2(n9623), .A3(n9622), .A4(n9621), .ZN(n14023)
         );
  NAND4_X1 U7603 ( .A1(n9588), .A2(n9587), .A3(n9586), .A4(n9585), .ZN(n14181)
         );
  NAND4_X1 U7604 ( .A1(n7309), .A2(n8651), .A3(n8650), .A4(n8652), .ZN(n15448)
         );
  AND4_X1 U7605 ( .A1(n8687), .A2(n8686), .A3(n8685), .A4(n8684), .ZN(n15424)
         );
  OR2_X1 U7606 ( .A1(n10888), .A2(n11607), .ZN(n7247) );
  OAI21_X1 U7607 ( .B1(n8758), .B2(n7411), .A(n7408), .ZN(n8780) );
  NAND2_X1 U7608 ( .A1(n6723), .A2(n6680), .ZN(n15142) );
  NOR2_X1 U7609 ( .A1(n12426), .A2(n14689), .ZN(n10106) );
  XNOR2_X1 U7610 ( .A(n14708), .B(n7123), .ZN(n14768) );
  NAND2_X1 U7611 ( .A1(n10177), .A2(n14188), .ZN(n6680) );
  INV_X1 U7612 ( .A(n6690), .ZN(n6668) );
  INV_X1 U7613 ( .A(n7875), .ZN(n7876) );
  INV_X1 U7615 ( .A(n6688), .ZN(n6669) );
  NAND2_X1 U7616 ( .A1(n10102), .A2(n10101), .ZN(n12426) );
  INV_X2 U7617 ( .A(n10639), .ZN(n8980) );
  AND2_X1 U7618 ( .A1(n10097), .A2(n10096), .ZN(n14690) );
  AND2_X1 U7619 ( .A1(n11695), .A2(n7913), .ZN(n11228) );
  MUX2_X1 U7620 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10100), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n10102) );
  XNOR2_X1 U7621 ( .A(n9549), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7588) );
  CLKBUF_X2 U7622 ( .A(n7913), .Z(n10188) );
  NAND2_X2 U7623 ( .A1(n10501), .A2(n12857), .ZN(n10639) );
  XNOR2_X1 U7624 ( .A(n9568), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14696) );
  OAI211_X1 U7625 ( .C1(n7869), .C2(n7622), .A(n7619), .B(n7617), .ZN(n9367)
         );
  AND2_X1 U7626 ( .A1(n7871), .A2(n7877), .ZN(n10187) );
  XNOR2_X1 U7627 ( .A(n8657), .B(n8656), .ZN(n10501) );
  OAI21_X1 U7628 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14764), .A(n14799), .ZN(
        n15933) );
  XNOR2_X1 U7629 ( .A(n9547), .B(n9546), .ZN(n12445) );
  XNOR2_X1 U7630 ( .A(n9566), .B(n9562), .ZN(n11674) );
  MUX2_X1 U7631 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9558), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n9560) );
  NAND2_X2 U7632 ( .A1(n10153), .A2(P2_U3088), .ZN(n13894) );
  MUX2_X1 U7633 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7870), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n7871) );
  OAI21_X1 U7634 ( .B1(n9354), .B2(n8643), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8657) );
  NAND2_X1 U7635 ( .A1(n9559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9557) );
  XNOR2_X1 U7636 ( .A(n7880), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U7637 ( .A1(n7343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7853) );
  XNOR2_X1 U7638 ( .A(n14702), .B(n7069), .ZN(n14756) );
  OAI21_X1 U7639 ( .B1(n7163), .B2(SI_1_), .A(n7807), .ZN(n7903) );
  INV_X2 U7640 ( .A(n11561), .ZN(n6670) );
  AND2_X2 U7641 ( .A1(n6683), .A2(n6894), .ZN(n9561) );
  NOR2_X1 U7642 ( .A1(n7952), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7956) );
  INV_X1 U7643 ( .A(n9757), .ZN(n6683) );
  NAND2_X1 U7644 ( .A1(n6684), .A2(n9603), .ZN(n9757) );
  NAND2_X1 U7645 ( .A1(n7102), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8680) );
  NOR2_X1 U7646 ( .A1(n9539), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6894) );
  NOR2_X1 U7647 ( .A1(n8142), .A2(n7939), .ZN(n7846) );
  NOR2_X1 U7648 ( .A1(n10092), .A2(n9542), .ZN(n9543) );
  NAND2_X1 U7649 ( .A1(n8678), .A2(n8679), .ZN(n8709) );
  AND3_X1 U7650 ( .A1(n7845), .A2(n7844), .A3(n7843), .ZN(n8144) );
  AND2_X1 U7651 ( .A1(n7290), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14759) );
  INV_X1 U7652 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9693) );
  NOR2_X1 U7653 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n9531) );
  INV_X1 U7654 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8173) );
  INV_X1 U7655 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7834) );
  NOR2_X1 U7656 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7836) );
  INV_X4 U7657 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U7658 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9579) );
  INV_X1 U7659 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9672) );
  INV_X1 U7660 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9822) );
  INV_X1 U7661 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8746) );
  INV_X1 U7662 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9562) );
  NOR2_X1 U7663 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7845) );
  NOR2_X1 U7664 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7844) );
  NOR2_X1 U7665 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7843) );
  INV_X1 U7666 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8140) );
  NOR2_X1 U7667 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8634) );
  INV_X1 U7668 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8014) );
  INV_X1 U7669 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7953) );
  INV_X4 U7670 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  XNOR2_X1 U7671 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n6861) );
  INV_X1 U7672 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7898) );
  OAI21_X1 U7673 ( .B1(n13940), .B2(n11488), .A(n10707), .ZN(n10708) );
  NAND2_X1 U7674 ( .A1(n11272), .A2(n11271), .ZN(n7380) );
  OAI21_X2 U7675 ( .B1(n14547), .B2(n6801), .A(n6671), .ZN(n14505) );
  NAND2_X1 U7676 ( .A1(n14582), .A2(n14319), .ZN(n14320) );
  NAND2_X1 U7677 ( .A1(n12244), .A2(n12246), .ZN(n6677) );
  XNOR2_X1 U7678 ( .A(n6679), .B(n11529), .ZN(n15153) );
  INV_X2 U7679 ( .A(n15142), .ZN(n11669) );
  AND2_X2 U7680 ( .A1(n9579), .A2(n9529), .ZN(n9603) );
  NAND4_X1 U7681 ( .A1(n9531), .A2(n9530), .A3(n9689), .A4(n9693), .ZN(n6685)
         );
  NOR2_X1 U7682 ( .A1(n10886), .A2(n10770), .ZN(n10885) );
  OAI21_X2 U7683 ( .B1(n8238), .B2(n7272), .A(n7269), .ZN(n8285) );
  NOR3_X4 U7684 ( .A1(n14481), .A2(n6905), .A3(n14437), .ZN(n14433) );
  NAND2_X1 U7685 ( .A1(n10107), .A2(n15020), .ZN(n6687) );
  NAND2_X1 U7686 ( .A1(n14684), .A2(n9550), .ZN(n6688) );
  OAI222_X1 U7687 ( .A1(P1_U3086), .A2(n14684), .B1(n14694), .B2(n14683), .C1(
        n14682), .C2(n14691), .ZN(P1_U3325) );
  BUF_X4 U7688 ( .A(n9886), .Z(n6689) );
  INV_X2 U7689 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n12470) );
  AND2_X1 U7690 ( .A1(n8189), .A2(n8188), .ZN(n8190) );
  AOI22_X1 U7691 ( .A1(n8165), .A2(n8164), .B1(n8163), .B2(n8162), .ZN(n8189)
         );
  XNOR2_X2 U7692 ( .A(n7851), .B(n7850), .ZN(n8626) );
  NOR2_X2 U7693 ( .A1(n8244), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8262) );
  INV_X1 U7694 ( .A(n8545), .ZN(n6692) );
  NOR2_X2 U7695 ( .A1(n15082), .A2(n15193), .ZN(n15081) );
  NAND2_X1 U7696 ( .A1(n9910), .A2(n10153), .ZN(n9878) );
  AND2_X4 U7697 ( .A1(n13492), .A2(n7008), .ZN(n9510) );
  INV_X1 U7698 ( .A(n8525), .ZN(n6693) );
  NAND2_X4 U7699 ( .A1(n9510), .A2(n10188), .ZN(n8525) );
  AOI21_X1 U7700 ( .B1(n14368), .B2(n15189), .A(n14367), .ZN(n14587) );
  INV_X1 U7701 ( .A(n9971), .ZN(n7518) );
  NAND2_X1 U7702 ( .A1(n8641), .A2(n7753), .ZN(n6948) );
  INV_X1 U7703 ( .A(n12461), .ZN(n7884) );
  OR2_X1 U7704 ( .A1(n13711), .A2(n13556), .ZN(n13521) );
  OR2_X1 U7705 ( .A1(n14963), .A2(n14294), .ZN(n14326) );
  OR2_X1 U7706 ( .A1(n11978), .A2(n10049), .ZN(n11834) );
  NAND2_X1 U7707 ( .A1(n8167), .A2(n8166), .ZN(n8170) );
  NAND2_X1 U7708 ( .A1(n7281), .A2(n7280), .ZN(n11715) );
  INV_X1 U7709 ( .A(n11441), .ZN(n7280) );
  OR2_X1 U7710 ( .A1(n9354), .A2(n7788), .ZN(n8655) );
  NAND2_X1 U7711 ( .A1(n7460), .A2(n7791), .ZN(n7788) );
  XNOR2_X1 U7712 ( .A(n12810), .B(n12824), .ZN(n12791) );
  NAND2_X1 U7713 ( .A1(n7057), .A2(n7056), .ZN(n9582) );
  NAND2_X1 U7714 ( .A1(n11487), .A2(n9660), .ZN(n7056) );
  NAND2_X1 U7715 ( .A1(n10051), .A2(n10544), .ZN(n7505) );
  NAND2_X1 U7716 ( .A1(n7681), .A2(n6745), .ZN(n7679) );
  NAND2_X1 U7717 ( .A1(n7646), .A2(n7645), .ZN(n7644) );
  NAND2_X1 U7718 ( .A1(n8304), .A2(n7658), .ZN(n7657) );
  INV_X1 U7719 ( .A(n9942), .ZN(n7513) );
  OR2_X1 U7720 ( .A1(n7513), .A2(n9944), .ZN(n7512) );
  NAND2_X1 U7721 ( .A1(n7269), .A2(n6920), .ZN(n6919) );
  AND2_X1 U7722 ( .A1(n7717), .A2(n7268), .ZN(n7267) );
  INV_X1 U7723 ( .A(n7797), .ZN(n6920) );
  NAND2_X1 U7724 ( .A1(n7772), .A2(n13097), .ZN(n6979) );
  AND2_X1 U7725 ( .A1(n6915), .A2(n6912), .ZN(n8557) );
  NAND2_X1 U7726 ( .A1(n6914), .A2(n6913), .ZN(n6912) );
  INV_X1 U7727 ( .A(n8601), .ZN(n6915) );
  NAND2_X1 U7728 ( .A1(n8555), .A2(n8554), .ZN(n6914) );
  NAND2_X1 U7729 ( .A1(n7516), .A2(n9983), .ZN(n7515) );
  NAND2_X1 U7730 ( .A1(n6701), .A2(n7517), .ZN(n7516) );
  INV_X1 U7731 ( .A(n9982), .ZN(n7105) );
  XNOR2_X1 U7732 ( .A(n13171), .B(n7140), .ZN(n12513) );
  INV_X1 U7733 ( .A(n11800), .ZN(n7438) );
  OR2_X1 U7734 ( .A1(n13183), .A2(n9162), .ZN(n9160) );
  NAND2_X1 U7735 ( .A1(n13243), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n6988) );
  OR2_X1 U7736 ( .A1(n12910), .A2(n12916), .ZN(n9341) );
  OR2_X1 U7737 ( .A1(n13125), .A2(n12956), .ZN(n9331) );
  OR2_X1 U7738 ( .A1(n13174), .A2(n13062), .ZN(n9293) );
  NAND3_X1 U7739 ( .A1(n6967), .A2(n6965), .A3(n12070), .ZN(n7752) );
  NAND2_X1 U7740 ( .A1(n10876), .A2(n10999), .ZN(n9222) );
  OAI21_X1 U7741 ( .B1(n7044), .B2(n12929), .A(n6787), .ZN(n7043) );
  AOI21_X1 U7742 ( .B1(n12942), .B2(n12900), .A(n12899), .ZN(n12928) );
  INV_X1 U7743 ( .A(n9464), .ZN(n9487) );
  AOI21_X1 U7744 ( .B1(n6707), .B2(n6695), .A(n6758), .ZN(n7161) );
  NAND2_X1 U7745 ( .A1(n7190), .A2(n7188), .ZN(n7187) );
  INV_X1 U7746 ( .A(n11991), .ZN(n7188) );
  NOR2_X1 U7747 ( .A1(n6744), .A2(n7347), .ZN(n7346) );
  INV_X1 U7748 ( .A(n12196), .ZN(n7347) );
  INV_X1 U7749 ( .A(n7190), .ZN(n7189) );
  INV_X1 U7750 ( .A(n11990), .ZN(n7148) );
  NAND2_X1 U7751 ( .A1(n12366), .A2(n12365), .ZN(n12377) );
  INV_X1 U7752 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7835) );
  AND2_X1 U7753 ( .A1(n7839), .A2(n7838), .ZN(n8613) );
  AND2_X1 U7754 ( .A1(n7624), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n7618) );
  NAND2_X1 U7755 ( .A1(n14461), .A2(n14337), .ZN(n7480) );
  XNOR2_X1 U7756 ( .A(n14461), .B(n14311), .ZN(n14338) );
  OR2_X1 U7757 ( .A1(n14512), .A2(n14109), .ZN(n9872) );
  NAND2_X1 U7758 ( .A1(n14512), .A2(n14109), .ZN(n14333) );
  OR2_X1 U7759 ( .A1(n14650), .A2(n14132), .ZN(n14329) );
  NOR2_X1 U7760 ( .A1(n11498), .A2(n7487), .ZN(n7486) );
  INV_X1 U7761 ( .A(n14179), .ZN(n6896) );
  INV_X1 U7762 ( .A(n11674), .ZN(n10728) );
  NAND2_X1 U7763 ( .A1(n7612), .A2(n7504), .ZN(n7611) );
  INV_X1 U7764 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7612) );
  INV_X1 U7765 ( .A(n8460), .ZN(n7737) );
  NAND2_X1 U7766 ( .A1(n6934), .A2(n6933), .ZN(n8529) );
  AND2_X1 U7767 ( .A1(n7259), .A2(n7735), .ZN(n6933) );
  INV_X1 U7768 ( .A(n8526), .ZN(n7259) );
  NAND2_X1 U7769 ( .A1(n7065), .A2(SI_20_), .ZN(n8372) );
  INV_X1 U7770 ( .A(n8332), .ZN(n7065) );
  NAND2_X1 U7771 ( .A1(n8134), .A2(n10148), .ZN(n8135) );
  XNOR2_X1 U7772 ( .A(n8168), .B(SI_12_), .ZN(n8166) );
  NAND2_X1 U7773 ( .A1(n14701), .A2(n7070), .ZN(n14702) );
  NAND2_X1 U7774 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7071), .ZN(n7070) );
  INV_X1 U7775 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7071) );
  NAND2_X1 U7776 ( .A1(n14706), .A2(n14707), .ZN(n14708) );
  AND2_X1 U7777 ( .A1(n14721), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n14749) );
  OAI21_X1 U7778 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14726), .A(n14725), .ZN(
        n14787) );
  OAI211_X1 U7779 ( .C1(n12570), .C2(n7427), .A(n7432), .B(n7425), .ZN(n7424)
         );
  NAND2_X1 U7780 ( .A1(n12568), .A2(n7430), .ZN(n7429) );
  NAND2_X1 U7781 ( .A1(n12664), .A2(n7434), .ZN(n7430) );
  NAND2_X1 U7782 ( .A1(n15426), .A2(n15444), .ZN(n10867) );
  AND2_X1 U7783 ( .A1(n6959), .A2(n10987), .ZN(n15457) );
  INV_X1 U7784 ( .A(n15448), .ZN(n6959) );
  XNOR2_X1 U7785 ( .A(n14863), .B(n7140), .ZN(n12432) );
  INV_X1 U7786 ( .A(n7442), .ZN(n7441) );
  OAI21_X1 U7787 ( .B1(n7445), .B2(n7443), .A(n12621), .ZN(n7442) );
  NAND2_X1 U7788 ( .A1(n12850), .A2(n11107), .ZN(n11583) );
  INV_X1 U7789 ( .A(n9123), .ZN(n9116) );
  NAND2_X1 U7790 ( .A1(n7086), .A2(n13243), .ZN(n9154) );
  NAND2_X1 U7791 ( .A1(n7283), .A2(n7282), .ZN(n10948) );
  OR2_X1 U7792 ( .A1(n11153), .A2(n11155), .ZN(n7211) );
  AND2_X1 U7793 ( .A1(n11715), .A2(n11714), .ZN(n11943) );
  NAND2_X1 U7794 ( .A1(n7279), .A2(n7278), .ZN(n12169) );
  INV_X1 U7795 ( .A(n11948), .ZN(n7278) );
  NAND2_X1 U7796 ( .A1(n7218), .A2(n7217), .ZN(n12790) );
  INV_X1 U7797 ( .A(n12765), .ZN(n7217) );
  AND2_X1 U7798 ( .A1(n9341), .A2(n9340), .ZN(n12903) );
  NOR2_X1 U7799 ( .A1(n13047), .A2(n6811), .ZN(n13030) );
  OR2_X1 U7800 ( .A1(n13163), .A2(n13061), .ZN(n13040) );
  AND2_X1 U7801 ( .A1(n9293), .A2(n9292), .ZN(n13087) );
  OR2_X1 U7802 ( .A1(n12325), .A2(n6733), .ZN(n6937) );
  AND4_X1 U7803 ( .A1(n8862), .A2(n8861), .A3(n8860), .A4(n8859), .ZN(n12870)
         );
  AOI21_X1 U7804 ( .B1(n11600), .B2(n7307), .A(n7306), .ZN(n7305) );
  INV_X1 U7805 ( .A(n9213), .ZN(n7306) );
  INV_X2 U7806 ( .A(n9014), .ZN(n9148) );
  NAND2_X1 U7807 ( .A1(n12928), .A2(n12929), .ZN(n12927) );
  AND2_X1 U7808 ( .A1(n15416), .A2(n13122), .ZN(n15466) );
  INV_X1 U7809 ( .A(n13238), .ZN(n6994) );
  NAND2_X1 U7810 ( .A1(n9080), .A2(n9079), .ZN(n9089) );
  NOR2_X1 U7811 ( .A1(n8785), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U7812 ( .A1(n8925), .A2(n8926), .ZN(n8928) );
  NAND2_X1 U7813 ( .A1(n8905), .A2(n8904), .ZN(n8920) );
  INV_X1 U7814 ( .A(n7792), .ZN(n7755) );
  INV_X1 U7815 ( .A(n7406), .ZN(n7405) );
  OAI21_X1 U7816 ( .B1(n8800), .B2(n7407), .A(n8818), .ZN(n7406) );
  INV_X1 U7817 ( .A(n8155), .ZN(n8537) );
  AND4_X1 U7818 ( .A1(n8159), .A2(n8158), .A3(n8157), .A4(n8156), .ZN(n11996)
         );
  INV_X1 U7819 ( .A(n7960), .ZN(n8474) );
  OR2_X1 U7820 ( .A1(n8155), .A2(n7892), .ZN(n7897) );
  XNOR2_X1 U7821 ( .A(n13764), .B(n13537), .ZN(n13611) );
  AOI21_X1 U7822 ( .B1(n7196), .B2(n13522), .A(n7195), .ZN(n7194) );
  NAND2_X1 U7823 ( .A1(n7182), .A2(n13530), .ZN(n13646) );
  NAND2_X1 U7824 ( .A1(n13510), .A2(n13509), .ZN(n7342) );
  OAI21_X1 U7825 ( .B1(n12358), .B2(n7698), .A(n7696), .ZN(n13552) );
  INV_X1 U7826 ( .A(n7699), .ZN(n7698) );
  AOI21_X1 U7827 ( .B1(n7697), .B2(n7699), .A(n13509), .ZN(n7696) );
  INV_X1 U7828 ( .A(n7700), .ZN(n7697) );
  NAND2_X1 U7829 ( .A1(n7145), .A2(n7144), .ZN(n14922) );
  AND2_X1 U7830 ( .A1(n14912), .A2(n6703), .ZN(n7144) );
  NAND2_X1 U7831 ( .A1(n11989), .A2(n7147), .ZN(n7145) );
  INV_X1 U7832 ( .A(n11989), .ZN(n7151) );
  NAND2_X1 U7833 ( .A1(n8579), .A2(n11762), .ZN(n11756) );
  XNOR2_X1 U7834 ( .A(n11228), .B(n9367), .ZN(n9368) );
  NAND2_X1 U7835 ( .A1(n10461), .A2(n10462), .ZN(n10464) );
  NAND2_X1 U7836 ( .A1(n13876), .A2(n8530), .ZN(n7029) );
  INV_X2 U7837 ( .A(n7938), .ZN(n8530) );
  INV_X1 U7838 ( .A(n11860), .ZN(n15382) );
  INV_X1 U7839 ( .A(n13806), .ZN(n14915) );
  NAND2_X1 U7840 ( .A1(n13877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7880) );
  AOI21_X1 U7841 ( .B1(n6706), .B2(n7365), .A(n7360), .ZN(n7359) );
  INV_X1 U7842 ( .A(n14010), .ZN(n7360) );
  OAI22_X1 U7843 ( .A1(n11488), .A2(n13941), .B1(n11669), .B2(n13942), .ZN(
        n10706) );
  NAND2_X1 U7844 ( .A1(n15058), .A2(n9799), .ZN(n15057) );
  XNOR2_X1 U7845 ( .A(n14258), .B(n14257), .ZN(n14250) );
  AND2_X1 U7846 ( .A1(n14420), .A2(n14341), .ZN(n7503) );
  AND2_X1 U7847 ( .A1(n6895), .A2(n7472), .ZN(n14429) );
  AOI21_X1 U7848 ( .B1(n7474), .B2(n7473), .A(n6776), .ZN(n7472) );
  OAI21_X1 U7849 ( .B1(n14553), .B2(n14552), .A(n14328), .ZN(n14537) );
  INV_X1 U7850 ( .A(n6690), .ZN(n10038) );
  OR2_X1 U7851 ( .A1(n10185), .A2(n6690), .ZN(n9723) );
  INV_X1 U7852 ( .A(n9997), .ZN(n10039) );
  NAND2_X1 U7853 ( .A1(n11736), .A2(n11735), .ZN(n11820) );
  AOI21_X1 U7854 ( .B1(n11744), .B2(n7591), .A(n6764), .ZN(n7590) );
  INV_X1 U7855 ( .A(n11641), .ZN(n7591) );
  NAND2_X2 U7856 ( .A1(n10107), .A2(n15020), .ZN(n9910) );
  INV_X1 U7857 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7290) );
  OAI22_X1 U7858 ( .A1(n12507), .A2(n12506), .B1(n12871), .B2(n12505), .ZN(
        n12541) );
  NOR2_X1 U7859 ( .A1(n11716), .A2(n8828), .ZN(n11944) );
  XNOR2_X1 U7860 ( .A(n7219), .B(n12714), .ZN(n12170) );
  NOR2_X1 U7861 ( .A1(n12170), .A2(n8877), .ZN(n12710) );
  OR2_X1 U7862 ( .A1(n12713), .A2(n12717), .ZN(n12737) );
  NOR2_X1 U7863 ( .A1(n12738), .A2(n12739), .ZN(n12761) );
  OAI21_X1 U7864 ( .B1(n12791), .B2(n6829), .A(n7220), .ZN(n12835) );
  INV_X1 U7865 ( .A(n12811), .ZN(n7222) );
  INV_X1 U7866 ( .A(n12852), .ZN(n7469) );
  NAND2_X1 U7867 ( .A1(n9102), .A2(n9201), .ZN(n12920) );
  INV_X1 U7868 ( .A(n12917), .ZN(n6975) );
  OR2_X1 U7869 ( .A1(n13541), .A2(n13806), .ZN(n13548) );
  NAND2_X1 U7870 ( .A1(n14631), .A2(n6694), .ZN(n14480) );
  NAND2_X1 U7871 ( .A1(n14631), .A2(n14310), .ZN(n14478) );
  OAI21_X1 U7872 ( .B1(n7977), .B2(n7976), .A(n7975), .ZN(n7999) );
  NAND2_X1 U7873 ( .A1(n7677), .A2(n6724), .ZN(n7672) );
  INV_X1 U7874 ( .A(n7679), .ZN(n7674) );
  NAND2_X1 U7875 ( .A1(n8086), .A2(n8087), .ZN(n7676) );
  NAND2_X1 U7876 ( .A1(n7680), .A2(n7679), .ZN(n7675) );
  NOR2_X1 U7877 ( .A1(n7681), .A2(n6745), .ZN(n7680) );
  NAND2_X1 U7878 ( .A1(n8116), .A2(n8115), .ZN(n7631) );
  NAND2_X1 U7879 ( .A1(n7027), .A2(n11580), .ZN(n7026) );
  INV_X1 U7880 ( .A(n9247), .ZN(n7027) );
  AOI21_X1 U7881 ( .B1(n8116), .B2(n7634), .A(n7633), .ZN(n7632) );
  INV_X1 U7882 ( .A(n8131), .ZN(n7633) );
  NOR2_X1 U7883 ( .A1(n8132), .A2(n8114), .ZN(n7634) );
  INV_X1 U7884 ( .A(n7637), .ZN(n7636) );
  NAND2_X1 U7885 ( .A1(n7630), .A2(n7628), .ZN(n7627) );
  INV_X1 U7886 ( .A(n7632), .ZN(n7628) );
  NOR2_X1 U7887 ( .A1(n8115), .A2(n8116), .ZN(n7637) );
  OAI22_X1 U7888 ( .A1(n9662), .A2(n6882), .B1(n9663), .B2(n6881), .ZN(n9679)
         );
  NOR2_X1 U7889 ( .A1(n9661), .A2(n9664), .ZN(n6882) );
  INV_X1 U7890 ( .A(n9661), .ZN(n6881) );
  OAI22_X1 U7891 ( .A1(n9645), .A2(n7529), .B1(n9644), .B2(n7528), .ZN(n9662)
         );
  OAI21_X1 U7892 ( .B1(n9679), .B2(n6702), .A(n7054), .ZN(n9701) );
  NOR2_X1 U7893 ( .A1(n9700), .A2(n7055), .ZN(n7054) );
  INV_X1 U7894 ( .A(n7507), .ZN(n7055) );
  NAND2_X1 U7895 ( .A1(n7641), .A2(n8231), .ZN(n7640) );
  NAND2_X1 U7896 ( .A1(n6705), .A2(n7642), .ZN(n7641) );
  OR2_X1 U7897 ( .A1(n8280), .A2(n8281), .ZN(n8282) );
  NAND2_X1 U7898 ( .A1(n7649), .A2(n7647), .ZN(n8279) );
  AOI21_X1 U7899 ( .B1(n7651), .B2(n7650), .A(n7648), .ZN(n7647) );
  OAI21_X1 U7900 ( .B1(n9762), .B2(n6868), .A(n6867), .ZN(n6869) );
  NAND2_X1 U7901 ( .A1(n9764), .A2(n9761), .ZN(n6867) );
  NOR2_X1 U7902 ( .A1(n9764), .A2(n9761), .ZN(n6868) );
  NAND2_X1 U7903 ( .A1(n14322), .A2(n6760), .ZN(n7098) );
  INV_X1 U7904 ( .A(n9776), .ZN(n7531) );
  NAND2_X1 U7905 ( .A1(n9778), .A2(n9776), .ZN(n7532) );
  NOR2_X1 U7906 ( .A1(n7666), .A2(n7671), .ZN(n7665) );
  INV_X1 U7907 ( .A(n8347), .ZN(n7670) );
  NAND2_X1 U7908 ( .A1(n7013), .A2(n7012), .ZN(n9873) );
  NAND2_X1 U7909 ( .A1(n14333), .A2(n9660), .ZN(n7012) );
  NAND2_X1 U7910 ( .A1(n9872), .A2(n10011), .ZN(n7013) );
  INV_X1 U7911 ( .A(n7665), .ZN(n7661) );
  INV_X1 U7912 ( .A(n8364), .ZN(n7664) );
  NAND2_X1 U7913 ( .A1(n7665), .A2(n6699), .ZN(n7663) );
  AOI21_X1 U7914 ( .B1(n6699), .B2(n7668), .A(n8363), .ZN(n7667) );
  NAND2_X1 U7915 ( .A1(n9326), .A2(n9063), .ZN(n7021) );
  OR3_X1 U7916 ( .A1(n9323), .A2(n12891), .A3(n9322), .ZN(n9325) );
  OAI22_X1 U7917 ( .A1(n9896), .A2(n6880), .B1(n9897), .B2(n6879), .ZN(n9913)
         );
  NOR2_X1 U7918 ( .A1(n9898), .A2(n9895), .ZN(n6880) );
  INV_X1 U7919 ( .A(n9895), .ZN(n6879) );
  NAND2_X1 U7920 ( .A1(n9571), .A2(n6870), .ZN(n6872) );
  AND2_X1 U7921 ( .A1(n10724), .A2(n10728), .ZN(n6870) );
  INV_X1 U7922 ( .A(n7269), .ZN(n6921) );
  INV_X1 U7923 ( .A(n7718), .ZN(n7717) );
  OAI21_X1 U7924 ( .B1(n8328), .B2(n7719), .A(n8327), .ZN(n7718) );
  NAND2_X1 U7925 ( .A1(n7720), .A2(n8288), .ZN(n7719) );
  NAND2_X1 U7926 ( .A1(n7722), .A2(n8288), .ZN(n7721) );
  INV_X1 U7927 ( .A(n8328), .ZN(n7722) );
  NAND2_X1 U7928 ( .A1(n7251), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7250) );
  NOR2_X1 U7929 ( .A1(n12896), .A2(n7771), .ZN(n7770) );
  OAI22_X1 U7930 ( .A1(n13659), .A2(n8545), .B1(n13288), .B2(n8565), .ZN(n8443) );
  OR2_X1 U7931 ( .A1(n9973), .A2(n7518), .ZN(n7517) );
  INV_X1 U7932 ( .A(n9983), .ZN(n7106) );
  OAI21_X1 U7933 ( .B1(n9943), .B2(n6696), .A(n6780), .ZN(n9958) );
  INV_X1 U7934 ( .A(n15088), .ZN(n11493) );
  OAI211_X1 U7935 ( .C1(n6911), .C2(n6909), .A(n6908), .B(n15613), .ZN(n8424)
         );
  NOR2_X1 U7936 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9538) );
  INV_X1 U7937 ( .A(n7800), .ZN(n7272) );
  AOI21_X1 U7938 ( .B1(n7800), .B2(n7271), .A(n7270), .ZN(n7269) );
  INV_X1 U7939 ( .A(n8237), .ZN(n7271) );
  INV_X1 U7940 ( .A(n8259), .ZN(n7270) );
  AND2_X1 U7941 ( .A1(n7706), .A2(n7265), .ZN(n7264) );
  NAND2_X1 U7942 ( .A1(n7825), .A2(n7826), .ZN(n7265) );
  INV_X1 U7943 ( .A(n7826), .ZN(n7266) );
  INV_X1 U7944 ( .A(n8117), .ZN(n7705) );
  XNOR2_X1 U7945 ( .A(n13157), .B(n7140), .ZN(n12518) );
  INV_X1 U7946 ( .A(n12640), .ZN(n7136) );
  INV_X1 U7947 ( .A(n7444), .ZN(n7443) );
  XNOR2_X1 U7948 ( .A(n12532), .B(n9248), .ZN(n12102) );
  AND2_X1 U7949 ( .A1(n13183), .A2(n9162), .ZN(n9347) );
  NOR2_X1 U7950 ( .A1(n7277), .A2(n6765), .ZN(n10788) );
  INV_X1 U7951 ( .A(n12695), .ZN(n7277) );
  NAND2_X1 U7952 ( .A1(n11167), .A2(n11166), .ZN(n7246) );
  NOR2_X1 U7953 ( .A1(n7091), .A2(n12807), .ZN(n7090) );
  INV_X1 U7954 ( .A(n12816), .ZN(n7091) );
  INV_X1 U7955 ( .A(n9076), .ZN(n7320) );
  INV_X1 U7956 ( .A(n7770), .ZN(n7765) );
  NOR2_X1 U7957 ( .A1(n12958), .A2(n7768), .ZN(n7767) );
  INV_X1 U7958 ( .A(n12895), .ZN(n7768) );
  NAND2_X1 U7959 ( .A1(n12983), .A2(n12891), .ZN(n12894) );
  OR2_X1 U7960 ( .A1(n12889), .A2(n13007), .ZN(n9178) );
  INV_X1 U7961 ( .A(n12886), .ZN(n7780) );
  INV_X1 U7962 ( .A(n12888), .ZN(n7777) );
  AND2_X1 U7963 ( .A1(n12889), .A2(n13007), .ZN(n9321) );
  OR2_X1 U7964 ( .A1(n7783), .A2(n8882), .ZN(n6983) );
  NOR2_X1 U7965 ( .A1(n7784), .A2(n14856), .ZN(n7783) );
  NAND2_X1 U7966 ( .A1(n7784), .A2(n14856), .ZN(n6982) );
  INV_X1 U7967 ( .A(n9263), .ZN(n6940) );
  INV_X1 U7968 ( .A(n7314), .ZN(n7313) );
  NAND2_X1 U7969 ( .A1(n12870), .A2(n14863), .ZN(n7787) );
  INV_X1 U7970 ( .A(n6957), .ZN(n6956) );
  OAI21_X1 U7971 ( .B1(n11772), .B2(n6958), .A(n11616), .ZN(n6957) );
  INV_X1 U7972 ( .A(n9244), .ZN(n6958) );
  INV_X1 U7973 ( .A(n15396), .ZN(n12073) );
  AND2_X1 U7974 ( .A1(n15411), .A2(n6969), .ZN(n6966) );
  AND2_X1 U7975 ( .A1(n11615), .A2(n11576), .ZN(n6969) );
  AND2_X1 U7976 ( .A1(n7758), .A2(n11614), .ZN(n7757) );
  NAND2_X1 U7977 ( .A1(n7761), .A2(n7759), .ZN(n7758) );
  NOR2_X1 U7978 ( .A1(n11600), .A2(n7762), .ZN(n7761) );
  INV_X1 U7979 ( .A(n11599), .ZN(n7762) );
  NAND2_X1 U7980 ( .A1(n11596), .A2(n11595), .ZN(n7763) );
  AND3_X1 U7981 ( .A1(n8683), .A2(n8682), .A3(n8681), .ZN(n10991) );
  OR2_X1 U7982 ( .A1(n8833), .A2(SI_2_), .ZN(n8683) );
  INV_X1 U7983 ( .A(n12881), .ZN(n7331) );
  NAND2_X1 U7984 ( .A1(n13045), .A2(n9297), .ZN(n6962) );
  NAND2_X1 U7985 ( .A1(n6999), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U7986 ( .A1(n8993), .A2(n8992), .ZN(n8994) );
  INV_X1 U7987 ( .A(n8954), .ZN(n7395) );
  NAND2_X1 U7988 ( .A1(n8864), .A2(n8863), .ZN(n6852) );
  INV_X1 U7989 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7756) );
  INV_X1 U7990 ( .A(n8776), .ZN(n7409) );
  NAND2_X1 U7991 ( .A1(n10158), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U7992 ( .A1(n10247), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U7993 ( .A1(n10164), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U7994 ( .A1(n13333), .A2(n9484), .ZN(n7585) );
  INV_X1 U7995 ( .A(n9486), .ZN(n7583) );
  NAND2_X1 U7996 ( .A1(n8563), .A2(n8562), .ZN(n7093) );
  NAND2_X1 U7997 ( .A1(n13528), .A2(n13530), .ZN(n7176) );
  NOR2_X1 U7998 ( .A1(n7158), .A2(n13633), .ZN(n7157) );
  INV_X1 U7999 ( .A(n13565), .ZN(n7158) );
  INV_X1 U8000 ( .A(n11762), .ZN(n7340) );
  AND2_X1 U8001 ( .A1(n11505), .A2(n8581), .ZN(n11378) );
  INV_X1 U8002 ( .A(n10900), .ZN(n7726) );
  INV_X1 U8003 ( .A(n7495), .ZN(n7490) );
  NAND2_X1 U8004 ( .A1(n14537), .A2(n14329), .ZN(n6886) );
  NOR2_X1 U8005 ( .A1(n7494), .A2(n7493), .ZN(n7492) );
  INV_X1 U8006 ( .A(n14333), .ZN(n7494) );
  INV_X1 U8007 ( .A(n14520), .ZN(n7493) );
  NOR2_X1 U8008 ( .A1(n14963), .A2(n14275), .ZN(n14557) );
  NOR2_X1 U8009 ( .A1(n12095), .A2(n14976), .ZN(n7089) );
  XNOR2_X1 U8010 ( .A(n14819), .B(n12042), .ZN(n12086) );
  NOR3_X1 U8011 ( .A1(n14384), .A2(n14583), .A3(n14576), .ZN(n6898) );
  NOR2_X1 U8012 ( .A1(n14527), .A2(n14512), .ZN(n14508) );
  OAI21_X1 U8013 ( .B1(n8500), .B2(n7746), .A(n7744), .ZN(n8493) );
  AOI21_X1 U8014 ( .B1(n7747), .B2(n7745), .A(n6825), .ZN(n7744) );
  INV_X1 U8015 ( .A(n7747), .ZN(n7746) );
  NAND2_X1 U8016 ( .A1(n7736), .A2(n15846), .ZN(n7735) );
  INV_X1 U8017 ( .A(n8459), .ZN(n7736) );
  OR2_X1 U8018 ( .A1(n8423), .A2(n15613), .ZN(n8448) );
  INV_X1 U8019 ( .A(n8375), .ZN(n6910) );
  NAND2_X1 U8020 ( .A1(n8424), .A2(n8448), .ZN(n7739) );
  OAI211_X1 U8021 ( .C1(n8372), .C2(n8371), .A(n8370), .B(n8369), .ZN(n8374)
         );
  INV_X1 U8022 ( .A(n8378), .ZN(n8377) );
  NAND2_X1 U8023 ( .A1(n9564), .A2(n9562), .ZN(n9567) );
  NAND2_X1 U8024 ( .A1(n7824), .A2(SI_8_), .ZN(n7826) );
  INV_X1 U8025 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9529) );
  INV_X1 U8026 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9602) );
  INV_X1 U8027 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8658) );
  INV_X1 U8028 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7123) );
  OAI21_X1 U8029 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n14713), .A(n14712), .ZN(
        n14714) );
  NOR2_X1 U8030 ( .A1(n14721), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n14748) );
  INV_X1 U8031 ( .A(n7428), .ZN(n7427) );
  OAI21_X1 U8032 ( .B1(n7429), .B2(n7434), .A(n7433), .ZN(n7428) );
  NAND2_X1 U8033 ( .A1(n12567), .A2(n12943), .ZN(n7433) );
  XNOR2_X1 U8034 ( .A(n12919), .B(n7140), .ZN(n12570) );
  OAI21_X1 U8035 ( .B1(n12608), .B2(n7436), .A(n7127), .ZN(n12576) );
  AOI21_X1 U8036 ( .B1(n7435), .B2(n6714), .A(n6774), .ZN(n7127) );
  XNOR2_X1 U8037 ( .A(n13010), .B(n7140), .ZN(n12524) );
  NOR2_X1 U8038 ( .A1(n12586), .A2(n7139), .ZN(n7138) );
  INV_X1 U8039 ( .A(n12523), .ZN(n7139) );
  XNOR2_X1 U8040 ( .A(n13139), .B(n7140), .ZN(n12551) );
  OAI21_X1 U8041 ( .B1(n12549), .B2(n7458), .A(n7456), .ZN(n12527) );
  NOR2_X1 U8042 ( .A1(n12547), .A2(n12985), .ZN(n7458) );
  INV_X1 U8043 ( .A(n7457), .ZN(n7456) );
  OAI21_X1 U8044 ( .B1(n12631), .B2(n12630), .A(n12525), .ZN(n7457) );
  NAND2_X1 U8045 ( .A1(n12599), .A2(n13094), .ZN(n7444) );
  NAND2_X1 U8046 ( .A1(n7446), .A2(n13062), .ZN(n7445) );
  INV_X1 U8047 ( .A(n12599), .ZN(n7446) );
  XNOR2_X1 U8048 ( .A(n14850), .B(n7140), .ZN(n12505) );
  AND2_X1 U8049 ( .A1(n7450), .A2(n12867), .ZN(n7448) );
  NAND2_X1 U8050 ( .A1(n12608), .A2(n12609), .ZN(n12607) );
  NAND2_X1 U8051 ( .A1(n12607), .A2(n6725), .ZN(n12106) );
  XNOR2_X1 U8052 ( .A(n14838), .B(n7140), .ZN(n12539) );
  NOR2_X1 U8053 ( .A1(n7329), .A2(n7325), .ZN(n7324) );
  AND4_X1 U8054 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), .ZN(n12107)
         );
  AND2_X1 U8055 ( .A1(n8665), .A2(n8664), .ZN(n7310) );
  INV_X1 U8056 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15864) );
  NAND2_X1 U8057 ( .A1(n7247), .A2(n6728), .ZN(n7462) );
  NAND2_X1 U8058 ( .A1(n10948), .A2(n6812), .ZN(n7212) );
  NAND2_X1 U8059 ( .A1(n7468), .A2(n7467), .ZN(n11167) );
  INV_X1 U8060 ( .A(n11007), .ZN(n7467) );
  XNOR2_X1 U8061 ( .A(n7246), .B(n11157), .ZN(n11168) );
  NOR2_X1 U8062 ( .A1(n11168), .A2(n12158), .ZN(n11431) );
  NAND2_X1 U8063 ( .A1(n7211), .A2(n6727), .ZN(n7281) );
  OR2_X1 U8064 ( .A1(n11728), .A2(n12336), .ZN(n7465) );
  XNOR2_X1 U8065 ( .A(n12721), .B(n7101), .ZN(n12185) );
  NOR3_X1 U8066 ( .A1(n12720), .A2(n12719), .A3(n12718), .ZN(n12745) );
  OR2_X1 U8067 ( .A1(n12782), .A2(n12781), .ZN(n12795) );
  NAND2_X1 U8068 ( .A1(n12790), .A2(n12789), .ZN(n12810) );
  OR2_X1 U8069 ( .A1(n12791), .A2(n12792), .ZN(n7224) );
  OR2_X1 U8070 ( .A1(n12828), .A2(n12827), .ZN(n7254) );
  AOI21_X1 U8071 ( .B1(n7318), .B2(n7320), .A(n7317), .ZN(n7316) );
  INV_X1 U8072 ( .A(n9332), .ZN(n7317) );
  OR2_X1 U8073 ( .A1(n9069), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U8074 ( .A1(n12968), .A2(n9206), .ZN(n12959) );
  NAND2_X1 U8075 ( .A1(n12959), .A2(n12958), .ZN(n12957) );
  INV_X1 U8076 ( .A(n12897), .ZN(n12970) );
  AOI21_X1 U8077 ( .B1(n12981), .B2(n12982), .A(n6757), .ZN(n12969) );
  OAI21_X1 U8078 ( .B1(n12998), .B2(n9321), .A(n9178), .ZN(n12981) );
  NAND2_X1 U8079 ( .A1(n6962), .A2(n6960), .ZN(n13023) );
  NOR2_X1 U8080 ( .A1(n13020), .A2(n6961), .ZN(n6960) );
  INV_X1 U8081 ( .A(n7330), .ZN(n6961) );
  AND2_X1 U8082 ( .A1(n9177), .A2(n12888), .ZN(n13008) );
  NAND2_X1 U8083 ( .A1(n13029), .A2(n12884), .ZN(n13016) );
  AND3_X1 U8084 ( .A1(n9005), .A2(n9004), .A3(n9003), .ZN(n13031) );
  NAND2_X1 U8085 ( .A1(n13030), .A2(n13041), .ZN(n13029) );
  NAND2_X1 U8086 ( .A1(n13069), .A2(n9296), .ZN(n13045) );
  NAND2_X1 U8087 ( .A1(n6821), .A2(n12875), .ZN(n13076) );
  AND2_X1 U8088 ( .A1(n12876), .A2(n12875), .ZN(n7772) );
  INV_X1 U8089 ( .A(n6939), .ZN(n6938) );
  OAI21_X1 U8090 ( .B1(n6733), .B2(n12334), .A(n7311), .ZN(n6939) );
  AOI21_X1 U8091 ( .B1(n7312), .B2(n7314), .A(n6741), .ZN(n7311) );
  INV_X1 U8092 ( .A(n14861), .ZN(n7312) );
  INV_X1 U8093 ( .A(n12334), .ZN(n12331) );
  AND2_X1 U8094 ( .A1(n9275), .A2(n9274), .ZN(n14861) );
  NAND2_X1 U8095 ( .A1(n12324), .A2(n9263), .ZN(n14862) );
  NAND2_X1 U8096 ( .A1(n14862), .A2(n14861), .ZN(n14860) );
  AOI21_X1 U8097 ( .B1(n7301), .B2(n9265), .A(n9262), .ZN(n7300) );
  INV_X1 U8098 ( .A(n8808), .ZN(n7301) );
  AND2_X1 U8099 ( .A1(n11581), .A2(n11580), .ZN(n15447) );
  NAND2_X1 U8100 ( .A1(n7761), .A2(n7763), .ZN(n11777) );
  AND4_X1 U8101 ( .A1(n8740), .A2(n8739), .A3(n8738), .A4(n8737), .ZN(n12613)
         );
  NAND2_X1 U8102 ( .A1(n6935), .A2(n9230), .ZN(n11566) );
  NAND2_X1 U8103 ( .A1(n11566), .A2(n7759), .ZN(n11568) );
  AND4_X1 U8104 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n15408)
         );
  OR2_X1 U8105 ( .A1(n9154), .A2(n10764), .ZN(n8700) );
  INV_X1 U8106 ( .A(n15447), .ZN(n15425) );
  OR2_X1 U8107 ( .A1(n9154), .A2(n10666), .ZN(n8672) );
  NAND2_X1 U8108 ( .A1(n10874), .A2(n11580), .ZN(n15450) );
  NAND2_X1 U8109 ( .A1(n12905), .A2(n15453), .ZN(n6986) );
  INV_X1 U8110 ( .A(n7043), .ZN(n7773) );
  AND2_X1 U8111 ( .A1(n9204), .A2(n9202), .ZN(n12919) );
  AND2_X1 U8112 ( .A1(n10198), .A2(n10604), .ZN(n10618) );
  OAI22_X1 U8113 ( .A1(n9131), .A2(n9130), .B1(P2_DATAO_REG_29__SCAN_IN), .B2(
        n12460), .ZN(n9145) );
  OR2_X1 U8114 ( .A1(n9145), .A2(n9144), .ZN(n9147) );
  NAND2_X1 U8115 ( .A1(n9024), .A2(n9023), .ZN(n9035) );
  AND2_X1 U8116 ( .A1(n9172), .A2(n9349), .ZN(n10860) );
  NAND2_X1 U8117 ( .A1(n8994), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U8118 ( .A1(n8975), .A2(n8974), .ZN(n8993) );
  NAND2_X1 U8119 ( .A1(n7397), .A2(n7398), .ZN(n8942) );
  AOI21_X1 U8120 ( .B1(n7400), .B2(n7402), .A(n7399), .ZN(n7398) );
  INV_X1 U8121 ( .A(n8938), .ZN(n7399) );
  INV_X1 U8122 ( .A(n7401), .ZN(n7400) );
  OAI21_X1 U8123 ( .B1(n8904), .B2(n7402), .A(n8922), .ZN(n7401) );
  INV_X1 U8124 ( .A(n8919), .ZN(n7402) );
  OR2_X1 U8125 ( .A1(n6852), .A2(n10457), .ZN(n8865) );
  NOR2_X1 U8126 ( .A1(n8785), .A2(n7754), .ZN(n8868) );
  NAND2_X1 U8127 ( .A1(n8840), .A2(n8839), .ZN(n8845) );
  INV_X1 U8128 ( .A(n8815), .ZN(n7407) );
  AND2_X1 U8129 ( .A1(n8815), .A2(n8799), .ZN(n8800) );
  NAND2_X1 U8130 ( .A1(n8801), .A2(n8800), .ZN(n8816) );
  NAND2_X1 U8131 ( .A1(n8780), .A2(n8779), .ZN(n8798) );
  NOR2_X1 U8132 ( .A1(n8761), .A2(n7413), .ZN(n7412) );
  INV_X1 U8133 ( .A(n8759), .ZN(n7413) );
  NAND2_X1 U8134 ( .A1(n8758), .A2(n8757), .ZN(n7414) );
  NAND2_X1 U8135 ( .A1(n6846), .A2(n8744), .ZN(n8758) );
  NAND2_X1 U8136 ( .A1(n8743), .A2(n8742), .ZN(n6846) );
  INV_X1 U8137 ( .A(n8741), .ZN(n8742) );
  INV_X1 U8138 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8711) );
  OR2_X1 U8139 ( .A1(n8709), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8710) );
  INV_X1 U8140 ( .A(n8688), .ZN(n6848) );
  INV_X1 U8141 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8679) );
  AND2_X1 U8142 ( .A1(n9432), .A2(n9431), .ZN(n7564) );
  OR2_X1 U8143 ( .A1(n9432), .A2(n7566), .ZN(n7565) );
  INV_X1 U8144 ( .A(n9431), .ZN(n7566) );
  OAI21_X1 U8145 ( .B1(n9442), .B2(n7552), .A(n13272), .ZN(n7551) );
  INV_X1 U8146 ( .A(n7561), .ZN(n7560) );
  AOI21_X1 U8147 ( .B1(n7561), .B2(n13305), .A(n6784), .ZN(n7559) );
  NOR2_X1 U8148 ( .A1(n13279), .A2(n7562), .ZN(n7561) );
  XNOR2_X1 U8149 ( .A(n9379), .B(n8585), .ZN(n10740) );
  NAND2_X1 U8150 ( .A1(n8295), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U8151 ( .A1(n6843), .A2(n9395), .ZN(n11120) );
  INV_X1 U8152 ( .A(n11228), .ZN(n9369) );
  NOR2_X1 U8153 ( .A1(n8601), .A2(n8600), .ZN(n8606) );
  AND2_X1 U8154 ( .A1(n8524), .A2(n8523), .ZN(n13573) );
  AND2_X1 U8155 ( .A1(n8544), .A2(n8543), .ZN(n13571) );
  AND3_X1 U8156 ( .A1(n8316), .A2(n8315), .A3(n8314), .ZN(n13555) );
  NAND2_X1 U8157 ( .A1(n8150), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U8158 ( .A1(n13618), .A2(n13570), .ZN(n7714) );
  NAND2_X1 U8159 ( .A1(n13636), .A2(n13568), .ZN(n13618) );
  NAND2_X1 U8160 ( .A1(n13566), .A2(n7157), .ZN(n13636) );
  NAND2_X1 U8161 ( .A1(n7183), .A2(n7184), .ZN(n7182) );
  INV_X1 U8162 ( .A(n13663), .ZN(n7183) );
  AND2_X1 U8163 ( .A1(n8410), .A2(n8409), .ZN(n13561) );
  INV_X1 U8164 ( .A(n13558), .ZN(n7730) );
  INV_X1 U8165 ( .A(n7197), .ZN(n7196) );
  OAI21_X1 U8166 ( .B1(n7198), .B2(n13522), .A(n13524), .ZN(n7197) );
  NOR2_X1 U8167 ( .A1(n7199), .A2(n13691), .ZN(n7198) );
  NAND2_X1 U8168 ( .A1(n7160), .A2(n7161), .ZN(n13690) );
  OR2_X1 U8169 ( .A1(n13733), .A2(n13747), .ZN(n13731) );
  OAI21_X1 U8170 ( .B1(n12377), .B2(n12376), .A(n12378), .ZN(n13510) );
  AOI21_X1 U8171 ( .B1(n7700), .B2(n12362), .A(n6770), .ZN(n7699) );
  AND2_X1 U8172 ( .A1(n12359), .A2(n7702), .ZN(n7700) );
  NAND2_X1 U8173 ( .A1(n7703), .A2(n12368), .ZN(n7702) );
  OR2_X1 U8174 ( .A1(n12358), .A2(n12362), .ZN(n7701) );
  NOR2_X1 U8175 ( .A1(n12193), .A2(n7191), .ZN(n7190) );
  INV_X1 U8176 ( .A(n11993), .ZN(n7191) );
  NAND2_X1 U8177 ( .A1(n12195), .A2(n12477), .ZN(n7152) );
  NAND2_X1 U8178 ( .A1(n7147), .A2(n11988), .ZN(n7146) );
  NAND2_X1 U8179 ( .A1(n11992), .A2(n11991), .ZN(n7192) );
  AOI21_X1 U8180 ( .B1(n7143), .B2(n11683), .A(n6817), .ZN(n7732) );
  INV_X1 U8181 ( .A(n6734), .ZN(n7143) );
  OR2_X1 U8182 ( .A1(n8079), .A2(n8078), .ZN(n8100) );
  OAI21_X1 U8183 ( .B1(n7339), .B2(n11073), .A(n11075), .ZN(n7338) );
  NOR2_X1 U8184 ( .A1(n7339), .A2(n7201), .ZN(n7200) );
  INV_X1 U8185 ( .A(n11070), .ZN(n7201) );
  OAI21_X1 U8186 ( .B1(n10400), .B2(n6697), .A(n10397), .ZN(n10462) );
  XNOR2_X1 U8187 ( .A(n13363), .B(n10469), .ZN(n10467) );
  XNOR2_X1 U8188 ( .A(n13364), .B(n8585), .ZN(n10400) );
  AND2_X1 U8189 ( .A1(n8532), .A2(n8531), .ZN(n13619) );
  OR2_X1 U8190 ( .A1(n11967), .A2(n7938), .ZN(n8381) );
  AND2_X1 U8191 ( .A1(n8336), .A2(n8335), .ZN(n13816) );
  OR2_X1 U8192 ( .A1(n11694), .A2(n7938), .ZN(n8336) );
  AND2_X1 U8193 ( .A1(n7749), .A2(n7852), .ZN(n7204) );
  INV_X1 U8194 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7852) );
  NOR2_X1 U8195 ( .A1(n7863), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n7840) );
  INV_X1 U8196 ( .A(n7620), .ZN(n7619) );
  OAI21_X1 U8197 ( .B1(n7624), .B2(n7622), .A(n7621), .ZN(n7620) );
  OR2_X1 U8198 ( .A1(n8073), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U8199 ( .A1(n7096), .A2(n7095), .ZN(n7952) );
  INV_X1 U8200 ( .A(n7939), .ZN(n7096) );
  AOI21_X1 U8201 ( .B1(n7375), .B2(n7377), .A(n6785), .ZN(n7371) );
  INV_X1 U8202 ( .A(n11889), .ZN(n7358) );
  NAND2_X1 U8203 ( .A1(n14108), .A2(n14107), .ZN(n7369) );
  INV_X1 U8204 ( .A(n14151), .ZN(n7385) );
  OR2_X1 U8205 ( .A1(n9683), .A2(n9682), .ZN(n9703) );
  AND2_X1 U8206 ( .A1(n7388), .A2(n7387), .ZN(n10550) );
  INV_X1 U8207 ( .A(n10545), .ZN(n7387) );
  NAND2_X1 U8208 ( .A1(n7369), .A2(n7368), .ZN(n14118) );
  OR2_X1 U8209 ( .A1(n9703), .A2(n10447), .ZN(n9734) );
  OR2_X1 U8210 ( .A1(n9945), .A2(n14068), .ZN(n9961) );
  AOI21_X1 U8211 ( .B1(n7527), .B2(n7521), .A(n7519), .ZN(n10084) );
  NAND2_X1 U8212 ( .A1(n7520), .A2(n7523), .ZN(n7519) );
  AND2_X1 U8213 ( .A1(n7522), .A2(n7525), .ZN(n7521) );
  OAI21_X1 U8214 ( .B1(n6878), .B2(n6877), .A(n6876), .ZN(n7527) );
  AND3_X1 U8215 ( .A1(n9857), .A2(n9856), .A3(n9855), .ZN(n14109) );
  AND4_X1 U8216 ( .A1(n9820), .A2(n9819), .A3(n9818), .A4(n9817), .ZN(n14132)
         );
  NAND2_X1 U8217 ( .A1(n10938), .A2(n10939), .ZN(n11247) );
  OR2_X1 U8218 ( .A1(n11252), .A2(n11251), .ZN(n6925) );
  NAND2_X1 U8219 ( .A1(n15057), .A2(n12020), .ZN(n12022) );
  OR2_X1 U8220 ( .A1(n12022), .A2(n12021), .ZN(n6930) );
  AND2_X1 U8221 ( .A1(n6930), .A2(n6929), .ZN(n14237) );
  NAND2_X1 U8222 ( .A1(n14234), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U8223 ( .A1(n10041), .A2(n10040), .ZN(n14284) );
  OR2_X1 U8224 ( .A1(n14370), .A2(n14361), .ZN(n7287) );
  XNOR2_X1 U8225 ( .A(n14576), .B(n10043), .ZN(n14348) );
  AND2_X1 U8226 ( .A1(n14379), .A2(n14318), .ZN(n7607) );
  NOR2_X1 U8227 ( .A1(n14417), .A2(n14596), .ZN(n14401) );
  NAND2_X1 U8228 ( .A1(n14407), .A2(n14342), .ZN(n7501) );
  NOR2_X1 U8229 ( .A1(n14407), .A2(n14342), .ZN(n7500) );
  NAND2_X1 U8230 ( .A1(n9954), .A2(n9953), .ZN(n14420) );
  NOR2_X1 U8231 ( .A1(n14412), .A2(n14413), .ZN(n14411) );
  NAND2_X1 U8232 ( .A1(n7046), .A2(n9932), .ZN(n14437) );
  NAND2_X1 U8233 ( .A1(n12424), .A2(n10038), .ZN(n7046) );
  OR2_X1 U8234 ( .A1(n6709), .A2(n7478), .ZN(n7477) );
  INV_X1 U8235 ( .A(n7480), .ZN(n7478) );
  NAND2_X1 U8236 ( .A1(n14490), .A2(n14335), .ZN(n14473) );
  NOR2_X1 U8237 ( .A1(n14332), .A2(n7496), .ZN(n7495) );
  INV_X1 U8238 ( .A(n14331), .ZN(n7496) );
  NAND2_X1 U8239 ( .A1(n6887), .A2(n10047), .ZN(n14539) );
  INV_X1 U8240 ( .A(n14537), .ZN(n6887) );
  NAND2_X1 U8241 ( .A1(n6888), .A2(n14326), .ZN(n14553) );
  AND2_X1 U8242 ( .A1(n11834), .A2(n10050), .ZN(n11747) );
  OR2_X1 U8243 ( .A1(n11820), .A2(n11821), .ZN(n11739) );
  NOR2_X1 U8244 ( .A1(n6667), .A2(n15071), .ZN(n7589) );
  OR2_X1 U8245 ( .A1(n10168), .A2(n6690), .ZN(n9697) );
  NAND2_X1 U8246 ( .A1(n11494), .A2(n11495), .ZN(n11539) );
  AND2_X1 U8247 ( .A1(n9880), .A2(n9879), .ZN(n14634) );
  OR2_X1 U8248 ( .A1(n11694), .A2(n6690), .ZN(n9880) );
  OR2_X1 U8249 ( .A1(n11523), .A2(n6690), .ZN(n9826) );
  NAND2_X1 U8250 ( .A1(n9815), .A2(n9814), .ZN(n14650) );
  NAND2_X1 U8251 ( .A1(n10091), .A2(n10090), .ZN(n15189) );
  INV_X1 U8252 ( .A(n15205), .ZN(n15143) );
  NAND2_X1 U8253 ( .A1(n10733), .A2(n11459), .ZN(n15192) );
  XNOR2_X1 U8254 ( .A(n8493), .B(n8489), .ZN(n13884) );
  NAND2_X1 U8255 ( .A1(n6772), .A2(n9561), .ZN(n9559) );
  INV_X1 U8256 ( .A(n7611), .ZN(n7609) );
  NAND2_X1 U8257 ( .A1(n6771), .A2(n9561), .ZN(n10104) );
  NAND2_X1 U8258 ( .A1(n8374), .A2(SI_22_), .ZN(n8399) );
  NAND2_X1 U8259 ( .A1(n7112), .A2(n8377), .ZN(n8400) );
  OR2_X1 U8260 ( .A1(n9567), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n10085) );
  XNOR2_X1 U8261 ( .A(n9563), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10540) );
  NAND2_X1 U8262 ( .A1(n9567), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9563) );
  XNOR2_X1 U8263 ( .A(n8352), .B(n8351), .ZN(n11900) );
  AND2_X1 U8264 ( .A1(n9809), .A2(n7389), .ZN(n9564) );
  AND2_X1 U8265 ( .A1(n7390), .A2(n9811), .ZN(n7389) );
  AND2_X1 U8266 ( .A1(n9822), .A2(n9569), .ZN(n7390) );
  OR2_X1 U8267 ( .A1(n8333), .A2(n8365), .ZN(n8348) );
  NOR2_X1 U8268 ( .A1(n9757), .A2(n9539), .ZN(n9809) );
  NAND2_X1 U8269 ( .A1(n8170), .A2(n8169), .ZN(n8196) );
  INV_X1 U8270 ( .A(n7707), .ZN(n7706) );
  OAI21_X1 U8271 ( .B1(n8089), .B2(n7708), .A(n7832), .ZN(n7707) );
  INV_X1 U8272 ( .A(n14759), .ZN(n7005) );
  INV_X1 U8273 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7069) );
  AND2_X1 U8274 ( .A1(n7291), .A2(n14810), .ZN(n14781) );
  OAI21_X1 U8275 ( .B1(n14812), .B2(n14811), .A(n7292), .ZN(n7291) );
  INV_X1 U8276 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7292) );
  OAI21_X1 U8277 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14724), .A(n14723), .ZN(
        n14785) );
  AOI22_X1 U8278 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14729), .B1(n14787), 
        .B2(n14728), .ZN(n14790) );
  AND3_X1 U8279 ( .A1(n8768), .A2(n8767), .A3(n8766), .ZN(n15496) );
  NAND2_X1 U8280 ( .A1(n9093), .A2(n9092), .ZN(n12933) );
  NAND2_X1 U8281 ( .A1(n10869), .A2(n10868), .ZN(n7419) );
  NAND2_X1 U8282 ( .A1(n10987), .A2(n15448), .ZN(n15445) );
  NAND2_X1 U8283 ( .A1(n9068), .A2(n9067), .ZN(n12960) );
  NAND2_X1 U8284 ( .A1(n12674), .A2(n12512), .ZN(n12601) );
  NAND2_X1 U8285 ( .A1(n8946), .A2(n8945), .ZN(n13171) );
  AND3_X1 U8286 ( .A1(n8717), .A2(n8716), .A3(n8715), .ZN(n11597) );
  NAND2_X1 U8287 ( .A1(n8999), .A2(n8998), .ZN(n13019) );
  OR2_X1 U8288 ( .A1(n11106), .A2(n9014), .ZN(n8999) );
  NAND2_X1 U8289 ( .A1(n12435), .A2(n12434), .ZN(n12507) );
  NAND2_X1 U8290 ( .A1(n7131), .A2(n7129), .ZN(n12655) );
  AOI21_X1 U8291 ( .B1(n7132), .B2(n7134), .A(n7130), .ZN(n7129) );
  AND2_X1 U8292 ( .A1(n7441), .A2(n7133), .ZN(n7132) );
  NAND2_X1 U8293 ( .A1(n12164), .A2(n9148), .ZN(n6845) );
  NAND4_X1 U8294 ( .A1(n8796), .A2(n8795), .A3(n8794), .A4(n8793), .ZN(n15397)
         );
  NAND2_X1 U8295 ( .A1(n7257), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7256) );
  OR2_X1 U8296 ( .A1(n11944), .A2(n11945), .ZN(n7279) );
  INV_X1 U8297 ( .A(n12752), .ZN(n12751) );
  NOR2_X1 U8298 ( .A1(n12710), .A2(n12711), .ZN(n12713) );
  INV_X1 U8299 ( .A(n7219), .ZN(n12709) );
  OR2_X1 U8300 ( .A1(n12761), .A2(n12762), .ZN(n7218) );
  AND2_X1 U8301 ( .A1(n12796), .A2(n13071), .ZN(n7032) );
  XNOR2_X1 U8302 ( .A(n7253), .B(n7252), .ZN(n7471) );
  INV_X1 U8303 ( .A(n12846), .ZN(n7252) );
  NAND2_X1 U8304 ( .A1(n7254), .A2(n12844), .ZN(n7253) );
  NOR2_X1 U8305 ( .A1(n12835), .A2(n12834), .ZN(n12836) );
  XNOR2_X1 U8306 ( .A(n12865), .B(n12903), .ZN(n13117) );
  INV_X1 U8307 ( .A(n12931), .ZN(n7082) );
  NAND2_X1 U8308 ( .A1(n6665), .A2(n15435), .ZN(n7083) );
  NAND2_X1 U8309 ( .A1(n8964), .A2(n8963), .ZN(n13163) );
  NAND2_X1 U8310 ( .A1(n8931), .A2(n8930), .ZN(n13174) );
  NAND2_X1 U8311 ( .A1(n8910), .A2(n8909), .ZN(n13178) );
  AND3_X1 U8312 ( .A1(n8825), .A2(n8824), .A3(n8823), .ZN(n12328) );
  NAND2_X1 U8313 ( .A1(n6973), .A2(n6976), .ZN(n6972) );
  NAND2_X1 U8314 ( .A1(n12915), .A2(n12919), .ZN(n6976) );
  AND2_X1 U8315 ( .A1(n12918), .A2(n15453), .ZN(n6973) );
  NAND2_X1 U8316 ( .A1(n12927), .A2(n12902), .ZN(n12915) );
  NAND2_X1 U8317 ( .A1(n7017), .A2(n6975), .ZN(n6971) );
  INV_X1 U8318 ( .A(n7018), .ZN(n7017) );
  OAI21_X1 U8319 ( .B1(n13121), .B2(n15466), .A(n13119), .ZN(n7018) );
  NOR2_X1 U8320 ( .A1(n13123), .A2(n7016), .ZN(n13191) );
  AND2_X1 U8321 ( .A1(n6665), .A2(n15509), .ZN(n7016) );
  NOR2_X1 U8322 ( .A1(n7789), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n6987) );
  INV_X1 U8323 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U8324 ( .A1(n8655), .A2(n8654), .ZN(n12857) );
  MUX2_X1 U8325 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8653), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8654) );
  NAND2_X1 U8326 ( .A1(n6947), .A2(n6946), .ZN(n6945) );
  XNOR2_X1 U8327 ( .A(n8979), .B(n8978), .ZN(n12850) );
  OAI21_X1 U8328 ( .B1(n8977), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8979) );
  INV_X1 U8329 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U8330 ( .A1(n8516), .A2(n8515), .ZN(n13764) );
  AND2_X1 U8331 ( .A1(n12484), .A2(n9426), .ZN(n6836) );
  NAND2_X1 U8332 ( .A1(n7579), .A2(n7578), .ZN(n7577) );
  OAI22_X1 U8333 ( .A1(n7580), .A2(n7576), .B1(n9489), .B2(n7579), .ZN(n7575)
         );
  XNOR2_X1 U8334 ( .A(n9372), .B(n10740), .ZN(n10661) );
  OR2_X1 U8335 ( .A1(n9385), .A2(n6698), .ZN(n7546) );
  NAND2_X1 U8336 ( .A1(n14900), .A2(n14898), .ZN(n6834) );
  NAND2_X1 U8337 ( .A1(n8429), .A2(n8428), .ZN(n13787) );
  NAND2_X1 U8338 ( .A1(n12424), .A2(n8530), .ZN(n8429) );
  NAND2_X1 U8339 ( .A1(n10112), .A2(n9385), .ZN(n10693) );
  NAND2_X1 U8340 ( .A1(n7613), .A2(n7273), .ZN(n8603) );
  INV_X1 U8341 ( .A(n13573), .ZN(n13537) );
  INV_X1 U8342 ( .A(n13288), .ZN(n13564) );
  AND4_X1 U8343 ( .A1(n7891), .A2(n7890), .A3(n7889), .A4(n7888), .ZN(n13354)
         );
  NAND4_X1 U8344 ( .A1(n7982), .A2(n7981), .A3(n7980), .A4(n7979), .ZN(n13362)
         );
  OR2_X1 U8345 ( .A1(n7914), .A2(n7978), .ZN(n7979) );
  AND2_X1 U8346 ( .A1(n13588), .A2(n13587), .ZN(n13760) );
  OR2_X1 U8347 ( .A1(n11523), .A2(n7938), .ZN(n8294) );
  NAND2_X1 U8348 ( .A1(n8201), .A2(n8200), .ZN(n14921) );
  OAI21_X1 U8349 ( .B1(n10185), .B2(n7938), .A(n7861), .ZN(n11860) );
  OR2_X1 U8350 ( .A1(n10194), .A2(n15365), .ZN(n13737) );
  NAND2_X1 U8351 ( .A1(n15389), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7352) );
  NAND2_X1 U8352 ( .A1(n13548), .A2(n6736), .ZN(n13847) );
  NAND2_X1 U8353 ( .A1(n12443), .A2(n8530), .ZN(n6917) );
  NAND2_X1 U8354 ( .A1(n7209), .A2(n13760), .ZN(n13849) );
  INV_X1 U8355 ( .A(n7210), .ZN(n7209) );
  OAI21_X1 U8356 ( .B1(n13761), .B2(n13842), .A(n13759), .ZN(n7210) );
  INV_X1 U8357 ( .A(n6686), .ZN(n12465) );
  OR2_X1 U8358 ( .A1(n10174), .A2(n6690), .ZN(n9677) );
  NAND2_X1 U8359 ( .A1(n9981), .A2(n9980), .ZN(n14589) );
  NOR2_X1 U8360 ( .A1(n7085), .A2(n6732), .ZN(n7084) );
  NOR2_X1 U8361 ( .A1(n9997), .A2(n10138), .ZN(n7085) );
  NAND2_X1 U8362 ( .A1(n7380), .A2(n11276), .ZN(n14020) );
  AND2_X1 U8363 ( .A1(n14032), .A2(n14030), .ZN(n7111) );
  INV_X1 U8364 ( .A(n14562), .ZN(n14656) );
  INV_X1 U8365 ( .A(n14165), .ZN(n14142) );
  NAND2_X1 U8366 ( .A1(n9979), .A2(n9978), .ZN(n14344) );
  OR2_X1 U8367 ( .A1(n10018), .A2(n10282), .ZN(n9639) );
  NAND2_X1 U8368 ( .A1(n10013), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9623) );
  NOR2_X1 U8369 ( .A1(n14260), .A2(n14259), .ZN(n14261) );
  NAND2_X1 U8370 ( .A1(n14308), .A2(n14307), .ZN(n14631) );
  INV_X1 U8371 ( .A(n7063), .ZN(n14308) );
  OAI22_X1 U8372 ( .A1(n10181), .A2(n10154), .B1(n10122), .B2(n10153), .ZN(
        n7481) );
  XNOR2_X1 U8373 ( .A(n9570), .B(n9569), .ZN(n14511) );
  NAND2_X1 U8374 ( .A1(n15930), .A2(n15931), .ZN(n15929) );
  NAND2_X1 U8375 ( .A1(n14781), .A2(n14782), .ZN(n14817) );
  NAND2_X1 U8376 ( .A1(n14817), .A2(n14818), .ZN(n14814) );
  NAND2_X1 U8377 ( .A1(n6854), .A2(n6853), .ZN(n14816) );
  INV_X1 U8378 ( .A(n14782), .ZN(n6853) );
  INV_X1 U8379 ( .A(n14781), .ZN(n6854) );
  AOI21_X1 U8380 ( .B1(n15918), .B2(n15919), .A(n6859), .ZN(n6858) );
  INV_X1 U8381 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n6859) );
  NOR2_X1 U8382 ( .A1(n15918), .A2(n15919), .ZN(n6860) );
  INV_X1 U8383 ( .A(n10053), .ZN(n10052) );
  AOI21_X1 U8384 ( .B1(n9235), .B2(n9234), .A(n9233), .ZN(n9243) );
  OAI21_X1 U8385 ( .B1(n8068), .B2(n7673), .A(n6777), .ZN(n8110) );
  NAND2_X1 U8386 ( .A1(n7677), .A2(n7675), .ZN(n7673) );
  OAI21_X1 U8387 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(n9628) );
  NOR2_X1 U8388 ( .A1(n7530), .A2(n9643), .ZN(n7529) );
  INV_X1 U8389 ( .A(n9644), .ZN(n7530) );
  INV_X1 U8390 ( .A(n9643), .ZN(n7528) );
  INV_X1 U8391 ( .A(n9678), .ZN(n7508) );
  NAND2_X1 U8392 ( .A1(n6702), .A2(n7507), .ZN(n7506) );
  NAND2_X1 U8393 ( .A1(n9679), .A2(n7507), .ZN(n7059) );
  OR2_X1 U8394 ( .A1(n9680), .A2(n7508), .ZN(n7507) );
  NOR2_X1 U8395 ( .A1(n6710), .A2(n12070), .ZN(n7024) );
  AOI22_X1 U8396 ( .A1(n7635), .A2(n7632), .B1(n7629), .B2(n7637), .ZN(n7626)
         );
  NAND2_X1 U8397 ( .A1(n7636), .A2(n7638), .ZN(n7635) );
  NAND2_X1 U8398 ( .A1(n9712), .A2(n9714), .ZN(n7099) );
  AND2_X1 U8399 ( .A1(n7644), .A2(n7643), .ZN(n7642) );
  INV_X1 U8400 ( .A(n8256), .ZN(n7652) );
  NAND2_X1 U8401 ( .A1(n7653), .A2(n7652), .ZN(n7650) );
  INV_X1 U8402 ( .A(n8281), .ZN(n7648) );
  NOR2_X1 U8403 ( .A1(n7653), .A2(n7652), .ZN(n7651) );
  NAND2_X1 U8404 ( .A1(n9746), .A2(n9748), .ZN(n7541) );
  OR3_X1 U8405 ( .A1(n9308), .A2(n9300), .A3(n7332), .ZN(n9310) );
  NAND2_X1 U8406 ( .A1(n8303), .A2(n7656), .ZN(n7655) );
  INV_X1 U8407 ( .A(n8304), .ZN(n7656) );
  AOI21_X1 U8408 ( .B1(n6869), .B2(n7532), .A(n7098), .ZN(n9808) );
  AND2_X1 U8409 ( .A1(n10047), .A2(n9849), .ZN(n7097) );
  NAND2_X1 U8410 ( .A1(n9873), .A2(n7536), .ZN(n7537) );
  NOR2_X1 U8411 ( .A1(n9873), .A2(n7536), .ZN(n7535) );
  AND2_X1 U8412 ( .A1(n9327), .A2(n12958), .ZN(n7020) );
  NAND2_X1 U8413 ( .A1(n7661), .A2(n6763), .ZN(n7660) );
  NAND2_X1 U8414 ( .A1(n9913), .A2(n9914), .ZN(n9912) );
  NAND2_X1 U8415 ( .A1(n7269), .A2(n7272), .ZN(n7268) );
  INV_X1 U8416 ( .A(n8284), .ZN(n7720) );
  OAI22_X1 U8417 ( .A1(n13865), .A2(n8565), .B1(n13561), .B2(n8545), .ZN(n8414) );
  NAND2_X1 U8418 ( .A1(n8552), .A2(n8551), .ZN(n6913) );
  INV_X1 U8419 ( .A(n9957), .ZN(n7107) );
  NAND2_X1 U8420 ( .A1(n6696), .A2(n7512), .ZN(n7511) );
  OAI21_X1 U8421 ( .B1(n6875), .B2(n6874), .A(n6873), .ZN(n9943) );
  NAND2_X1 U8422 ( .A1(n9929), .A2(n9931), .ZN(n6873) );
  NOR2_X1 U8423 ( .A1(n9931), .A2(n9929), .ZN(n6874) );
  NAND2_X1 U8424 ( .A1(n9918), .A2(n9917), .ZN(n6875) );
  NAND2_X1 U8425 ( .A1(n9571), .A2(n10724), .ZN(n10027) );
  NAND2_X1 U8426 ( .A1(n9339), .A2(n12903), .ZN(n9342) );
  MUX2_X1 U8427 ( .A(n11580), .B(n9205), .S(n9204), .Z(n9338) );
  OAI22_X1 U8428 ( .A1(n13580), .A2(n8545), .B1(n9514), .B2(n6692), .ZN(n8552)
         );
  INV_X1 U8429 ( .A(n10029), .ZN(n7524) );
  INV_X1 U8430 ( .A(n10030), .ZN(n7526) );
  INV_X1 U8431 ( .A(n7590), .ZN(n7227) );
  OR2_X1 U8432 ( .A1(n11496), .A2(n7595), .ZN(n7594) );
  INV_X1 U8433 ( .A(n11477), .ZN(n7595) );
  AOI21_X1 U8434 ( .B1(n8499), .B2(n8470), .A(n7748), .ZN(n7747) );
  INV_X1 U8435 ( .A(n8483), .ZN(n7748) );
  INV_X1 U8436 ( .A(n8470), .ZN(n7745) );
  AOI21_X1 U8437 ( .B1(n8399), .B2(n7693), .A(n6820), .ZN(n7692) );
  NOR2_X1 U8438 ( .A1(n8421), .A2(n8377), .ZN(n7693) );
  AND2_X1 U8439 ( .A1(n8399), .A2(n7694), .ZN(n6911) );
  INV_X1 U8440 ( .A(n8421), .ZN(n7694) );
  NAND2_X1 U8441 ( .A1(n6922), .A2(n7715), .ZN(n8332) );
  AOI21_X1 U8442 ( .B1(n7717), .B2(n7721), .A(n6819), .ZN(n7715) );
  OAI21_X1 U8443 ( .B1(n8236), .B2(n6921), .A(n6786), .ZN(n6922) );
  NAND2_X1 U8444 ( .A1(n8170), .A2(n7742), .ZN(n7741) );
  NOR2_X1 U8445 ( .A1(n8195), .A2(n7743), .ZN(n7742) );
  INV_X1 U8446 ( .A(n8169), .ZN(n7743) );
  INV_X1 U8447 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9533) );
  INV_X1 U8448 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9530) );
  INV_X1 U8449 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7258) );
  NAND2_X1 U8450 ( .A1(n6856), .A2(n14704), .ZN(n14705) );
  NAND2_X1 U8451 ( .A1(n14756), .A2(n14703), .ZN(n6856) );
  INV_X1 U8452 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15887) );
  INV_X1 U8453 ( .A(n12609), .ZN(n7128) );
  INV_X1 U8454 ( .A(n12105), .ZN(n7437) );
  XNOR2_X1 U8455 ( .A(n12159), .B(n12532), .ZN(n12114) );
  INV_X1 U8456 ( .A(n9204), .ZN(n7325) );
  NAND2_X1 U8457 ( .A1(n10782), .A2(n7275), .ZN(n10785) );
  NOR2_X1 U8458 ( .A1(n10783), .A2(n7276), .ZN(n7275) );
  INV_X1 U8459 ( .A(n10781), .ZN(n7276) );
  NAND2_X1 U8460 ( .A1(n11953), .A2(n7251), .ZN(n7249) );
  NAND2_X1 U8461 ( .A1(n12795), .A2(n12794), .ZN(n12825) );
  NAND2_X1 U8462 ( .A1(n12894), .A2(n7770), .ZN(n7769) );
  OR2_X1 U8463 ( .A1(n13171), .A2(n12656), .ZN(n9296) );
  AOI21_X1 U8464 ( .B1(n13091), .B2(n7772), .A(n6978), .ZN(n6977) );
  NAND2_X1 U8465 ( .A1(n6979), .A2(n12877), .ZN(n6978) );
  OR2_X1 U8466 ( .A1(n13178), .A2(n14833), .ZN(n9291) );
  NOR2_X1 U8467 ( .A1(n9278), .A2(n7315), .ZN(n7314) );
  INV_X1 U8468 ( .A(n9274), .ZN(n7315) );
  INV_X1 U8469 ( .A(n8807), .ZN(n7299) );
  INV_X1 U8470 ( .A(n7757), .ZN(n6968) );
  NOR2_X1 U8471 ( .A1(n11595), .A2(n7308), .ZN(n7304) );
  INV_X1 U8472 ( .A(n11600), .ZN(n7308) );
  NAND2_X1 U8473 ( .A1(n15422), .A2(n9225), .ZN(n15407) );
  INV_X1 U8474 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9350) );
  NOR2_X1 U8475 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8636) );
  INV_X1 U8476 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9169) );
  NAND2_X1 U8477 ( .A1(n8926), .A2(n6704), .ZN(n8960) );
  AND2_X1 U8478 ( .A1(n7334), .A2(n7333), .ZN(n7792) );
  NOR2_X1 U8479 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7334) );
  NOR2_X1 U8480 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7333) );
  OR2_X1 U8481 ( .A1(n13252), .A2(n7587), .ZN(n7586) );
  INV_X1 U8482 ( .A(n9484), .ZN(n7587) );
  INV_X1 U8483 ( .A(n9457), .ZN(n7562) );
  NAND2_X1 U8484 ( .A1(n6916), .A2(n8566), .ZN(n8601) );
  NAND2_X1 U8485 ( .A1(n7041), .A2(n13344), .ZN(n6916) );
  INV_X1 U8486 ( .A(n7157), .ZN(n7154) );
  AND2_X1 U8487 ( .A1(n7711), .A2(n13568), .ZN(n7156) );
  OR2_X1 U8488 ( .A1(n7712), .A2(n13570), .ZN(n7710) );
  NAND2_X1 U8489 ( .A1(n7713), .A2(n13572), .ZN(n7712) );
  INV_X1 U8490 ( .A(n13611), .ZN(n7713) );
  INV_X1 U8491 ( .A(n13677), .ZN(n7195) );
  NAND2_X1 U8492 ( .A1(n13659), .A2(n7234), .ZN(n7233) );
  INV_X1 U8493 ( .A(n7235), .ZN(n7234) );
  NAND2_X1 U8494 ( .A1(n13865), .A2(n7236), .ZN(n7235) );
  INV_X1 U8495 ( .A(n13518), .ZN(n7199) );
  NAND2_X1 U8496 ( .A1(n7241), .A2(n13550), .ZN(n7240) );
  INV_X1 U8497 ( .A(n7242), .ZN(n7241) );
  NAND2_X1 U8498 ( .A1(n12383), .A2(n7703), .ZN(n7242) );
  INV_X1 U8499 ( .A(n11758), .ZN(n7733) );
  NAND2_X1 U8500 ( .A1(n7232), .A2(n12066), .ZN(n7231) );
  AND2_X1 U8501 ( .A1(n11501), .A2(n7687), .ZN(n7686) );
  NAND2_X1 U8502 ( .A1(n11087), .A2(n11371), .ZN(n7687) );
  INV_X1 U8503 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8001) );
  NOR2_X1 U8504 ( .A1(n7231), .A2(n7230), .ZN(n11995) );
  INV_X1 U8505 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U8506 ( .A1(n7874), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n7621) );
  NAND2_X1 U8507 ( .A1(n7623), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7622) );
  INV_X1 U8508 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7623) );
  AND2_X1 U8509 ( .A1(n7867), .A2(n7868), .ZN(n7624) );
  NOR2_X1 U8510 ( .A1(n7863), .A2(n7866), .ZN(n7572) );
  AND2_X1 U8511 ( .A1(n11702), .A2(n7376), .ZN(n7375) );
  NAND2_X1 U8512 ( .A1(n11280), .A2(n6991), .ZN(n11281) );
  NAND2_X1 U8513 ( .A1(n14026), .A2(n6666), .ZN(n6991) );
  INV_X1 U8514 ( .A(n10725), .ZN(n10544) );
  INV_X1 U8515 ( .A(n14116), .ZN(n7370) );
  OAI21_X1 U8516 ( .B1(n9972), .B2(n6701), .A(n6779), .ZN(n9984) );
  NOR2_X1 U8517 ( .A1(n10001), .A2(n10002), .ZN(n6877) );
  NAND2_X1 U8518 ( .A1(n10002), .A2(n10001), .ZN(n6876) );
  OR2_X1 U8519 ( .A1(n7524), .A2(n7526), .ZN(n7522) );
  NAND2_X1 U8520 ( .A1(n10031), .A2(n10032), .ZN(n7525) );
  NAND2_X1 U8521 ( .A1(n10034), .A2(n10033), .ZN(n7523) );
  NAND2_X1 U8522 ( .A1(n12017), .A2(n6923), .ZN(n12019) );
  OR2_X1 U8523 ( .A1(n12018), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8524 ( .A1(n14613), .A2(n6906), .ZN(n6905) );
  INV_X1 U8525 ( .A(n6721), .ZN(n7473) );
  INV_X1 U8526 ( .A(n14296), .ZN(n7597) );
  NAND2_X1 U8527 ( .A1(n7089), .A2(n7088), .ZN(n14275) );
  NAND2_X1 U8528 ( .A1(n8529), .A2(n8463), .ZN(n7682) );
  INV_X1 U8529 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10094) );
  INV_X1 U8530 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10086) );
  NAND2_X1 U8531 ( .A1(n7716), .A2(n8288), .ZN(n8329) );
  INV_X1 U8532 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9537) );
  INV_X1 U8533 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U8534 ( .A1(n8236), .A2(n7797), .ZN(n8238) );
  NAND3_X1 U8535 ( .A1(n7262), .A2(n7263), .A3(n7704), .ZN(n8137) );
  AOI21_X1 U8536 ( .B1(n7706), .B2(n7708), .A(n7705), .ZN(n7704) );
  XNOR2_X1 U8537 ( .A(n8133), .B(SI_11_), .ZN(n8136) );
  NAND2_X1 U8538 ( .A1(n7830), .A2(SI_10_), .ZN(n8117) );
  OR2_X1 U8539 ( .A1(n9720), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9742) );
  AND2_X1 U8540 ( .A1(n9673), .A2(n9672), .ZN(n9690) );
  NOR2_X1 U8541 ( .A1(n9655), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U8542 ( .A1(n7261), .A2(SI_5_), .ZN(n7817) );
  OR2_X1 U8543 ( .A1(n9631), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9655) );
  XNOR2_X1 U8544 ( .A(n14705), .B(n15887), .ZN(n14755) );
  NAND2_X1 U8545 ( .A1(n9222), .A2(n15457), .ZN(n10869) );
  NAND2_X1 U8546 ( .A1(n15426), .A2(n10876), .ZN(n15428) );
  AND2_X1 U8547 ( .A1(n12345), .A2(n12343), .ZN(n7452) );
  XNOR2_X1 U8548 ( .A(n12974), .B(n7140), .ZN(n12631) );
  INV_X1 U8549 ( .A(n9055), .ZN(n9054) );
  OR2_X1 U8550 ( .A1(n11322), .A2(n11321), .ZN(n11793) );
  NAND2_X1 U8551 ( .A1(n12576), .A2(n12577), .ZN(n12112) );
  XNOR2_X1 U8552 ( .A(n13019), .B(n7140), .ZN(n12521) );
  OAI21_X1 U8553 ( .B1(n12641), .B2(n7137), .A(n7135), .ZN(n12549) );
  INV_X1 U8554 ( .A(n7138), .ZN(n7137) );
  AOI21_X1 U8555 ( .B1(n7138), .B2(n7136), .A(n6773), .ZN(n7135) );
  NAND2_X1 U8556 ( .A1(n12346), .A2(n7451), .ZN(n7450) );
  INV_X1 U8557 ( .A(n12343), .ZN(n7451) );
  OR2_X1 U8558 ( .A1(n12344), .A2(n12345), .ZN(n7449) );
  NAND2_X1 U8559 ( .A1(n12344), .A2(n7452), .ZN(n7447) );
  INV_X1 U8560 ( .A(n12512), .ZN(n7134) );
  OR2_X1 U8561 ( .A1(n12675), .A2(n7134), .ZN(n7133) );
  INV_X1 U8562 ( .A(n7439), .ZN(n7130) );
  AOI21_X1 U8563 ( .B1(n7441), .B2(n7443), .A(n6762), .ZN(n7439) );
  XNOR2_X1 U8564 ( .A(n13163), .B(n7140), .ZN(n12514) );
  XNOR2_X1 U8565 ( .A(n13178), .B(n7140), .ZN(n12511) );
  AND2_X1 U8566 ( .A1(n9158), .A2(n9143), .ZN(n9162) );
  AND2_X1 U8567 ( .A1(n9363), .A2(n10604), .ZN(n10627) );
  NAND2_X1 U8568 ( .A1(n7034), .A2(n7033), .ZN(n10518) );
  NAND2_X1 U8569 ( .A1(n12840), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7034) );
  NAND2_X1 U8570 ( .A1(n12814), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7033) );
  OAI21_X1 U8571 ( .B1(n10854), .B2(n10853), .A(n10852), .ZN(n12687) );
  XNOR2_X1 U8572 ( .A(n10788), .B(n10894), .ZN(n10886) );
  INV_X1 U8573 ( .A(n7247), .ZN(n10887) );
  OAI21_X1 U8574 ( .B1(n12689), .B2(n10882), .A(n10881), .ZN(n10880) );
  NAND2_X1 U8575 ( .A1(n7462), .A2(n7461), .ZN(n10966) );
  INV_X1 U8576 ( .A(n10756), .ZN(n7461) );
  NOR2_X1 U8577 ( .A1(n10967), .A2(n10951), .ZN(n11004) );
  OAI21_X1 U8578 ( .B1(n10958), .B2(n10957), .A(n10956), .ZN(n11016) );
  AND2_X1 U8579 ( .A1(n7216), .A2(n7215), .ZN(n11024) );
  AND2_X1 U8580 ( .A1(n10948), .A2(n10947), .ZN(n11018) );
  NOR2_X1 U8581 ( .A1(n11432), .A2(n11431), .ZN(n11434) );
  INV_X1 U8582 ( .A(n7246), .ZN(n11430) );
  NOR2_X1 U8583 ( .A1(n11720), .A2(n11719), .ZN(n11722) );
  NOR2_X1 U8584 ( .A1(n11722), .A2(n11721), .ZN(n11960) );
  NAND2_X1 U8585 ( .A1(n12169), .A2(n12168), .ZN(n7219) );
  XNOR2_X1 U8586 ( .A(n12825), .B(n12824), .ZN(n12796) );
  INV_X1 U8587 ( .A(n7223), .ZN(n7221) );
  NAND2_X1 U8588 ( .A1(n12810), .A2(n12824), .ZN(n7223) );
  NOR2_X1 U8589 ( .A1(n9117), .A2(n7328), .ZN(n7327) );
  INV_X1 U8590 ( .A(n9201), .ZN(n7328) );
  OAI21_X1 U8591 ( .B1(n12959), .B2(n6951), .A(n6950), .ZN(n9102) );
  AOI21_X1 U8592 ( .B1(n7316), .B2(n7319), .A(n12929), .ZN(n6950) );
  INV_X1 U8593 ( .A(n7316), .ZN(n6951) );
  INV_X1 U8594 ( .A(n7767), .ZN(n7766) );
  AOI21_X1 U8595 ( .B1(n7767), .B2(n7765), .A(n6775), .ZN(n7764) );
  NAND2_X1 U8596 ( .A1(n7769), .A2(n7767), .ZN(n12952) );
  INV_X1 U8597 ( .A(n12966), .ZN(n9063) );
  OR2_X1 U8598 ( .A1(n9027), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9039) );
  INV_X1 U8599 ( .A(n7779), .ZN(n7778) );
  AOI21_X1 U8600 ( .B1(n7779), .B2(n9006), .A(n7777), .ZN(n7776) );
  NOR2_X1 U8601 ( .A1(n12887), .A2(n7780), .ZN(n7779) );
  NAND2_X1 U8602 ( .A1(n7321), .A2(n9313), .ZN(n12998) );
  NOR2_X1 U8603 ( .A1(n9315), .A2(n7323), .ZN(n7322) );
  INV_X1 U8604 ( .A(n9007), .ZN(n7323) );
  OR2_X1 U8605 ( .A1(n9320), .A2(n9321), .ZN(n12999) );
  OR2_X1 U8606 ( .A1(n9000), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9019) );
  NOR2_X1 U8607 ( .A1(n13048), .A2(n13049), .ZN(n13047) );
  OR2_X1 U8608 ( .A1(n13045), .A2(n7332), .ZN(n13039) );
  NAND2_X1 U8609 ( .A1(n8947), .A2(n15625), .ZN(n8965) );
  INV_X1 U8610 ( .A(n8948), .ZN(n8947) );
  NAND2_X1 U8611 ( .A1(n8912), .A2(n8911), .ZN(n8932) );
  OR2_X1 U8612 ( .A1(n8932), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U8613 ( .A1(n6941), .A2(n9283), .ZN(n13098) );
  NAND2_X1 U8614 ( .A1(n6937), .A2(n6936), .ZN(n6941) );
  AND2_X1 U8615 ( .A1(n6938), .A2(n9179), .ZN(n6936) );
  AND2_X1 U8616 ( .A1(n6983), .A2(n6982), .ZN(n6981) );
  NOR2_X1 U8617 ( .A1(n14856), .A2(n14850), .ZN(n6984) );
  NAND2_X1 U8618 ( .A1(n12869), .A2(n7785), .ZN(n6985) );
  NOR2_X1 U8619 ( .A1(n8856), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8874) );
  OR2_X1 U8620 ( .A1(n8826), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8856) );
  AND2_X1 U8621 ( .A1(n8855), .A2(n8854), .ZN(n14863) );
  AND2_X1 U8622 ( .A1(n9263), .A2(n9267), .ZN(n12334) );
  NAND2_X1 U8623 ( .A1(n12325), .A2(n12334), .ZN(n12324) );
  NAND2_X1 U8624 ( .A1(n8791), .A2(n8790), .ZN(n8809) );
  NAND2_X1 U8625 ( .A1(n12154), .A2(n12075), .ZN(n12327) );
  AOI21_X1 U8626 ( .B1(n6956), .B2(n6958), .A(n6953), .ZN(n6952) );
  INV_X1 U8627 ( .A(n9249), .ZN(n6953) );
  INV_X1 U8628 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11027) );
  AND2_X1 U8629 ( .A1(n9253), .A2(n9254), .ZN(n15396) );
  NAND2_X1 U8630 ( .A1(n7752), .A2(n12072), .ZN(n15395) );
  NOR2_X1 U8631 ( .A1(n8751), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8769) );
  AND4_X1 U8632 ( .A1(n8775), .A2(n8774), .A3(n8773), .A4(n8772), .ZN(n12497)
         );
  OAI21_X1 U8633 ( .B1(n11596), .B2(n7760), .A(n7757), .ZN(n11778) );
  OR2_X1 U8634 ( .A1(n8735), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U8635 ( .A1(n7763), .A2(n11599), .ZN(n11601) );
  NOR2_X1 U8636 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8719) );
  AND2_X1 U8637 ( .A1(n15412), .A2(n15410), .ZN(n11573) );
  INV_X1 U8638 ( .A(n10991), .ZN(n15437) );
  NAND2_X1 U8639 ( .A1(n10869), .A2(n10867), .ZN(n15423) );
  OR2_X1 U8640 ( .A1(n9154), .A2(n10759), .ZN(n8684) );
  AND2_X1 U8641 ( .A1(n12859), .A2(n12906), .ZN(n13184) );
  NAND2_X1 U8642 ( .A1(n12927), .A2(n7774), .ZN(n12918) );
  NAND2_X1 U8643 ( .A1(n6962), .A2(n7330), .ZN(n13021) );
  NAND2_X1 U8644 ( .A1(n14860), .A2(n9274), .ZN(n14849) );
  OR2_X1 U8645 ( .A1(n10920), .A2(n10807), .ZN(n10918) );
  AND2_X1 U8646 ( .A1(n8656), .A2(n8644), .ZN(n7791) );
  OAI21_X1 U8647 ( .B1(n9119), .B2(n9118), .A(n9120), .ZN(n9131) );
  AND2_X1 U8648 ( .A1(n8782), .A2(n6942), .ZN(n6946) );
  NOR2_X1 U8649 ( .A1(n7459), .A2(n6943), .ZN(n6942) );
  NAND2_X1 U8650 ( .A1(n8642), .A2(n8783), .ZN(n6943) );
  NAND2_X1 U8651 ( .A1(n7460), .A2(n8656), .ZN(n7459) );
  INV_X1 U8652 ( .A(n6948), .ZN(n6947) );
  NAND2_X1 U8653 ( .A1(n9065), .A2(n9051), .ZN(n9064) );
  OR2_X1 U8654 ( .A1(n9175), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U8655 ( .A1(n9009), .A2(n9008), .ZN(n9012) );
  NAND2_X1 U8656 ( .A1(n8868), .A2(n7028), .ZN(n9173) );
  INV_X1 U8657 ( .A(n9167), .ZN(n7028) );
  NAND2_X1 U8658 ( .A1(n9170), .A2(n9169), .ZN(n9175) );
  INV_X1 U8659 ( .A(n9173), .ZN(n9170) );
  AND2_X1 U8660 ( .A1(n6704), .A2(n8961), .ZN(n7141) );
  AOI21_X1 U8661 ( .B1(n8957), .B2(n7395), .A(n7394), .ZN(n7393) );
  INV_X1 U8662 ( .A(n8957), .ZN(n7396) );
  INV_X1 U8663 ( .A(n8971), .ZN(n7394) );
  INV_X1 U8664 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8925) );
  AND2_X1 U8665 ( .A1(n8868), .A2(n8907), .ZN(n8926) );
  AND2_X1 U8666 ( .A1(n8863), .A2(n8846), .ZN(n8847) );
  NAND2_X1 U8667 ( .A1(n8848), .A2(n8847), .ZN(n8864) );
  NAND2_X1 U8668 ( .A1(n6847), .A2(n7403), .ZN(n8840) );
  AOI21_X1 U8669 ( .B1(n7405), .B2(n7407), .A(n7404), .ZN(n7403) );
  NAND2_X1 U8670 ( .A1(n8801), .A2(n7405), .ZN(n6847) );
  INV_X1 U8671 ( .A(n8836), .ZN(n7404) );
  AND2_X1 U8672 ( .A1(n8844), .A2(n8838), .ZN(n8839) );
  INV_X1 U8673 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8783) );
  AOI21_X1 U8674 ( .B1(n7412), .B2(n7410), .A(n7409), .ZN(n7408) );
  INV_X1 U8675 ( .A(n7412), .ZN(n7411) );
  INV_X1 U8676 ( .A(n8757), .ZN(n7410) );
  AND2_X1 U8677 ( .A1(n8797), .A2(n8778), .ZN(n8779) );
  NAND2_X1 U8678 ( .A1(n7391), .A2(n8729), .ZN(n8743) );
  INV_X1 U8679 ( .A(n8726), .ZN(n8727) );
  NAND2_X1 U8680 ( .A1(n6850), .A2(n8677), .ZN(n8689) );
  NAND2_X1 U8681 ( .A1(n8676), .A2(n6851), .ZN(n6850) );
  NAND2_X1 U8682 ( .A1(n8690), .A2(n6849), .ZN(n8688) );
  NAND2_X1 U8683 ( .A1(n10129), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6849) );
  OR2_X1 U8684 ( .A1(n8534), .A2(n8484), .ZN(n8535) );
  NAND2_X1 U8685 ( .A1(n13315), .A2(n13314), .ZN(n6844) );
  NOR2_X1 U8686 ( .A1(n7586), .A2(n7578), .ZN(n7574) );
  NAND2_X1 U8687 ( .A1(n7583), .A2(n7582), .ZN(n7581) );
  OR2_X1 U8688 ( .A1(n13252), .A2(n7585), .ZN(n7584) );
  INV_X1 U8689 ( .A(n9485), .ZN(n7582) );
  AND2_X1 U8690 ( .A1(n7586), .A2(n7578), .ZN(n7576) );
  INV_X1 U8691 ( .A(n9489), .ZN(n7578) );
  INV_X1 U8692 ( .A(n11856), .ZN(n6838) );
  AOI21_X1 U8693 ( .B1(n11857), .B2(n9415), .A(n6781), .ZN(n7557) );
  INV_X1 U8694 ( .A(n9415), .ZN(n7558) );
  NOR2_X1 U8695 ( .A1(n13295), .A2(n7544), .ZN(n7543) );
  INV_X1 U8696 ( .A(n9468), .ZN(n7544) );
  AND2_X1 U8697 ( .A1(n8223), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8268) );
  AND2_X1 U8698 ( .A1(n6841), .A2(n11404), .ZN(n7569) );
  INV_X1 U8699 ( .A(n9401), .ZN(n6842) );
  INV_X1 U8700 ( .A(n9396), .ZN(n7570) );
  NAND2_X1 U8701 ( .A1(n9456), .A2(n9455), .ZN(n13302) );
  INV_X1 U8702 ( .A(n12239), .ZN(n7064) );
  INV_X1 U8703 ( .A(n12238), .ZN(n6837) );
  OR2_X1 U8704 ( .A1(n8355), .A2(n13281), .ZN(n8383) );
  NOR2_X1 U8705 ( .A1(n8002), .A2(n8001), .ZN(n8037) );
  AOI21_X1 U8706 ( .B1(n10652), .B2(n6698), .A(n6778), .ZN(n7547) );
  NAND2_X1 U8707 ( .A1(n8457), .A2(n8458), .ZN(n7614) );
  OR2_X1 U8708 ( .A1(n8559), .A2(n8558), .ZN(n7061) );
  AND2_X1 U8709 ( .A1(n8344), .A2(n8343), .ZN(n13556) );
  AND3_X1 U8710 ( .A1(n8301), .A2(n8300), .A3(n8299), .ZN(n13553) );
  AND3_X1 U8711 ( .A1(n8277), .A2(n8276), .A3(n8275), .ZN(n13549) );
  OR2_X1 U8712 ( .A1(n15268), .A2(n15267), .ZN(n15265) );
  AOI21_X1 U8713 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n10564), .A(n10563), .ZN(
        n10567) );
  AOI21_X1 U8714 ( .B1(n10831), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10827), .ZN(
        n10830) );
  AOI21_X1 U8715 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n13456), .A(n13447), .ZN(
        n15280) );
  NOR2_X1 U8716 ( .A1(n13451), .A2(n15289), .ZN(n13453) );
  OR2_X1 U8717 ( .A1(n13453), .A2(n13452), .ZN(n13483) );
  AND2_X1 U8718 ( .A1(n15301), .A2(n15300), .ZN(n15302) );
  INV_X1 U8719 ( .A(n13577), .ZN(n12448) );
  AND2_X1 U8720 ( .A1(n8512), .A2(n8511), .ZN(n13545) );
  OAI211_X1 U8721 ( .C1(n13566), .C2(n7155), .A(n7709), .B(n7153), .ZN(n13591)
         );
  AND2_X1 U8722 ( .A1(n7710), .A2(n6809), .ZN(n7709) );
  INV_X1 U8723 ( .A(n7156), .ZN(n7155) );
  NAND2_X1 U8724 ( .A1(n7156), .A2(n7154), .ZN(n7153) );
  AOI21_X1 U8725 ( .B1(n13601), .B2(n13611), .A(n6726), .ZN(n13586) );
  INV_X1 U8726 ( .A(n7712), .ZN(n7711) );
  NOR2_X1 U8727 ( .A1(n13694), .A2(n7233), .ZN(n13653) );
  NOR2_X1 U8728 ( .A1(n13694), .A2(n7235), .ZN(n13670) );
  NOR2_X1 U8729 ( .A1(n13694), .A2(n13802), .ZN(n13680) );
  AOI21_X1 U8730 ( .B1(n7729), .B2(n13689), .A(n6740), .ZN(n7728) );
  NAND2_X1 U8731 ( .A1(n13519), .A2(n13518), .ZN(n13706) );
  NOR2_X1 U8732 ( .A1(n7238), .A2(n14927), .ZN(n13735) );
  NAND2_X1 U8733 ( .A1(n13744), .A2(n7239), .ZN(n7238) );
  INV_X1 U8734 ( .A(n7240), .ZN(n7239) );
  NOR2_X1 U8735 ( .A1(n14927), .A2(n7240), .ZN(n13734) );
  NOR2_X1 U8736 ( .A1(n14927), .A2(n7242), .ZN(n12388) );
  NOR2_X1 U8737 ( .A1(n14927), .A2(n12364), .ZN(n12371) );
  AND2_X1 U8738 ( .A1(n7346), .A2(n7187), .ZN(n7186) );
  OR2_X1 U8739 ( .A1(n14921), .A2(n14926), .ZN(n14927) );
  NAND2_X1 U8740 ( .A1(n11995), .A2(n12195), .ZN(n14926) );
  NOR2_X1 U8741 ( .A1(n8152), .A2(n8151), .ZN(n8179) );
  INV_X1 U8742 ( .A(n7169), .ZN(n11928) );
  AOI21_X1 U8743 ( .B1(n11681), .B2(n6738), .A(n7170), .ZN(n7169) );
  OAI21_X1 U8744 ( .B1(n11683), .B2(n7340), .A(n11761), .ZN(n7170) );
  INV_X1 U8745 ( .A(n7231), .ZN(n11937) );
  INV_X1 U8746 ( .A(n7232), .ZN(n11766) );
  INV_X1 U8747 ( .A(n11756), .ZN(n11683) );
  NAND2_X1 U8748 ( .A1(n11681), .A2(n11680), .ZN(n11682) );
  NAND2_X1 U8749 ( .A1(n11682), .A2(n11683), .ZN(n11763) );
  NOR2_X1 U8750 ( .A1(n8100), .A2(n8099), .ZN(n8098) );
  NAND2_X1 U8751 ( .A1(n7684), .A2(n7683), .ZN(n11676) );
  AOI21_X1 U8752 ( .B1(n7686), .B2(n7688), .A(n6769), .ZN(n7683) );
  NAND2_X1 U8753 ( .A1(n11370), .A2(n7686), .ZN(n7684) );
  INV_X1 U8754 ( .A(n11371), .ZN(n7688) );
  OR2_X1 U8755 ( .A1(n8058), .A2(n8057), .ZN(n8079) );
  NOR2_X1 U8756 ( .A1(n7338), .A2(n6783), .ZN(n7336) );
  NAND2_X1 U8757 ( .A1(n7685), .A2(n11371), .ZN(n11502) );
  NAND2_X1 U8758 ( .A1(n11370), .A2(n11369), .ZN(n7685) );
  AND4_X1 U8759 ( .A1(n8085), .A2(n8084), .A3(n8083), .A4(n8082), .ZN(n11503)
         );
  OR2_X1 U8760 ( .A1(n9519), .A2(n10320), .ZN(n13326) );
  OAI21_X1 U8761 ( .B1(n10898), .B2(n7724), .A(n7723), .ZN(n11109) );
  INV_X1 U8762 ( .A(n7725), .ZN(n7724) );
  NOR2_X1 U8763 ( .A1(n11082), .A2(n7726), .ZN(n7725) );
  NAND2_X1 U8764 ( .A1(n10905), .A2(n11240), .ZN(n11110) );
  NAND2_X1 U8765 ( .A1(n7349), .A2(n7993), .ZN(n7350) );
  OR2_X1 U8766 ( .A1(n13593), .A2(n13592), .ZN(n13759) );
  AND2_X1 U8767 ( .A1(n11695), .A2(n11968), .ZN(n7008) );
  NAND2_X1 U8768 ( .A1(n11074), .A2(n11073), .ZN(n11113) );
  NAND2_X1 U8769 ( .A1(n11071), .A2(n11070), .ZN(n11074) );
  INV_X1 U8770 ( .A(n7956), .ZN(n8146) );
  OR2_X1 U8771 ( .A1(n8146), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8013) );
  INV_X1 U8772 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9665) );
  OR2_X1 U8773 ( .A1(n9666), .A2(n9665), .ZN(n9683) );
  NAND2_X1 U8774 ( .A1(n11274), .A2(n11275), .ZN(n11276) );
  INV_X4 U8775 ( .A(n13942), .ZN(n14042) );
  OR2_X1 U8776 ( .A1(n9837), .A2(n9836), .ZN(n9839) );
  NAND2_X1 U8777 ( .A1(n11886), .A2(n7356), .ZN(n11915) );
  NAND2_X1 U8778 ( .A1(n10703), .A2(n10550), .ZN(n10705) );
  NAND2_X1 U8779 ( .A1(n9765), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U8780 ( .A1(n7364), .A2(n7370), .ZN(n7363) );
  INV_X1 U8781 ( .A(n7366), .ZN(n7364) );
  AOI21_X1 U8782 ( .B1(n7368), .B2(n7367), .A(n13953), .ZN(n7366) );
  INV_X1 U8783 ( .A(n14107), .ZN(n7367) );
  NAND2_X1 U8784 ( .A1(n7368), .A2(n7370), .ZN(n7365) );
  NAND2_X1 U8785 ( .A1(n12221), .A2(n12220), .ZN(n12272) );
  OR2_X1 U8786 ( .A1(n11408), .A2(n11407), .ZN(n7376) );
  AND2_X1 U8787 ( .A1(n11408), .A2(n11407), .ZN(n7377) );
  INV_X1 U8788 ( .A(n9961), .ZN(n9960) );
  NAND2_X1 U8789 ( .A1(n13915), .A2(n13916), .ZN(n14152) );
  NAND2_X1 U8790 ( .A1(n14152), .A2(n14151), .ZN(n7383) );
  INV_X1 U8791 ( .A(n10082), .ZN(n6866) );
  AND4_X1 U8792 ( .A1(n9844), .A2(n9843), .A3(n9842), .A4(n9841), .ZN(n14298)
         );
  NOR2_X1 U8793 ( .A1(n15035), .A2(n6813), .ZN(n10378) );
  NAND2_X1 U8794 ( .A1(n10378), .A2(n10377), .ZN(n10376) );
  NAND2_X1 U8795 ( .A1(n10376), .A2(n6926), .ZN(n10283) );
  OR2_X1 U8796 ( .A1(n10293), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6926) );
  NOR2_X1 U8797 ( .A1(n10283), .A2(n10284), .ZN(n10357) );
  NOR2_X1 U8798 ( .A1(n10413), .A2(n6928), .ZN(n10417) );
  AND2_X1 U8799 ( .A1(n10414), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6928) );
  NAND2_X1 U8800 ( .A1(n10417), .A2(n10416), .ZN(n10436) );
  NOR2_X1 U8801 ( .A1(n10592), .A2(n6931), .ZN(n10596) );
  AND2_X1 U8802 ( .A1(n10593), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U8803 ( .A1(n10596), .A2(n10595), .ZN(n10936) );
  NAND2_X1 U8804 ( .A1(n10936), .A2(n6989), .ZN(n10938) );
  OR2_X1 U8805 ( .A1(n10937), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6989) );
  AND2_X1 U8806 ( .A1(n6925), .A2(n6924), .ZN(n11340) );
  NAND2_X1 U8807 ( .A1(n11339), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U8808 ( .A1(n11340), .A2(n11341), .ZN(n12017) );
  NOR2_X1 U8809 ( .A1(n14248), .A2(n6832), .ZN(n14258) );
  NOR2_X1 U8810 ( .A1(n14250), .A2(n14251), .ZN(n14260) );
  AOI21_X1 U8811 ( .B1(n7607), .B2(n14317), .A(n6768), .ZN(n7606) );
  NAND2_X1 U8812 ( .A1(n14319), .A2(n10045), .ZN(n14375) );
  OR2_X1 U8813 ( .A1(n14583), .A2(n14346), .ZN(n10045) );
  NAND2_X1 U8814 ( .A1(n14433), .A2(n14418), .ZN(n14417) );
  NOR2_X1 U8815 ( .A1(n14428), .A2(n7602), .ZN(n7601) );
  INV_X1 U8816 ( .A(n14314), .ZN(n7602) );
  NAND2_X1 U8817 ( .A1(n14427), .A2(n14340), .ZN(n14412) );
  INV_X1 U8818 ( .A(n14424), .ZN(n14413) );
  INV_X1 U8819 ( .A(n14437), .ZN(n14435) );
  INV_X1 U8820 ( .A(n14432), .ZN(n14428) );
  AOI21_X1 U8821 ( .B1(n6694), .B2(n14500), .A(n6767), .ZN(n7604) );
  NOR2_X1 U8822 ( .A1(n14481), .A2(n14461), .ZN(n14460) );
  NAND2_X1 U8823 ( .A1(n14546), .A2(n14329), .ZN(n6885) );
  NAND2_X1 U8824 ( .A1(n7286), .A2(n14529), .ZN(n14527) );
  NAND2_X1 U8825 ( .A1(n9795), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9837) );
  INV_X1 U8826 ( .A(n9797), .ZN(n9795) );
  OR2_X1 U8827 ( .A1(n9784), .A2(n9783), .ZN(n9797) );
  NAND2_X1 U8828 ( .A1(n6889), .A2(n14324), .ZN(n14952) );
  INV_X1 U8829 ( .A(n7089), .ZN(n12255) );
  NAND2_X1 U8830 ( .A1(n9736), .A2(n9735), .ZN(n9750) );
  AND3_X1 U8831 ( .A1(n7087), .A2(n15081), .A3(n6903), .ZN(n11844) );
  NOR2_X1 U8832 ( .A1(n11978), .A2(n11879), .ZN(n6903) );
  AND2_X1 U8833 ( .A1(n11844), .A2(n14984), .ZN(n12096) );
  INV_X1 U8834 ( .A(n11834), .ZN(n7499) );
  NAND2_X1 U8835 ( .A1(n15081), .A2(n15201), .ZN(n11827) );
  NAND2_X1 U8836 ( .A1(n7285), .A2(n7284), .ZN(n15082) );
  AOI21_X1 U8837 ( .B1(n7486), .B2(n11496), .A(n6735), .ZN(n7485) );
  NAND2_X1 U8838 ( .A1(n6902), .A2(n6900), .ZN(n11550) );
  NOR2_X1 U8839 ( .A1(n14026), .A2(n6901), .ZN(n6900) );
  NOR2_X1 U8840 ( .A1(n15100), .A2(n14026), .ZN(n15101) );
  OR2_X1 U8841 ( .A1(n10018), .A2(n9572), .ZN(n9574) );
  NAND2_X1 U8842 ( .A1(n10013), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U8843 ( .A1(n6897), .A2(n7287), .ZN(n6899) );
  XNOR2_X1 U8844 ( .A(n8496), .B(n8495), .ZN(n13876) );
  AND2_X1 U8845 ( .A1(n9543), .A2(n7610), .ZN(n7608) );
  NOR2_X1 U8846 ( .A1(n7611), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n7610) );
  XNOR2_X1 U8847 ( .A(n6918), .B(n8483), .ZN(n12443) );
  OAI21_X1 U8848 ( .B1(n8500), .B2(n8499), .A(n8470), .ZN(n6918) );
  AND2_X1 U8849 ( .A1(n8529), .A2(n8528), .ZN(n13887) );
  NAND2_X1 U8850 ( .A1(n6934), .A2(n7735), .ZN(n8527) );
  NAND2_X1 U8851 ( .A1(n8448), .A2(n7740), .ZN(n8461) );
  NOR2_X1 U8852 ( .A1(n10093), .A2(n10092), .ZN(n10098) );
  AND2_X1 U8853 ( .A1(n8449), .A2(n8427), .ZN(n12424) );
  NAND2_X1 U8854 ( .A1(n9561), .A2(n9822), .ZN(n10093) );
  INV_X1 U8855 ( .A(n9561), .ZN(n9821) );
  AND2_X1 U8856 ( .A1(n9690), .A2(n9689), .ZN(n9694) );
  INV_X1 U8857 ( .A(n7260), .ZN(n8009) );
  OAI21_X1 U8858 ( .B1(SI_5_), .B2(n7261), .A(n7817), .ZN(n7260) );
  NOR2_X1 U8859 ( .A1(n9590), .A2(n9603), .ZN(n10289) );
  INV_X1 U8860 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15861) );
  OAI21_X1 U8861 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n15864), .A(n14700), .ZN(
        n14758) );
  XNOR2_X1 U8862 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14757) );
  XNOR2_X1 U8863 ( .A(n14755), .B(n15052), .ZN(n14766) );
  NAND2_X1 U8864 ( .A1(n14711), .A2(n14710), .ZN(n14773) );
  NOR2_X1 U8865 ( .A1(n14803), .A2(n14776), .ZN(n14778) );
  OAI21_X1 U8866 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15822), .A(n14718), .ZN(
        n14752) );
  NOR2_X1 U8867 ( .A1(n14749), .A2(n14722), .ZN(n14747) );
  AND2_X1 U8868 ( .A1(n7288), .A2(n14998), .ZN(n14789) );
  INV_X1 U8869 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7289) );
  OAI21_X1 U8870 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14731), .A(n14730), .ZN(
        n14744) );
  NAND2_X1 U8871 ( .A1(n12106), .A2(n12105), .ZN(n12493) );
  AOI21_X1 U8872 ( .B1(n12921), .B2(n9116), .A(n9115), .ZN(n12930) );
  INV_X1 U8873 ( .A(n12986), .ZN(n12630) );
  NAND2_X1 U8874 ( .A1(n9038), .A2(n9037), .ZN(n13139) );
  OR2_X1 U8875 ( .A1(n12570), .A2(n7429), .ZN(n7426) );
  INV_X1 U8876 ( .A(n7424), .ZN(n7423) );
  NAND2_X1 U8877 ( .A1(n11570), .A2(n6828), .ZN(n10871) );
  NAND2_X1 U8878 ( .A1(n12639), .A2(n12523), .ZN(n12585) );
  INV_X1 U8879 ( .A(n7125), .ZN(n12431) );
  OAI22_X1 U8880 ( .A1(n12344), .A2(n7126), .B1(n7452), .B2(n7448), .ZN(n7125)
         );
  AND2_X1 U8881 ( .A1(n7448), .A2(n12345), .ZN(n7126) );
  AND4_X1 U8882 ( .A1(n8970), .A2(n8969), .A3(n8968), .A4(n8967), .ZN(n13061)
         );
  NAND2_X1 U8883 ( .A1(n7440), .A2(n7444), .ZN(n12620) );
  NAND2_X1 U8884 ( .A1(n12601), .A2(n7445), .ZN(n7440) );
  OR2_X1 U8885 ( .A1(n12135), .A2(n12134), .ZN(n12137) );
  NAND2_X1 U8886 ( .A1(n12641), .A2(n12640), .ZN(n12639) );
  NAND2_X1 U8887 ( .A1(n9026), .A2(n9025), .ZN(n12889) );
  AND4_X1 U8888 ( .A1(n8814), .A2(n8813), .A3(n8812), .A4(n8811), .ZN(n12353)
         );
  AND2_X1 U8889 ( .A1(n8843), .A2(n8842), .ZN(n12355) );
  XNOR2_X1 U8890 ( .A(n12532), .B(n10876), .ZN(n10992) );
  INV_X1 U8891 ( .A(n12677), .ZN(n12657) );
  NAND2_X1 U8892 ( .A1(n12607), .A2(n11797), .ZN(n11799) );
  AND2_X1 U8893 ( .A1(n10642), .A2(n10983), .ZN(n12670) );
  INV_X1 U8894 ( .A(n7453), .ZN(n12676) );
  OAI21_X1 U8895 ( .B1(n12541), .B2(n12508), .A(n12510), .ZN(n7453) );
  NAND2_X1 U8896 ( .A1(n12676), .A2(n12675), .ZN(n12674) );
  XNOR2_X1 U8897 ( .A(n6996), .B(n12850), .ZN(n9199) );
  NAND2_X1 U8898 ( .A1(n6997), .A2(n6743), .ZN(n6996) );
  NAND2_X1 U8899 ( .A1(n7045), .A2(n15455), .ZN(n7081) );
  AND2_X1 U8900 ( .A1(n9158), .A2(n9128), .ZN(n12916) );
  NAND2_X1 U8901 ( .A1(n9087), .A2(n9086), .ZN(n12898) );
  INV_X1 U8902 ( .A(n12870), .ZN(n14844) );
  INV_X1 U8903 ( .A(n12353), .ZN(n12342) );
  INV_X1 U8904 ( .A(n12497), .ZN(n12110) );
  INV_X1 U8905 ( .A(n12107), .ZN(n15399) );
  INV_X1 U8906 ( .A(n12613), .ZN(n12104) );
  INV_X1 U8907 ( .A(n15408), .ZN(n11598) );
  INV_X1 U8908 ( .A(n15426), .ZN(n10999) );
  NAND2_X1 U8909 ( .A1(n9138), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7309) );
  AND2_X1 U8910 ( .A1(n7040), .A2(n7039), .ZN(n10520) );
  NAND2_X1 U8911 ( .A1(n10518), .A2(n10524), .ZN(n7039) );
  NAND2_X1 U8912 ( .A1(n10520), .A2(n11056), .ZN(n10673) );
  AOI21_X1 U8913 ( .B1(n10673), .B2(n7040), .A(n10672), .ZN(n10854) );
  AOI21_X1 U8914 ( .B1(n12687), .B2(n12686), .A(n12685), .ZN(n12689) );
  INV_X1 U8915 ( .A(n7462), .ZN(n10757) );
  AOI21_X1 U8916 ( .B1(n11016), .B2(n11015), .A(n11014), .ZN(n11162) );
  INV_X1 U8917 ( .A(n7468), .ZN(n11008) );
  INV_X1 U8918 ( .A(n7211), .ZN(n11439) );
  OAI21_X1 U8919 ( .B1(n11162), .B2(n11161), .A(n11160), .ZN(n11428) );
  INV_X1 U8920 ( .A(n7281), .ZN(n11442) );
  AOI21_X1 U8921 ( .B1(n11428), .B2(n11427), .A(n11426), .ZN(n11720) );
  INV_X1 U8922 ( .A(n7465), .ZN(n11952) );
  XNOR2_X1 U8923 ( .A(n12760), .B(n12775), .ZN(n12738) );
  INV_X1 U8924 ( .A(n7254), .ZN(n12845) );
  NAND2_X1 U8925 ( .A1(n12817), .A2(n12818), .ZN(n7036) );
  NAND2_X1 U8926 ( .A1(n6949), .A2(n7316), .ZN(n12926) );
  NAND2_X1 U8927 ( .A1(n12959), .A2(n7318), .ZN(n6949) );
  NAND2_X1 U8928 ( .A1(n12957), .A2(n9076), .ZN(n12939) );
  NAND2_X1 U8929 ( .A1(n7781), .A2(n12886), .ZN(n13005) );
  NAND2_X1 U8930 ( .A1(n13016), .A2(n13020), .ZN(n7781) );
  NAND2_X1 U8931 ( .A1(n13023), .A2(n9007), .ZN(n13009) );
  NAND2_X1 U8932 ( .A1(n8982), .A2(n8981), .ZN(n13157) );
  NAND2_X1 U8933 ( .A1(n6821), .A2(n7772), .ZN(n13080) );
  NAND2_X1 U8934 ( .A1(n6937), .A2(n6938), .ZN(n14837) );
  NAND2_X1 U8935 ( .A1(n12869), .A2(n12868), .ZN(n14855) );
  INV_X1 U8936 ( .A(n15460), .ZN(n14864) );
  NAND2_X1 U8937 ( .A1(n7302), .A2(n8808), .ZN(n12080) );
  NAND2_X1 U8938 ( .A1(n12150), .A2(n8807), .ZN(n7302) );
  NAND2_X1 U8939 ( .A1(n6955), .A2(n9244), .ZN(n11612) );
  NAND2_X1 U8940 ( .A1(n11773), .A2(n11772), .ZN(n6955) );
  NAND2_X1 U8941 ( .A1(n11568), .A2(n9212), .ZN(n11594) );
  NAND3_X1 U8942 ( .A1(n7454), .A2(n8661), .A3(n7455), .ZN(n10987) );
  NAND2_X1 U8943 ( .A1(n10639), .A2(n6815), .ZN(n7455) );
  NAND2_X1 U8944 ( .A1(n8666), .A2(SI_0_), .ZN(n7454) );
  INV_X1 U8945 ( .A(n13104), .ZN(n13085) );
  INV_X1 U8946 ( .A(n15458), .ZN(n15442) );
  NAND2_X1 U8947 ( .A1(n9150), .A2(n9149), .ZN(n13111) );
  INV_X1 U8948 ( .A(n13111), .ZN(n13189) );
  OAI211_X1 U8949 ( .C1(n13117), .C2(n15466), .A(n6986), .B(n6756), .ZN(n13190) );
  NAND2_X1 U8950 ( .A1(n12910), .A2(n15495), .ZN(n7050) );
  OR2_X1 U8951 ( .A1(n13173), .A2(n13172), .ZN(n13231) );
  OR3_X1 U8952 ( .A1(n13182), .A2(n13181), .A3(n13180), .ZN(n13233) );
  INV_X1 U8953 ( .A(n10987), .ZN(n10927) );
  AND2_X1 U8954 ( .A1(n10606), .A2(n10605), .ZN(n13234) );
  AND2_X1 U8955 ( .A1(n10609), .A2(n10608), .ZN(n13236) );
  NAND2_X1 U8956 ( .A1(n9147), .A2(n9133), .ZN(n9135) );
  OR2_X1 U8957 ( .A1(n6994), .A2(n8645), .ZN(n8647) );
  NOR2_X1 U8958 ( .A1(n6994), .A2(n6993), .ZN(n6992) );
  OR2_X1 U8959 ( .A1(n8648), .A2(n7790), .ZN(n6995) );
  NOR2_X1 U8960 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6993) );
  XNOR2_X1 U8961 ( .A(n9089), .B(n9081), .ZN(n12164) );
  XNOR2_X1 U8962 ( .A(n9200), .B(P3_IR_REG_22__SCAN_IN), .ZN(n13115) );
  NAND2_X1 U8963 ( .A1(n9349), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9200) );
  INV_X1 U8964 ( .A(n10860), .ZN(n11565) );
  NAND2_X1 U8965 ( .A1(n8995), .A2(n9008), .ZN(n8996) );
  NAND2_X1 U8966 ( .A1(n8958), .A2(n8957), .ZN(n8972) );
  NAND2_X1 U8967 ( .A1(n8955), .A2(n8954), .ZN(n8958) );
  OAI21_X1 U8968 ( .B1(n8905), .B2(n7402), .A(n7400), .ZN(n8939) );
  NAND2_X1 U8969 ( .A1(n8920), .A2(n8919), .ZN(n8923) );
  NAND2_X1 U8970 ( .A1(n8883), .A2(n8865), .ZN(n8866) );
  INV_X1 U8971 ( .A(n8868), .ZN(n9168) );
  OAI21_X1 U8972 ( .B1(n8801), .B2(n7407), .A(n7405), .ZN(n8837) );
  NAND2_X1 U8973 ( .A1(n8816), .A2(n8815), .ZN(n8819) );
  INV_X1 U8974 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U8975 ( .A1(n7414), .A2(n7412), .ZN(n8777) );
  NAND2_X1 U8976 ( .A1(n7414), .A2(n8759), .ZN(n8762) );
  NAND2_X2 U8977 ( .A1(n8714), .A2(n8713), .ZN(n10787) );
  INV_X1 U8978 ( .A(n8678), .ZN(n7102) );
  NAND2_X1 U8979 ( .A1(n7568), .A2(n11119), .ZN(n11391) );
  NAND2_X1 U8980 ( .A1(n7108), .A2(n9396), .ZN(n7568) );
  NAND2_X1 U8981 ( .A1(n13331), .A2(n9484), .ZN(n13253) );
  XNOR2_X1 U8982 ( .A(n9486), .B(n9485), .ZN(n13252) );
  NAND2_X1 U8983 ( .A1(n13324), .A2(n9445), .ZN(n13273) );
  INV_X1 U8984 ( .A(n11504), .ZN(n15372) );
  NAND2_X1 U8985 ( .A1(n13302), .A2(n9457), .ZN(n13280) );
  NAND2_X1 U8986 ( .A1(n7556), .A2(n7554), .ZN(n11874) );
  AOI21_X1 U8987 ( .B1(n7557), .B2(n7558), .A(n7555), .ZN(n7554) );
  NAND2_X1 U8988 ( .A1(n6838), .A2(n7557), .ZN(n7556) );
  INV_X1 U8989 ( .A(n11868), .ZN(n7555) );
  NAND2_X1 U8990 ( .A1(n7567), .A2(n7564), .ZN(n7563) );
  NAND2_X1 U8991 ( .A1(n7545), .A2(n9468), .ZN(n13296) );
  OAI21_X1 U8992 ( .B1(n7108), .B2(n7571), .A(n7569), .ZN(n11400) );
  NAND2_X1 U8993 ( .A1(n7049), .A2(n13271), .ZN(n13304) );
  INV_X1 U8994 ( .A(n7551), .ZN(n7550) );
  NAND2_X1 U8995 ( .A1(n11809), .A2(n9415), .ZN(n11866) );
  NAND2_X1 U8996 ( .A1(n7553), .A2(n9442), .ZN(n13324) );
  INV_X1 U8997 ( .A(n13323), .ZN(n7553) );
  CLKBUF_X1 U8998 ( .A(n11120), .Z(n7108) );
  XNOR2_X1 U8999 ( .A(n7567), .B(n9432), .ZN(n12291) );
  INV_X1 U9000 ( .A(n13545), .ZN(n13538) );
  OR2_X1 U9001 ( .A1(n7914), .A2(n10476), .ZN(n7963) );
  OR2_X1 U9002 ( .A1(n7930), .A2(n7961), .ZN(n7962) );
  NAND4_X1 U9003 ( .A1(n7934), .A2(n7933), .A3(n7932), .A4(n7931), .ZN(n13363)
         );
  OR2_X1 U9004 ( .A1(n7914), .A2(n7928), .ZN(n7934) );
  OR2_X1 U9005 ( .A1(n7930), .A2(n7893), .ZN(n7896) );
  OR2_X1 U9006 ( .A1(n7914), .A2(n10264), .ZN(n7895) );
  NAND2_X1 U9007 ( .A1(n7960), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7918) );
  OR2_X1 U9008 ( .A1(n7930), .A2(n12469), .ZN(n7915) );
  OR2_X1 U9009 ( .A1(n8155), .A2(n12473), .ZN(n7916) );
  AND2_X1 U9010 ( .A1(n8075), .A2(n8093), .ZN(n13438) );
  INV_X1 U9011 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13497) );
  XNOR2_X1 U9012 ( .A(n13487), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13489) );
  INV_X1 U9013 ( .A(n13764), .ZN(n13609) );
  NAND2_X1 U9014 ( .A1(n7714), .A2(n13572), .ZN(n13612) );
  NAND2_X1 U9015 ( .A1(n7714), .A2(n7711), .ZN(n13766) );
  NAND2_X1 U9016 ( .A1(n13663), .A2(n7177), .ZN(n7178) );
  NAND2_X1 U9017 ( .A1(n13566), .A2(n13565), .ZN(n13634) );
  NAND2_X1 U9018 ( .A1(n7182), .A2(n7177), .ZN(n13649) );
  NAND2_X1 U9019 ( .A1(n7731), .A2(n13558), .ZN(n13676) );
  NAND2_X1 U9020 ( .A1(n13690), .A2(n13692), .ZN(n7731) );
  OAI21_X1 U9021 ( .B1(n13519), .B2(n13522), .A(n7196), .ZN(n13675) );
  NAND2_X1 U9022 ( .A1(n8354), .A2(n8353), .ZN(n13699) );
  INV_X1 U9023 ( .A(n13816), .ZN(n13711) );
  NAND2_X1 U9024 ( .A1(n7162), .A2(n6700), .ZN(n13704) );
  OR2_X1 U9025 ( .A1(n13727), .A2(n6695), .ZN(n7162) );
  AND2_X1 U9026 ( .A1(n8310), .A2(n8309), .ZN(n13725) );
  NAND2_X1 U9027 ( .A1(n7342), .A2(n13512), .ZN(n13746) );
  NAND2_X1 U9028 ( .A1(n7695), .A2(n7699), .ZN(n12386) );
  NAND2_X1 U9029 ( .A1(n12358), .A2(n7700), .ZN(n7695) );
  NAND2_X1 U9030 ( .A1(n7701), .A2(n7700), .ZN(n12384) );
  NAND2_X1 U9031 ( .A1(n7701), .A2(n7702), .ZN(n12360) );
  NAND2_X1 U9032 ( .A1(n12197), .A2(n12196), .ZN(n14913) );
  NAND2_X1 U9033 ( .A1(n7192), .A2(n7190), .ZN(n12197) );
  NAND2_X1 U9034 ( .A1(n7145), .A2(n6703), .ZN(n14924) );
  NAND2_X1 U9035 ( .A1(n7149), .A2(n11990), .ZN(n12191) );
  NAND2_X1 U9036 ( .A1(n7151), .A2(n7150), .ZN(n7149) );
  NAND2_X1 U9037 ( .A1(n7192), .A2(n11993), .ZN(n12194) );
  NAND2_X1 U9038 ( .A1(n7734), .A2(n11758), .ZN(n11925) );
  NAND2_X1 U9039 ( .A1(n11757), .A2(n11756), .ZN(n7734) );
  NAND2_X1 U9040 ( .A1(n7335), .A2(n7337), .ZN(n11374) );
  INV_X1 U9041 ( .A(n7338), .ZN(n7337) );
  NOR2_X1 U9042 ( .A1(n14919), .A2(n11090), .ZN(n14932) );
  NAND2_X1 U9043 ( .A1(n7727), .A2(n10900), .ZN(n11083) );
  NAND2_X1 U9044 ( .A1(n10898), .A2(n10897), .ZN(n7727) );
  INV_X1 U9045 ( .A(n13741), .ZN(n14919) );
  INV_X1 U9046 ( .A(n13743), .ZN(n14920) );
  INV_X1 U9047 ( .A(n13713), .ZN(n14931) );
  INV_X1 U9048 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7207) );
  NAND2_X1 U9049 ( .A1(n8097), .A2(n8096), .ZN(n11677) );
  INV_X1 U9050 ( .A(n13619), .ZN(n13854) );
  NAND2_X1 U9051 ( .A1(n8036), .A2(n8035), .ZN(n11211) );
  OR2_X1 U9052 ( .A1(n10250), .A2(n10249), .ZN(n15386) );
  AND2_X1 U9053 ( .A1(n7204), .A2(n7203), .ZN(n7202) );
  AND2_X1 U9054 ( .A1(n7850), .A2(n7882), .ZN(n7203) );
  INV_X1 U9055 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10356) );
  INV_X1 U9056 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10186) );
  INV_X1 U9057 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10170) );
  INV_X1 U9058 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10169) );
  INV_X1 U9059 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10175) );
  INV_X1 U9060 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10161) );
  INV_X1 U9061 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10158) );
  INV_X1 U9062 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10164) );
  NOR2_X2 U9063 ( .A1(n7957), .A2(n7956), .ZN(n13386) );
  INV_X1 U9064 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10167) );
  AOI21_X1 U9065 ( .B1(n11914), .B2(n7357), .A(n6711), .ZN(n7354) );
  INV_X1 U9066 ( .A(n11914), .ZN(n7355) );
  NAND2_X1 U9067 ( .A1(n11886), .A2(n11885), .ZN(n11888) );
  AND2_X1 U9068 ( .A1(n7369), .A2(n6737), .ZN(n14055) );
  AND2_X1 U9069 ( .A1(n7384), .A2(n7382), .ZN(n7381) );
  OR2_X1 U9070 ( .A1(n14073), .A2(n7385), .ZN(n7384) );
  OR2_X1 U9071 ( .A1(n14073), .A2(n13916), .ZN(n7382) );
  AND2_X1 U9072 ( .A1(n7383), .A2(n7386), .ZN(n14074) );
  XNOR2_X1 U9073 ( .A(n11350), .B(n11348), .ZN(n11288) );
  NAND2_X1 U9074 ( .A1(n11915), .A2(n11914), .ZN(n11973) );
  NAND2_X1 U9075 ( .A1(n13934), .A2(n7110), .ZN(n7109) );
  INV_X1 U9076 ( .A(n13939), .ZN(n7110) );
  NAND2_X1 U9077 ( .A1(n7362), .A2(n7363), .ZN(n14120) );
  OR2_X1 U9078 ( .A1(n14108), .A2(n7365), .ZN(n7362) );
  NAND2_X1 U9079 ( .A1(n7374), .A2(n7373), .ZN(n11703) );
  INV_X1 U9080 ( .A(n7377), .ZN(n7373) );
  NAND2_X1 U9081 ( .A1(n11409), .A2(n7376), .ZN(n7374) );
  NAND2_X1 U9082 ( .A1(n10551), .A2(n10543), .ZN(n14165) );
  INV_X1 U9083 ( .A(n7383), .ZN(n14154) );
  AND2_X1 U9084 ( .A1(n14062), .A2(n15192), .ZN(n14163) );
  AND2_X1 U9085 ( .A1(n10179), .A2(n14197), .ZN(n14521) );
  NAND2_X1 U9086 ( .A1(n10078), .A2(n6866), .ZN(n6865) );
  AND4_X1 U9087 ( .A1(n9803), .A2(n9802), .A3(n9801), .A4(n9800), .ZN(n14294)
         );
  AND4_X1 U9088 ( .A1(n9789), .A2(n9788), .A3(n9787), .A4(n9786), .ZN(n14155)
         );
  INV_X1 U9089 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10247) );
  OR2_X1 U9090 ( .A1(n10018), .A2(n15019), .ZN(n9552) );
  OAI21_X1 U9091 ( .B1(n10280), .B2(n14208), .A(n14200), .ZN(n14212) );
  AOI21_X1 U9092 ( .B1(n10358), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10357), .ZN(
        n10361) );
  NAND2_X1 U9093 ( .A1(n10436), .A2(n6927), .ZN(n10438) );
  NAND2_X1 U9094 ( .A1(n10441), .A2(n10415), .ZN(n6927) );
  NAND2_X1 U9095 ( .A1(n10438), .A2(n10439), .ZN(n10481) );
  INV_X1 U9096 ( .A(n6925), .ZN(n11338) );
  INV_X1 U9097 ( .A(n6930), .ZN(n14233) );
  NOR2_X1 U9098 ( .A1(n14276), .A2(n14349), .ZN(n14277) );
  AOI22_X1 U9099 ( .A1(n13884), .A2(n10038), .B1(n10039), .B2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n14573) );
  OAI22_X1 U9100 ( .A1(n14365), .A2(n14347), .B1(n14358), .B2(n14583), .ZN(
        n6884) );
  OR3_X1 U9101 ( .A1(n14370), .A2(n14369), .A3(n15205), .ZN(n14586) );
  NAND2_X1 U9102 ( .A1(n14396), .A2(n14318), .ZN(n14390) );
  INV_X1 U9103 ( .A(n7502), .ZN(n14395) );
  NAND2_X1 U9104 ( .A1(n7476), .A2(n7477), .ZN(n14443) );
  NAND2_X1 U9105 ( .A1(n14473), .A2(n6721), .ZN(n7476) );
  AND2_X1 U9106 ( .A1(n7479), .A2(n6739), .ZN(n14457) );
  NAND2_X1 U9107 ( .A1(n14473), .A2(n14477), .ZN(n7479) );
  INV_X1 U9108 ( .A(n14634), .ZN(n14499) );
  NAND2_X1 U9109 ( .A1(n7495), .A2(n7497), .ZN(n14506) );
  NAND2_X1 U9110 ( .A1(n14519), .A2(n14520), .ZN(n7497) );
  NAND2_X1 U9111 ( .A1(n7599), .A2(n14301), .ZN(n14518) );
  NAND2_X1 U9112 ( .A1(n14960), .A2(n14296), .ZN(n7598) );
  AND2_X1 U9113 ( .A1(n9848), .A2(n9847), .ZN(n14562) );
  NAND2_X1 U9114 ( .A1(n9793), .A2(n9792), .ZN(n14963) );
  NAND2_X1 U9115 ( .A1(n9775), .A2(n9774), .ZN(n14976) );
  NAND2_X1 U9116 ( .A1(n9760), .A2(n9759), .ZN(n14819) );
  NAND2_X1 U9117 ( .A1(n11739), .A2(n11738), .ZN(n11835) );
  NAND2_X1 U9118 ( .A1(n7589), .A2(n15072), .ZN(n7226) );
  NAND2_X1 U9119 ( .A1(n15072), .A2(n11640), .ZN(n7592) );
  NAND2_X1 U9120 ( .A1(n7488), .A2(n11497), .ZN(n11545) );
  NAND2_X1 U9121 ( .A1(n11539), .A2(n11538), .ZN(n7488) );
  NAND2_X1 U9122 ( .A1(n7593), .A2(n11477), .ZN(n11543) );
  NAND2_X1 U9123 ( .A1(n11533), .A2(n11496), .ZN(n7593) );
  INV_X1 U9124 ( .A(n15098), .ZN(n14958) );
  OR2_X1 U9125 ( .A1(n15108), .A2(n11459), .ZN(n15098) );
  NAND2_X1 U9126 ( .A1(n14353), .A2(n15094), .ZN(n14532) );
  XNOR2_X1 U9127 ( .A(n11486), .B(n11669), .ZN(n15144) );
  INV_X1 U9128 ( .A(n14564), .ZN(n14967) );
  INV_X1 U9129 ( .A(n15233), .ZN(n15231) );
  NAND2_X1 U9130 ( .A1(n14568), .A2(n7121), .ZN(n14660) );
  INV_X1 U9131 ( .A(n7122), .ZN(n7121) );
  OAI21_X1 U9132 ( .B1(n14569), .B2(n15213), .A(n14571), .ZN(n7122) );
  OR2_X1 U9133 ( .A1(n14629), .A2(n14628), .ZN(n14670) );
  OR2_X1 U9134 ( .A1(n14636), .A2(n14635), .ZN(n14671) );
  NAND2_X1 U9135 ( .A1(n10104), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U9136 ( .A1(n8399), .A2(n8400), .ZN(n8422) );
  NAND2_X1 U9137 ( .A1(n10085), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9568) );
  INV_X1 U9138 ( .A(n10540), .ZN(n11905) );
  NAND2_X1 U9139 ( .A1(n9565), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U9140 ( .A1(n8348), .A2(n8334), .ZN(n11694) );
  NAND2_X1 U9141 ( .A1(n8306), .A2(n8291), .ZN(n11523) );
  INV_X1 U9142 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10235) );
  INV_X1 U9143 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10184) );
  OAI21_X1 U9144 ( .B1(n8090), .B2(n7708), .A(n7706), .ZN(n8118) );
  NAND2_X1 U9145 ( .A1(n8092), .A2(n7004), .ZN(n7833) );
  NOR2_X1 U9146 ( .A1(n7832), .A2(n7708), .ZN(n7004) );
  INV_X1 U9147 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10171) );
  INV_X1 U9148 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10152) );
  INV_X1 U9149 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10150) );
  INV_X1 U9150 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10141) );
  INV_X1 U9151 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10130) );
  INV_X1 U9152 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10131) );
  INV_X1 U9153 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10138) );
  OAI22_X1 U9154 ( .A1(n9603), .A2(n6932), .B1(P1_IR_REG_3__SCAN_IN), .B2(
        P1_IR_REG_31__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U9155 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6932) );
  NOR2_X1 U9156 ( .A1(n9580), .A2(n9579), .ZN(n14188) );
  INV_X1 U9157 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7804) );
  NOR2_X1 U9158 ( .A1(n14763), .A2(n15936), .ZN(n14800) );
  AOI21_X1 U9159 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14765), .A(n15932), .ZN(
        n15924) );
  XNOR2_X1 U9160 ( .A(n14766), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15923) );
  XNOR2_X1 U9161 ( .A(n14769), .B(n7294), .ZN(n15927) );
  NAND2_X1 U9162 ( .A1(n15927), .A2(n15926), .ZN(n15925) );
  XNOR2_X1 U9163 ( .A(n14775), .B(n14774), .ZN(n14804) );
  NOR2_X1 U9164 ( .A1(n14805), .A2(n14804), .ZN(n14803) );
  XNOR2_X1 U9165 ( .A(n14778), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15930) );
  OAI21_X1 U9166 ( .B1(n14780), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n14806), .ZN(
        n14812) );
  NAND2_X1 U9167 ( .A1(n14812), .A2(n14811), .ZN(n14810) );
  NAND2_X1 U9168 ( .A1(n14814), .A2(n14816), .ZN(n14995) );
  NOR2_X1 U9169 ( .A1(n14995), .A2(n14996), .ZN(n14994) );
  NOR2_X1 U9170 ( .A1(n14789), .A2(n14788), .ZN(n15003) );
  OAI21_X1 U9171 ( .B1(n14792), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n15007), .ZN(
        n15013) );
  NAND2_X1 U9172 ( .A1(n15013), .A2(n15012), .ZN(n15011) );
  NAND2_X1 U9173 ( .A1(n6855), .A2(n15011), .ZN(n15017) );
  OAI21_X1 U9174 ( .B1(n15013), .B2(n15012), .A(n7293), .ZN(n6855) );
  NOR2_X1 U9175 ( .A1(n15017), .A2(n15016), .ZN(n15015) );
  INV_X1 U9176 ( .A(n7279), .ZN(n11949) );
  INV_X1 U9177 ( .A(n12737), .ZN(n12736) );
  INV_X1 U9178 ( .A(n7218), .ZN(n12764) );
  OAI21_X1 U9179 ( .B1(n12808), .B2(n12855), .A(n7030), .ZN(P3_U3199) );
  NOR2_X1 U9180 ( .A1(n12806), .A2(n7031), .ZN(n7030) );
  OR2_X1 U9181 ( .A1(n12805), .A2(n6824), .ZN(n7031) );
  NAND2_X1 U9182 ( .A1(n7471), .A2(n12702), .ZN(n6990) );
  AND2_X1 U9183 ( .A1(n6972), .A2(n6975), .ZN(n13120) );
  NAND2_X1 U9184 ( .A1(n6963), .A2(n6823), .ZN(P3_U3487) );
  OAI21_X1 U9185 ( .B1(n6971), .B2(n6964), .A(n15532), .ZN(n6963) );
  INV_X1 U9186 ( .A(n6972), .ZN(n6964) );
  OAI211_X1 U9187 ( .C1(n6972), .C2(n15517), .A(n6970), .B(n6974), .ZN(
        P3_U3455) );
  NAND2_X1 U9188 ( .A1(n15517), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U9189 ( .A1(n6971), .A2(n15519), .ZN(n6970) );
  OAI21_X1 U9190 ( .B1(n13191), .B2(n15517), .A(n7052), .ZN(P3_U3454) );
  INV_X1 U9191 ( .A(n7053), .ZN(n7052) );
  OAI22_X1 U9192 ( .A1(n13193), .A2(n13229), .B1(n15519), .B2(n13192), .ZN(
        n7053) );
  NAND2_X1 U9193 ( .A1(n9513), .A2(n6814), .ZN(n9527) );
  OAI211_X1 U9194 ( .C1(n10112), .C2(n6698), .A(n10652), .B(n7546), .ZN(n10657) );
  OAI21_X1 U9195 ( .B1(n8603), .B2(n8571), .A(n8607), .ZN(n8632) );
  AND2_X1 U9196 ( .A1(n8603), .A2(n7796), .ZN(n8633) );
  INV_X1 U9197 ( .A(n7351), .ZN(n7074) );
  OAI21_X1 U9198 ( .B1(n13580), .B2(n7353), .A(n7352), .ZN(n7351) );
  NAND2_X1 U9199 ( .A1(n7208), .A2(n7205), .ZN(P2_U3527) );
  NAND2_X1 U9200 ( .A1(n13849), .A2(n15391), .ZN(n7208) );
  NOR2_X1 U9201 ( .A1(n15391), .A2(n7207), .ZN(n7206) );
  AOI21_X1 U9202 ( .B1(n13848), .B2(n13873), .A(n7244), .ZN(n7243) );
  NOR2_X1 U9203 ( .A1(n15387), .A2(n8487), .ZN(n7244) );
  NAND2_X1 U9204 ( .A1(n7168), .A2(n7166), .ZN(P2_U3495) );
  AOI21_X1 U9205 ( .B1(n13850), .B2(n13873), .A(n7167), .ZN(n7166) );
  NAND2_X1 U9206 ( .A1(n13849), .A2(n15387), .ZN(n7168) );
  NOR2_X1 U9207 ( .A1(n15387), .A2(n8509), .ZN(n7167) );
  MUX2_X1 U9208 ( .A(n14272), .B(n14271), .S(n14511), .Z(n14274) );
  NAND2_X1 U9209 ( .A1(n7120), .A2(n7119), .ZN(P1_U3559) );
  OR2_X1 U9210 ( .A1(n15233), .A2(n10016), .ZN(n7119) );
  NAND2_X1 U9211 ( .A1(n14660), .A2(n15233), .ZN(n7120) );
  INV_X1 U9212 ( .A(n14816), .ZN(n14815) );
  XNOR2_X1 U9213 ( .A(n7072), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9214 ( .A1(n7295), .A2(n7073), .ZN(n7072) );
  INV_X1 U9215 ( .A(n6860), .ZN(n7295) );
  NOR2_X1 U9216 ( .A1(n6860), .A2(n6858), .ZN(n6857) );
  AND2_X1 U9217 ( .A1(n7605), .A2(n14310), .ZN(n6694) );
  AND2_X1 U9218 ( .A1(n13725), .A2(n13555), .ZN(n6695) );
  NAND2_X1 U9219 ( .A1(n7350), .A2(n6759), .ZN(n8585) );
  INV_X1 U9220 ( .A(n11737), .ZN(n11821) );
  AND2_X1 U9221 ( .A1(n9944), .A2(n7513), .ZN(n6696) );
  INV_X1 U9222 ( .A(n15444), .ZN(n10876) );
  AND2_X1 U9223 ( .A1(n8582), .A2(n10428), .ZN(n6697) );
  NAND2_X1 U9224 ( .A1(n7029), .A2(n8497), .ZN(n13498) );
  INV_X1 U9225 ( .A(n12251), .ZN(n14322) );
  AND2_X1 U9226 ( .A1(n10650), .A2(n9387), .ZN(n6698) );
  INV_X1 U9227 ( .A(n11637), .ZN(n7284) );
  AND2_X1 U9228 ( .A1(n8345), .A2(n7670), .ZN(n6699) );
  OR2_X1 U9229 ( .A1(n13725), .A2(n13555), .ZN(n6700) );
  NAND2_X1 U9230 ( .A1(n6917), .A2(n6830), .ZN(n13848) );
  INV_X1 U9231 ( .A(n13848), .ZN(n13580) );
  AND2_X1 U9232 ( .A1(n9973), .A2(n7518), .ZN(n6701) );
  AND2_X1 U9233 ( .A1(n9680), .A2(n7508), .ZN(n6702) );
  NAND2_X1 U9234 ( .A1(n8222), .A2(n8221), .ZN(n12364) );
  INV_X1 U9235 ( .A(n12364), .ZN(n7703) );
  AND2_X1 U9236 ( .A1(n7146), .A2(n7152), .ZN(n6703) );
  AND2_X1 U9237 ( .A1(n8925), .A2(n7142), .ZN(n6704) );
  AND2_X1 U9238 ( .A1(n8212), .A2(n8210), .ZN(n6705) );
  AND2_X1 U9239 ( .A1(n7363), .A2(n13963), .ZN(n6706) );
  AND2_X1 U9240 ( .A1(n6700), .A2(n6746), .ZN(n6707) );
  NAND2_X1 U9241 ( .A1(n9970), .A2(n9969), .ZN(n14596) );
  AND2_X1 U9242 ( .A1(n11304), .A2(n9403), .ZN(n6708) );
  AND2_X1 U9243 ( .A1(n14338), .A2(n6739), .ZN(n6709) );
  AND3_X1 U9244 ( .A1(n12104), .A2(n9248), .A3(n11580), .ZN(n6710) );
  AND2_X1 U9245 ( .A1(n11972), .A2(n11971), .ZN(n6711) );
  AND2_X1 U9246 ( .A1(n14444), .A2(n14314), .ZN(n6712) );
  OR2_X1 U9247 ( .A1(n8560), .A2(n6761), .ZN(n6713) );
  OR2_X1 U9248 ( .A1(n7437), .A2(n7128), .ZN(n6714) );
  NAND2_X1 U9249 ( .A1(n8347), .A2(n7669), .ZN(n7668) );
  INV_X1 U9250 ( .A(n7668), .ZN(n7666) );
  INV_X1 U9251 ( .A(n12195), .ZN(n12242) );
  AND2_X1 U9252 ( .A1(n8178), .A2(n8177), .ZN(n12195) );
  INV_X1 U9253 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8656) );
  INV_X1 U9254 ( .A(n9194), .ZN(n12929) );
  XNOR2_X1 U9255 ( .A(n12933), .B(n12901), .ZN(n9194) );
  NAND2_X1 U9256 ( .A1(n9122), .A2(n9121), .ZN(n12910) );
  INV_X1 U9257 ( .A(n9712), .ZN(n7539) );
  OR2_X1 U9258 ( .A1(n7001), .A2(n7000), .ZN(n6715) );
  AND2_X1 U9259 ( .A1(n7214), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6716) );
  AND2_X1 U9260 ( .A1(n9433), .A2(n7565), .ZN(n6717) );
  OR2_X1 U9261 ( .A1(n6984), .A2(n7786), .ZN(n6718) );
  AND2_X1 U9262 ( .A1(n14329), .A2(n9861), .ZN(n10047) );
  INV_X1 U9263 ( .A(n12182), .ZN(n7251) );
  AND2_X1 U9264 ( .A1(n7257), .A2(n6833), .ZN(n6719) );
  NAND2_X1 U9265 ( .A1(n8782), .A2(n8783), .ZN(n8785) );
  XOR2_X1 U9266 ( .A(n14284), .B(n10074), .Z(n6720) );
  AND2_X1 U9267 ( .A1(n8403), .A2(n8402), .ZN(n13865) );
  INV_X1 U9268 ( .A(n13865), .ZN(n7237) );
  NAND2_X1 U9269 ( .A1(n14539), .A2(n14329), .ZN(n14519) );
  NAND2_X1 U9270 ( .A1(n10639), .A2(n10123), .ZN(n9014) );
  NAND4_X1 U9271 ( .A1(n7965), .A2(n7964), .A3(n7963), .A4(n7962), .ZN(n8584)
         );
  NAND2_X1 U9272 ( .A1(n13248), .A2(n13243), .ZN(n7001) );
  NAND2_X1 U9273 ( .A1(n6947), .A2(n6944), .ZN(n9354) );
  NAND2_X1 U9274 ( .A1(n13885), .A2(n7884), .ZN(n7930) );
  INV_X1 U9275 ( .A(n11108), .ZN(n7339) );
  OR2_X1 U9276 ( .A1(n10518), .A2(n10524), .ZN(n7040) );
  INV_X1 U9277 ( .A(n8458), .ZN(n7615) );
  NAND2_X1 U9278 ( .A1(n8798), .A2(n8797), .ZN(n8801) );
  NAND4_X1 U9279 ( .A1(n7918), .A2(n7917), .A3(n7916), .A4(n7915), .ZN(n8582)
         );
  INV_X1 U9280 ( .A(n8087), .ZN(n7678) );
  AND2_X1 U9281 ( .A1(n7480), .A2(n14477), .ZN(n6721) );
  XNOR2_X1 U9282 ( .A(n12355), .B(n7140), .ZN(n12345) );
  OR2_X1 U9283 ( .A1(n8785), .A2(n7755), .ZN(n6722) );
  AND2_X1 U9284 ( .A1(n13040), .A2(n9303), .ZN(n13049) );
  NAND2_X1 U9285 ( .A1(n6687), .A2(n7481), .ZN(n6723) );
  AND4_X1 U9286 ( .A1(n8671), .A2(n8673), .A3(n8674), .A4(n8672), .ZN(n15451)
         );
  AND2_X1 U9287 ( .A1(n7675), .A2(n7674), .ZN(n6724) );
  INV_X1 U9288 ( .A(n7863), .ZN(n7864) );
  AND2_X1 U9289 ( .A1(n7438), .A2(n11797), .ZN(n6725) );
  INV_X1 U9290 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14676) );
  NOR2_X1 U9291 ( .A1(n13609), .A2(n13537), .ZN(n6726) );
  OR2_X1 U9292 ( .A1(n11438), .A2(n11437), .ZN(n6727) );
  OR2_X1 U9293 ( .A1(n10894), .A2(n10754), .ZN(n6728) );
  INV_X1 U9294 ( .A(n8210), .ZN(n7645) );
  NAND2_X1 U9295 ( .A1(n14646), .A2(n14330), .ZN(n6729) );
  NAND2_X1 U9296 ( .A1(n13744), .A2(n13513), .ZN(n6730) );
  MUX2_X1 U9297 ( .A(n14437), .B(n14169), .S(n10075), .Z(n9944) );
  INV_X1 U9298 ( .A(n14442), .ZN(n7475) );
  NAND2_X1 U9299 ( .A1(n14435), .A2(n14315), .ZN(n6731) );
  AND2_X1 U9300 ( .A1(n10177), .A2(n14218), .ZN(n6732) );
  OR2_X1 U9301 ( .A1(n7313), .A2(n6940), .ZN(n6733) );
  OR2_X1 U9302 ( .A1(n11924), .A2(n7733), .ZN(n6734) );
  INV_X1 U9303 ( .A(n11595), .ZN(n7759) );
  INV_X1 U9304 ( .A(n9212), .ZN(n7307) );
  NAND2_X1 U9305 ( .A1(n9782), .A2(n9781), .ZN(n14292) );
  INV_X1 U9306 ( .A(n14292), .ZN(n7088) );
  INV_X1 U9307 ( .A(n10894), .ZN(n7463) );
  INV_X1 U9308 ( .A(n13647), .ZN(n7174) );
  AND2_X1 U9309 ( .A1(n14178), .A2(n11552), .ZN(n6735) );
  INV_X1 U9310 ( .A(n9882), .ZN(n7536) );
  XNOR2_X1 U9311 ( .A(n13019), .B(n13031), .ZN(n13020) );
  NAND2_X1 U9312 ( .A1(n6995), .A2(n6992), .ZN(n13248) );
  AND3_X1 U9313 ( .A1(n13758), .A2(n13757), .A3(n13547), .ZN(n6736) );
  NOR2_X1 U9314 ( .A1(n6948), .A2(n8785), .ZN(n9357) );
  NOR2_X1 U9315 ( .A1(n14182), .A2(n11480), .ZN(n11487) );
  INV_X1 U9316 ( .A(n11487), .ZN(n7058) );
  NAND2_X1 U9317 ( .A1(n13944), .A2(n13945), .ZN(n6737) );
  AND2_X1 U9318 ( .A1(n11762), .A2(n11680), .ZN(n6738) );
  NAND2_X1 U9319 ( .A1(n14627), .A2(n14336), .ZN(n6739) );
  AND2_X1 U9320 ( .A1(n13802), .A2(n13559), .ZN(n6740) );
  AND2_X1 U9321 ( .A1(n8882), .A2(n14856), .ZN(n6741) );
  INV_X1 U9322 ( .A(n8132), .ZN(n7638) );
  AND2_X1 U9323 ( .A1(n8451), .A2(n8450), .ZN(n13639) );
  INV_X1 U9324 ( .A(n13639), .ZN(n13858) );
  AND2_X1 U9325 ( .A1(n9340), .A2(n11580), .ZN(n6742) );
  INV_X1 U9326 ( .A(n9908), .ZN(n7112) );
  NOR2_X1 U9327 ( .A1(n9347), .A2(n9164), .ZN(n6743) );
  NOR2_X1 U9328 ( .A1(n14921), .A2(n12198), .ZN(n6744) );
  INV_X1 U9329 ( .A(n7319), .ZN(n7318) );
  OAI21_X1 U9330 ( .B1(n12958), .B2(n7320), .A(n9331), .ZN(n7319) );
  INV_X1 U9331 ( .A(n8303), .ZN(n7658) );
  INV_X1 U9332 ( .A(n8345), .ZN(n7669) );
  AND2_X1 U9333 ( .A1(n8066), .A2(n8065), .ZN(n6745) );
  OR2_X1 U9334 ( .A1(n13816), .A2(n13556), .ZN(n6746) );
  AND2_X1 U9335 ( .A1(n13361), .A2(n11084), .ZN(n6747) );
  AND3_X1 U9336 ( .A1(n9619), .A2(n9618), .A3(n9617), .ZN(n15167) );
  INV_X1 U9337 ( .A(n15167), .ZN(n6901) );
  NAND2_X1 U9338 ( .A1(n7174), .A2(n13530), .ZN(n7181) );
  INV_X1 U9339 ( .A(n7181), .ZN(n7177) );
  AND2_X1 U9340 ( .A1(n14396), .A2(n7607), .ZN(n6748) );
  OR2_X1 U9341 ( .A1(n7999), .A2(n7998), .ZN(n6749) );
  AND2_X1 U9342 ( .A1(n8266), .A2(n8265), .ZN(n13550) );
  INV_X1 U9343 ( .A(n13550), .ZN(n14907) );
  OR2_X1 U9344 ( .A1(n7045), .A2(n11583), .ZN(n6750) );
  NAND2_X1 U9345 ( .A1(n7827), .A2(SI_9_), .ZN(n7829) );
  INV_X1 U9346 ( .A(n7829), .ZN(n7708) );
  AND2_X1 U9347 ( .A1(n10004), .A2(n10003), .ZN(n14361) );
  INV_X1 U9348 ( .A(n14361), .ZN(n14576) );
  NOR2_X1 U9349 ( .A1(n12190), .A2(n7148), .ZN(n7147) );
  AND2_X1 U9350 ( .A1(n7497), .A2(n14331), .ZN(n6751) );
  INV_X1 U9351 ( .A(n12070), .ZN(n11616) );
  AND2_X1 U9352 ( .A1(n12639), .A2(n7138), .ZN(n6752) );
  AND2_X1 U9353 ( .A1(n7731), .A2(n7729), .ZN(n6753) );
  NAND2_X1 U9354 ( .A1(n8397), .A2(n8396), .ZN(n6754) );
  INV_X1 U9355 ( .A(n7357), .ZN(n7356) );
  NAND2_X1 U9356 ( .A1(n7358), .A2(n11885), .ZN(n7357) );
  AND2_X1 U9357 ( .A1(n14413), .A2(n6731), .ZN(n6755) );
  AND2_X1 U9358 ( .A1(n7050), .A2(n12909), .ZN(n6756) );
  NOR2_X1 U9359 ( .A1(n13139), .A2(n12997), .ZN(n6757) );
  AND2_X1 U9360 ( .A1(n13816), .A2(n13556), .ZN(n6758) );
  NAND3_X1 U9361 ( .A1(n12458), .A2(n8626), .A3(n13373), .ZN(n6759) );
  AND2_X1 U9362 ( .A1(n9291), .A2(n9285), .ZN(n13097) );
  INV_X1 U9363 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U9364 ( .A1(n9777), .A2(n7531), .ZN(n6760) );
  AND2_X1 U9365 ( .A1(n7616), .A2(n7615), .ZN(n6761) );
  INV_X1 U9366 ( .A(n11988), .ZN(n7150) );
  AND2_X1 U9367 ( .A1(n12513), .A2(n12656), .ZN(n6762) );
  OR2_X1 U9368 ( .A1(n7664), .A2(n7666), .ZN(n6763) );
  NOR2_X1 U9369 ( .A1(n11879), .A2(n14175), .ZN(n6764) );
  AND2_X1 U9370 ( .A1(n10787), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6765) );
  AND2_X1 U9371 ( .A1(n7476), .A2(n7474), .ZN(n6766) );
  NOR2_X1 U9372 ( .A1(n14484), .A2(n14336), .ZN(n6767) );
  NOR2_X1 U9373 ( .A1(n14589), .A2(n14344), .ZN(n6768) );
  NOR2_X1 U9374 ( .A1(n11504), .A2(n11503), .ZN(n6769) );
  NOR2_X1 U9375 ( .A1(n12383), .A2(n12382), .ZN(n6770) );
  INV_X1 U9376 ( .A(n8363), .ZN(n7671) );
  AND2_X1 U9377 ( .A1(n9543), .A2(n7504), .ZN(n6771) );
  AND2_X1 U9378 ( .A1(n9543), .A2(n7609), .ZN(n6772) );
  AND2_X1 U9379 ( .A1(n12524), .A2(n13018), .ZN(n6773) );
  AND2_X1 U9380 ( .A1(n15399), .A2(n12108), .ZN(n6774) );
  AND2_X1 U9381 ( .A1(n12960), .A2(n12897), .ZN(n6775) );
  AND2_X1 U9382 ( .A1(n14452), .A2(n14339), .ZN(n6776) );
  INV_X1 U9383 ( .A(n7436), .ZN(n7435) );
  OAI21_X1 U9384 ( .B1(n6725), .B2(n7437), .A(n12494), .ZN(n7436) );
  INV_X1 U9385 ( .A(n14026), .ZN(n15159) );
  NAND2_X1 U9386 ( .A1(n9606), .A2(n7084), .ZN(n14026) );
  AND2_X1 U9387 ( .A1(n7672), .A2(n7676), .ZN(n6777) );
  AND2_X1 U9388 ( .A1(n9390), .A2(n9389), .ZN(n6778) );
  AND2_X1 U9389 ( .A1(n7517), .A2(n7106), .ZN(n6779) );
  AND2_X1 U9390 ( .A1(n7512), .A2(n7107), .ZN(n6780) );
  AND2_X1 U9391 ( .A1(n9417), .A2(n9416), .ZN(n6781) );
  NAND2_X1 U9392 ( .A1(n7603), .A2(n6731), .ZN(n6782) );
  INV_X1 U9393 ( .A(n7580), .ZN(n7579) );
  NAND2_X1 U9394 ( .A1(n7584), .A2(n7581), .ZN(n7580) );
  INV_X1 U9395 ( .A(n12919), .ZN(n7775) );
  AND2_X1 U9396 ( .A1(n11375), .A2(n11392), .ZN(n6783) );
  NOR2_X1 U9397 ( .A1(n9459), .A2(n9458), .ZN(n6784) );
  OR2_X1 U9398 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n8643) );
  INV_X1 U9399 ( .A(n8643), .ZN(n7460) );
  AND2_X1 U9400 ( .A1(n11706), .A2(n11705), .ZN(n6785) );
  INV_X1 U9401 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9811) );
  AND2_X1 U9402 ( .A1(n7267), .A2(n6919), .ZN(n6786) );
  INV_X1 U9403 ( .A(n11953), .ZN(n7464) );
  NAND2_X1 U9404 ( .A1(n13118), .A2(n12908), .ZN(n6787) );
  AND2_X1 U9405 ( .A1(n8248), .A2(n8247), .ZN(n12383) );
  INV_X1 U9406 ( .A(n12383), .ZN(n14893) );
  INV_X1 U9407 ( .A(n10047), .ZN(n14546) );
  XOR2_X1 U9408 ( .A(n15921), .B(n15920), .Z(n6788) );
  AND2_X1 U9409 ( .A1(n7769), .A2(n12895), .ZN(n6789) );
  AND2_X1 U9410 ( .A1(n14054), .A2(n6737), .ZN(n7368) );
  INV_X1 U9411 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8642) );
  INV_X1 U9412 ( .A(n7630), .ZN(n7629) );
  NAND2_X1 U9413 ( .A1(n7631), .A2(n8132), .ZN(n7630) );
  INV_X1 U9414 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U9415 ( .A1(n14026), .A2(n6896), .ZN(n11494) );
  XNOR2_X1 U9416 ( .A(n14589), .B(n10044), .ZN(n14379) );
  INV_X1 U9417 ( .A(n12359), .ZN(n12367) );
  OR2_X1 U9418 ( .A1(n8048), .A2(n8047), .ZN(n6790) );
  OR2_X1 U9419 ( .A1(n7810), .A2(SI_2_), .ZN(n6791) );
  AND2_X1 U9420 ( .A1(n6899), .A2(n14577), .ZN(n6792) );
  AND3_X1 U9421 ( .A1(n14586), .A2(n14584), .A3(n14585), .ZN(n6793) );
  AND2_X1 U9422 ( .A1(n8872), .A2(n8871), .ZN(n14850) );
  NOR2_X1 U9423 ( .A1(n13677), .A2(n7730), .ZN(n7729) );
  AND2_X1 U9424 ( .A1(n6720), .A2(n10042), .ZN(n6794) );
  INV_X1 U9425 ( .A(n9445), .ZN(n7552) );
  AND2_X1 U9426 ( .A1(n8194), .A2(n15873), .ZN(n6795) );
  NAND2_X1 U9427 ( .A1(n13910), .A2(n13909), .ZN(n6796) );
  OR2_X1 U9428 ( .A1(n9881), .A2(n9882), .ZN(n6797) );
  AND2_X1 U9429 ( .A1(n9591), .A2(n9592), .ZN(n6798) );
  AND2_X1 U9430 ( .A1(n12073), .A2(n12072), .ZN(n6799) );
  AND2_X1 U9431 ( .A1(n6730), .A2(n13512), .ZN(n6800) );
  AND2_X1 U9432 ( .A1(n7470), .A2(n7469), .ZN(n6802) );
  AND2_X1 U9433 ( .A1(n7506), .A2(n9700), .ZN(n6803) );
  AND2_X1 U9434 ( .A1(n13548), .A2(n13547), .ZN(n6804) );
  AND2_X1 U9435 ( .A1(n7655), .A2(n8319), .ZN(n6805) );
  AND2_X1 U9436 ( .A1(n7224), .A2(n7223), .ZN(n6806) );
  OAI21_X1 U9437 ( .B1(n7667), .B2(n7664), .A(n7663), .ZN(n7662) );
  NAND2_X1 U9438 ( .A1(n7539), .A2(n9713), .ZN(n6807) );
  NAND2_X1 U9439 ( .A1(n7542), .A2(n9747), .ZN(n6808) );
  OR2_X1 U9440 ( .A1(n13609), .A2(n13573), .ZN(n6809) );
  INV_X1 U9441 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9569) );
  INV_X1 U9442 ( .A(n7786), .ZN(n7785) );
  NAND2_X1 U9443 ( .A1(n7787), .A2(n12868), .ZN(n7786) );
  AND2_X1 U9444 ( .A1(n7475), .A2(n7477), .ZN(n7474) );
  INV_X1 U9445 ( .A(n7044), .ZN(n7774) );
  NAND2_X1 U9446 ( .A1(n7775), .A2(n12902), .ZN(n7044) );
  INV_X1 U9447 ( .A(n7750), .ZN(n7749) );
  NAND2_X1 U9448 ( .A1(n7849), .A2(n7751), .ZN(n7750) );
  OR2_X1 U9449 ( .A1(n13248), .A2(n6988), .ZN(n6810) );
  INV_X1 U9450 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7095) );
  INV_X1 U9451 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7142) );
  INV_X1 U9452 ( .A(n7798), .ZN(n12389) );
  INV_X1 U9453 ( .A(SI_3_), .ZN(n7067) );
  INV_X1 U9454 ( .A(n14477), .ZN(n7605) );
  AND2_X1 U9455 ( .A1(n8149), .A2(n8148), .ZN(n14945) );
  INV_X1 U9456 ( .A(n14945), .ZN(n7230) );
  NAND2_X1 U9457 ( .A1(n8381), .A2(n8380), .ZN(n13802) );
  INV_X1 U9458 ( .A(n13802), .ZN(n7236) );
  NAND2_X1 U9459 ( .A1(n8610), .A2(n7849), .ZN(n8608) );
  NOR2_X1 U9460 ( .A1(n13163), .A2(n12880), .ZN(n6811) );
  AND2_X1 U9461 ( .A1(n10947), .A2(n11019), .ZN(n6812) );
  AND2_X1 U9462 ( .A1(n15038), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6813) );
  INV_X1 U9463 ( .A(n13596), .ZN(n13850) );
  AND2_X1 U9464 ( .A1(n8502), .A2(n8501), .ZN(n13596) );
  NAND2_X1 U9465 ( .A1(n8658), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8675) );
  AND2_X1 U9466 ( .A1(n13596), .A2(n14903), .ZN(n6814) );
  AND3_X1 U9467 ( .A1(n8806), .A2(n8805), .A3(n8804), .ZN(n12131) );
  AND2_X1 U9468 ( .A1(n7848), .A2(n7847), .ZN(n8610) );
  AND2_X1 U9469 ( .A1(n10123), .A2(n10134), .ZN(n6815) );
  AND4_X1 U9470 ( .A1(n8185), .A2(n8184), .A3(n8183), .A4(n8182), .ZN(n12477)
         );
  INV_X1 U9471 ( .A(n14461), .ZN(n6906) );
  NAND2_X1 U9472 ( .A1(n12332), .A2(n12331), .ZN(n12869) );
  AND3_X1 U9473 ( .A1(n7449), .A2(n7448), .A3(n7447), .ZN(n6816) );
  INV_X1 U9474 ( .A(n7286), .ZN(n14541) );
  NOR2_X1 U9475 ( .A1(n14558), .A2(n14650), .ZN(n7286) );
  NOR2_X1 U9476 ( .A1(n12064), .A2(n13353), .ZN(n6817) );
  AND2_X1 U9477 ( .A1(n12291), .A2(n9431), .ZN(n6818) );
  AND2_X1 U9478 ( .A1(n8331), .A2(n15895), .ZN(n6819) );
  AND2_X1 U9479 ( .A1(n8420), .A2(n15662), .ZN(n6820) );
  INV_X1 U9480 ( .A(n7784), .ZN(n7782) );
  NOR2_X1 U9481 ( .A1(n12870), .A2(n14863), .ZN(n7784) );
  OR2_X1 U9482 ( .A1(n13091), .A2(n13097), .ZN(n6821) );
  INV_X1 U9483 ( .A(n6904), .ZN(n14447) );
  NOR2_X1 U9484 ( .A1(n14481), .A2(n6905), .ZN(n6904) );
  INV_X1 U9485 ( .A(n9746), .ZN(n7542) );
  AND2_X1 U9486 ( .A1(n7465), .A2(n7464), .ZN(n6822) );
  OR2_X1 U9487 ( .A1(n13915), .A2(n13916), .ZN(n7386) );
  INV_X1 U9488 ( .A(n12867), .ZN(n14857) );
  AND4_X1 U9489 ( .A1(n8832), .A2(n8831), .A3(n8830), .A4(n8829), .ZN(n12867)
         );
  INV_X1 U9490 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7790) );
  INV_X1 U9491 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10232) );
  INV_X1 U9492 ( .A(n14935), .ZN(n13741) );
  INV_X1 U9493 ( .A(n12775), .ZN(n7038) );
  INV_X1 U9494 ( .A(n12672), .ZN(n7432) );
  INV_X1 U9495 ( .A(n11912), .ZN(n7087) );
  INV_X1 U9496 ( .A(n12714), .ZN(n7101) );
  AND2_X2 U9497 ( .A1(n10982), .A2(n10824), .ZN(n15532) );
  INV_X1 U9498 ( .A(n15532), .ZN(n15530) );
  NAND2_X1 U9499 ( .A1(n15411), .A2(n11576), .ZN(n11596) );
  NAND2_X1 U9500 ( .A1(n7226), .A2(n7590), .ZN(n11818) );
  NAND2_X1 U9501 ( .A1(n6954), .A2(n6952), .ZN(n15393) );
  NAND2_X1 U9502 ( .A1(n7592), .A2(n11641), .ZN(n11745) );
  INV_X1 U9503 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7751) );
  OR2_X1 U9504 ( .A1(n15532), .A2(n9114), .ZN(n6823) );
  AND2_X1 U9505 ( .A1(n12822), .A2(n12807), .ZN(n6824) );
  INV_X1 U9506 ( .A(n7285), .ZN(n11551) );
  NOR2_X1 U9507 ( .A1(n11550), .A2(n11556), .ZN(n7285) );
  AND2_X1 U9508 ( .A1(n8472), .A2(n15597), .ZN(n6825) );
  OR2_X1 U9509 ( .A1(n15532), .A2(n9126), .ZN(n6826) );
  AND2_X1 U9510 ( .A1(n6985), .A2(n7782), .ZN(n6827) );
  NAND2_X1 U9511 ( .A1(n10111), .A2(n10627), .ZN(n11368) );
  NOR2_X1 U9512 ( .A1(n15389), .A2(n15381), .ZN(n13837) );
  INV_X1 U9513 ( .A(n14181), .ZN(n7011) );
  NAND2_X1 U9514 ( .A1(n11579), .A2(n11578), .ZN(n15453) );
  NAND2_X1 U9515 ( .A1(n10819), .A2(n11565), .ZN(n15512) );
  INV_X1 U9516 ( .A(n12850), .ZN(n11577) );
  AND2_X1 U9517 ( .A1(n10870), .A2(n7140), .ZN(n6828) );
  INV_X1 U9518 ( .A(n15100), .ZN(n6902) );
  OR2_X1 U9519 ( .A1(n12811), .A2(n12792), .ZN(n6829) );
  INV_X1 U9520 ( .A(n11119), .ZN(n7571) );
  AND2_X1 U9521 ( .A1(n11587), .A2(n11586), .ZN(n15416) );
  INV_X1 U9522 ( .A(n15416), .ZN(n15435) );
  OR2_X1 U9523 ( .A1(n7990), .A2(n12460), .ZN(n6830) );
  NOR2_X1 U9524 ( .A1(n7990), .A2(n13886), .ZN(n6831) );
  AND2_X1 U9525 ( .A1(n14249), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6832) );
  OR2_X1 U9526 ( .A1(n10885), .A2(n10789), .ZN(n7283) );
  INV_X1 U9527 ( .A(n10790), .ZN(n7282) );
  AND2_X1 U9528 ( .A1(n12699), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6833) );
  INV_X1 U9529 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7690) );
  INV_X1 U9530 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7000) );
  INV_X1 U9531 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7293) );
  XNOR2_X1 U9532 ( .A(n11003), .B(n11019), .ZN(n10967) );
  OR2_X1 U9533 ( .A1(n10947), .A2(n11019), .ZN(n7214) );
  OR2_X1 U9534 ( .A1(n10948), .A2(n11019), .ZN(n7213) );
  OR2_X1 U9535 ( .A1(n10195), .A2(n10249), .ZN(n15389) );
  AOI21_X1 U9536 ( .B1(n13850), .B2(n13837), .A(n7206), .ZN(n7205) );
  INV_X1 U9537 ( .A(n13837), .ZN(n7353) );
  NAND2_X2 U9538 ( .A1(n11933), .A2(n9369), .ZN(n9379) );
  NAND2_X1 U9539 ( .A1(n11874), .A2(n9421), .ZN(n12238) );
  NAND2_X1 U9540 ( .A1(n6838), .A2(n9413), .ZN(n11809) );
  NAND2_X1 U9541 ( .A1(n6840), .A2(n6839), .ZN(n9404) );
  AOI21_X1 U9542 ( .B1(n7569), .B2(n7571), .A(n6708), .ZN(n6839) );
  NAND2_X1 U9543 ( .A1(n11120), .A2(n7569), .ZN(n6840) );
  AOI21_X1 U9544 ( .B1(n11119), .B2(n7570), .A(n6842), .ZN(n6841) );
  INV_X1 U9545 ( .A(n11036), .ZN(n6843) );
  NAND2_X1 U9546 ( .A1(n6844), .A2(n9463), .ZN(n13260) );
  XNOR2_X1 U9547 ( .A(n9462), .B(n9460), .ZN(n13315) );
  INV_X2 U9548 ( .A(n8615), .ZN(n7869) );
  NAND2_X2 U9549 ( .A1(n7847), .A2(n7572), .ZN(n8615) );
  NAND2_X1 U9550 ( .A1(n7869), .A2(n7867), .ZN(n7877) );
  NAND2_X1 U9551 ( .A1(n8689), .A2(n6848), .ZN(n8691) );
  NAND2_X1 U9552 ( .A1(n10167), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8690) );
  INV_X1 U9553 ( .A(n8675), .ZN(n6851) );
  NAND3_X1 U9554 ( .A1(n8995), .A2(n9008), .A3(n11673), .ZN(n9009) );
  NAND3_X1 U9555 ( .A1(n8865), .A2(P1_DATAO_REG_13__SCAN_IN), .A3(n8883), .ZN(
        n8884) );
  NAND2_X1 U9556 ( .A1(n6852), .A2(n10457), .ZN(n8883) );
  XNOR2_X1 U9557 ( .A(n6857), .B(n6788), .ZN(SUB_1596_U4) );
  OAI21_X2 U9558 ( .B1(n14797), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n14827), .ZN(
        n15918) );
  NAND2_X1 U9559 ( .A1(n6861), .A2(n14759), .ZN(n14700) );
  XNOR2_X1 U9560 ( .A(n7005), .B(n6861), .ZN(n14761) );
  NAND2_X1 U9561 ( .A1(n6862), .A2(n10109), .ZN(P1_U3242) );
  NAND2_X1 U9562 ( .A1(n6863), .A2(n10089), .ZN(n6862) );
  OAI211_X1 U9563 ( .C1(n10084), .C2(n6865), .A(n6864), .B(n7794), .ZN(n6863)
         );
  NAND2_X1 U9564 ( .A1(n10084), .A2(n6794), .ZN(n6864) );
  AND2_X2 U9565 ( .A1(n6872), .A2(n6871), .ZN(n9858) );
  NAND2_X1 U9566 ( .A1(n10027), .A2(n11905), .ZN(n6871) );
  NAND2_X1 U9567 ( .A1(n9985), .A2(n9984), .ZN(n6878) );
  NAND2_X1 U9568 ( .A1(n7103), .A2(n6883), .ZN(n14662) );
  NAND2_X1 U9569 ( .A1(n14579), .A2(n15189), .ZN(n6883) );
  XNOR2_X1 U9570 ( .A(n6884), .B(n14348), .ZN(n14579) );
  NAND3_X1 U9571 ( .A1(n6886), .A2(n6885), .A3(n7492), .ZN(n7491) );
  NAND2_X1 U9572 ( .A1(n14952), .A2(n14325), .ZN(n6888) );
  NAND2_X1 U9573 ( .A1(n14323), .A2(n14322), .ZN(n6889) );
  OAI211_X1 U9574 ( .C1(n11820), .C2(n6891), .A(n6890), .B(n12036), .ZN(n12040) );
  NAND2_X1 U9575 ( .A1(n7498), .A2(n6893), .ZN(n6890) );
  INV_X1 U9576 ( .A(n7498), .ZN(n6891) );
  NAND2_X1 U9577 ( .A1(n6892), .A2(n7498), .ZN(n12037) );
  NAND2_X1 U9578 ( .A1(n11820), .A2(n11738), .ZN(n6892) );
  INV_X1 U9579 ( .A(n11738), .ZN(n6893) );
  AOI21_X2 U9580 ( .B1(n7502), .B2(n7501), .A(n7500), .ZN(n14380) );
  NAND3_X1 U9581 ( .A1(n7474), .A2(n14490), .A3(n14335), .ZN(n6895) );
  NAND2_X1 U9582 ( .A1(n7801), .A2(n14500), .ZN(n14490) );
  NAND2_X1 U9583 ( .A1(n9610), .A2(n11494), .ZN(n15088) );
  NAND2_X1 U9584 ( .A1(n10128), .A2(n6668), .ZN(n9593) );
  NAND2_X1 U9585 ( .A1(n14349), .A2(n7287), .ZN(n14578) );
  INV_X1 U9586 ( .A(n6898), .ZN(n14349) );
  NOR2_X1 U9587 ( .A1(n6898), .A2(n15205), .ZN(n6897) );
  NOR2_X1 U9588 ( .A1(n14384), .A2(n14583), .ZN(n14370) );
  NAND3_X1 U9589 ( .A1(n7087), .A2(n15081), .A3(n15201), .ZN(n11843) );
  NAND2_X1 U9590 ( .A1(n6907), .A2(n7692), .ZN(n8423) );
  NAND2_X1 U9591 ( .A1(n6911), .A2(n6910), .ZN(n6907) );
  NAND2_X1 U9592 ( .A1(n8375), .A2(n7692), .ZN(n6908) );
  INV_X1 U9593 ( .A(n7692), .ZN(n6909) );
  NAND2_X1 U9594 ( .A1(n8375), .A2(n8399), .ZN(n9908) );
  NAND3_X1 U9595 ( .A1(n7740), .A2(n8448), .A3(n7737), .ZN(n6934) );
  NAND2_X1 U9596 ( .A1(n7304), .A2(n11566), .ZN(n7303) );
  NAND2_X1 U9597 ( .A1(n15407), .A2(n8698), .ZN(n6935) );
  NAND2_X1 U9598 ( .A1(n6945), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U9599 ( .A1(n11773), .A2(n6956), .ZN(n6954) );
  AND2_X2 U9600 ( .A1(n10639), .A2(n10154), .ZN(n8666) );
  AND2_X1 U9601 ( .A1(n6967), .A2(n6965), .ZN(n12071) );
  NAND2_X1 U9602 ( .A1(n7761), .A2(n6966), .ZN(n6965) );
  NAND2_X1 U9603 ( .A1(n6968), .A2(n11615), .ZN(n6967) );
  INV_X1 U9604 ( .A(n6977), .ZN(n13059) );
  INV_X1 U9605 ( .A(n12869), .ZN(n6980) );
  OAI21_X1 U9606 ( .B1(n6980), .B2(n6718), .A(n6981), .ZN(n14832) );
  NAND2_X1 U9607 ( .A1(n6986), .A2(n12909), .ZN(n13114) );
  AND3_X2 U9608 ( .A1(n7310), .A2(n6810), .A3(n6715), .ZN(n15426) );
  NAND2_X1 U9609 ( .A1(n9357), .A2(n6987), .ZN(n13238) );
  NAND2_X1 U9610 ( .A1(n12151), .A2(n12074), .ZN(n12154) );
  INV_X1 U9611 ( .A(n7740), .ZN(n7738) );
  XNOR2_X1 U9612 ( .A(n12019), .B(n12027), .ZN(n15058) );
  NAND2_X1 U9613 ( .A1(n7511), .A2(n9957), .ZN(n7510) );
  OAI21_X1 U9614 ( .B1(n13016), .B2(n7778), .A(n7776), .ZN(n12995) );
  OR2_X1 U9615 ( .A1(n7514), .A2(n7105), .ZN(n9985) );
  NAND2_X1 U9616 ( .A1(n8563), .A2(n8546), .ZN(n8560) );
  OAI211_X1 U9617 ( .C1(n8560), .C2(n7061), .A(n7093), .B(n7094), .ZN(n7014)
         );
  INV_X1 U9618 ( .A(n7014), .ZN(n8568) );
  NAND2_X2 U9619 ( .A1(n7361), .A2(n7359), .ZN(n14097) );
  NAND2_X1 U9620 ( .A1(n14128), .A2(n7111), .ZN(n14031) );
  INV_X2 U9621 ( .A(n7048), .ZN(n13915) );
  OAI21_X2 U9622 ( .B1(n14099), .B2(n14065), .A(n14064), .ZN(n14063) );
  AOI21_X2 U9623 ( .B1(n14097), .B2(n14096), .A(n14095), .ZN(n14099) );
  NAND2_X1 U9624 ( .A1(n14140), .A2(n14141), .ZN(n14139) );
  OAI211_X1 U9625 ( .C1(n12856), .C2(n12855), .A(n6802), .B(n6990), .ZN(
        P3_U3201) );
  NAND2_X1 U9626 ( .A1(n7326), .A2(n9204), .ZN(n12865) );
  MUX2_X1 U9627 ( .A(n13190), .B(P3_REG0_REG_29__SCAN_IN), .S(n15517), .Z(
        P3_U3456) );
  INV_X1 U9628 ( .A(n11571), .ZN(n15429) );
  AOI21_X1 U9629 ( .B1(n7332), .B2(n9297), .A(n7331), .ZN(n7330) );
  NAND2_X1 U9630 ( .A1(n7303), .A2(n7305), .ZN(n11773) );
  NAND2_X1 U9631 ( .A1(n10423), .A2(n15437), .ZN(n9226) );
  XNOR2_X1 U9632 ( .A(n11281), .B(n11282), .ZN(n14019) );
  OAI21_X1 U9633 ( .B1(n13907), .B2(n13908), .A(n6796), .ZN(n7048) );
  OAI22_X2 U9634 ( .A1(n13915), .A2(n7381), .B1(n13916), .B2(n7384), .ZN(
        n14086) );
  NAND2_X1 U9635 ( .A1(n7297), .A2(n7300), .ZN(n12325) );
  OAI21_X2 U9636 ( .B1(n14086), .B2(n14085), .A(n14084), .ZN(n14083) );
  NAND2_X1 U9637 ( .A1(n11352), .A2(n11351), .ZN(n11409) );
  NAND2_X2 U9638 ( .A1(n10106), .A2(n14690), .ZN(n10546) );
  NAND2_X1 U9639 ( .A1(n14083), .A2(n13930), .ZN(n14129) );
  NAND2_X1 U9640 ( .A1(n12969), .A2(n9063), .ZN(n12968) );
  NAND2_X1 U9641 ( .A1(n8887), .A2(n8886), .ZN(n8902) );
  NAND2_X1 U9642 ( .A1(n12407), .A2(n12406), .ZN(n13907) );
  NAND2_X1 U9643 ( .A1(n7415), .A2(n9348), .ZN(n7045) );
  NAND2_X1 U9644 ( .A1(n12219), .A2(n12218), .ZN(n12223) );
  NAND2_X1 U9645 ( .A1(n7021), .A2(n7020), .ZN(n9330) );
  NAND2_X1 U9646 ( .A1(n11697), .A2(n10038), .ZN(n7015) );
  OAI22_X2 U9647 ( .A1(n14380), .A2(n14379), .B1(n14389), .B2(n14344), .ZN(
        n14365) );
  NAND2_X1 U9648 ( .A1(n14333), .A2(n7490), .ZN(n7489) );
  NAND2_X1 U9649 ( .A1(n7113), .A2(n8323), .ZN(n8306) );
  NAND2_X1 U9650 ( .A1(n14587), .A2(n6793), .ZN(n14663) );
  NAND2_X1 U9651 ( .A1(n7112), .A2(n10153), .ZN(n9909) );
  NAND2_X1 U9652 ( .A1(n7042), .A2(n11696), .ZN(n8995) );
  NAND2_X1 U9653 ( .A1(n9165), .A2(n9166), .ZN(n6997) );
  OAI22_X1 U9654 ( .A1(n9199), .A2(n11578), .B1(n6998), .B2(n10862), .ZN(n9353) );
  XNOR2_X1 U9655 ( .A(n9198), .B(n11577), .ZN(n6998) );
  INV_X1 U9656 ( .A(n9050), .ZN(n6999) );
  INV_X1 U9657 ( .A(n8994), .ZN(n7042) );
  OAI22_X1 U9658 ( .A1(n12995), .A2(n12890), .B1(n13007), .B2(n13213), .ZN(
        n12983) );
  NAND2_X1 U9659 ( .A1(n11572), .A2(n11571), .ZN(n15432) );
  NAND2_X1 U9660 ( .A1(n12874), .A2(n12873), .ZN(n13091) );
  NAND2_X1 U9661 ( .A1(n12330), .A2(n12329), .ZN(n12333) );
  OR2_X1 U9662 ( .A1(n9123), .A2(n15459), .ZN(n8664) );
  NAND2_X1 U9663 ( .A1(n7752), .A2(n6799), .ZN(n12151) );
  NAND2_X1 U9664 ( .A1(n11570), .A2(n15445), .ZN(n15427) );
  NAND2_X1 U9665 ( .A1(n7002), .A2(n12879), .ZN(n13048) );
  NAND2_X1 U9666 ( .A1(n13059), .A2(n12878), .ZN(n7002) );
  NAND2_X1 U9667 ( .A1(n10867), .A2(n9222), .ZN(n11570) );
  INV_X1 U9669 ( .A(n7761), .ZN(n7760) );
  OAI21_X1 U9670 ( .B1(n12928), .B2(n7044), .A(n7773), .ZN(n12904) );
  NAND2_X1 U9671 ( .A1(n8072), .A2(n7826), .ZN(n8090) );
  NAND2_X1 U9672 ( .A1(n12044), .A2(n12043), .ZN(n12248) );
  NAND2_X1 U9673 ( .A1(n7491), .A2(n7489), .ZN(n7801) );
  AND2_X2 U9674 ( .A1(n9238), .A2(n9213), .ZN(n11600) );
  INV_X1 U9675 ( .A(n11497), .ZN(n7487) );
  INV_X1 U9676 ( .A(n7486), .ZN(n7483) );
  NAND2_X1 U9677 ( .A1(n15004), .A2(n15002), .ZN(n15009) );
  OAI21_X1 U9678 ( .B1(n11628), .B2(n11627), .A(n11626), .ZN(n15070) );
  AOI21_X1 U9679 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(n14783), .A(n14994), .ZN(
        n15000) );
  NOR2_X1 U9680 ( .A1(n9266), .A2(n7299), .ZN(n7298) );
  NOR2_X1 U9681 ( .A1(n9167), .A2(n8640), .ZN(n8641) );
  NAND2_X1 U9682 ( .A1(n9225), .A2(n9226), .ZN(n11571) );
  NAND2_X1 U9683 ( .A1(n13098), .A2(n13097), .ZN(n13100) );
  NAND2_X1 U9684 ( .A1(n8789), .A2(n9253), .ZN(n12150) );
  NAND2_X1 U9685 ( .A1(n7007), .A2(n7627), .ZN(n7625) );
  NAND2_X1 U9686 ( .A1(n7009), .A2(n8111), .ZN(n7007) );
  AOI21_X1 U9687 ( .B1(n8346), .B2(n7660), .A(n7662), .ZN(n8397) );
  OAI21_X1 U9688 ( .B1(n8257), .B2(n7651), .A(n7650), .ZN(n8280) );
  INV_X1 U9689 ( .A(n7077), .ZN(n7076) );
  OR2_X1 U9690 ( .A1(n8113), .A2(n8112), .ZN(n7009) );
  NOR2_X2 U9691 ( .A1(n8175), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n8219) );
  AOI21_X2 U9692 ( .B1(n6693), .B2(n8585), .A(n7171), .ZN(n7910) );
  NAND2_X1 U9693 ( .A1(n14300), .A2(n14299), .ZN(n14547) );
  XNOR2_X2 U9694 ( .A(n14320), .B(n14348), .ZN(n14580) );
  INV_X1 U9695 ( .A(n11542), .ZN(n11544) );
  NAND4_X1 U9696 ( .A1(n6797), .A2(n7060), .A3(n9870), .A4(n7538), .ZN(n7533)
         );
  NAND3_X1 U9697 ( .A1(n9850), .A2(n14520), .A3(n7097), .ZN(n7060) );
  NAND2_X1 U9698 ( .A1(n7059), .A2(n6803), .ZN(n9699) );
  NAND2_X1 U9699 ( .A1(n10137), .A2(n6668), .ZN(n9606) );
  NAND2_X2 U9700 ( .A1(n7015), .A2(n9851), .ZN(n14512) );
  AOI21_X1 U9701 ( .B1(n9943), .B2(n7512), .A(n7510), .ZN(n7509) );
  NAND2_X1 U9702 ( .A1(n15432), .A2(n11573), .ZN(n15411) );
  NAND2_X1 U9703 ( .A1(n7019), .A2(n9366), .ZN(P3_U3296) );
  OAI21_X1 U9704 ( .B1(n7080), .B2(n9353), .A(n9352), .ZN(n7019) );
  AOI21_X2 U9705 ( .B1(n13884), .B2(n8530), .A(n6831), .ZN(n13504) );
  NAND2_X1 U9706 ( .A1(n7022), .A2(n13097), .ZN(n9290) );
  NAND2_X1 U9707 ( .A1(n9282), .A2(n7023), .ZN(n7022) );
  OR2_X1 U9708 ( .A1(n9283), .A2(n10820), .ZN(n7023) );
  NAND2_X1 U9709 ( .A1(n7025), .A2(n7024), .ZN(n9252) );
  NAND2_X1 U9710 ( .A1(n9246), .A2(n7026), .ZN(n7025) );
  NOR2_X1 U9711 ( .A1(n12776), .A2(n12777), .ZN(n12782) );
  NOR2_X1 U9712 ( .A1(n12823), .A2(n7032), .ZN(n12799) );
  XNOR2_X1 U9713 ( .A(n12767), .B(n7038), .ZN(n12747) );
  AND2_X1 U9714 ( .A1(n12767), .A2(n7038), .ZN(n7035) );
  NAND2_X1 U9715 ( .A1(n7792), .A2(n7756), .ZN(n7754) );
  AOI21_X1 U9716 ( .B1(n10880), .B2(n10778), .A(n10777), .ZN(n10958) );
  NOR2_X1 U9717 ( .A1(n12745), .A2(n12744), .ZN(n12767) );
  CLKBUF_X3 U9718 ( .A(n10501), .Z(n12814) );
  AOI21_X1 U9719 ( .B1(n7037), .B2(n7036), .A(n12819), .ZN(n12820) );
  INV_X1 U9720 ( .A(n12837), .ZN(n7037) );
  INV_X1 U9721 ( .A(n13498), .ZN(n7041) );
  NAND2_X1 U9722 ( .A1(n7047), .A2(n9338), .ZN(n9339) );
  NAND2_X1 U9723 ( .A1(n9337), .A2(n12919), .ZN(n7047) );
  INV_X1 U9724 ( .A(n8561), .ZN(n7094) );
  NAND2_X1 U9725 ( .A1(n8070), .A2(n7264), .ZN(n7262) );
  NAND2_X1 U9726 ( .A1(n8448), .A2(n7738), .ZN(n8449) );
  NAND2_X1 U9727 ( .A1(n11288), .A2(n11287), .ZN(n11352) );
  NAND2_X1 U9728 ( .A1(n14021), .A2(n11283), .ZN(n11350) );
  NAND2_X1 U9729 ( .A1(n8052), .A2(n7823), .ZN(n8070) );
  NAND2_X1 U9730 ( .A1(n14501), .A2(n6694), .ZN(n7092) );
  NAND2_X1 U9731 ( .A1(n7549), .A2(n7550), .ZN(n7049) );
  NAND2_X1 U9732 ( .A1(n8070), .A2(n8069), .ZN(n8072) );
  NAND2_X1 U9733 ( .A1(n8050), .A2(n8049), .ZN(n8052) );
  OAI21_X2 U9734 ( .B1(n9456), .B2(n7560), .A(n7559), .ZN(n9462) );
  NAND2_X1 U9735 ( .A1(n7092), .A2(n7604), .ZN(n14469) );
  INV_X1 U9736 ( .A(n7104), .ZN(n7103) );
  NAND2_X1 U9737 ( .A1(n14960), .A2(n7596), .ZN(n14300) );
  NAND2_X1 U9738 ( .A1(n14306), .A2(n14305), .ZN(n14501) );
  NAND2_X1 U9739 ( .A1(n7066), .A2(n7986), .ZN(n7946) );
  NAND2_X1 U9740 ( .A1(n8089), .A2(n8090), .ZN(n8092) );
  NAND2_X1 U9741 ( .A1(n7051), .A2(n6826), .ZN(P3_U3488) );
  NAND2_X1 U9742 ( .A1(n13088), .A2(n13087), .ZN(n13086) );
  NAND2_X1 U9743 ( .A1(n13190), .A2(n15532), .ZN(n7051) );
  NAND3_X1 U9744 ( .A1(n7505), .A2(n9858), .A3(n7058), .ZN(n7057) );
  OAI21_X1 U9745 ( .B1(n7793), .B2(n9609), .A(n9608), .ZN(n9615) );
  NAND2_X1 U9746 ( .A1(n9959), .A2(n9958), .ZN(n9972) );
  NAND2_X1 U9747 ( .A1(n7100), .A2(n7099), .ZN(n9726) );
  AND2_X2 U9748 ( .A1(n13602), .A2(n13596), .ZN(n13593) );
  AND2_X2 U9749 ( .A1(n13621), .A2(n13609), .ZN(n13602) );
  NAND2_X1 U9750 ( .A1(n14469), .A2(n14468), .ZN(n7225) );
  NAND2_X1 U9751 ( .A1(n7062), .A2(n11474), .ZN(n15086) );
  NOR2_X2 U9752 ( .A1(n13500), .A2(n12389), .ZN(n13753) );
  NAND2_X1 U9753 ( .A1(n7548), .A2(n7547), .ZN(n11036) );
  INV_X1 U9754 ( .A(n10192), .ZN(n11227) );
  OAI21_X1 U9755 ( .B1(n7567), .B2(n6717), .A(n7563), .ZN(n14889) );
  NAND2_X1 U9756 ( .A1(n7682), .A2(n8464), .ZN(n8467) );
  NAND2_X1 U9757 ( .A1(n7068), .A2(n7067), .ZN(n7066) );
  INV_X1 U9758 ( .A(n7946), .ZN(n7114) );
  INV_X1 U9759 ( .A(n7809), .ZN(n7068) );
  NOR2_X1 U9760 ( .A1(n14808), .A2(n14807), .ZN(n14780) );
  NAND2_X1 U9761 ( .A1(n15918), .A2(n15919), .ZN(n7073) );
  NAND2_X1 U9762 ( .A1(n7075), .A2(n7074), .ZN(P2_U3528) );
  NAND2_X1 U9763 ( .A1(n13847), .A2(n15391), .ZN(n7075) );
  NAND2_X1 U9764 ( .A1(n13847), .A2(n15387), .ZN(n7245) );
  NAND2_X1 U9765 ( .A1(n7076), .A2(n6790), .ZN(n8068) );
  AOI21_X1 U9766 ( .B1(n8048), .B2(n8047), .A(n8046), .ZN(n7077) );
  NAND2_X1 U9767 ( .A1(n8302), .A2(n7657), .ZN(n7654) );
  NAND2_X1 U9768 ( .A1(n7654), .A2(n7655), .ZN(n8320) );
  OAI21_X1 U9769 ( .B1(n8110), .B2(n8109), .A(n8108), .ZN(n8111) );
  NAND2_X1 U9770 ( .A1(n7078), .A2(n7925), .ZN(n7926) );
  NAND2_X1 U9771 ( .A1(n7910), .A2(n7911), .ZN(n7078) );
  NAND2_X1 U9772 ( .A1(n7659), .A2(n8318), .ZN(n8322) );
  NAND2_X1 U9773 ( .A1(n12932), .A2(n15453), .ZN(n7115) );
  NOR2_X1 U9774 ( .A1(n6693), .A2(n7172), .ZN(n7171) );
  NAND2_X1 U9775 ( .A1(n8845), .A2(n8844), .ZN(n8848) );
  NAND2_X1 U9776 ( .A1(n7418), .A2(n7417), .ZN(n7416) );
  NAND2_X1 U9777 ( .A1(n7416), .A2(n9345), .ZN(n7415) );
  NAND2_X1 U9778 ( .A1(n7081), .A2(n6750), .ZN(n7080) );
  NAND3_X1 U9779 ( .A1(n7083), .A2(n7115), .A3(n7082), .ZN(n13123) );
  NAND2_X1 U9780 ( .A1(n9102), .A2(n7327), .ZN(n7326) );
  NAND2_X1 U9781 ( .A1(n12854), .A2(n12853), .ZN(n7470) );
  NAND2_X1 U9782 ( .A1(n7264), .A2(n7266), .ZN(n7263) );
  NAND3_X1 U9783 ( .A1(n13497), .A2(n7258), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7691) );
  NAND2_X2 U9784 ( .A1(n12470), .A2(n7898), .ZN(n7939) );
  AOI21_X2 U9785 ( .B1(n15309), .B2(P2_REG1_REG_17__SCAN_IN), .A(n15302), .ZN(
        n13485) );
  AOI21_X2 U9786 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n15284), .A(n15279), .ZN(
        n13450) );
  OAI21_X2 U9787 ( .B1(n7950), .B2(n7814), .A(n7813), .ZN(n7988) );
  INV_X1 U9788 ( .A(n8290), .ZN(n7113) );
  NAND2_X1 U9789 ( .A1(n8091), .A2(n8092), .ZN(n10172) );
  NAND3_X1 U9790 ( .A1(n9701), .A2(n9702), .A3(n6807), .ZN(n7100) );
  NAND2_X1 U9791 ( .A1(n7245), .A2(n7243), .ZN(P2_U3496) );
  OAI211_X1 U9792 ( .C1(n13663), .C2(n7175), .A(n13633), .B(n7179), .ZN(n13629) );
  INV_X1 U9793 ( .A(n7175), .ZN(n7180) );
  AND3_X2 U9794 ( .A1(n7248), .A2(n12184), .A3(n7249), .ZN(n12721) );
  NOR2_X1 U9795 ( .A1(n12755), .A2(n12754), .ZN(n12776) );
  NOR2_X1 U9796 ( .A1(n12722), .A2(n12723), .ZN(n12725) );
  NOR2_X1 U9797 ( .A1(n12823), .A2(n7255), .ZN(n12828) );
  OAI21_X1 U9798 ( .B1(n14580), .B2(n15176), .A(n6792), .ZN(n7104) );
  AOI21_X1 U9799 ( .B1(n11738), .B2(n11821), .A(n7499), .ZN(n7498) );
  AOI21_X1 U9800 ( .B1(n7537), .B2(n9881), .A(n7535), .ZN(n7534) );
  NAND2_X1 U9801 ( .A1(n7114), .A2(n6791), .ZN(n7812) );
  NAND2_X1 U9802 ( .A1(n8373), .A2(n15660), .ZN(n8375) );
  NAND2_X1 U9803 ( .A1(n7545), .A2(n7543), .ZN(n9474) );
  NAND2_X1 U9804 ( .A1(n9370), .A2(n10661), .ZN(n10741) );
  OAI21_X1 U9805 ( .B1(n9630), .B2(n9629), .A(n9628), .ZN(n9645) );
  NAND2_X1 U9806 ( .A1(n9343), .A2(n10820), .ZN(n7418) );
  NAND2_X1 U9807 ( .A1(n9078), .A2(n9077), .ZN(n9080) );
  XNOR2_X1 U9808 ( .A(n9119), .B(n9106), .ZN(n12491) );
  NAND2_X1 U9809 ( .A1(n7392), .A2(n8707), .ZN(n8728) );
  NAND2_X1 U9810 ( .A1(n8691), .A2(n8690), .ZN(n8706) );
  NAND2_X1 U9811 ( .A1(n9047), .A2(n9046), .ZN(n9049) );
  NAND2_X1 U9812 ( .A1(n9049), .A2(n9048), .ZN(n9050) );
  NOR2_X1 U9813 ( .A1(n12796), .A2(n13071), .ZN(n12823) );
  AOI21_X1 U9814 ( .B1(n7256), .B2(n12699), .A(n10753), .ZN(n12704) );
  NOR2_X1 U9815 ( .A1(n12185), .A2(n8876), .ZN(n12722) );
  XNOR2_X1 U9816 ( .A(n10754), .B(n10894), .ZN(n10888) );
  NAND2_X2 U9817 ( .A1(n10546), .A2(n10725), .ZN(n13942) );
  NAND2_X2 U9818 ( .A1(n14031), .A2(n7109), .ZN(n14108) );
  NAND2_X1 U9819 ( .A1(n8285), .A2(n8284), .ZN(n7716) );
  NAND3_X1 U9820 ( .A1(n7804), .A2(n7803), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7689) );
  INV_X1 U9821 ( .A(n7812), .ZN(n7948) );
  NAND2_X1 U9822 ( .A1(n8568), .A2(n7274), .ZN(n7273) );
  NAND2_X1 U9823 ( .A1(n14832), .A2(n14836), .ZN(n12874) );
  NAND2_X1 U9824 ( .A1(n7118), .A2(n7116), .ZN(P3_U3486) );
  INV_X1 U9825 ( .A(n7117), .ZN(n7116) );
  NAND2_X1 U9826 ( .A1(n14508), .A2(n14634), .ZN(n14495) );
  INV_X1 U9827 ( .A(n14770), .ZN(n7294) );
  OAI21_X1 U9828 ( .B1(n15000), .B2(n14999), .A(n7289), .ZN(n7288) );
  NOR2_X1 U9829 ( .A1(n12837), .A2(n7124), .ZN(n12843) );
  AND2_X1 U9830 ( .A1(n12839), .A2(n12838), .ZN(n7124) );
  NOR2_X4 U9831 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8678) );
  NOR2_X2 U9832 ( .A1(n8709), .A2(n8635), .ZN(n8782) );
  NAND2_X1 U9833 ( .A1(n12676), .A2(n7132), .ZN(n7131) );
  NAND2_X1 U9834 ( .A1(n8926), .A2(n7141), .ZN(n8977) );
  NAND2_X1 U9835 ( .A1(n13727), .A2(n6707), .ZN(n7160) );
  NAND2_X1 U9836 ( .A1(n7159), .A2(n7728), .ZN(n13667) );
  NAND3_X1 U9837 ( .A1(n7160), .A2(n7161), .A3(n7729), .ZN(n7159) );
  NAND2_X1 U9838 ( .A1(n7163), .A2(SI_1_), .ZN(n7807) );
  MUX2_X1 U9839 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n7816), .Z(n7163) );
  NAND2_X2 U9840 ( .A1(n7165), .A2(n7164), .ZN(n7816) );
  NAND2_X1 U9841 ( .A1(n7689), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U9842 ( .A1(n7691), .A2(n7690), .ZN(n7165) );
  NAND2_X1 U9843 ( .A1(n6693), .A2(n13364), .ZN(n7907) );
  INV_X1 U9844 ( .A(n13364), .ZN(n7172) );
  NAND4_X2 U9845 ( .A1(n7896), .A2(n7895), .A3(n7897), .A4(n7894), .ZN(n13364)
         );
  OAI21_X1 U9846 ( .B1(n13647), .B2(n7176), .A(n13531), .ZN(n7175) );
  NAND2_X1 U9847 ( .A1(n7178), .A2(n7180), .ZN(n13630) );
  NAND2_X1 U9848 ( .A1(n7180), .A2(n7181), .ZN(n7179) );
  INV_X1 U9849 ( .A(n13528), .ZN(n7184) );
  OR2_X1 U9850 ( .A1(n11992), .A2(n7189), .ZN(n7185) );
  NAND2_X1 U9851 ( .A1(n7185), .A2(n7186), .ZN(n7345) );
  NAND2_X1 U9852 ( .A1(n13519), .A2(n7196), .ZN(n7193) );
  NAND2_X1 U9853 ( .A1(n7193), .A2(n7194), .ZN(n13527) );
  NAND2_X1 U9854 ( .A1(n11071), .A2(n7200), .ZN(n7335) );
  NAND2_X1 U9855 ( .A1(n7336), .A2(n7335), .ZN(n11377) );
  AND4_X1 U9856 ( .A1(n7847), .A2(n7848), .A3(n7850), .A4(n7204), .ZN(n7881)
         );
  NAND3_X1 U9857 ( .A1(n7847), .A2(n7848), .A3(n7202), .ZN(n13877) );
  NAND3_X1 U9858 ( .A1(n7847), .A2(n7848), .A3(n7204), .ZN(n7879) );
  AND2_X2 U9859 ( .A1(n11152), .A2(n11151), .ZN(n11437) );
  NAND3_X1 U9860 ( .A1(n7213), .A2(n7214), .A3(n7212), .ZN(n10949) );
  NAND3_X1 U9861 ( .A1(n7213), .A2(n6716), .A3(n7212), .ZN(n7216) );
  INV_X1 U9862 ( .A(n7216), .ZN(n11020) );
  INV_X1 U9863 ( .A(n11021), .ZN(n7215) );
  NAND2_X1 U9864 ( .A1(n7221), .A2(n7222), .ZN(n7220) );
  INV_X1 U9865 ( .A(n7224), .ZN(n12809) );
  NAND3_X1 U9866 ( .A1(n7229), .A2(n7228), .A3(n11478), .ZN(n11636) );
  NAND3_X1 U9867 ( .A1(n11544), .A2(n7594), .A3(n7595), .ZN(n7228) );
  NAND3_X1 U9868 ( .A1(n11544), .A2(n7594), .A3(n11533), .ZN(n7229) );
  NAND2_X2 U9869 ( .A1(n9560), .A2(n9559), .ZN(n15020) );
  NOR2_X2 U9870 ( .A1(n11688), .A2(n11860), .ZN(n7232) );
  OR2_X2 U9871 ( .A1(n12725), .A2(n12724), .ZN(n12752) );
  AND2_X1 U9872 ( .A1(n12825), .A2(n12824), .ZN(n7255) );
  NAND2_X1 U9873 ( .A1(n7257), .A2(n12699), .ZN(n10843) );
  INV_X4 U9874 ( .A(n10123), .ZN(n10154) );
  MUX2_X1 U9875 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n10123), .Z(n7261) );
  NAND2_X1 U9876 ( .A1(n8238), .A2(n8237), .ZN(n8258) );
  NAND2_X1 U9877 ( .A1(n10782), .A2(n10781), .ZN(n10784) );
  XNOR2_X2 U9878 ( .A(n11943), .B(n11951), .ZN(n11716) );
  NAND2_X1 U9879 ( .A1(n15000), .A2(n14999), .ZN(n14998) );
  NOR2_X2 U9880 ( .A1(n15922), .A2(n14767), .ZN(n14769) );
  NAND2_X1 U9881 ( .A1(n12150), .A2(n7298), .ZN(n7297) );
  NAND2_X1 U9882 ( .A1(n13023), .A2(n7322), .ZN(n7321) );
  NAND2_X1 U9883 ( .A1(n7326), .A2(n7324), .ZN(n9166) );
  INV_X1 U9884 ( .A(n9341), .ZN(n7329) );
  INV_X1 U9885 ( .A(n13049), .ZN(n7332) );
  INV_X1 U9886 ( .A(n11761), .ZN(n7341) );
  NAND2_X1 U9887 ( .A1(n7342), .A2(n6800), .ZN(n13515) );
  INV_X2 U9888 ( .A(n7862), .ZN(n7847) );
  NAND2_X1 U9889 ( .A1(n7848), .A2(n7344), .ZN(n7343) );
  NOR2_X1 U9890 ( .A1(n7862), .A2(n7750), .ZN(n7344) );
  AND3_X2 U9891 ( .A1(n7841), .A2(n8613), .A3(n7840), .ZN(n7848) );
  NAND2_X1 U9892 ( .A1(n7345), .A2(n12199), .ZN(n12363) );
  NAND2_X1 U9893 ( .A1(n10153), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7348) );
  OAI21_X1 U9894 ( .B1(n10181), .B2(n10153), .A(n7348), .ZN(n7349) );
  NAND2_X2 U9895 ( .A1(n12458), .A2(n8626), .ZN(n7993) );
  OAI21_X2 U9896 ( .B1(n11886), .B2(n7355), .A(n7354), .ZN(n12214) );
  NAND2_X1 U9897 ( .A1(n14108), .A2(n6706), .ZN(n7361) );
  NAND2_X1 U9898 ( .A1(n11409), .A2(n7375), .ZN(n7372) );
  INV_X1 U9899 ( .A(n11276), .ZN(n7379) );
  NOR2_X1 U9900 ( .A1(n14019), .A2(n7379), .ZN(n7378) );
  NAND3_X1 U9901 ( .A1(n14042), .A2(n15205), .A3(n14182), .ZN(n7388) );
  NAND2_X1 U9902 ( .A1(n8728), .A2(n8727), .ZN(n7391) );
  NAND2_X1 U9903 ( .A1(n8706), .A2(n8705), .ZN(n7392) );
  NAND2_X1 U9904 ( .A1(n8905), .A2(n7400), .ZN(n7397) );
  NAND2_X1 U9905 ( .A1(n8884), .A2(n8883), .ZN(n8887) );
  OAI21_X2 U9906 ( .B1(n9104), .B2(n9103), .A(n9105), .ZN(n9119) );
  NAND2_X1 U9907 ( .A1(n10872), .A2(n7419), .ZN(n10994) );
  OAI21_X1 U9908 ( .B1(n12663), .B2(n12664), .A(n7434), .ZN(n12569) );
  NAND2_X1 U9909 ( .A1(n7421), .A2(n7420), .ZN(n7431) );
  NAND3_X1 U9910 ( .A1(n12663), .A2(n12570), .A3(n7427), .ZN(n7420) );
  INV_X1 U9911 ( .A(n7422), .ZN(n7421) );
  OAI21_X1 U9912 ( .B1(n12663), .B2(n7426), .A(n7423), .ZN(n7422) );
  NAND3_X1 U9913 ( .A1(n7427), .A2(n12570), .A3(n7429), .ZN(n7425) );
  NAND2_X1 U9914 ( .A1(n7431), .A2(n12575), .ZN(P3_U3160) );
  OR2_X1 U9915 ( .A1(n12533), .A2(n12898), .ZN(n7434) );
  NAND3_X1 U9916 ( .A1(n7449), .A2(n7450), .A3(n7447), .ZN(n12347) );
  NAND2_X1 U9917 ( .A1(n12312), .A2(n12311), .ZN(n12402) );
  INV_X1 U9918 ( .A(n12223), .ZN(n12221) );
  NAND2_X1 U9919 ( .A1(n10780), .A2(n10667), .ZN(n7466) );
  XNOR2_X2 U9920 ( .A(n8680), .B(n8679), .ZN(n10780) );
  OAI21_X1 U9921 ( .B1(n10780), .B2(n10667), .A(n7466), .ZN(n10682) );
  NAND2_X1 U9922 ( .A1(n10681), .A2(n10682), .ZN(n10751) );
  NAND2_X1 U9923 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  NAND2_X1 U9924 ( .A1(n11495), .A2(n7482), .ZN(n7484) );
  NOR2_X1 U9925 ( .A1(n7483), .A2(n9611), .ZN(n7482) );
  NAND2_X1 U9926 ( .A1(n7484), .A2(n7485), .ZN(n11628) );
  NAND2_X1 U9927 ( .A1(n9561), .A2(n9543), .ZN(n10096) );
  INV_X1 U9928 ( .A(n7509), .ZN(n9956) );
  AOI21_X1 U9929 ( .B1(n9972), .B2(n7517), .A(n7515), .ZN(n7514) );
  NAND3_X1 U9930 ( .A1(n7524), .A2(n7526), .A3(n7525), .ZN(n7520) );
  NAND2_X1 U9931 ( .A1(n7533), .A2(n7534), .ZN(n9896) );
  AND2_X1 U9932 ( .A1(n14507), .A2(n9871), .ZN(n7538) );
  INV_X1 U9933 ( .A(n9726), .ZN(n9729) );
  NAND3_X1 U9934 ( .A1(n9731), .A2(n9730), .A3(n6808), .ZN(n7540) );
  NAND2_X1 U9935 ( .A1(n7540), .A2(n7541), .ZN(n9762) );
  NAND3_X1 U9936 ( .A1(n10112), .A2(n9385), .A3(n10652), .ZN(n7548) );
  NAND2_X1 U9937 ( .A1(n13323), .A2(n9445), .ZN(n7549) );
  NAND2_X1 U9938 ( .A1(n7865), .A2(n7864), .ZN(n8175) );
  NAND2_X1 U9939 ( .A1(n8615), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U9940 ( .A1(n13334), .A2(n7574), .ZN(n7573) );
  OAI211_X1 U9941 ( .C1(n13334), .C2(n7577), .A(n7575), .B(n7573), .ZN(n9512)
         );
  NOR2_X1 U9942 ( .A1(n14297), .A2(n7597), .ZN(n7596) );
  XNOR2_X1 U9943 ( .A(n7598), .B(n14563), .ZN(n14659) );
  NAND4_X2 U9945 ( .A1(n9573), .A2(n9574), .A3(n9575), .A4(n9576), .ZN(n11661)
         );
  NAND2_X1 U9946 ( .A1(n11661), .A2(n15142), .ZN(n10053) );
  NAND2_X1 U9947 ( .A1(n14398), .A2(n14397), .ZN(n14396) );
  NAND2_X1 U9948 ( .A1(n9561), .A2(n7608), .ZN(n9545) );
  INV_X1 U9949 ( .A(n8457), .ZN(n7616) );
  NAND2_X1 U9950 ( .A1(n7869), .A2(n7624), .ZN(n8572) );
  NAND2_X1 U9951 ( .A1(n7869), .A2(n7618), .ZN(n7617) );
  NAND2_X1 U9952 ( .A1(n7625), .A2(n7626), .ZN(n8160) );
  OAI21_X1 U9953 ( .B1(n8211), .B2(n6705), .A(n7644), .ZN(n8233) );
  INV_X1 U9954 ( .A(n7639), .ZN(n8235) );
  AOI21_X1 U9955 ( .B1(n8211), .B2(n7642), .A(n7640), .ZN(n7639) );
  INV_X1 U9956 ( .A(n8232), .ZN(n7643) );
  INV_X1 U9957 ( .A(n8212), .ZN(n7646) );
  NAND2_X1 U9958 ( .A1(n8257), .A2(n7650), .ZN(n7649) );
  INV_X1 U9959 ( .A(n8255), .ZN(n7653) );
  NAND2_X1 U9960 ( .A1(n7654), .A2(n6805), .ZN(n7659) );
  NAND2_X1 U9961 ( .A1(n8088), .A2(n7678), .ZN(n7677) );
  INV_X1 U9962 ( .A(n8067), .ZN(n7681) );
  XNOR2_X1 U9963 ( .A(n7682), .B(n8514), .ZN(n12457) );
  AOI21_X1 U9964 ( .B1(n10901), .B2(n7725), .A(n6747), .ZN(n7723) );
  OAI21_X1 U9965 ( .B1(n11757), .B2(n6734), .A(n7732), .ZN(n11989) );
  NAND2_X1 U9966 ( .A1(n8424), .A2(n8425), .ZN(n7740) );
  NAND2_X1 U9967 ( .A1(n8198), .A2(n8213), .ZN(n8215) );
  NAND2_X1 U9968 ( .A1(n7741), .A2(n6795), .ZN(n8213) );
  NAND2_X1 U9969 ( .A1(n7741), .A2(n8194), .ZN(n8197) );
  INV_X1 U9970 ( .A(n7754), .ZN(n7753) );
  NAND2_X1 U9971 ( .A1(n12894), .A2(n12893), .ZN(n12967) );
  INV_X1 U9972 ( .A(n12893), .ZN(n7771) );
  NAND3_X1 U9973 ( .A1(n7460), .A2(n7791), .A3(n7790), .ZN(n7789) );
  NAND2_X1 U9974 ( .A1(n9916), .A2(n9915), .ZN(n9917) );
  OAI21_X1 U9975 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9850) );
  NAND2_X1 U9976 ( .A1(n9545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9547) );
  AND2_X1 U9977 ( .A1(n7951), .A2(n7987), .ZN(n10137) );
  OR2_X1 U9978 ( .A1(n11295), .A2(n9014), .ZN(n9016) );
  NAND2_X1 U9979 ( .A1(n7879), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7851) );
  OR2_X1 U9980 ( .A1(n6688), .A2(n10280), .ZN(n9586) );
  AND2_X2 U9981 ( .A1(n7885), .A2(n12461), .ZN(n7960) );
  AND2_X1 U9982 ( .A1(n9584), .A2(n9583), .ZN(n7793) );
  NOR2_X1 U9983 ( .A1(n10081), .A2(n10080), .ZN(n7794) );
  INV_X1 U9984 ( .A(n7885), .ZN(n13885) );
  XOR2_X1 U9985 ( .A(n6822), .B(n12182), .Z(n7795) );
  OR2_X1 U9986 ( .A1(n12465), .A2(n8569), .ZN(n7796) );
  INV_X1 U9987 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8790) );
  INV_X1 U9988 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8720) );
  INV_X1 U9989 ( .A(n11563), .ZN(n9352) );
  AND2_X1 U9990 ( .A1(n8237), .A2(n8218), .ZN(n7797) );
  INV_X1 U9991 ( .A(n12142), .ZN(n10089) );
  AND2_X1 U9992 ( .A1(n11227), .A2(n11695), .ZN(n7798) );
  AND3_X1 U9993 ( .A1(n8606), .A2(n8605), .A3(n12465), .ZN(n7799) );
  AND2_X1 U9994 ( .A1(n8259), .A2(n8241), .ZN(n7800) );
  AND2_X1 U9995 ( .A1(n8550), .A2(n8549), .ZN(n7802) );
  AND4_X1 U9996 ( .A1(n8881), .A2(n8880), .A3(n8879), .A4(n8878), .ZN(n12871)
         );
  INV_X1 U9997 ( .A(n11529), .ZN(n9609) );
  AND2_X1 U9998 ( .A1(n10428), .A2(n9369), .ZN(n7920) );
  NOR2_X1 U9999 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  INV_X1 U10000 ( .A(n7911), .ZN(n7908) );
  OAI21_X1 U10001 ( .B1(n11240), .B2(n8525), .A(n8021), .ZN(n8022) );
  INV_X1 U10002 ( .A(n8086), .ZN(n8088) );
  OAI22_X1 U10003 ( .A1(n13550), .A2(n8545), .B1(n13549), .B2(n6692), .ZN(
        n8278) );
  OAI22_X1 U10004 ( .A1(n13744), .A2(n8545), .B1(n13553), .B2(n6692), .ZN(
        n8303) );
  NAND2_X1 U10005 ( .A1(n8320), .A2(n8317), .ZN(n8321) );
  OAI22_X1 U10006 ( .A1(n13816), .A2(n8545), .B1(n13556), .B2(n6692), .ZN(
        n8345) );
  OAI22_X1 U10007 ( .A1(n13865), .A2(n8545), .B1(n13561), .B2(n6692), .ZN(
        n8411) );
  INV_X1 U10008 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9532) );
  INV_X1 U10009 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9535) );
  AND2_X1 U10010 ( .A1(n13183), .A2(n9346), .ZN(n9164) );
  INV_X1 U10011 ( .A(n9019), .ZN(n9018) );
  NAND3_X1 U10012 ( .A1(n8368), .A2(n8367), .A3(n8366), .ZN(n8370) );
  INV_X1 U10013 ( .A(n8913), .ZN(n8912) );
  OR2_X1 U10014 ( .A1(n9095), .A2(n9094), .ZN(n9110) );
  NAND2_X1 U10015 ( .A1(n9018), .A2(n9017), .ZN(n9027) );
  INV_X1 U10016 ( .A(n13020), .ZN(n9006) );
  INV_X1 U10017 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7803) );
  INV_X1 U10018 ( .A(n8297), .ZN(n8295) );
  INV_X1 U10019 ( .A(n8431), .ZN(n8430) );
  INV_X1 U10020 ( .A(n8383), .ZN(n8382) );
  INV_X1 U10021 ( .A(n10428), .ZN(n7919) );
  INV_X1 U10022 ( .A(n9767), .ZN(n9765) );
  NOR2_X1 U10023 ( .A1(n9839), .A2(n14091), .ZN(n9827) );
  INV_X1 U10024 ( .A(n15397), .ZN(n12113) );
  INV_X1 U10025 ( .A(n8987), .ZN(n8986) );
  OR2_X1 U10026 ( .A1(n9039), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9055) );
  OR2_X1 U10027 ( .A1(n9123), .A2(n8670), .ZN(n8674) );
  INV_X1 U10028 ( .A(n12891), .ZN(n12982) );
  INV_X1 U10029 ( .A(n12878), .ZN(n13066) );
  NAND2_X1 U10030 ( .A1(n8874), .A2(n8873), .ZN(n8892) );
  OR2_X1 U10031 ( .A1(n8809), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8826) );
  OR2_X1 U10032 ( .A1(n8312), .A2(n8311), .ZN(n8337) );
  INV_X1 U10033 ( .A(n14888), .ZN(n9434) );
  OR2_X1 U10034 ( .A1(n8337), .A2(n13308), .ZN(n8355) );
  AND2_X1 U10035 ( .A1(n8179), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U10036 ( .A1(n8430), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8534) );
  OR2_X1 U10037 ( .A1(n15284), .A2(n13459), .ZN(n15275) );
  AND2_X1 U10038 ( .A1(n8506), .A2(n8505), .ZN(n13594) );
  NAND2_X1 U10039 ( .A1(n8382), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8404) );
  OR2_X1 U10040 ( .A1(n8124), .A2(n8123), .ZN(n8152) );
  INV_X1 U10041 ( .A(n11378), .ZN(n11501) );
  INV_X1 U10042 ( .A(n9884), .ZN(n9883) );
  INV_X1 U10043 ( .A(n12224), .ZN(n12220) );
  OR2_X1 U10044 ( .A1(n9989), .A2(n9988), .ZN(n14355) );
  NAND2_X1 U10045 ( .A1(n9960), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9989) );
  OR2_X1 U10046 ( .A1(n9853), .A2(n9852), .ZN(n9874) );
  INV_X1 U10047 ( .A(n14507), .ZN(n14332) );
  OR2_X1 U10048 ( .A1(n9750), .A2(n9749), .ZN(n9767) );
  INV_X1 U10049 ( .A(n14511), .ZN(n14448) );
  NAND2_X1 U10050 ( .A1(n8197), .A2(SI_14_), .ZN(n8198) );
  NOR2_X1 U10051 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14748), .ZN(n14722) );
  NAND2_X1 U10052 ( .A1(n8986), .A2(n8985), .ZN(n9000) );
  NAND2_X1 U10053 ( .A1(n9054), .A2(n15847), .ZN(n9069) );
  OR2_X1 U10054 ( .A1(n8965), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8987) );
  OR2_X1 U10055 ( .A1(n13235), .A2(n10627), .ZN(n10920) );
  AND4_X1 U10056 ( .A1(n8937), .A2(n8936), .A3(n8935), .A4(n8934), .ZN(n13062)
         );
  INV_X1 U10057 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15894) );
  INV_X1 U10058 ( .A(n15392), .ZN(n12813) );
  AND2_X1 U10059 ( .A1(n9101), .A2(n9100), .ZN(n12943) );
  INV_X1 U10060 ( .A(n12898), .ZN(n12956) );
  AND3_X1 U10061 ( .A1(n8991), .A2(n8990), .A3(n8989), .ZN(n13051) );
  INV_X1 U10062 ( .A(n13087), .ZN(n12876) );
  OR2_X1 U10063 ( .A1(n8892), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8913) );
  AND2_X1 U10064 ( .A1(n8769), .A2(n11027), .ZN(n8791) );
  INV_X1 U10065 ( .A(n15438), .ZN(n15455) );
  INV_X1 U10066 ( .A(n13115), .ZN(n10819) );
  INV_X1 U10067 ( .A(n15453), .ZN(n15430) );
  AND2_X1 U10068 ( .A1(n8836), .A2(n8817), .ZN(n8818) );
  AND2_X1 U10069 ( .A1(n8202), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8223) );
  INV_X1 U10070 ( .A(n11857), .ZN(n9413) );
  OR2_X1 U10071 ( .A1(n11142), .A2(n11140), .ZN(n13458) );
  OR2_X1 U10072 ( .A1(n8404), .A2(n13264), .ZN(n8431) );
  INV_X1 U10073 ( .A(n13744), .ZN(n13828) );
  OR2_X1 U10074 ( .A1(n9919), .A2(n14015), .ZN(n9934) );
  NAND2_X1 U10075 ( .A1(n9883), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U10076 ( .A1(n15143), .A2(n14448), .ZN(n10733) );
  AND2_X1 U10077 ( .A1(n9990), .A2(n14355), .ZN(n14371) );
  OR2_X1 U10078 ( .A1(n9874), .A2(n14111), .ZN(n9884) );
  INV_X1 U10079 ( .A(n14156), .ZN(n14281) );
  NAND2_X1 U10080 ( .A1(n11454), .A2(n11453), .ZN(n15094) );
  INV_X1 U10081 ( .A(n14317), .ZN(n14397) );
  INV_X1 U10082 ( .A(n14521), .ZN(n14357) );
  AND2_X1 U10083 ( .A1(n9045), .A2(n9044), .ZN(n12997) );
  OR2_X1 U10084 ( .A1(n11058), .A2(n9352), .ZN(n12666) );
  OR2_X1 U10085 ( .A1(n12860), .A2(n9123), .ZN(n9158) );
  INV_X1 U10086 ( .A(n12851), .ZN(n12822) );
  INV_X1 U10087 ( .A(n12871), .ZN(n14856) );
  INV_X1 U10088 ( .A(n11774), .ZN(n15419) );
  NAND2_X1 U10089 ( .A1(n10983), .A2(n15455), .ZN(n15458) );
  INV_X1 U10090 ( .A(n15512), .ZN(n15495) );
  AND2_X1 U10091 ( .A1(n10823), .A2(n10822), .ZN(n10824) );
  INV_X1 U10092 ( .A(n15466), .ZN(n15515) );
  INV_X1 U10093 ( .A(n13122), .ZN(n15509) );
  INV_X1 U10094 ( .A(n15450), .ZN(n15398) );
  INV_X1 U10095 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8693) );
  INV_X1 U10096 ( .A(n13725), .ZN(n13822) );
  NAND2_X1 U10097 ( .A1(n8268), .A2(n8267), .ZN(n8297) );
  INV_X1 U10098 ( .A(n13339), .ZN(n14905) );
  AND2_X1 U10099 ( .A1(n9518), .A2(n9509), .ZN(n14903) );
  INV_X1 U10100 ( .A(n8628), .ZN(n8629) );
  AND2_X1 U10101 ( .A1(n8438), .A2(n8437), .ZN(n13288) );
  AND2_X1 U10102 ( .A1(n10342), .A2(n10341), .ZN(n15306) );
  AND2_X1 U10103 ( .A1(n10190), .A2(n10189), .ZN(n13806) );
  INV_X1 U10104 ( .A(n14941), .ZN(n13842) );
  AND2_X1 U10105 ( .A1(n9492), .A2(n9491), .ZN(n15332) );
  AND2_X1 U10106 ( .A1(n8618), .A2(n8617), .ZN(n9493) );
  INV_X1 U10107 ( .A(n14133), .ZN(n14159) );
  INV_X1 U10108 ( .A(n15036), .ZN(n15059) );
  INV_X1 U10109 ( .A(n15055), .ZN(n15046) );
  INV_X1 U10110 ( .A(n15192), .ZN(n15213) );
  AND2_X1 U10111 ( .A1(n15187), .A2(n15197), .ZN(n15176) );
  INV_X1 U10112 ( .A(n15176), .ZN(n15218) );
  NOR2_X1 U10113 ( .A1(n11452), .A2(n11454), .ZN(n12303) );
  NOR2_X1 U10114 ( .A1(n10244), .A2(n10176), .ZN(n11453) );
  AND2_X1 U10115 ( .A1(n10506), .A2(n10505), .ZN(n15392) );
  AND2_X1 U10116 ( .A1(n12992), .A2(n12081), .ZN(n15460) );
  OR2_X1 U10117 ( .A1(n15517), .A2(n15512), .ZN(n13229) );
  NAND2_X1 U10118 ( .A1(n10497), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13235) );
  INV_X1 U10119 ( .A(SI_12_), .ZN(n15814) );
  INV_X1 U10120 ( .A(n9525), .ZN(n9526) );
  NOR2_X1 U10121 ( .A1(n7799), .A2(n8629), .ZN(n8630) );
  INV_X1 U10122 ( .A(n13571), .ZN(n13569) );
  INV_X1 U10123 ( .A(n13555), .ZN(n13517) );
  AND2_X1 U10124 ( .A1(n11081), .A2(n13737), .ZN(n14935) );
  CLKBUF_X1 U10125 ( .A(n15360), .Z(n15364) );
  INV_X1 U10126 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11105) );
  INV_X1 U10127 ( .A(n14124), .ZN(n14161) );
  NAND2_X1 U10128 ( .A1(n9996), .A2(n9995), .ZN(n14346) );
  OR2_X1 U10129 ( .A1(n10244), .A2(n10546), .ZN(n14180) );
  OR2_X1 U10130 ( .A1(n15030), .A2(n14197), .ZN(n15064) );
  AND2_X1 U10131 ( .A1(n14431), .A2(n14430), .ZN(n14610) );
  INV_X1 U10132 ( .A(n14532), .ZN(n15096) );
  OR2_X1 U10133 ( .A1(n15108), .A2(n11455), .ZN(n14564) );
  INV_X1 U10134 ( .A(n15221), .ZN(n15219) );
  INV_X1 U10135 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10354) );
  INV_X1 U10136 ( .A(n14180), .ZN(P1_U4016) );
  INV_X1 U10137 ( .A(n7903), .ZN(n7806) );
  INV_X1 U10138 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8659) );
  MUX2_X1 U10139 ( .A(n8659), .B(n8658), .S(n7816), .Z(n7805) );
  INV_X1 U10140 ( .A(SI_0_), .ZN(n10135) );
  NOR2_X1 U10141 ( .A1(n7805), .A2(n10135), .ZN(n7901) );
  INV_X1 U10142 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10129) );
  MUX2_X1 U10143 ( .A(n10129), .B(n10167), .S(n7816), .Z(n7935) );
  INV_X1 U10144 ( .A(SI_2_), .ZN(n10144) );
  NOR2_X1 U10145 ( .A1(n7935), .A2(n10144), .ZN(n7949) );
  INV_X1 U10146 ( .A(n7949), .ZN(n7808) );
  MUX2_X1 U10147 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7816), .Z(n7809) );
  NAND2_X1 U10148 ( .A1(n7808), .A2(n7986), .ZN(n7814) );
  INV_X1 U10149 ( .A(n7935), .ZN(n7810) );
  MUX2_X1 U10150 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7816), .Z(n7811) );
  NAND2_X1 U10151 ( .A1(n7811), .A2(SI_4_), .ZN(n7815) );
  OAI21_X1 U10152 ( .B1(SI_4_), .B2(n7811), .A(n7815), .ZN(n7985) );
  NAND2_X1 U10153 ( .A1(n7988), .A2(n7815), .ZN(n8010) );
  INV_X1 U10154 ( .A(n7816), .ZN(n10123) );
  NAND2_X1 U10155 ( .A1(n8010), .A2(n8009), .ZN(n8012) );
  NAND2_X1 U10156 ( .A1(n8012), .A2(n7817), .ZN(n8031) );
  MUX2_X1 U10157 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10154), .Z(n7818) );
  NAND2_X1 U10158 ( .A1(n7818), .A2(SI_6_), .ZN(n7820) );
  OAI21_X1 U10159 ( .B1(SI_6_), .B2(n7818), .A(n7820), .ZN(n7819) );
  INV_X1 U10160 ( .A(n7819), .ZN(n8030) );
  NAND2_X1 U10161 ( .A1(n8031), .A2(n8030), .ZN(n8033) );
  NAND2_X1 U10162 ( .A1(n8033), .A2(n7820), .ZN(n8050) );
  MUX2_X1 U10163 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10154), .Z(n7821) );
  NAND2_X1 U10164 ( .A1(n7821), .A2(SI_7_), .ZN(n7823) );
  OAI21_X1 U10165 ( .B1(n7821), .B2(SI_7_), .A(n7823), .ZN(n7822) );
  INV_X1 U10166 ( .A(n7822), .ZN(n8049) );
  MUX2_X1 U10167 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10154), .Z(n7824) );
  OAI21_X1 U10168 ( .B1(SI_8_), .B2(n7824), .A(n7826), .ZN(n7825) );
  INV_X1 U10169 ( .A(n7825), .ZN(n8069) );
  MUX2_X1 U10170 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10154), .Z(n7827) );
  OAI21_X1 U10171 ( .B1(SI_9_), .B2(n7827), .A(n7829), .ZN(n7828) );
  INV_X1 U10172 ( .A(n7828), .ZN(n8089) );
  MUX2_X1 U10173 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10154), .Z(n7830) );
  OAI21_X1 U10174 ( .B1(SI_10_), .B2(n7830), .A(n8117), .ZN(n7831) );
  INV_X1 U10175 ( .A(n7831), .ZN(n7832) );
  NOR2_X1 U10176 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n7837) );
  NAND4_X1 U10177 ( .A1(n7837), .A2(n7836), .A3(n7835), .A4(n7834), .ZN(n7866)
         );
  INV_X1 U10178 ( .A(n7866), .ZN(n7841) );
  NAND3_X1 U10179 ( .A1(n7953), .A2(n7095), .A3(n8173), .ZN(n7863) );
  NOR2_X1 U10180 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n7839) );
  NOR2_X1 U10181 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n7838) );
  INV_X1 U10182 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7842) );
  NAND3_X1 U10183 ( .A1(n8014), .A2(n7842), .A3(n8140), .ZN(n8142) );
  NAND2_X1 U10184 ( .A1(n7846), .A2(n8144), .ZN(n7862) );
  XNOR2_X2 U10185 ( .A(n7853), .B(n7852), .ZN(n12458) );
  INV_X2 U10186 ( .A(n7993), .ZN(n8623) );
  INV_X1 U10187 ( .A(n8139), .ZN(n7855) );
  INV_X1 U10188 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U10189 ( .A1(n7855), .A2(n7854), .ZN(n8053) );
  INV_X1 U10190 ( .A(n8053), .ZN(n7857) );
  INV_X1 U10191 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10192 ( .A1(n7857), .A2(n7856), .ZN(n8073) );
  INV_X1 U10193 ( .A(n8093), .ZN(n7859) );
  INV_X1 U10194 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10195 ( .A1(n7859), .A2(n7858), .ZN(n8119) );
  NAND2_X1 U10196 ( .A1(n8119), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7860) );
  XNOR2_X1 U10197 ( .A(n7860), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10564) );
  INV_X2 U10198 ( .A(n7990), .ZN(n8308) );
  AOI22_X1 U10199 ( .A1(n8623), .A2(n10564), .B1(n8308), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n7861) );
  INV_X1 U10200 ( .A(n7862), .ZN(n7865) );
  INV_X1 U10201 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7867) );
  INV_X1 U10202 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7868) );
  INV_X1 U10203 ( .A(n9367), .ZN(n11968) );
  INV_X1 U10204 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7872) );
  INV_X1 U10205 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7873) );
  INV_X1 U10206 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7874) );
  AOI21_X1 U10207 ( .B1(n8262), .B2(n7834), .A(n7874), .ZN(n7875) );
  NAND2_X1 U10208 ( .A1(n7877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7878) );
  XNOR2_X1 U10209 ( .A(n7878), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7913) );
  INV_X1 U10210 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U10211 ( .A1(n8538), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7891) );
  INV_X1 U10212 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11687) );
  OR2_X1 U10213 ( .A1(n8474), .A2(n11687), .ZN(n7890) );
  NAND2_X2 U10214 ( .A1(n7885), .A2(n7884), .ZN(n8155) );
  NAND2_X1 U10215 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8002) );
  NAND2_X1 U10216 ( .A1(n8037), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8058) );
  INV_X1 U10217 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8057) );
  INV_X1 U10218 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8078) );
  INV_X1 U10219 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10220 ( .A1(n8098), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8124) );
  OR2_X1 U10221 ( .A1(n8098), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U10222 ( .A1(n8124), .A2(n7886), .ZN(n11854) );
  OR2_X1 U10223 ( .A1(n8155), .A2(n11854), .ZN(n7889) );
  NAND2_X2 U10224 ( .A1(n13885), .A2(n12461), .ZN(n7914) );
  INV_X1 U10225 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7887) );
  OR2_X1 U10226 ( .A1(n7914), .A2(n7887), .ZN(n7888) );
  OAI22_X1 U10227 ( .A1(n15382), .A2(n8565), .B1(n13354), .B2(n8525), .ZN(
        n8116) );
  INV_X1 U10228 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7892) );
  INV_X1 U10229 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7893) );
  NAND2_X1 U10230 ( .A1(n7960), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U10231 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7899) );
  MUX2_X1 U10232 ( .A(n7899), .B(P2_IR_REG_31__SCAN_IN), .S(n7898), .Z(n7900)
         );
  NAND2_X1 U10233 ( .A1(n7900), .A2(n7939), .ZN(n13368) );
  INV_X1 U10234 ( .A(n7901), .ZN(n7902) );
  NAND2_X1 U10235 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  NAND2_X1 U10236 ( .A1(n7905), .A2(n7904), .ZN(n10181) );
  INV_X1 U10237 ( .A(n7910), .ZN(n7909) );
  NAND2_X1 U10238 ( .A1(n8525), .A2(n8585), .ZN(n7906) );
  NAND2_X1 U10239 ( .A1(n7907), .A2(n7906), .ZN(n7911) );
  NAND2_X1 U10240 ( .A1(n7909), .A2(n7908), .ZN(n7927) );
  NAND2_X1 U10241 ( .A1(n10154), .A2(SI_0_), .ZN(n7912) );
  XNOR2_X1 U10242 ( .A(n7912), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13895) );
  MUX2_X1 U10243 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13895), .S(n7993), .Z(n10428)
         );
  INV_X1 U10244 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n12473) );
  INV_X1 U10245 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n12469) );
  OAI211_X1 U10246 ( .C1(n7919), .C2(n9369), .A(n8582), .B(n7079), .ZN(n7924)
         );
  NAND2_X1 U10247 ( .A1(n8582), .A2(n7919), .ZN(n8583) );
  INV_X1 U10248 ( .A(n9510), .ZN(n15377) );
  AND2_X1 U10249 ( .A1(n11228), .A2(n15377), .ZN(n7921) );
  NAND2_X1 U10250 ( .A1(n8583), .A2(n7922), .ZN(n7923) );
  NAND2_X1 U10251 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U10252 ( .A1(n7927), .A2(n7926), .ZN(n7972) );
  INV_X1 U10253 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7928) );
  INV_X1 U10254 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7929) );
  OR2_X1 U10255 ( .A1(n8155), .A2(n7929), .ZN(n7933) );
  NAND2_X1 U10256 ( .A1(n7960), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7932) );
  INV_X1 U10257 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10305) );
  OR2_X1 U10258 ( .A1(n7930), .A2(n10305), .ZN(n7931) );
  INV_X1 U10259 ( .A(n8565), .ZN(n8456) );
  NAND2_X1 U10260 ( .A1(n13363), .A2(n7079), .ZN(n7944) );
  NAND2_X1 U10261 ( .A1(n7950), .A2(SI_2_), .ZN(n7945) );
  OAI21_X1 U10262 ( .B1(n7950), .B2(SI_2_), .A(n7945), .ZN(n7936) );
  OR2_X1 U10263 ( .A1(n7936), .A2(n7935), .ZN(n7947) );
  NAND2_X1 U10264 ( .A1(n7936), .A2(n7935), .ZN(n7937) );
  AND2_X1 U10265 ( .A1(n7947), .A2(n7937), .ZN(n10128) );
  NAND2_X1 U10266 ( .A1(n10128), .A2(n8530), .ZN(n7942) );
  NAND2_X1 U10267 ( .A1(n7939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7940) );
  XNOR2_X1 U10268 ( .A(n7940), .B(P2_IR_REG_2__SCAN_IN), .ZN(n15239) );
  AOI22_X1 U10269 ( .A1(n8308), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n8623), .B2(
        n15239), .ZN(n7941) );
  NAND2_X1 U10270 ( .A1(n10469), .A2(n7173), .ZN(n7943) );
  NAND2_X1 U10271 ( .A1(n7944), .A2(n7943), .ZN(n7971) );
  NAND3_X1 U10272 ( .A1(n7947), .A2(n7946), .A3(n7945), .ZN(n7951) );
  OAI21_X1 U10273 ( .B1(n7950), .B2(n7949), .A(n7948), .ZN(n7987) );
  NAND2_X1 U10274 ( .A1(n10137), .A2(n8530), .ZN(n7959) );
  NAND2_X1 U10275 ( .A1(n7952), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7954) );
  MUX2_X1 U10276 ( .A(n7954), .B(P2_IR_REG_31__SCAN_IN), .S(n7953), .Z(n7955)
         );
  INV_X1 U10277 ( .A(n7955), .ZN(n7957) );
  AOI22_X1 U10278 ( .A1(n8308), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n13386), 
        .B2(n8623), .ZN(n7958) );
  NAND2_X1 U10279 ( .A1(n7079), .A2(n10580), .ZN(n7967) );
  NAND2_X1 U10280 ( .A1(n7960), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7965) );
  OR2_X1 U10281 ( .A1(n8155), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7964) );
  INV_X1 U10282 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U10283 ( .A1(n8584), .A2(n6693), .ZN(n7966) );
  AND2_X1 U10284 ( .A1(n7967), .A2(n7966), .ZN(n7974) );
  NAND2_X1 U10285 ( .A1(n10580), .A2(n7173), .ZN(n7969) );
  NAND2_X1 U10286 ( .A1(n8584), .A2(n7079), .ZN(n7968) );
  NAND2_X1 U10287 ( .A1(n7969), .A2(n7968), .ZN(n7973) );
  OAI22_X1 U10288 ( .A1(n7972), .A2(n7971), .B1(n7974), .B2(n7973), .ZN(n7977)
         );
  AOI22_X1 U10289 ( .A1(n8565), .A2(n13363), .B1(n7079), .B2(n10469), .ZN(
        n7970) );
  AOI21_X1 U10290 ( .B1(n7972), .B2(n7971), .A(n7970), .ZN(n7976) );
  NAND2_X1 U10291 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  NAND2_X1 U10292 ( .A1(n8538), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7982) );
  INV_X1 U10293 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11199) );
  OR2_X1 U10294 ( .A1(n8474), .A2(n11199), .ZN(n7981) );
  OAI21_X1 U10295 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8002), .ZN(n11200) );
  OR2_X1 U10296 ( .A1(n8155), .A2(n11200), .ZN(n7980) );
  INV_X1 U10297 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7978) );
  NAND2_X1 U10298 ( .A1(n13362), .A2(n7079), .ZN(n7995) );
  NAND2_X1 U10299 ( .A1(n8146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7983) );
  MUX2_X1 U10300 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7983), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7984) );
  NAND2_X1 U10301 ( .A1(n7984), .A2(n8013), .ZN(n15249) );
  NAND3_X1 U10302 ( .A1(n7987), .A2(n7986), .A3(n7985), .ZN(n7989) );
  NAND2_X1 U10303 ( .A1(n7989), .A2(n7988), .ZN(n10155) );
  OR2_X1 U10304 ( .A1(n10155), .A2(n7938), .ZN(n7992) );
  OR2_X1 U10305 ( .A1(n7990), .A2(n10247), .ZN(n7991) );
  OAI211_X1 U10306 ( .C1(n7993), .C2(n15249), .A(n7992), .B(n7991), .ZN(n10899) );
  NAND2_X1 U10307 ( .A1(n10899), .A2(n8565), .ZN(n7994) );
  NAND2_X1 U10308 ( .A1(n7995), .A2(n7994), .ZN(n7998) );
  AOI22_X1 U10309 ( .A1(n8565), .A2(n13362), .B1(n7079), .B2(n10899), .ZN(
        n7996) );
  AOI21_X1 U10310 ( .B1(n7999), .B2(n7998), .A(n7996), .ZN(n7997) );
  INV_X1 U10311 ( .A(n7997), .ZN(n8000) );
  NAND2_X1 U10312 ( .A1(n8000), .A2(n6749), .ZN(n8024) );
  NAND2_X1 U10313 ( .A1(n8538), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8008) );
  INV_X1 U10314 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10329) );
  OR2_X1 U10315 ( .A1(n8474), .A2(n10329), .ZN(n8007) );
  AND2_X1 U10316 ( .A1(n8002), .A2(n8001), .ZN(n8003) );
  OR2_X1 U10317 ( .A1(n8003), .A2(n8037), .ZN(n11239) );
  OR2_X1 U10318 ( .A1(n8155), .A2(n11239), .ZN(n8006) );
  INV_X1 U10319 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8004) );
  OR2_X1 U10320 ( .A1(n7914), .A2(n8004), .ZN(n8005) );
  NAND4_X1 U10321 ( .A1(n8008), .A2(n8007), .A3(n8006), .A4(n8005), .ZN(n13361) );
  NAND2_X1 U10322 ( .A1(n13361), .A2(n8565), .ZN(n8020) );
  OR2_X1 U10323 ( .A1(n8010), .A2(n8009), .ZN(n8011) );
  NAND2_X1 U10324 ( .A1(n8012), .A2(n8011), .ZN(n10157) );
  OR2_X1 U10325 ( .A1(n10157), .A2(n7938), .ZN(n8018) );
  NAND2_X1 U10326 ( .A1(n8013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8015) );
  MUX2_X1 U10327 ( .A(n8015), .B(P2_IR_REG_31__SCAN_IN), .S(n8014), .Z(n8016)
         );
  AOI22_X1 U10328 ( .A1(n8308), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8623), .B2(
        n13399), .ZN(n8017) );
  NAND2_X1 U10329 ( .A1(n8018), .A2(n8017), .ZN(n11084) );
  NAND2_X1 U10330 ( .A1(n8456), .A2(n11084), .ZN(n8019) );
  NAND2_X1 U10331 ( .A1(n8020), .A2(n8019), .ZN(n8025) );
  NAND2_X1 U10332 ( .A1(n8024), .A2(n8025), .ZN(n8023) );
  INV_X1 U10333 ( .A(n11084), .ZN(n11240) );
  NAND2_X1 U10334 ( .A1(n13361), .A2(n8525), .ZN(n8021) );
  NAND2_X1 U10335 ( .A1(n8023), .A2(n8022), .ZN(n8029) );
  INV_X1 U10336 ( .A(n8024), .ZN(n8027) );
  INV_X1 U10337 ( .A(n8025), .ZN(n8026) );
  NAND2_X1 U10338 ( .A1(n8027), .A2(n8026), .ZN(n8028) );
  NAND2_X1 U10339 ( .A1(n8029), .A2(n8028), .ZN(n8048) );
  OR2_X1 U10340 ( .A1(n8031), .A2(n8030), .ZN(n8032) );
  NAND2_X1 U10341 ( .A1(n8033), .A2(n8032), .ZN(n10160) );
  OR2_X1 U10342 ( .A1(n10160), .A2(n7938), .ZN(n8036) );
  NAND2_X1 U10343 ( .A1(n8139), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8034) );
  AOI22_X1 U10344 ( .A1(n8308), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8623), .B2(
        n13410), .ZN(n8035) );
  NAND2_X1 U10345 ( .A1(n11211), .A2(n8565), .ZN(n8045) );
  NAND2_X1 U10346 ( .A1(n8538), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8043) );
  INV_X1 U10347 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11210) );
  OR2_X1 U10348 ( .A1(n8474), .A2(n11210), .ZN(n8042) );
  OR2_X1 U10349 ( .A1(n8037), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10350 ( .A1(n8058), .A2(n8038), .ZN(n11212) );
  OR2_X1 U10351 ( .A1(n8155), .A2(n11212), .ZN(n8041) );
  INV_X1 U10352 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8039) );
  OR2_X1 U10353 ( .A1(n7914), .A2(n8039), .ZN(n8040) );
  NAND4_X1 U10354 ( .A1(n8043), .A2(n8042), .A3(n8041), .A4(n8040), .ZN(n13360) );
  NAND2_X1 U10355 ( .A1(n13360), .A2(n8525), .ZN(n8044) );
  NAND2_X1 U10356 ( .A1(n8045), .A2(n8044), .ZN(n8047) );
  AOI22_X1 U10357 ( .A1(n11211), .A2(n8525), .B1(n8565), .B2(n13360), .ZN(
        n8046) );
  OR2_X1 U10358 ( .A1(n8050), .A2(n8049), .ZN(n8051) );
  NAND2_X1 U10359 ( .A1(n8052), .A2(n8051), .ZN(n10174) );
  OR2_X1 U10360 ( .A1(n10174), .A2(n7938), .ZN(n8056) );
  NAND2_X1 U10361 ( .A1(n8053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8054) );
  XNOR2_X1 U10362 ( .A(n8054), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U10363 ( .A1(n8308), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8623), .B2(
        n13424), .ZN(n8055) );
  NAND2_X2 U10364 ( .A1(n8056), .A2(n8055), .ZN(n11375) );
  NAND2_X1 U10365 ( .A1(n11375), .A2(n8456), .ZN(n8066) );
  NAND2_X1 U10366 ( .A1(n8538), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8064) );
  INV_X1 U10367 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11097) );
  OR2_X1 U10368 ( .A1(n8474), .A2(n11097), .ZN(n8063) );
  NAND2_X1 U10369 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  NAND2_X1 U10370 ( .A1(n8079), .A2(n8059), .ZN(n11125) );
  OR2_X1 U10371 ( .A1(n8155), .A2(n11125), .ZN(n8062) );
  INV_X1 U10372 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8060) );
  OR2_X1 U10373 ( .A1(n7914), .A2(n8060), .ZN(n8061) );
  NAND4_X1 U10374 ( .A1(n8064), .A2(n8063), .A3(n8062), .A4(n8061), .ZN(n13359) );
  NAND2_X1 U10375 ( .A1(n13359), .A2(n8565), .ZN(n8065) );
  AOI22_X1 U10376 ( .A1(n11375), .A2(n8565), .B1(n13359), .B2(n8456), .ZN(
        n8067) );
  OR2_X1 U10377 ( .A1(n8070), .A2(n8069), .ZN(n8071) );
  NAND2_X1 U10378 ( .A1(n8072), .A2(n8071), .ZN(n10168) );
  OR2_X1 U10379 ( .A1(n10168), .A2(n7938), .ZN(n8077) );
  NAND2_X1 U10380 ( .A1(n8073), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8074) );
  MUX2_X1 U10381 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8074), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8075) );
  AOI22_X1 U10382 ( .A1(n8308), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8623), .B2(
        n13438), .ZN(n8076) );
  NAND2_X1 U10383 ( .A1(n8538), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8085) );
  INV_X1 U10384 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11383) );
  OR2_X1 U10385 ( .A1(n8474), .A2(n11383), .ZN(n8084) );
  NAND2_X1 U10386 ( .A1(n8079), .A2(n8078), .ZN(n8080) );
  NAND2_X1 U10387 ( .A1(n8100), .A2(n8080), .ZN(n11399) );
  OR2_X1 U10388 ( .A1(n8155), .A2(n11399), .ZN(n8083) );
  INV_X1 U10389 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8081) );
  OR2_X1 U10390 ( .A1(n7914), .A2(n8081), .ZN(n8082) );
  OAI22_X1 U10391 ( .A1(n11504), .A2(n8525), .B1(n11503), .B2(n8565), .ZN(
        n8087) );
  INV_X1 U10392 ( .A(n11503), .ZN(n13358) );
  AOI22_X1 U10393 ( .A1(n15372), .A2(n8525), .B1(n8565), .B2(n13358), .ZN(
        n8086) );
  INV_X1 U10394 ( .A(n8110), .ZN(n8113) );
  OR2_X1 U10395 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  OR2_X1 U10396 ( .A1(n10172), .A2(n7938), .ZN(n8097) );
  NAND2_X1 U10397 ( .A1(n8093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8094) );
  MUX2_X1 U10398 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8094), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8095) );
  NAND2_X1 U10399 ( .A1(n8095), .A2(n8119), .ZN(n10339) );
  INV_X1 U10400 ( .A(n10339), .ZN(n15259) );
  AOI22_X1 U10401 ( .A1(n8308), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n15259), 
        .B2(n8623), .ZN(n8096) );
  NAND2_X1 U10402 ( .A1(n8538), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8107) );
  INV_X1 U10403 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11515) );
  OR2_X1 U10404 ( .A1(n8474), .A2(n11515), .ZN(n8106) );
  INV_X1 U10405 ( .A(n8098), .ZN(n8102) );
  NAND2_X1 U10406 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  NAND2_X1 U10407 ( .A1(n8102), .A2(n8101), .ZN(n11514) );
  OR2_X1 U10408 ( .A1(n8155), .A2(n11514), .ZN(n8105) );
  INV_X1 U10409 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8103) );
  OR2_X1 U10410 ( .A1(n7914), .A2(n8103), .ZN(n8104) );
  NAND4_X1 U10411 ( .A1(n8107), .A2(n8106), .A3(n8105), .A4(n8104), .ZN(n13357) );
  AOI22_X1 U10412 ( .A1(n11677), .A2(n8545), .B1(n8565), .B2(n13357), .ZN(
        n8109) );
  INV_X1 U10413 ( .A(n8109), .ZN(n8112) );
  INV_X1 U10414 ( .A(n11677), .ZN(n11653) );
  INV_X1 U10415 ( .A(n13357), .ZN(n11684) );
  OAI22_X1 U10416 ( .A1(n11653), .A2(n8545), .B1(n11684), .B2(n8565), .ZN(
        n8108) );
  OAI22_X1 U10417 ( .A1(n15382), .A2(n8525), .B1(n13354), .B2(n8565), .ZN(
        n8114) );
  INV_X1 U10418 ( .A(n8114), .ZN(n8115) );
  MUX2_X1 U10419 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10154), .Z(n8133) );
  XNOR2_X1 U10420 ( .A(n8137), .B(n8136), .ZN(n10234) );
  NAND2_X1 U10421 ( .A1(n10234), .A2(n8530), .ZN(n8122) );
  OAI21_X1 U10422 ( .B1(n8119), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8120) );
  XNOR2_X1 U10423 ( .A(n8120), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U10424 ( .A1(n10831), .A2(n8623), .B1(n8308), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U10425 ( .A1(n8538), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8130) );
  INV_X1 U10426 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11767) );
  OR2_X1 U10427 ( .A1(n8474), .A2(n11767), .ZN(n8129) );
  INV_X1 U10428 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10429 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  NAND2_X1 U10430 ( .A1(n8152), .A2(n8125), .ZN(n11808) );
  OR2_X1 U10431 ( .A1(n8155), .A2(n11808), .ZN(n8128) );
  INV_X1 U10432 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8126) );
  OR2_X1 U10433 ( .A1(n7914), .A2(n8126), .ZN(n8127) );
  NAND4_X1 U10434 ( .A1(n8130), .A2(n8129), .A3(n8128), .A4(n8127), .ZN(n13353) );
  AOI22_X1 U10435 ( .A1(n12064), .A2(n8525), .B1(n8565), .B2(n13353), .ZN(
        n8132) );
  INV_X1 U10436 ( .A(n12064), .ZN(n12066) );
  INV_X1 U10437 ( .A(n13353), .ZN(n11926) );
  OAI22_X1 U10438 ( .A1(n12066), .A2(n8545), .B1(n11926), .B2(n8565), .ZN(
        n8131) );
  INV_X1 U10439 ( .A(n8133), .ZN(n8134) );
  INV_X1 U10440 ( .A(SI_11_), .ZN(n10148) );
  OAI21_X2 U10441 ( .B1(n8137), .B2(n8136), .A(n8135), .ZN(n8167) );
  MUX2_X1 U10442 ( .A(n10354), .B(n10356), .S(n10154), .Z(n8168) );
  XNOR2_X1 U10443 ( .A(n8167), .B(n8166), .ZN(n10353) );
  NAND2_X1 U10444 ( .A1(n10353), .A2(n8530), .ZN(n8149) );
  INV_X1 U10445 ( .A(n8144), .ZN(n8138) );
  OAI21_X1 U10446 ( .B1(n8139), .B2(n8138), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8141) );
  MUX2_X1 U10447 ( .A(n8141), .B(P2_IR_REG_31__SCAN_IN), .S(n8140), .Z(n8147)
         );
  INV_X1 U10448 ( .A(n8142), .ZN(n8143) );
  NAND2_X1 U10449 ( .A1(n8144), .A2(n8143), .ZN(n8145) );
  OR2_X1 U10450 ( .A1(n8146), .A2(n8145), .ZN(n8172) );
  NAND2_X1 U10451 ( .A1(n8147), .A2(n8172), .ZN(n11135) );
  INV_X1 U10452 ( .A(n11135), .ZN(n11132) );
  AOI22_X1 U10453 ( .A1(n8308), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8623), 
        .B2(n11132), .ZN(n8148) );
  NAND2_X1 U10454 ( .A1(n8150), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8159) );
  INV_X1 U10455 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10828) );
  OR2_X1 U10456 ( .A1(n7930), .A2(n10828), .ZN(n8158) );
  INV_X1 U10457 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11935) );
  OR2_X1 U10458 ( .A1(n8474), .A2(n11935), .ZN(n8157) );
  INV_X1 U10459 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8151) );
  INV_X1 U10460 ( .A(n8179), .ZN(n8154) );
  NAND2_X1 U10461 ( .A1(n8152), .A2(n8151), .ZN(n8153) );
  NAND2_X1 U10462 ( .A1(n8154), .A2(n8153), .ZN(n11934) );
  OR2_X1 U10463 ( .A1(n8155), .A2(n11934), .ZN(n8156) );
  OAI22_X1 U10464 ( .A1(n14945), .A2(n8545), .B1(n11996), .B2(n8565), .ZN(
        n8161) );
  NAND2_X1 U10465 ( .A1(n8160), .A2(n8161), .ZN(n8165) );
  OAI22_X1 U10466 ( .A1(n14945), .A2(n8565), .B1(n11996), .B2(n8545), .ZN(
        n8164) );
  INV_X1 U10467 ( .A(n8160), .ZN(n8163) );
  INV_X1 U10468 ( .A(n8161), .ZN(n8162) );
  INV_X1 U10469 ( .A(n8189), .ZN(n8186) );
  NAND2_X1 U10470 ( .A1(n8168), .A2(n15814), .ZN(n8169) );
  MUX2_X1 U10471 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10154), .Z(n8193) );
  INV_X1 U10472 ( .A(SI_13_), .ZN(n10182) );
  XNOR2_X1 U10473 ( .A(n8193), .B(n10182), .ZN(n8171) );
  XNOR2_X1 U10474 ( .A(n8196), .B(n8171), .ZN(n10455) );
  NAND2_X1 U10475 ( .A1(n10455), .A2(n8530), .ZN(n8178) );
  NAND2_X1 U10476 ( .A1(n8172), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8174) );
  MUX2_X1 U10477 ( .A(n8174), .B(P2_IR_REG_31__SCAN_IN), .S(n8173), .Z(n8176)
         );
  NAND2_X1 U10478 ( .A1(n8176), .A2(n8175), .ZN(n11148) );
  INV_X1 U10479 ( .A(n11148), .ZN(n13456) );
  AOI22_X1 U10480 ( .A1(n8308), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8623), 
        .B2(n13456), .ZN(n8177) );
  NAND2_X1 U10481 ( .A1(n8538), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8185) );
  INV_X1 U10482 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11139) );
  OR2_X1 U10483 ( .A1(n8474), .A2(n11139), .ZN(n8184) );
  NOR2_X1 U10484 ( .A1(n8179), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8180) );
  OR2_X1 U10485 ( .A1(n8202), .A2(n8180), .ZN(n12236) );
  OR2_X1 U10486 ( .A1(n8155), .A2(n12236), .ZN(n8183) );
  INV_X1 U10487 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8181) );
  OR2_X1 U10488 ( .A1(n7914), .A2(n8181), .ZN(n8182) );
  OAI22_X1 U10489 ( .A1(n12195), .A2(n6692), .B1(n12477), .B2(n8545), .ZN(
        n8187) );
  NAND2_X1 U10490 ( .A1(n8186), .A2(n8187), .ZN(n8192) );
  OAI22_X1 U10491 ( .A1(n12195), .A2(n8545), .B1(n12477), .B2(n6692), .ZN(
        n8191) );
  INV_X1 U10492 ( .A(n8187), .ZN(n8188) );
  NOR2_X1 U10493 ( .A1(n8193), .A2(SI_13_), .ZN(n8195) );
  NAND2_X1 U10494 ( .A1(n8193), .A2(SI_13_), .ZN(n8194) );
  MUX2_X1 U10495 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10154), .Z(n8214) );
  XNOR2_X1 U10496 ( .A(n8215), .B(n8214), .ZN(n10913) );
  NAND2_X1 U10497 ( .A1(n10913), .A2(n8530), .ZN(n8201) );
  NAND2_X1 U10498 ( .A1(n8175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8199) );
  XNOR2_X1 U10499 ( .A(n8199), .B(P2_IR_REG_14__SCAN_IN), .ZN(n15284) );
  AOI22_X1 U10500 ( .A1(n8308), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8623), 
        .B2(n15284), .ZN(n8200) );
  NOR2_X1 U10501 ( .A1(n8202), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8203) );
  OR2_X1 U10502 ( .A1(n8223), .A2(n8203), .ZN(n12481) );
  INV_X1 U10503 ( .A(n12481), .ZN(n14917) );
  NAND2_X1 U10504 ( .A1(n8537), .A2(n14917), .ZN(n8209) );
  INV_X1 U10505 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8204) );
  OR2_X1 U10506 ( .A1(n8474), .A2(n8204), .ZN(n8208) );
  INV_X1 U10507 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8205) );
  OR2_X1 U10508 ( .A1(n7914), .A2(n8205), .ZN(n8207) );
  INV_X1 U10509 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13448) );
  OR2_X1 U10510 ( .A1(n7930), .A2(n13448), .ZN(n8206) );
  NAND4_X1 U10511 ( .A1(n8209), .A2(n8208), .A3(n8207), .A4(n8206), .ZN(n13350) );
  AOI22_X1 U10512 ( .A1(n14921), .A2(n6692), .B1(n13350), .B2(n8545), .ZN(
        n8210) );
  INV_X1 U10513 ( .A(n14921), .ZN(n14937) );
  INV_X1 U10514 ( .A(n13350), .ZN(n12198) );
  OAI22_X1 U10515 ( .A1(n14937), .A2(n8565), .B1(n12198), .B2(n8545), .ZN(
        n8212) );
  OAI21_X2 U10516 ( .B1(n8215), .B2(n8214), .A(n8213), .ZN(n8236) );
  INV_X1 U10517 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11103) );
  MUX2_X1 U10518 ( .A(n11103), .B(n11105), .S(n10154), .Z(n8216) );
  INV_X1 U10519 ( .A(SI_15_), .ZN(n15875) );
  NAND2_X1 U10520 ( .A1(n8216), .A2(n15875), .ZN(n8237) );
  INV_X1 U10521 ( .A(n8216), .ZN(n8217) );
  NAND2_X1 U10522 ( .A1(n8217), .A2(SI_15_), .ZN(n8218) );
  XNOR2_X1 U10523 ( .A(n8236), .B(n7797), .ZN(n11102) );
  NAND2_X1 U10524 ( .A1(n11102), .A2(n8530), .ZN(n8222) );
  OR2_X1 U10525 ( .A1(n8219), .A2(n7874), .ZN(n8220) );
  XNOR2_X1 U10526 ( .A(n8220), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15293) );
  AOI22_X1 U10527 ( .A1(n8308), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8623), 
        .B2(n15293), .ZN(n8221) );
  NOR2_X1 U10528 ( .A1(n8223), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8224) );
  OR2_X1 U10529 ( .A1(n8268), .A2(n8224), .ZN(n12292) );
  INV_X1 U10530 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8225) );
  OR2_X1 U10531 ( .A1(n7930), .A2(n8225), .ZN(n8228) );
  INV_X1 U10532 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8226) );
  OR2_X1 U10533 ( .A1(n8474), .A2(n8226), .ZN(n8227) );
  AND2_X1 U10534 ( .A1(n8228), .A2(n8227), .ZN(n8230) );
  NAND2_X1 U10535 ( .A1(n8150), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8229) );
  OAI211_X1 U10536 ( .C1(n12292), .C2(n8155), .A(n8230), .B(n8229), .ZN(n13349) );
  AOI22_X1 U10537 ( .A1(n12364), .A2(n8545), .B1(n8565), .B2(n13349), .ZN(
        n8232) );
  INV_X1 U10538 ( .A(n13349), .ZN(n12368) );
  OAI22_X1 U10539 ( .A1(n7703), .A2(n8545), .B1(n12368), .B2(n8565), .ZN(n8231) );
  NAND2_X1 U10540 ( .A1(n8233), .A2(n8232), .ZN(n8234) );
  NAND2_X1 U10541 ( .A1(n8235), .A2(n8234), .ZN(n8257) );
  INV_X1 U10542 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11195) );
  INV_X1 U10543 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11196) );
  MUX2_X1 U10544 ( .A(n11195), .B(n11196), .S(n10154), .Z(n8239) );
  INV_X1 U10545 ( .A(SI_16_), .ZN(n15595) );
  NAND2_X1 U10546 ( .A1(n8239), .A2(n15595), .ZN(n8259) );
  INV_X1 U10547 ( .A(n8239), .ZN(n8240) );
  NAND2_X1 U10548 ( .A1(n8240), .A2(SI_16_), .ZN(n8241) );
  XNOR2_X1 U10549 ( .A(n8258), .B(n7800), .ZN(n11194) );
  NAND2_X1 U10550 ( .A1(n11194), .A2(n8530), .ZN(n8248) );
  NOR2_X1 U10551 ( .A1(n8242), .A2(n7874), .ZN(n8243) );
  MUX2_X1 U10552 ( .A(n7874), .B(n8243), .S(P2_IR_REG_16__SCAN_IN), .Z(n8246)
         );
  INV_X1 U10553 ( .A(n8244), .ZN(n8245) );
  NOR2_X1 U10554 ( .A1(n8246), .A2(n8245), .ZN(n13481) );
  AOI22_X1 U10555 ( .A1(n8308), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8623), 
        .B2(n13481), .ZN(n8247) );
  XNOR2_X1 U10556 ( .A(n8268), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n14896) );
  OR2_X1 U10557 ( .A1(n14896), .A2(n8155), .ZN(n8254) );
  INV_X1 U10558 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8251) );
  NAND2_X1 U10559 ( .A1(n7960), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U10560 ( .A1(n8538), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8249) );
  OAI211_X1 U10561 ( .C1(n7914), .C2(n8251), .A(n8250), .B(n8249), .ZN(n8252)
         );
  INV_X1 U10562 ( .A(n8252), .ZN(n8253) );
  AND2_X1 U10563 ( .A1(n8254), .A2(n8253), .ZN(n12382) );
  OAI22_X1 U10564 ( .A1(n12383), .A2(n8545), .B1(n12382), .B2(n6692), .ZN(
        n8256) );
  INV_X1 U10565 ( .A(n12382), .ZN(n13348) );
  AOI22_X1 U10566 ( .A1(n14893), .A2(n8545), .B1(n8565), .B2(n13348), .ZN(
        n8255) );
  MUX2_X1 U10567 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10154), .Z(n8286) );
  INV_X1 U10568 ( .A(SI_17_), .ZN(n10459) );
  XNOR2_X1 U10569 ( .A(n8286), .B(n10459), .ZN(n8260) );
  XNOR2_X1 U10570 ( .A(n8285), .B(n8260), .ZN(n11310) );
  NAND2_X1 U10571 ( .A1(n11310), .A2(n8530), .ZN(n8266) );
  NAND2_X1 U10572 ( .A1(n8244), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8261) );
  MUX2_X1 U10573 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8261), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8264) );
  INV_X1 U10574 ( .A(n8262), .ZN(n8263) );
  AND2_X1 U10575 ( .A1(n8264), .A2(n8263), .ZN(n15309) );
  AOI22_X1 U10576 ( .A1(n8308), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8623), 
        .B2(n15309), .ZN(n8265) );
  AND2_X1 U10577 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n8267) );
  INV_X1 U10578 ( .A(n8268), .ZN(n8271) );
  INV_X1 U10579 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8270) );
  INV_X1 U10580 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8269) );
  OAI21_X1 U10581 ( .B1(n8271), .B2(n8270), .A(n8269), .ZN(n8272) );
  NAND2_X1 U10582 ( .A1(n8297), .A2(n8272), .ZN(n14910) );
  OR2_X1 U10583 ( .A1(n14910), .A2(n8155), .ZN(n8277) );
  NAND2_X1 U10584 ( .A1(n8150), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U10585 ( .A1(n8538), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8273) );
  AND2_X1 U10586 ( .A1(n8274), .A2(n8273), .ZN(n8276) );
  NAND2_X1 U10587 ( .A1(n7960), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8275) );
  OAI22_X1 U10588 ( .A1(n13550), .A2(n6692), .B1(n13549), .B2(n8545), .ZN(
        n8281) );
  NAND2_X1 U10589 ( .A1(n8279), .A2(n8278), .ZN(n8283) );
  NAND2_X1 U10590 ( .A1(n8283), .A2(n8282), .ZN(n8302) );
  NAND2_X1 U10591 ( .A1(n8286), .A2(SI_17_), .ZN(n8284) );
  INV_X1 U10592 ( .A(n8286), .ZN(n8287) );
  NAND2_X1 U10593 ( .A1(n8287), .A2(n10459), .ZN(n8288) );
  INV_X1 U10594 ( .A(SI_18_), .ZN(n10495) );
  NAND2_X1 U10595 ( .A1(n8329), .A2(n10495), .ZN(n8289) );
  NAND2_X1 U10596 ( .A1(n8305), .A2(n8289), .ZN(n8290) );
  INV_X1 U10597 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11522) );
  INV_X1 U10598 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11521) );
  MUX2_X1 U10599 ( .A(n11522), .B(n11521), .S(n10154), .Z(n8324) );
  NAND2_X1 U10600 ( .A1(n8290), .A2(n8324), .ZN(n8291) );
  NAND2_X1 U10601 ( .A1(n8263), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8292) );
  XNOR2_X1 U10602 ( .A(n8292), .B(P2_IR_REG_18__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U10603 ( .A1(n8308), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8623), 
        .B2(n11520), .ZN(n8293) );
  INV_X1 U10604 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10605 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U10606 ( .A1(n8312), .A2(n8298), .ZN(n13738) );
  OR2_X1 U10607 ( .A1(n13738), .A2(n8155), .ZN(n8301) );
  AOI22_X1 U10608 ( .A1(n8538), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n7960), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U10609 ( .A1(n8150), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8299) );
  OAI22_X1 U10610 ( .A1(n13744), .A2(n8565), .B1(n13553), .B2(n8545), .ZN(
        n8304) );
  NAND2_X1 U10611 ( .A1(n8306), .A2(n8305), .ZN(n8307) );
  MUX2_X1 U10612 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10154), .Z(n8330) );
  XNOR2_X1 U10613 ( .A(n8330), .B(SI_19_), .ZN(n8326) );
  XNOR2_X2 U10614 ( .A(n8307), .B(n8326), .ZN(n11697) );
  NAND2_X1 U10615 ( .A1(n11697), .A2(n8530), .ZN(n8310) );
  AOI22_X1 U10616 ( .A1(n8308), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6686), 
        .B2(n8623), .ZN(n8309) );
  INV_X1 U10617 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8311) );
  NAND2_X1 U10618 ( .A1(n8312), .A2(n8311), .ZN(n8313) );
  NAND2_X1 U10619 ( .A1(n8337), .A2(n8313), .ZN(n13722) );
  OR2_X1 U10620 ( .A1(n13722), .A2(n8155), .ZN(n8316) );
  AOI22_X1 U10621 ( .A1(n8150), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n7960), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10622 ( .A1(n8538), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8314) );
  OAI22_X1 U10623 ( .A1(n13725), .A2(n6692), .B1(n13555), .B2(n8545), .ZN(
        n8319) );
  INV_X1 U10624 ( .A(n8319), .ZN(n8317) );
  OAI22_X1 U10625 ( .A1(n13725), .A2(n8545), .B1(n13555), .B2(n8565), .ZN(
        n8318) );
  NAND2_X1 U10626 ( .A1(n8322), .A2(n8321), .ZN(n8346) );
  INV_X1 U10627 ( .A(n8324), .ZN(n8323) );
  NOR2_X1 U10628 ( .A1(n8323), .A2(SI_18_), .ZN(n8328) );
  NOR2_X1 U10629 ( .A1(n8324), .A2(n10495), .ZN(n8325) );
  NOR2_X1 U10630 ( .A1(n8326), .A2(n8325), .ZN(n8327) );
  INV_X1 U10631 ( .A(n8330), .ZN(n8331) );
  INV_X1 U10632 ( .A(SI_19_), .ZN(n15895) );
  INV_X1 U10633 ( .A(SI_20_), .ZN(n15844) );
  NAND2_X1 U10634 ( .A1(n8332), .A2(n15844), .ZN(n8368) );
  NAND2_X1 U10635 ( .A1(n8372), .A2(n8368), .ZN(n8333) );
  INV_X1 U10636 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11673) );
  INV_X1 U10637 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11696) );
  MUX2_X1 U10638 ( .A(n11673), .B(n11696), .S(n10154), .Z(n8365) );
  NAND2_X1 U10639 ( .A1(n8333), .A2(n8365), .ZN(n8334) );
  OR2_X1 U10640 ( .A1(n7990), .A2(n11696), .ZN(n8335) );
  INV_X1 U10641 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13308) );
  NAND2_X1 U10642 ( .A1(n8337), .A2(n13308), .ZN(n8338) );
  NAND2_X1 U10643 ( .A1(n8355), .A2(n8338), .ZN(n13306) );
  INV_X1 U10644 ( .A(n13306), .ZN(n13708) );
  NAND2_X1 U10645 ( .A1(n13708), .A2(n8537), .ZN(n8344) );
  INV_X1 U10646 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10647 ( .A1(n7960), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10648 ( .A1(n8538), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8339) );
  OAI211_X1 U10649 ( .C1(n8341), .C2(n7914), .A(n8340), .B(n8339), .ZN(n8342)
         );
  INV_X1 U10650 ( .A(n8342), .ZN(n8343) );
  OAI22_X1 U10651 ( .A1(n13816), .A2(n6692), .B1(n13556), .B2(n8545), .ZN(
        n8347) );
  NAND2_X1 U10652 ( .A1(n8348), .A2(n8372), .ZN(n8352) );
  INV_X1 U10653 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11903) );
  INV_X1 U10654 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11902) );
  MUX2_X1 U10655 ( .A(n11903), .B(n11902), .S(n10154), .Z(n8349) );
  INV_X1 U10656 ( .A(SI_21_), .ZN(n11296) );
  NAND2_X1 U10657 ( .A1(n8349), .A2(n11296), .ZN(n8366) );
  INV_X1 U10658 ( .A(n8349), .ZN(n8350) );
  NAND2_X1 U10659 ( .A1(n8350), .A2(SI_21_), .ZN(n8369) );
  NAND2_X1 U10660 ( .A1(n8366), .A2(n8369), .ZN(n8351) );
  NAND2_X1 U10661 ( .A1(n11900), .A2(n8530), .ZN(n8354) );
  OR2_X1 U10662 ( .A1(n7990), .A2(n11902), .ZN(n8353) );
  INV_X1 U10663 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13281) );
  NAND2_X1 U10664 ( .A1(n8355), .A2(n13281), .ZN(n8356) );
  AND2_X1 U10665 ( .A1(n8383), .A2(n8356), .ZN(n13696) );
  NAND2_X1 U10666 ( .A1(n13696), .A2(n8537), .ZN(n8362) );
  INV_X1 U10667 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U10668 ( .A1(n7960), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10669 ( .A1(n8538), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8357) );
  OAI211_X1 U10670 ( .C1(n8359), .C2(n7914), .A(n8358), .B(n8357), .ZN(n8360)
         );
  INV_X1 U10671 ( .A(n8360), .ZN(n8361) );
  NAND2_X1 U10672 ( .A1(n8362), .A2(n8361), .ZN(n13557) );
  AOI22_X1 U10673 ( .A1(n13699), .A2(n8545), .B1(n8565), .B2(n13557), .ZN(
        n8363) );
  INV_X1 U10674 ( .A(n13699), .ZN(n13809) );
  INV_X1 U10675 ( .A(n13557), .ZN(n13523) );
  OAI22_X1 U10676 ( .A1(n13809), .A2(n8545), .B1(n13523), .B2(n8565), .ZN(
        n8364) );
  INV_X1 U10677 ( .A(n8397), .ZN(n8392) );
  INV_X1 U10678 ( .A(n8366), .ZN(n8371) );
  INV_X1 U10679 ( .A(n8365), .ZN(n8367) );
  INV_X1 U10680 ( .A(n8374), .ZN(n8373) );
  INV_X1 U10681 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8376) );
  INV_X1 U10682 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11969) );
  MUX2_X1 U10683 ( .A(n8376), .B(n11969), .S(n10154), .Z(n8378) );
  NAND2_X1 U10684 ( .A1(n9908), .A2(n8378), .ZN(n8379) );
  NAND2_X1 U10685 ( .A1(n8400), .A2(n8379), .ZN(n11967) );
  OR2_X1 U10686 ( .A1(n7990), .A2(n11969), .ZN(n8380) );
  INV_X1 U10687 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13318) );
  NAND2_X1 U10688 ( .A1(n8383), .A2(n13318), .ZN(n8384) );
  NAND2_X1 U10689 ( .A1(n8404), .A2(n8384), .ZN(n13682) );
  OR2_X1 U10690 ( .A1(n13682), .A2(n8155), .ZN(n8390) );
  INV_X1 U10691 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10692 ( .A1(n7960), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10693 ( .A1(n8538), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8385) );
  OAI211_X1 U10694 ( .C1(n7914), .C2(n8387), .A(n8386), .B(n8385), .ZN(n8388)
         );
  INV_X1 U10695 ( .A(n8388), .ZN(n8389) );
  NAND2_X1 U10696 ( .A1(n8390), .A2(n8389), .ZN(n13559) );
  AOI22_X1 U10697 ( .A1(n13802), .A2(n6692), .B1(n13559), .B2(n8545), .ZN(
        n8396) );
  INV_X1 U10698 ( .A(n8396), .ZN(n8391) );
  NAND2_X1 U10699 ( .A1(n8392), .A2(n8391), .ZN(n8395) );
  AOI22_X1 U10700 ( .A1(n13802), .A2(n8545), .B1(n6692), .B2(n13559), .ZN(
        n8393) );
  INV_X1 U10701 ( .A(n8393), .ZN(n8394) );
  NAND2_X1 U10702 ( .A1(n8395), .A2(n8394), .ZN(n8398) );
  NAND2_X1 U10703 ( .A1(n8398), .A2(n6754), .ZN(n8413) );
  MUX2_X1 U10704 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10154), .Z(n8419) );
  XNOR2_X1 U10705 ( .A(n8419), .B(SI_23_), .ZN(n8401) );
  NAND2_X1 U10706 ( .A1(n12146), .A2(n8530), .ZN(n8403) );
  INV_X1 U10707 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12149) );
  OR2_X1 U10708 ( .A1(n7990), .A2(n12149), .ZN(n8402) );
  INV_X1 U10709 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13264) );
  NAND2_X1 U10710 ( .A1(n8404), .A2(n13264), .ZN(n8405) );
  AND2_X1 U10711 ( .A1(n8431), .A2(n8405), .ZN(n13666) );
  NAND2_X1 U10712 ( .A1(n13666), .A2(n8537), .ZN(n8410) );
  INV_X1 U10713 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13862) );
  NAND2_X1 U10714 ( .A1(n7960), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U10715 ( .A1(n8538), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8406) );
  OAI211_X1 U10716 ( .C1(n7914), .C2(n13862), .A(n8407), .B(n8406), .ZN(n8408)
         );
  INV_X1 U10717 ( .A(n8408), .ZN(n8409) );
  NAND2_X1 U10718 ( .A1(n8413), .A2(n8414), .ZN(n8412) );
  NAND2_X1 U10719 ( .A1(n8412), .A2(n8411), .ZN(n8418) );
  INV_X1 U10720 ( .A(n8413), .ZN(n8416) );
  INV_X1 U10721 ( .A(n8414), .ZN(n8415) );
  NAND2_X1 U10722 ( .A1(n8416), .A2(n8415), .ZN(n8417) );
  NAND2_X1 U10723 ( .A1(n8418), .A2(n8417), .ZN(n8442) );
  INV_X1 U10724 ( .A(n8419), .ZN(n8420) );
  INV_X1 U10725 ( .A(SI_23_), .ZN(n15662) );
  NOR2_X1 U10726 ( .A1(n8420), .A2(n15662), .ZN(n8421) );
  INV_X1 U10727 ( .A(SI_24_), .ZN(n15613) );
  MUX2_X1 U10728 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10154), .Z(n8425) );
  INV_X1 U10729 ( .A(n8425), .ZN(n8426) );
  NAND2_X1 U10730 ( .A1(n7739), .A2(n8426), .ZN(n8427) );
  INV_X1 U10731 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12427) );
  OR2_X1 U10732 ( .A1(n7990), .A2(n12427), .ZN(n8428) );
  INV_X1 U10733 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13297) );
  NAND2_X1 U10734 ( .A1(n8431), .A2(n13297), .ZN(n8432) );
  NAND2_X1 U10735 ( .A1(n8534), .A2(n8432), .ZN(n13655) );
  OR2_X1 U10736 ( .A1(n13655), .A2(n8155), .ZN(n8438) );
  INV_X1 U10737 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10738 ( .A1(n7960), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U10739 ( .A1(n8538), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8433) );
  OAI211_X1 U10740 ( .C1(n8435), .C2(n7914), .A(n8434), .B(n8433), .ZN(n8436)
         );
  INV_X1 U10741 ( .A(n8436), .ZN(n8437) );
  NAND2_X1 U10742 ( .A1(n8442), .A2(n8443), .ZN(n8441) );
  AOI22_X1 U10743 ( .A1(n13787), .A2(n8545), .B1(n6692), .B2(n13564), .ZN(
        n8439) );
  INV_X1 U10744 ( .A(n8439), .ZN(n8440) );
  NAND2_X1 U10745 ( .A1(n8441), .A2(n8440), .ZN(n8447) );
  INV_X1 U10746 ( .A(n8442), .ZN(n8445) );
  INV_X1 U10747 ( .A(n8443), .ZN(n8444) );
  NAND2_X1 U10748 ( .A1(n8445), .A2(n8444), .ZN(n8446) );
  MUX2_X1 U10749 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10154), .Z(n8459) );
  XNOR2_X1 U10750 ( .A(n8459), .B(SI_25_), .ZN(n8460) );
  XNOR2_X1 U10751 ( .A(n8461), .B(n8460), .ZN(n13890) );
  NAND2_X1 U10752 ( .A1(n13890), .A2(n8530), .ZN(n8451) );
  INV_X1 U10753 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13893) );
  OR2_X1 U10754 ( .A1(n7990), .A2(n13893), .ZN(n8450) );
  XNOR2_X1 U10755 ( .A(n8534), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n13637) );
  INV_X1 U10756 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U10757 ( .A1(n7960), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10758 ( .A1(n8538), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8452) );
  OAI211_X1 U10759 ( .C1(n7914), .C2(n8454), .A(n8453), .B(n8452), .ZN(n8455)
         );
  AOI21_X1 U10760 ( .B1(n13637), .B2(n8537), .A(n8455), .ZN(n13567) );
  OAI22_X1 U10761 ( .A1(n13639), .A2(n6692), .B1(n13567), .B2(n8545), .ZN(
        n8458) );
  INV_X1 U10762 ( .A(n13567), .ZN(n13532) );
  AOI22_X1 U10763 ( .A1(n13858), .A2(n6693), .B1(n13532), .B2(n8545), .ZN(
        n8457) );
  MUX2_X1 U10764 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10154), .Z(n8462) );
  NAND2_X1 U10765 ( .A1(n8462), .A2(SI_26_), .ZN(n8463) );
  OAI21_X1 U10766 ( .B1(SI_26_), .B2(n8462), .A(n8463), .ZN(n8526) );
  INV_X1 U10767 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14685) );
  INV_X1 U10768 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12459) );
  MUX2_X1 U10769 ( .A(n14685), .B(n12459), .S(n10154), .Z(n8465) );
  INV_X1 U10770 ( .A(SI_27_), .ZN(n12262) );
  NAND2_X1 U10771 ( .A1(n8465), .A2(n12262), .ZN(n8464) );
  INV_X1 U10772 ( .A(n8465), .ZN(n8513) );
  NAND2_X1 U10773 ( .A1(n8513), .A2(SI_27_), .ZN(n8466) );
  MUX2_X1 U10774 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10154), .Z(n8468) );
  XNOR2_X1 U10775 ( .A(n8468), .B(SI_28_), .ZN(n8499) );
  INV_X1 U10776 ( .A(n8468), .ZN(n8469) );
  INV_X1 U10777 ( .A(SI_28_), .ZN(n15799) );
  NAND2_X1 U10778 ( .A1(n8469), .A2(n15799), .ZN(n8470) );
  MUX2_X1 U10779 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n10154), .Z(n8471) );
  INV_X1 U10780 ( .A(SI_29_), .ZN(n15597) );
  XNOR2_X1 U10781 ( .A(n8471), .B(n15597), .ZN(n8483) );
  INV_X1 U10782 ( .A(n8471), .ZN(n8472) );
  MUX2_X1 U10783 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10154), .Z(n8490) );
  INV_X1 U10784 ( .A(SI_30_), .ZN(n13245) );
  XNOR2_X1 U10785 ( .A(n8490), .B(n13245), .ZN(n8489) );
  INV_X1 U10786 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13886) );
  INV_X1 U10787 ( .A(n13504), .ZN(n8576) );
  INV_X1 U10788 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n12455) );
  OR2_X1 U10789 ( .A1(n7930), .A2(n12455), .ZN(n8477) );
  INV_X1 U10790 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8473) );
  OR2_X1 U10791 ( .A1(n8474), .A2(n8473), .ZN(n8476) );
  INV_X1 U10792 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n12452) );
  OR2_X1 U10793 ( .A1(n7914), .A2(n12452), .ZN(n8475) );
  AND3_X1 U10794 ( .A1(n8477), .A2(n8476), .A3(n8475), .ZN(n13543) );
  INV_X1 U10795 ( .A(n13543), .ZN(n13345) );
  AOI22_X1 U10796 ( .A1(n8576), .A2(n8545), .B1(n8565), .B2(n13345), .ZN(n8555) );
  INV_X1 U10797 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13845) );
  NAND2_X1 U10798 ( .A1(n7960), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U10799 ( .A1(n8538), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8478) );
  OAI211_X1 U10800 ( .C1(n7914), .C2(n13845), .A(n8479), .B(n8478), .ZN(n13344) );
  NAND2_X1 U10801 ( .A1(n6686), .A2(n9367), .ZN(n10190) );
  OR2_X1 U10802 ( .A1(n10190), .A2(n10187), .ZN(n8480) );
  NAND2_X1 U10803 ( .A1(n12465), .A2(n11695), .ZN(n9522) );
  NAND3_X1 U10804 ( .A1(n8480), .A2(n10188), .A3(n9522), .ZN(n8481) );
  AOI21_X1 U10805 ( .B1(n13344), .B2(n8545), .A(n8481), .ZN(n8482) );
  OAI22_X1 U10806 ( .A1(n13504), .A2(n8545), .B1(n13543), .B2(n8482), .ZN(
        n8554) );
  INV_X1 U10807 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12460) );
  NAND2_X1 U10808 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n8484) );
  INV_X1 U10809 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13254) );
  NOR2_X1 U10810 ( .A1(n8535), .A2(n13254), .ZN(n8503) );
  AND2_X1 U10811 ( .A1(n8503), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13578) );
  INV_X1 U10812 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U10813 ( .A1(n8538), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10814 ( .A1(n7960), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8485) );
  OAI211_X1 U10815 ( .C1(n8487), .C2(n7914), .A(n8486), .B(n8485), .ZN(n8488)
         );
  AOI21_X1 U10816 ( .B1(n13578), .B2(n8537), .A(n8488), .ZN(n9514) );
  INV_X1 U10817 ( .A(n9514), .ZN(n13346) );
  AOI22_X1 U10818 ( .A1(n13848), .A2(n8545), .B1(n6692), .B2(n13346), .ZN(
        n8551) );
  INV_X1 U10819 ( .A(n8489), .ZN(n8492) );
  NAND2_X1 U10820 ( .A1(n8490), .A2(SI_30_), .ZN(n8491) );
  MUX2_X1 U10821 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10154), .Z(n8494) );
  XNOR2_X1 U10822 ( .A(n8494), .B(SI_31_), .ZN(n8495) );
  INV_X1 U10823 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13879) );
  OR2_X1 U10824 ( .A1(n7990), .A2(n13879), .ZN(n8497) );
  INV_X1 U10825 ( .A(n13344), .ZN(n8498) );
  NAND2_X1 U10826 ( .A1(n13498), .A2(n8498), .ZN(n8566) );
  NAND2_X1 U10827 ( .A1(n12446), .A2(n8530), .ZN(n8502) );
  INV_X1 U10828 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n12464) );
  OR2_X1 U10829 ( .A1(n7990), .A2(n12464), .ZN(n8501) );
  INV_X1 U10830 ( .A(n13578), .ZN(n8506) );
  INV_X1 U10831 ( .A(n8503), .ZN(n8518) );
  INV_X1 U10832 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U10833 ( .A1(n8518), .A2(n8504), .ZN(n8505) );
  NAND2_X1 U10834 ( .A1(n13594), .A2(n8537), .ZN(n8512) );
  INV_X1 U10835 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U10836 ( .A1(n8538), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10837 ( .A1(n7960), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8507) );
  OAI211_X1 U10838 ( .C1(n8509), .C2(n7914), .A(n8508), .B(n8507), .ZN(n8510)
         );
  INV_X1 U10839 ( .A(n8510), .ZN(n8511) );
  AOI22_X1 U10840 ( .A1(n13850), .A2(n8545), .B1(n8565), .B2(n13538), .ZN(
        n8550) );
  OAI22_X1 U10841 ( .A1(n13596), .A2(n8545), .B1(n13545), .B2(n6692), .ZN(
        n8549) );
  XNOR2_X1 U10842 ( .A(n8513), .B(SI_27_), .ZN(n8514) );
  NAND2_X1 U10843 ( .A1(n12457), .A2(n8530), .ZN(n8516) );
  OR2_X1 U10844 ( .A1(n7990), .A2(n12459), .ZN(n8515) );
  NAND2_X1 U10845 ( .A1(n8535), .A2(n13254), .ZN(n8517) );
  NAND2_X1 U10846 ( .A1(n8518), .A2(n8517), .ZN(n13604) );
  OR2_X1 U10847 ( .A1(n13604), .A2(n8155), .ZN(n8524) );
  INV_X1 U10848 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U10849 ( .A1(n8538), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U10850 ( .A1(n7960), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8519) );
  OAI211_X1 U10851 ( .C1(n8521), .C2(n7914), .A(n8520), .B(n8519), .ZN(n8522)
         );
  INV_X1 U10852 ( .A(n8522), .ZN(n8523) );
  OAI22_X1 U10853 ( .A1(n13609), .A2(n8545), .B1(n13573), .B2(n6692), .ZN(
        n8548) );
  AOI22_X1 U10854 ( .A1(n13764), .A2(n8545), .B1(n8565), .B2(n13537), .ZN(
        n8547) );
  NAND2_X1 U10855 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  NAND2_X1 U10856 ( .A1(n13887), .A2(n8530), .ZN(n8532) );
  INV_X1 U10857 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13888) );
  OR2_X1 U10858 ( .A1(n7990), .A2(n13888), .ZN(n8531) );
  INV_X1 U10859 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13289) );
  INV_X1 U10860 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8533) );
  OAI21_X1 U10861 ( .B1(n8534), .B2(n13289), .A(n8533), .ZN(n8536) );
  AND2_X1 U10862 ( .A1(n8536), .A2(n8535), .ZN(n13622) );
  NAND2_X1 U10863 ( .A1(n13622), .A2(n8537), .ZN(n8544) );
  INV_X1 U10864 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U10865 ( .A1(n8538), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U10866 ( .A1(n7960), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8539) );
  OAI211_X1 U10867 ( .C1(n8541), .C2(n7914), .A(n8540), .B(n8539), .ZN(n8542)
         );
  INV_X1 U10868 ( .A(n8542), .ZN(n8543) );
  AOI22_X1 U10869 ( .A1(n13854), .A2(n8545), .B1(n8565), .B2(n13569), .ZN(
        n8559) );
  OAI22_X1 U10870 ( .A1(n13619), .A2(n8545), .B1(n13571), .B2(n6692), .ZN(
        n8558) );
  AOI22_X1 U10871 ( .A1(n8548), .A2(n8547), .B1(n8559), .B2(n8558), .ZN(n8546)
         );
  NOR2_X1 U10872 ( .A1(n8548), .A2(n8547), .ZN(n8562) );
  OAI22_X1 U10873 ( .A1(n8552), .A2(n8551), .B1(n8550), .B2(n8549), .ZN(n8553)
         );
  NOR2_X1 U10874 ( .A1(n8601), .A2(n8553), .ZN(n8556) );
  OAI22_X1 U10875 ( .A1(n8557), .A2(n8556), .B1(n8555), .B2(n8554), .ZN(n8561)
         );
  NAND2_X1 U10876 ( .A1(n6692), .A2(n13344), .ZN(n8564) );
  OAI22_X1 U10877 ( .A1(n8566), .A2(n8565), .B1(n8564), .B2(n13498), .ZN(n8567) );
  INV_X1 U10878 ( .A(n10188), .ZN(n11901) );
  MUX2_X1 U10879 ( .A(n11901), .B(n11968), .S(n11695), .Z(n8569) );
  NAND2_X1 U10880 ( .A1(n12465), .A2(n10188), .ZN(n8570) );
  OAI211_X1 U10881 ( .C1(n9367), .C2(n9369), .A(n9522), .B(n8570), .ZN(n8571)
         );
  OAI21_X1 U10882 ( .B1(n8572), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8574) );
  INV_X1 U10883 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8573) );
  XNOR2_X1 U10884 ( .A(n8574), .B(n8573), .ZN(n8622) );
  INV_X1 U10885 ( .A(n8622), .ZN(n8575) );
  AND2_X1 U10886 ( .A1(n8575), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U10887 ( .A(n8576), .B(n13345), .ZN(n8599) );
  NAND2_X1 U10888 ( .A1(n13850), .A2(n13538), .ZN(n13574) );
  OR2_X1 U10889 ( .A1(n13850), .A2(n13538), .ZN(n8577) );
  NAND2_X1 U10890 ( .A1(n13574), .A2(n8577), .ZN(n13585) );
  NAND2_X1 U10891 ( .A1(n13659), .A2(n13564), .ZN(n8578) );
  NAND2_X1 U10892 ( .A1(n13787), .A2(n13288), .ZN(n13531) );
  NAND2_X1 U10893 ( .A1(n8578), .A2(n13531), .ZN(n13647) );
  XNOR2_X1 U10894 ( .A(n7237), .B(n13561), .ZN(n13668) );
  XNOR2_X1 U10895 ( .A(n13802), .B(n13559), .ZN(n13677) );
  NAND2_X1 U10896 ( .A1(n13711), .A2(n13556), .ZN(n13520) );
  NAND2_X1 U10897 ( .A1(n13521), .A2(n13520), .ZN(n13703) );
  INV_X1 U10898 ( .A(n13553), .ZN(n13513) );
  XNOR2_X1 U10899 ( .A(n13828), .B(n13513), .ZN(n13747) );
  XNOR2_X1 U10900 ( .A(n14893), .B(n12382), .ZN(n12359) );
  XNOR2_X1 U10901 ( .A(n12364), .B(n12368), .ZN(n12200) );
  XNOR2_X1 U10902 ( .A(n14921), .B(n12198), .ZN(n14912) );
  XNOR2_X1 U10903 ( .A(n12242), .B(n12477), .ZN(n11994) );
  INV_X1 U10904 ( .A(n11996), .ZN(n13352) );
  XNOR2_X1 U10905 ( .A(n7230), .B(n13352), .ZN(n11929) );
  NAND2_X1 U10906 ( .A1(n11860), .A2(n13354), .ZN(n11762) );
  OR2_X1 U10907 ( .A1(n11860), .A2(n13354), .ZN(n8579) );
  NAND2_X1 U10908 ( .A1(n11677), .A2(n11684), .ZN(n11680) );
  OR2_X1 U10909 ( .A1(n11677), .A2(n11684), .ZN(n8580) );
  NAND2_X1 U10910 ( .A1(n11680), .A2(n8580), .ZN(n11675) );
  NAND2_X1 U10911 ( .A1(n15372), .A2(n11503), .ZN(n11505) );
  OR2_X1 U10912 ( .A1(n15372), .A2(n11503), .ZN(n8581) );
  OR2_X1 U10913 ( .A1(n8582), .A2(n7919), .ZN(n10258) );
  AND2_X1 U10914 ( .A1(n10258), .A2(n8583), .ZN(n11230) );
  XNOR2_X1 U10915 ( .A(n13362), .B(n10899), .ZN(n10901) );
  XNOR2_X1 U10916 ( .A(n13361), .B(n11084), .ZN(n11070) );
  NAND4_X1 U10917 ( .A1(n11230), .A2(n10187), .A3(n10901), .A4(n11070), .ZN(
        n8587) );
  XNOR2_X1 U10918 ( .A(n8584), .B(n10580), .ZN(n10578) );
  NAND3_X1 U10919 ( .A1(n10578), .A2(n10467), .A3(n10400), .ZN(n8586) );
  NOR2_X1 U10920 ( .A1(n8587), .A2(n8586), .ZN(n8588) );
  XNOR2_X1 U10921 ( .A(n11375), .B(n13359), .ZN(n11087) );
  XNOR2_X1 U10922 ( .A(n11211), .B(n13360), .ZN(n11108) );
  NAND4_X1 U10923 ( .A1(n11378), .A2(n8588), .A3(n11087), .A4(n11108), .ZN(
        n8589) );
  NOR2_X1 U10924 ( .A1(n11675), .A2(n8589), .ZN(n8590) );
  XNOR2_X1 U10925 ( .A(n12064), .B(n13353), .ZN(n11761) );
  NAND4_X1 U10926 ( .A1(n11929), .A2(n11683), .A3(n8590), .A4(n11761), .ZN(
        n8591) );
  OR4_X1 U10927 ( .A1(n12200), .A2(n14912), .A3(n11994), .A4(n8591), .ZN(n8592) );
  NOR2_X1 U10928 ( .A1(n12359), .A2(n8592), .ZN(n8593) );
  INV_X1 U10929 ( .A(n13549), .ZN(n13511) );
  XNOR2_X1 U10930 ( .A(n14907), .B(n13511), .ZN(n13509) );
  NAND3_X1 U10931 ( .A1(n13747), .A2(n8593), .A3(n13509), .ZN(n8594) );
  NOR2_X1 U10932 ( .A1(n13703), .A2(n8594), .ZN(n8595) );
  XNOR2_X1 U10933 ( .A(n13699), .B(n13557), .ZN(n13689) );
  XNOR2_X1 U10934 ( .A(n13822), .B(n13517), .ZN(n13726) );
  NAND4_X1 U10935 ( .A1(n13677), .A2(n8595), .A3(n13689), .A4(n13726), .ZN(
        n8596) );
  NOR3_X1 U10936 ( .A1(n13647), .A2(n13668), .A3(n8596), .ZN(n8597) );
  XNOR2_X1 U10937 ( .A(n13858), .B(n13532), .ZN(n13633) );
  XNOR2_X1 U10938 ( .A(n13854), .B(n13569), .ZN(n13616) );
  AND4_X1 U10939 ( .A1(n13585), .A2(n8597), .A3(n13633), .A4(n13616), .ZN(
        n8598) );
  XNOR2_X1 U10940 ( .A(n13848), .B(n13346), .ZN(n13575) );
  NAND4_X1 U10941 ( .A1(n8599), .A2(n8598), .A3(n13575), .A4(n13611), .ZN(
        n8600) );
  NAND2_X1 U10942 ( .A1(n8607), .A2(n11901), .ZN(n8604) );
  NOR3_X1 U10943 ( .A1(n8606), .A2(n12465), .A3(n8604), .ZN(n8602) );
  INV_X1 U10944 ( .A(n8604), .ZN(n8605) );
  INV_X1 U10945 ( .A(n8607), .ZN(n12147) );
  NAND2_X1 U10946 ( .A1(n8608), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8609) );
  XNOR2_X1 U10947 ( .A(n8609), .B(n7751), .ZN(n13889) );
  INV_X1 U10948 ( .A(n8610), .ZN(n8617) );
  NAND2_X1 U10949 ( .A1(n8617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8611) );
  MUX2_X1 U10950 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8611), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8612) );
  NAND2_X1 U10951 ( .A1(n8612), .A2(n8608), .ZN(n13891) );
  NOR2_X1 U10952 ( .A1(n13889), .A2(n13891), .ZN(n8619) );
  INV_X1 U10953 ( .A(n8613), .ZN(n8614) );
  OAI21_X1 U10954 ( .B1(n8615), .B2(n8614), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8616) );
  MUX2_X1 U10955 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8616), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8618) );
  NAND2_X1 U10956 ( .A1(n8619), .A2(n9493), .ZN(n8620) );
  NAND2_X1 U10957 ( .A1(n8622), .A2(n8620), .ZN(n9520) );
  NAND2_X1 U10958 ( .A1(n9367), .A2(n10188), .ZN(n9519) );
  OR2_X1 U10959 ( .A1(n9520), .A2(n9519), .ZN(n8625) );
  INV_X1 U10960 ( .A(n8620), .ZN(n8621) );
  NAND2_X1 U10961 ( .A1(n8622), .A2(n8621), .ZN(n10110) );
  NAND2_X1 U10962 ( .A1(n10110), .A2(n8623), .ZN(n8624) );
  NAND2_X1 U10963 ( .A1(n8625), .A2(n8624), .ZN(n10317) );
  AND2_X1 U10964 ( .A1(n10317), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15328) );
  INV_X1 U10965 ( .A(n12458), .ZN(n10341) );
  INV_X1 U10966 ( .A(n8626), .ZN(n10320) );
  INV_X1 U10967 ( .A(n9522), .ZN(n9517) );
  NAND4_X1 U10968 ( .A1(n15328), .A2(n10341), .A3(n10320), .A4(n9517), .ZN(
        n8627) );
  OAI211_X1 U10969 ( .C1(n9367), .C2(n12147), .A(n8627), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8628) );
  OAI211_X1 U10970 ( .C1(n8633), .C2(n8632), .A(n8631), .B(n8630), .ZN(
        P2_U3328) );
  NAND4_X1 U10971 ( .A1(n8634), .A2(n8711), .A3(n8746), .A4(n8693), .ZN(n8635)
         );
  NOR2_X1 U10972 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), 
        .ZN(n8637) );
  NAND4_X1 U10973 ( .A1(n8637), .A2(n8636), .A3(n7142), .A4(n8925), .ZN(n9167)
         );
  INV_X1 U10974 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8639) );
  INV_X1 U10975 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8638) );
  NAND4_X1 U10976 ( .A1(n8639), .A2(n8638), .A3(n9169), .A4(n9350), .ZN(n8640)
         );
  INV_X1 U10977 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8644) );
  INV_X1 U10978 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U10979 ( .A1(n8655), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U10980 ( .A1(n9151), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8652) );
  INV_X1 U10981 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11046) );
  OR2_X1 U10982 ( .A1(n9123), .A2(n11046), .ZN(n8651) );
  INV_X1 U10983 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10519) );
  OR2_X1 U10984 ( .A1(n9154), .A2(n10519), .ZN(n8650) );
  INV_X1 U10985 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U10986 ( .A1(n8659), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U10987 ( .A1(n8675), .A2(n8660), .ZN(n10134) );
  NAND2_X1 U10988 ( .A1(n8980), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8661) );
  INV_X1 U10989 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n8662) );
  OR2_X1 U10990 ( .A1(n9139), .A2(n8662), .ZN(n8665) );
  INV_X1 U10991 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15459) );
  INV_X1 U10992 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8663) );
  XNOR2_X1 U10993 ( .A(n8676), .B(n8675), .ZN(n10146) );
  NAND2_X1 U10994 ( .A1(n8666), .A2(SI_1_), .ZN(n8669) );
  NAND2_X1 U10995 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8667) );
  XNOR2_X1 U10996 ( .A(n8667), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U10997 ( .A1(n8980), .A2(n10508), .ZN(n8668) );
  OAI211_X1 U10998 ( .C1(n9014), .C2(n10146), .A(n8669), .B(n8668), .ZN(n15444) );
  INV_X1 U10999 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n8670) );
  INV_X1 U11000 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10667) );
  OR2_X1 U11001 ( .A1(n9139), .A2(n10667), .ZN(n8673) );
  INV_X1 U11002 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U11003 ( .A1(n9138), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11004 ( .A1(n10232), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8677) );
  XNOR2_X1 U11005 ( .A(n8689), .B(n8688), .ZN(n10145) );
  NAND2_X1 U11006 ( .A1(n9148), .A2(n10145), .ZN(n8682) );
  NAND2_X1 U11007 ( .A1(n8980), .A2(n10780), .ZN(n8681) );
  NAND2_X1 U11008 ( .A1(n15451), .A2(n10991), .ZN(n9225) );
  INV_X1 U11009 ( .A(n15451), .ZN(n10423) );
  NAND2_X1 U11010 ( .A1(n15423), .A2(n15429), .ZN(n15422) );
  NAND2_X1 U11011 ( .A1(n9138), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8687) );
  OR2_X1 U11012 ( .A1(n9123), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8686) );
  INV_X1 U11013 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10760) );
  OR2_X1 U11014 ( .A1(n9139), .A2(n10760), .ZN(n8685) );
  INV_X1 U11015 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U11016 ( .A1(n8666), .A2(n7067), .ZN(n8697) );
  NAND2_X1 U11017 ( .A1(n10138), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U11018 ( .A1(n8707), .A2(n8692), .ZN(n8704) );
  XNOR2_X1 U11019 ( .A(n8706), .B(n8704), .ZN(n10142) );
  NAND2_X1 U11020 ( .A1(n9148), .A2(n10142), .ZN(n8696) );
  NAND2_X1 U11021 ( .A1(n8709), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8694) );
  XNOR2_X1 U11022 ( .A(n8694), .B(n8693), .ZN(n10783) );
  NAND2_X1 U11023 ( .A1(n8980), .A2(n10783), .ZN(n8695) );
  NAND2_X1 U11024 ( .A1(n15424), .A2(n11574), .ZN(n9230) );
  INV_X1 U11025 ( .A(n11574), .ZN(n15418) );
  NAND2_X1 U11026 ( .A1(n11575), .A2(n15418), .ZN(n9231) );
  NAND2_X1 U11027 ( .A1(n9230), .A2(n9231), .ZN(n15412) );
  INV_X1 U11028 ( .A(n15412), .ZN(n8698) );
  NAND2_X1 U11029 ( .A1(n9138), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8703) );
  INV_X1 U11030 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10765) );
  OR2_X1 U11031 ( .A1(n9139), .A2(n10765), .ZN(n8702) );
  AND2_X1 U11032 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8699) );
  NOR2_X1 U11033 ( .A1(n8719), .A2(n8699), .ZN(n11569) );
  OR2_X1 U11034 ( .A1(n9123), .A2(n11569), .ZN(n8701) );
  INV_X1 U11035 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10764) );
  INV_X1 U11036 ( .A(SI_4_), .ZN(n15586) );
  NAND2_X1 U11037 ( .A1(n8666), .A2(n15586), .ZN(n8717) );
  INV_X1 U11038 ( .A(n8704), .ZN(n8705) );
  NAND2_X1 U11039 ( .A1(n10131), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11040 ( .A1(n8729), .A2(n8708), .ZN(n8726) );
  XNOR2_X1 U11041 ( .A(n8728), .B(n8726), .ZN(n10143) );
  NAND2_X1 U11042 ( .A1(n9148), .A2(n10143), .ZN(n8716) );
  NOR2_X2 U11043 ( .A1(n8710), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8747) );
  INV_X1 U11044 ( .A(n8747), .ZN(n8714) );
  NAND2_X1 U11045 ( .A1(n8710), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8712) );
  MUX2_X1 U11046 ( .A(n8712), .B(P3_IR_REG_31__SCAN_IN), .S(n8711), .Z(n8713)
         );
  NAND2_X1 U11047 ( .A1(n8980), .A2(n10787), .ZN(n8715) );
  NAND2_X1 U11048 ( .A1(n15408), .A2(n11597), .ZN(n9212) );
  INV_X1 U11049 ( .A(n11597), .ZN(n8718) );
  NAND2_X1 U11050 ( .A1(n11598), .A2(n8718), .ZN(n9236) );
  NAND2_X1 U11051 ( .A1(n9212), .A2(n9236), .ZN(n11595) );
  NAND2_X1 U11052 ( .A1(n9138), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8725) );
  INV_X1 U11053 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11607) );
  OR2_X1 U11054 ( .A1(n9139), .A2(n11607), .ZN(n8724) );
  NAND2_X1 U11055 ( .A1(n8719), .A2(n8720), .ZN(n8735) );
  OR2_X1 U11056 ( .A1(n8720), .A2(n8719), .ZN(n8721) );
  AND2_X1 U11057 ( .A1(n8735), .A2(n8721), .ZN(n11608) );
  OR2_X1 U11058 ( .A1(n9123), .A2(n11608), .ZN(n8723) );
  INV_X1 U11059 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10770) );
  OR2_X1 U11060 ( .A1(n9154), .A2(n10770), .ZN(n8722) );
  INV_X1 U11061 ( .A(SI_5_), .ZN(n15867) );
  NAND2_X1 U11062 ( .A1(n8666), .A2(n15867), .ZN(n8734) );
  NAND2_X1 U11063 ( .A1(n10130), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8730) );
  NAND2_X1 U11064 ( .A1(n8744), .A2(n8730), .ZN(n8741) );
  XNOR2_X1 U11065 ( .A(n8743), .B(n8741), .ZN(n10127) );
  NAND2_X1 U11066 ( .A1(n9148), .A2(n10127), .ZN(n8733) );
  OR2_X1 U11067 ( .A1(n8747), .A2(n8645), .ZN(n8731) );
  XNOR2_X1 U11068 ( .A(n8731), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10894) );
  NAND2_X1 U11069 ( .A1(n8980), .A2(n7463), .ZN(n8732) );
  NAND2_X1 U11070 ( .A1(n11795), .A2(n12612), .ZN(n9213) );
  INV_X1 U11071 ( .A(n11795), .ZN(n10265) );
  INV_X1 U11072 ( .A(n12612), .ZN(n11613) );
  NAND2_X1 U11073 ( .A1(n10265), .A2(n11613), .ZN(n9238) );
  NAND2_X1 U11074 ( .A1(n9138), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8740) );
  INV_X1 U11075 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10963) );
  OR2_X1 U11076 ( .A1(n9139), .A2(n10963), .ZN(n8739) );
  NAND2_X1 U11077 ( .A1(n8735), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8736) );
  AND2_X1 U11078 ( .A1(n8751), .A2(n8736), .ZN(n11787) );
  OR2_X1 U11079 ( .A1(n9123), .A2(n11787), .ZN(n8738) );
  INV_X1 U11080 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10946) );
  OR2_X1 U11081 ( .A1(n9154), .A2(n10946), .ZN(n8737) );
  INV_X1 U11082 ( .A(SI_6_), .ZN(n15843) );
  XNOR2_X1 U11083 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8745) );
  XNOR2_X1 U11084 ( .A(n8758), .B(n8745), .ZN(n10132) );
  NAND2_X1 U11085 ( .A1(n9148), .A2(n10132), .ZN(n8750) );
  NAND2_X1 U11086 ( .A1(n8747), .A2(n8746), .ZN(n8764) );
  NAND2_X1 U11087 ( .A1(n8764), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8748) );
  XNOR2_X1 U11088 ( .A(n8748), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10964) );
  NAND2_X1 U11089 ( .A1(n8980), .A2(n10964), .ZN(n8749) );
  OAI211_X1 U11090 ( .C1(n8833), .C2(n15843), .A(n8750), .B(n8749), .ZN(n11791) );
  NAND2_X1 U11091 ( .A1(n12613), .A2(n11791), .ZN(n9244) );
  INV_X1 U11092 ( .A(n11791), .ZN(n9248) );
  NAND2_X1 U11093 ( .A1(n12104), .A2(n9248), .ZN(n9237) );
  NAND2_X1 U11094 ( .A1(n9244), .A2(n9237), .ZN(n11775) );
  INV_X1 U11095 ( .A(n11775), .ZN(n11772) );
  NAND2_X1 U11096 ( .A1(n9138), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8756) );
  INV_X1 U11097 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10951) );
  OR2_X1 U11098 ( .A1(n9139), .A2(n10951), .ZN(n8755) );
  AND2_X1 U11099 ( .A1(n8751), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8752) );
  NOR2_X1 U11100 ( .A1(n8769), .A2(n8752), .ZN(n12499) );
  OR2_X1 U11101 ( .A1(n9123), .A2(n12499), .ZN(n8754) );
  OR2_X1 U11102 ( .A1(n9154), .A2(n15526), .ZN(n8753) );
  INV_X1 U11103 ( .A(SI_7_), .ZN(n10125) );
  NAND2_X1 U11104 ( .A1(n8666), .A2(n10125), .ZN(n8768) );
  NAND2_X1 U11105 ( .A1(n10141), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U11106 ( .A1(n10161), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U11107 ( .A1(n10150), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11108 ( .A1(n10175), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U11109 ( .A1(n8776), .A2(n8760), .ZN(n8761) );
  NAND2_X1 U11110 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  NAND2_X1 U11111 ( .A1(n8777), .A2(n8763), .ZN(n10126) );
  NAND2_X1 U11112 ( .A1(n9148), .A2(n10126), .ZN(n8767) );
  OAI21_X1 U11113 ( .B1(n8764), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8765) );
  XNOR2_X1 U11114 ( .A(n8765), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11019) );
  INV_X1 U11115 ( .A(n11019), .ZN(n10953) );
  NAND2_X1 U11116 ( .A1(n8980), .A2(n10953), .ZN(n8766) );
  NAND2_X1 U11117 ( .A1(n12107), .A2(n15496), .ZN(n9249) );
  INV_X1 U11118 ( .A(n15496), .ZN(n11621) );
  NAND2_X1 U11119 ( .A1(n15399), .A2(n11621), .ZN(n9250) );
  NAND2_X1 U11120 ( .A1(n9249), .A2(n9250), .ZN(n12070) );
  NAND2_X1 U11121 ( .A1(n9138), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8775) );
  INV_X1 U11122 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11009) );
  OR2_X1 U11123 ( .A1(n9139), .A2(n11009), .ZN(n8774) );
  NOR2_X1 U11124 ( .A1(n8769), .A2(n11027), .ZN(n8770) );
  OR2_X1 U11125 ( .A1(n8791), .A2(n8770), .ZN(n15404) );
  INV_X1 U11126 ( .A(n15404), .ZN(n8771) );
  OR2_X1 U11127 ( .A1(n9123), .A2(n8771), .ZN(n8773) );
  INV_X1 U11128 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11022) );
  OR2_X1 U11129 ( .A1(n9154), .A2(n11022), .ZN(n8772) );
  NAND2_X1 U11130 ( .A1(n10152), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U11131 ( .A1(n10169), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8778) );
  OR2_X1 U11132 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  NAND2_X1 U11133 ( .A1(n8798), .A2(n8781), .ZN(n10140) );
  NAND2_X1 U11134 ( .A1(n8666), .A2(SI_8_), .ZN(n8788) );
  OR2_X1 U11135 ( .A1(n8782), .A2(n8645), .ZN(n8784) );
  MUX2_X1 U11136 ( .A(n8784), .B(P3_IR_REG_31__SCAN_IN), .S(n8783), .Z(n8786)
         );
  NAND2_X1 U11137 ( .A1(n8786), .A2(n8785), .ZN(n11165) );
  INV_X1 U11138 ( .A(n11165), .ZN(n11010) );
  NAND2_X1 U11139 ( .A1(n8980), .A2(n11010), .ZN(n8787) );
  OAI211_X1 U11140 ( .C1(n9014), .C2(n10140), .A(n8788), .B(n8787), .ZN(n12580) );
  NAND2_X1 U11141 ( .A1(n12497), .A2(n12580), .ZN(n9253) );
  INV_X1 U11142 ( .A(n12580), .ZN(n15403) );
  NAND2_X1 U11143 ( .A1(n12110), .A2(n15403), .ZN(n9254) );
  NAND2_X1 U11144 ( .A1(n15393), .A2(n15396), .ZN(n8789) );
  NAND2_X1 U11145 ( .A1(n9138), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8796) );
  INV_X1 U11146 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12158) );
  OR2_X1 U11147 ( .A1(n9139), .A2(n12158), .ZN(n8795) );
  OR2_X1 U11148 ( .A1(n8791), .A2(n8790), .ZN(n8792) );
  AND2_X1 U11149 ( .A1(n8809), .A2(n8792), .ZN(n12129) );
  OR2_X1 U11150 ( .A1(n9123), .A2(n12129), .ZN(n8794) );
  INV_X1 U11151 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11155) );
  OR2_X1 U11152 ( .A1(n9154), .A2(n11155), .ZN(n8793) );
  NAND2_X1 U11153 ( .A1(n10171), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U11154 ( .A1(n10170), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8799) );
  OR2_X1 U11155 ( .A1(n8801), .A2(n8800), .ZN(n8802) );
  NAND2_X1 U11156 ( .A1(n8816), .A2(n8802), .ZN(n10124) );
  NAND2_X1 U11157 ( .A1(n9148), .A2(n10124), .ZN(n8806) );
  INV_X1 U11158 ( .A(SI_9_), .ZN(n15789) );
  NAND2_X1 U11159 ( .A1(n8666), .A2(n15789), .ZN(n8805) );
  NAND2_X1 U11160 ( .A1(n8785), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8803) );
  XNOR2_X1 U11161 ( .A(n8803), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11438) );
  INV_X1 U11162 ( .A(n11438), .ZN(n11157) );
  NAND2_X1 U11163 ( .A1(n8980), .A2(n11157), .ZN(n8804) );
  INV_X1 U11164 ( .A(n12131), .ZN(n12159) );
  NAND2_X1 U11165 ( .A1(n15397), .A2(n12159), .ZN(n8807) );
  NAND2_X1 U11166 ( .A1(n12113), .A2(n12131), .ZN(n8808) );
  NAND2_X1 U11167 ( .A1(n9138), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8814) );
  INV_X1 U11168 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12077) );
  OR2_X1 U11169 ( .A1(n9139), .A2(n12077), .ZN(n8813) );
  NAND2_X1 U11170 ( .A1(n8809), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8810) );
  AND2_X1 U11171 ( .A1(n8826), .A2(n8810), .ZN(n12121) );
  OR2_X1 U11172 ( .A1(n9123), .A2(n12121), .ZN(n8812) );
  INV_X1 U11173 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11440) );
  OR2_X1 U11174 ( .A1(n7003), .A2(n11440), .ZN(n8811) );
  NAND2_X1 U11175 ( .A1(n10184), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U11176 ( .A1(n10186), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8817) );
  OR2_X1 U11177 ( .A1(n8819), .A2(n8818), .ZN(n8820) );
  NAND2_X1 U11178 ( .A1(n8837), .A2(n8820), .ZN(n10147) );
  NAND2_X1 U11179 ( .A1(n9148), .A2(n10147), .ZN(n8825) );
  INV_X1 U11180 ( .A(SI_10_), .ZN(n15823) );
  NAND2_X1 U11181 ( .A1(n8666), .A2(n15823), .ZN(n8824) );
  OR2_X1 U11182 ( .A1(n8785), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U11183 ( .A1(n8834), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8822) );
  XNOR2_X1 U11184 ( .A(n8822), .B(n8821), .ZN(n11727) );
  NAND2_X1 U11185 ( .A1(n8980), .A2(n11727), .ZN(n8823) );
  INV_X1 U11186 ( .A(n12328), .ZN(n15513) );
  NAND2_X1 U11187 ( .A1(n12342), .A2(n15513), .ZN(n9265) );
  NAND2_X1 U11188 ( .A1(n12353), .A2(n12328), .ZN(n9261) );
  NAND2_X1 U11189 ( .A1(n9138), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8832) );
  INV_X1 U11190 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12336) );
  OR2_X1 U11191 ( .A1(n9139), .A2(n12336), .ZN(n8831) );
  NAND2_X1 U11192 ( .A1(n8826), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8827) );
  AND2_X1 U11193 ( .A1(n8856), .A2(n8827), .ZN(n12349) );
  OR2_X1 U11194 ( .A1(n9123), .A2(n12349), .ZN(n8830) );
  INV_X1 U11195 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8828) );
  OR2_X1 U11196 ( .A1(n7003), .A2(n8828), .ZN(n8829) );
  OR2_X1 U11197 ( .A1(n8834), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U11198 ( .A1(n8850), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8835) );
  XNOR2_X1 U11199 ( .A(n8835), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11951) );
  INV_X1 U11200 ( .A(n11951), .ZN(n11957) );
  AOI22_X1 U11201 ( .A1(n8666), .A2(n10148), .B1(n8980), .B2(n11957), .ZN(
        n8843) );
  NAND2_X1 U11202 ( .A1(n10235), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8844) );
  INV_X1 U11203 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U11204 ( .A1(n10237), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8838) );
  OR2_X1 U11205 ( .A1(n8840), .A2(n8839), .ZN(n8841) );
  NAND2_X1 U11206 ( .A1(n8845), .A2(n8841), .ZN(n10149) );
  NAND2_X1 U11207 ( .A1(n10149), .A2(n9148), .ZN(n8842) );
  NAND2_X1 U11208 ( .A1(n12867), .A2(n12355), .ZN(n9263) );
  INV_X1 U11209 ( .A(n12355), .ZN(n12866) );
  NAND2_X1 U11210 ( .A1(n14857), .A2(n12866), .ZN(n9267) );
  NAND2_X1 U11211 ( .A1(n10354), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8863) );
  NAND2_X1 U11212 ( .A1(n10356), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8846) );
  OR2_X1 U11213 ( .A1(n8848), .A2(n8847), .ZN(n8849) );
  NAND2_X1 U11214 ( .A1(n8864), .A2(n8849), .ZN(n10151) );
  OR2_X1 U11215 ( .A1(n10151), .A2(n9014), .ZN(n8855) );
  OAI21_X1 U11216 ( .B1(n8850), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8852) );
  MUX2_X1 U11217 ( .A(n8852), .B(P3_IR_REG_31__SCAN_IN), .S(n8851), .Z(n8853)
         );
  NAND2_X1 U11218 ( .A1(n8853), .A2(n6722), .ZN(n12183) );
  INV_X1 U11219 ( .A(n12183), .ZN(n12173) );
  AOI22_X1 U11220 ( .A1(n8666), .A2(SI_12_), .B1(n8980), .B2(n12173), .ZN(
        n8854) );
  NAND2_X1 U11221 ( .A1(n9151), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8862) );
  AND2_X1 U11222 ( .A1(n8856), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8857) );
  OR2_X1 U11223 ( .A1(n8857), .A2(n8874), .ZN(n14859) );
  INV_X1 U11224 ( .A(n14859), .ZN(n12419) );
  OR2_X1 U11225 ( .A1(n9123), .A2(n12419), .ZN(n8861) );
  INV_X1 U11226 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11946) );
  OR2_X1 U11227 ( .A1(n7003), .A2(n11946), .ZN(n8860) );
  INV_X1 U11228 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8858) );
  OR2_X1 U11229 ( .A1(n7001), .A2(n8858), .ZN(n8859) );
  NAND2_X1 U11230 ( .A1(n14863), .A2(n14844), .ZN(n9275) );
  INV_X1 U11231 ( .A(n14863), .ZN(n12421) );
  NAND2_X1 U11232 ( .A1(n12870), .A2(n12421), .ZN(n9274) );
  INV_X1 U11233 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10457) );
  INV_X1 U11234 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10456) );
  NAND2_X1 U11235 ( .A1(n8866), .A2(n10456), .ZN(n8867) );
  NAND2_X1 U11236 ( .A1(n8884), .A2(n8867), .ZN(n10183) );
  NAND2_X1 U11237 ( .A1(n10183), .A2(n9148), .ZN(n8872) );
  NAND2_X1 U11238 ( .A1(n6722), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8869) );
  MUX2_X1 U11239 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8869), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8870) );
  NAND2_X1 U11240 ( .A1(n9168), .A2(n8870), .ZN(n12714) );
  AOI22_X1 U11241 ( .A1(n8666), .A2(n10182), .B1(n8980), .B2(n12714), .ZN(
        n8871) );
  INV_X1 U11242 ( .A(n14850), .ZN(n8882) );
  NAND2_X1 U11243 ( .A1(n9138), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8881) );
  INV_X1 U11244 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8873) );
  OR2_X1 U11245 ( .A1(n8874), .A2(n8873), .ZN(n8875) );
  AND2_X1 U11246 ( .A1(n8875), .A2(n8892), .ZN(n14847) );
  OR2_X1 U11247 ( .A1(n9123), .A2(n14847), .ZN(n8880) );
  INV_X1 U11248 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8876) );
  OR2_X1 U11249 ( .A1(n9139), .A2(n8876), .ZN(n8879) );
  INV_X1 U11250 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8877) );
  OR2_X1 U11251 ( .A1(n7003), .A2(n8877), .ZN(n8878) );
  NOR2_X1 U11252 ( .A1(n8882), .A2(n14856), .ZN(n9278) );
  INV_X1 U11253 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10916) );
  NAND2_X1 U11254 ( .A1(n10916), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8901) );
  INV_X1 U11255 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10914) );
  NAND2_X1 U11256 ( .A1(n10914), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8885) );
  AND2_X1 U11257 ( .A1(n8901), .A2(n8885), .ZN(n8886) );
  OR2_X1 U11258 ( .A1(n8887), .A2(n8886), .ZN(n8888) );
  NAND2_X1 U11259 ( .A1(n8902), .A2(n8888), .ZN(n10231) );
  NAND2_X1 U11260 ( .A1(n10231), .A2(n9148), .ZN(n8891) );
  INV_X1 U11261 ( .A(SI_14_), .ZN(n15873) );
  OR2_X1 U11262 ( .A1(n8868), .A2(n8645), .ZN(n8889) );
  INV_X1 U11263 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8907) );
  XNOR2_X1 U11264 ( .A(n8889), .B(n8907), .ZN(n12729) );
  AOI22_X1 U11265 ( .A1(n8666), .A2(n15873), .B1(n8980), .B2(n12729), .ZN(
        n8890) );
  NAND2_X1 U11266 ( .A1(n8891), .A2(n8890), .ZN(n14838) );
  NAND2_X1 U11267 ( .A1(n9151), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11268 ( .A1(n8892), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8893) );
  NAND2_X1 U11269 ( .A1(n8913), .A2(n8893), .ZN(n14835) );
  INV_X1 U11270 ( .A(n14835), .ZN(n8894) );
  OR2_X1 U11271 ( .A1(n9123), .A2(n8894), .ZN(n8899) );
  INV_X1 U11272 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n8895) );
  OR2_X1 U11273 ( .A1(n7001), .A2(n8895), .ZN(n8898) );
  INV_X1 U11274 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n8896) );
  OR2_X1 U11275 ( .A1(n7003), .A2(n8896), .ZN(n8897) );
  NAND4_X1 U11276 ( .A1(n8900), .A2(n8899), .A3(n8898), .A4(n8897), .ZN(n14843) );
  NAND2_X1 U11277 ( .A1(n14838), .A2(n14843), .ZN(n9179) );
  INV_X1 U11278 ( .A(n9179), .ZN(n9284) );
  OR2_X1 U11279 ( .A1(n14838), .A2(n14843), .ZN(n9283) );
  NAND2_X1 U11280 ( .A1(n11103), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U11281 ( .A1(n11105), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8903) );
  AND2_X1 U11282 ( .A1(n8919), .A2(n8903), .ZN(n8904) );
  OR2_X1 U11283 ( .A1(n8905), .A2(n8904), .ZN(n8906) );
  NAND2_X1 U11284 ( .A1(n8920), .A2(n8906), .ZN(n10255) );
  NAND2_X1 U11285 ( .A1(n10255), .A2(n9148), .ZN(n8910) );
  OR2_X1 U11286 ( .A1(n8926), .A2(n8645), .ZN(n8908) );
  XNOR2_X1 U11287 ( .A(n8908), .B(n8925), .ZN(n12775) );
  AOI22_X1 U11288 ( .A1(n8666), .A2(n15875), .B1(n8980), .B2(n12775), .ZN(
        n8909) );
  NAND2_X1 U11289 ( .A1(n9138), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8918) );
  INV_X1 U11290 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12755) );
  OR2_X1 U11291 ( .A1(n9139), .A2(n12755), .ZN(n8917) );
  INV_X1 U11292 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U11293 ( .A1(n8913), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8914) );
  AND2_X1 U11294 ( .A1(n8932), .A2(n8914), .ZN(n13101) );
  OR2_X1 U11295 ( .A1(n9123), .A2(n13101), .ZN(n8916) );
  INV_X1 U11296 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12739) );
  OR2_X1 U11297 ( .A1(n7003), .A2(n12739), .ZN(n8915) );
  NAND4_X1 U11298 ( .A1(n8918), .A2(n8917), .A3(n8916), .A4(n8915), .ZN(n14833) );
  NAND2_X1 U11299 ( .A1(n13178), .A2(n14833), .ZN(n9285) );
  NAND2_X1 U11300 ( .A1(n13100), .A2(n9291), .ZN(n13088) );
  NAND2_X1 U11301 ( .A1(n11195), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11302 ( .A1(n11196), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8921) );
  AND2_X1 U11303 ( .A1(n8938), .A2(n8921), .ZN(n8922) );
  OR2_X1 U11304 ( .A1(n8923), .A2(n8922), .ZN(n8924) );
  NAND2_X1 U11305 ( .A1(n8939), .A2(n8924), .ZN(n10302) );
  OR2_X1 U11306 ( .A1(n10302), .A2(n9014), .ZN(n8931) );
  NAND2_X1 U11307 ( .A1(n8928), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8927) );
  MUX2_X1 U11308 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8927), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8929) );
  AND2_X1 U11309 ( .A1(n8929), .A2(n8960), .ZN(n12778) );
  AOI22_X1 U11310 ( .A1(n8666), .A2(SI_16_), .B1(n8980), .B2(n12778), .ZN(
        n8930) );
  NAND2_X1 U11311 ( .A1(n9138), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8937) );
  INV_X1 U11312 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13083) );
  OR2_X1 U11313 ( .A1(n9139), .A2(n13083), .ZN(n8936) );
  NAND2_X1 U11314 ( .A1(n8932), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8933) );
  AND2_X1 U11315 ( .A1(n8948), .A2(n8933), .ZN(n13082) );
  OR2_X1 U11316 ( .A1(n9123), .A2(n13082), .ZN(n8935) );
  INV_X1 U11317 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12768) );
  OR2_X1 U11318 ( .A1(n7003), .A2(n12768), .ZN(n8934) );
  NAND2_X1 U11319 ( .A1(n13174), .A2(n13062), .ZN(n9292) );
  NAND2_X1 U11320 ( .A1(n13086), .A2(n9292), .ZN(n13067) );
  INV_X1 U11321 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11311) );
  NAND2_X1 U11322 ( .A1(n11311), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8954) );
  INV_X1 U11323 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U11324 ( .A1(n11313), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8940) );
  AND2_X1 U11325 ( .A1(n8954), .A2(n8940), .ZN(n8941) );
  OR2_X1 U11326 ( .A1(n8942), .A2(n8941), .ZN(n8943) );
  NAND2_X1 U11327 ( .A1(n8955), .A2(n8943), .ZN(n10460) );
  NAND2_X1 U11328 ( .A1(n10460), .A2(n9148), .ZN(n8946) );
  NAND2_X1 U11329 ( .A1(n8960), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8944) );
  XNOR2_X1 U11330 ( .A(n8944), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12807) );
  INV_X1 U11331 ( .A(n12807), .ZN(n12824) );
  AOI22_X1 U11332 ( .A1(n8666), .A2(n10459), .B1(n8980), .B2(n12824), .ZN(
        n8945) );
  NAND2_X1 U11333 ( .A1(n9138), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8953) );
  INV_X1 U11334 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15625) );
  NAND2_X1 U11335 ( .A1(n8948), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8949) );
  AND2_X1 U11336 ( .A1(n8965), .A2(n8949), .ZN(n13070) );
  OR2_X1 U11337 ( .A1(n9123), .A2(n13070), .ZN(n8952) );
  INV_X1 U11338 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13071) );
  OR2_X1 U11339 ( .A1(n9139), .A2(n13071), .ZN(n8951) );
  INV_X1 U11340 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12792) );
  OR2_X1 U11341 ( .A1(n7003), .A2(n12792), .ZN(n8950) );
  NAND4_X1 U11342 ( .A1(n8953), .A2(n8952), .A3(n8951), .A4(n8950), .ZN(n12656) );
  NAND2_X1 U11343 ( .A1(n13171), .A2(n12656), .ZN(n9301) );
  NAND2_X1 U11344 ( .A1(n9296), .A2(n9301), .ZN(n12878) );
  NAND2_X1 U11345 ( .A1(n13067), .A2(n13066), .ZN(n13069) );
  NAND2_X1 U11346 ( .A1(n11522), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U11347 ( .A1(n11521), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8956) );
  AND2_X1 U11348 ( .A1(n8971), .A2(n8956), .ZN(n8957) );
  OR2_X1 U11349 ( .A1(n8958), .A2(n8957), .ZN(n8959) );
  NAND2_X1 U11350 ( .A1(n8972), .A2(n8959), .ZN(n10496) );
  OR2_X1 U11351 ( .A1(n10496), .A2(n9014), .ZN(n8964) );
  INV_X1 U11352 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U11353 ( .A1(n8977), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8962) );
  XNOR2_X1 U11354 ( .A(n8962), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U11355 ( .A1(n8666), .A2(SI_18_), .B1(n8980), .B2(n12838), .ZN(
        n8963) );
  NAND2_X1 U11356 ( .A1(n8965), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11357 ( .A1(n8987), .A2(n8966), .ZN(n13052) );
  NAND2_X1 U11358 ( .A1(n9116), .A2(n13052), .ZN(n8970) );
  INV_X1 U11359 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13054) );
  OR2_X1 U11360 ( .A1(n9139), .A2(n13054), .ZN(n8969) );
  INV_X1 U11361 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13227) );
  OR2_X1 U11362 ( .A1(n7001), .A2(n13227), .ZN(n8968) );
  INV_X1 U11363 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13166) );
  OR2_X1 U11364 ( .A1(n7003), .A2(n13166), .ZN(n8967) );
  NAND2_X1 U11365 ( .A1(n13163), .A2(n13061), .ZN(n9303) );
  INV_X1 U11366 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11698) );
  NAND2_X1 U11367 ( .A1(n11698), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8992) );
  INV_X1 U11368 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12467) );
  NAND2_X1 U11369 ( .A1(n12467), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8973) );
  AND2_X1 U11370 ( .A1(n8992), .A2(n8973), .ZN(n8974) );
  OR2_X1 U11371 ( .A1(n8975), .A2(n8974), .ZN(n8976) );
  NAND2_X1 U11372 ( .A1(n8993), .A2(n8976), .ZN(n10702) );
  OR2_X1 U11373 ( .A1(n10702), .A2(n9014), .ZN(n8982) );
  INV_X1 U11374 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8978) );
  AOI22_X1 U11375 ( .A1(n8666), .A2(SI_19_), .B1(n11577), .B2(n8980), .ZN(
        n8981) );
  INV_X1 U11376 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13037) );
  OR2_X1 U11377 ( .A1(n9139), .A2(n13037), .ZN(n8984) );
  INV_X1 U11378 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13222) );
  OR2_X1 U11379 ( .A1(n7001), .A2(n13222), .ZN(n8983) );
  AND2_X1 U11380 ( .A1(n8984), .A2(n8983), .ZN(n8991) );
  INV_X1 U11381 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11382 ( .A1(n8987), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U11383 ( .A1(n9000), .A2(n8988), .ZN(n13035) );
  NAND2_X1 U11384 ( .A1(n13035), .A2(n9116), .ZN(n8990) );
  INV_X1 U11385 ( .A(n7003), .ZN(n9002) );
  NAND2_X1 U11386 ( .A1(n9002), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8989) );
  OR2_X1 U11387 ( .A1(n13157), .A2(n13051), .ZN(n12882) );
  AND2_X1 U11388 ( .A1(n12882), .A2(n13040), .ZN(n9297) );
  NAND2_X1 U11389 ( .A1(n13157), .A2(n13051), .ZN(n12881) );
  NAND2_X1 U11390 ( .A1(n8996), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U11391 ( .A1(n9009), .A2(n8997), .ZN(n11106) );
  NAND2_X1 U11392 ( .A1(n8666), .A2(SI_20_), .ZN(n8998) );
  NAND2_X1 U11393 ( .A1(n9000), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9001) );
  NAND2_X1 U11394 ( .A1(n9019), .A2(n9001), .ZN(n13024) );
  NAND2_X1 U11395 ( .A1(n13024), .A2(n9116), .ZN(n9005) );
  AOI22_X1 U11396 ( .A1(n9151), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n9138), .B2(
        P3_REG0_REG_20__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11397 ( .A1(n9002), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9003) );
  OR2_X1 U11398 ( .A1(n13019), .A2(n13031), .ZN(n9007) );
  NAND2_X1 U11399 ( .A1(n11903), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U11400 ( .A1(n11902), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9010) );
  AND2_X1 U11401 ( .A1(n9023), .A2(n9010), .ZN(n9011) );
  OR2_X1 U11402 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  NAND2_X1 U11403 ( .A1(n9024), .A2(n9013), .ZN(n11295) );
  NAND2_X1 U11404 ( .A1(n8666), .A2(SI_21_), .ZN(n9015) );
  INV_X1 U11405 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13151) );
  INV_X1 U11406 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U11407 ( .A1(n9019), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U11408 ( .A1(n9027), .A2(n9020), .ZN(n13011) );
  NAND2_X1 U11409 ( .A1(n13011), .A2(n9116), .ZN(n9022) );
  AOI22_X1 U11410 ( .A1(n9151), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n9138), .B2(
        P3_REG0_REG_21__SCAN_IN), .ZN(n9021) );
  OAI211_X1 U11411 ( .C1(n7003), .C2(n13151), .A(n9022), .B(n9021), .ZN(n12648) );
  INV_X1 U11412 ( .A(n12648), .ZN(n13018) );
  NOR2_X1 U11413 ( .A1(n13010), .A2(n13018), .ZN(n9315) );
  NAND2_X1 U11414 ( .A1(n13010), .A2(n13018), .ZN(n9313) );
  XNOR2_X1 U11415 ( .A(n11969), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9034) );
  XNOR2_X1 U11416 ( .A(n9035), .B(n9034), .ZN(n11328) );
  NAND2_X1 U11417 ( .A1(n11328), .A2(n9148), .ZN(n9026) );
  NAND2_X1 U11418 ( .A1(n8666), .A2(SI_22_), .ZN(n9025) );
  NAND2_X1 U11419 ( .A1(n9027), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11420 ( .A1(n9039), .A2(n9028), .ZN(n13000) );
  NAND2_X1 U11421 ( .A1(n13000), .A2(n9116), .ZN(n9033) );
  INV_X1 U11422 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13147) );
  NAND2_X1 U11423 ( .A1(n9138), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9030) );
  NAND2_X1 U11424 ( .A1(n9151), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9029) );
  OAI211_X1 U11425 ( .C1(n13147), .C2(n7003), .A(n9030), .B(n9029), .ZN(n9031)
         );
  INV_X1 U11426 ( .A(n9031), .ZN(n9032) );
  NAND2_X1 U11427 ( .A1(n9033), .A2(n9032), .ZN(n12985) );
  NAND2_X1 U11428 ( .A1(n11969), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9036) );
  XNOR2_X1 U11429 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9046) );
  XNOR2_X1 U11430 ( .A(n9047), .B(n9046), .ZN(n11562) );
  NAND2_X1 U11431 ( .A1(n11562), .A2(n9148), .ZN(n9038) );
  NAND2_X1 U11432 ( .A1(n8666), .A2(SI_23_), .ZN(n9037) );
  NAND2_X1 U11433 ( .A1(n9039), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9040) );
  NAND2_X1 U11434 ( .A1(n9055), .A2(n9040), .ZN(n12989) );
  NAND2_X1 U11435 ( .A1(n12989), .A2(n9116), .ZN(n9045) );
  INV_X1 U11436 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13143) );
  NAND2_X1 U11437 ( .A1(n9138), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U11438 ( .A1(n9151), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9041) );
  OAI211_X1 U11439 ( .C1(n13143), .C2(n7003), .A(n9042), .B(n9041), .ZN(n9043)
         );
  INV_X1 U11440 ( .A(n9043), .ZN(n9044) );
  XNOR2_X1 U11441 ( .A(n13139), .B(n12997), .ZN(n12891) );
  NAND2_X1 U11442 ( .A1(n12149), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11443 ( .A1(n9050), .A2(n12427), .ZN(n9051) );
  INV_X1 U11444 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12425) );
  XNOR2_X1 U11445 ( .A(n9064), .B(n12425), .ZN(n11897) );
  NAND2_X1 U11446 ( .A1(n11897), .A2(n9148), .ZN(n9053) );
  NAND2_X1 U11447 ( .A1(n8666), .A2(SI_24_), .ZN(n9052) );
  INV_X1 U11448 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15847) );
  NAND2_X1 U11449 ( .A1(n9055), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11450 ( .A1(n9069), .A2(n9056), .ZN(n12975) );
  NAND2_X1 U11451 ( .A1(n12975), .A2(n9116), .ZN(n9061) );
  INV_X1 U11452 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13137) );
  NAND2_X1 U11453 ( .A1(n9138), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U11454 ( .A1(n9151), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9057) );
  OAI211_X1 U11455 ( .C1(n13137), .C2(n7003), .A(n9058), .B(n9057), .ZN(n9059)
         );
  INV_X1 U11456 ( .A(n9059), .ZN(n9060) );
  NAND2_X1 U11457 ( .A1(n9061), .A2(n9060), .ZN(n12986) );
  NAND2_X1 U11458 ( .A1(n12974), .A2(n12630), .ZN(n9206) );
  OR2_X1 U11459 ( .A1(n12974), .A2(n12630), .ZN(n9062) );
  NAND2_X1 U11460 ( .A1(n9206), .A2(n9062), .ZN(n12966) );
  XNOR2_X1 U11461 ( .A(n13893), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9066) );
  XNOR2_X1 U11462 ( .A(n9078), .B(n9066), .ZN(n12013) );
  NAND2_X1 U11463 ( .A1(n12013), .A2(n9148), .ZN(n9068) );
  NAND2_X1 U11464 ( .A1(n8666), .A2(SI_25_), .ZN(n9067) );
  NAND2_X1 U11465 ( .A1(n9069), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U11466 ( .A1(n9095), .A2(n9070), .ZN(n12961) );
  NAND2_X1 U11467 ( .A1(n12961), .A2(n9116), .ZN(n9075) );
  INV_X1 U11468 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13133) );
  NAND2_X1 U11469 ( .A1(n9138), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11470 ( .A1(n9151), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9071) );
  OAI211_X1 U11471 ( .C1(n13133), .C2(n7003), .A(n9072), .B(n9071), .ZN(n9073)
         );
  INV_X1 U11472 ( .A(n9073), .ZN(n9074) );
  NAND2_X1 U11473 ( .A1(n9075), .A2(n9074), .ZN(n12897) );
  NAND2_X1 U11474 ( .A1(n12960), .A2(n12970), .ZN(n9076) );
  NAND2_X1 U11475 ( .A1(n13893), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9077) );
  INV_X1 U11476 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14692) );
  NAND2_X1 U11477 ( .A1(n14692), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9079) );
  XNOR2_X1 U11478 ( .A(n13888), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U11479 ( .A1(n8666), .A2(SI_26_), .ZN(n9082) );
  XNOR2_X1 U11480 ( .A(n9095), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n12947) );
  NAND2_X1 U11481 ( .A1(n12947), .A2(n9116), .ZN(n9087) );
  INV_X1 U11482 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U11483 ( .A1(n9138), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11484 ( .A1(n9151), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9083) );
  OAI211_X1 U11485 ( .C1(n13129), .C2(n7003), .A(n9084), .B(n9083), .ZN(n9085)
         );
  INV_X1 U11486 ( .A(n9085), .ZN(n9086) );
  NAND2_X1 U11487 ( .A1(n13125), .A2(n12956), .ZN(n9332) );
  NOR2_X1 U11488 ( .A1(n13888), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9088) );
  NAND2_X1 U11489 ( .A1(n13888), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9090) );
  XNOR2_X1 U11490 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9091) );
  XNOR2_X1 U11491 ( .A(n9104), .B(n9091), .ZN(n12261) );
  NAND2_X1 U11492 ( .A1(n12261), .A2(n9148), .ZN(n9093) );
  NAND2_X1 U11493 ( .A1(n8666), .A2(SI_27_), .ZN(n9092) );
  OAI21_X1 U11494 ( .B1(n9095), .B2(P3_REG3_REG_26__SCAN_IN), .A(
        P3_REG3_REG_27__SCAN_IN), .ZN(n9096) );
  INV_X1 U11495 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15653) );
  INV_X1 U11496 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15812) );
  NAND2_X1 U11497 ( .A1(n15653), .A2(n15812), .ZN(n9094) );
  NAND2_X1 U11498 ( .A1(n9096), .A2(n9110), .ZN(n12934) );
  NAND2_X1 U11499 ( .A1(n12934), .A2(n9116), .ZN(n9101) );
  INV_X1 U11500 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13124) );
  NAND2_X1 U11501 ( .A1(n9138), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U11502 ( .A1(n9151), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9097) );
  OAI211_X1 U11503 ( .C1(n13124), .C2(n7003), .A(n9098), .B(n9097), .ZN(n9099)
         );
  INV_X1 U11504 ( .A(n9099), .ZN(n9100) );
  NAND2_X1 U11505 ( .A1(n12933), .A2(n12943), .ZN(n9201) );
  AND2_X1 U11506 ( .A1(n12459), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11507 ( .A1(n14685), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9105) );
  XNOR2_X1 U11508 ( .A(n12464), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U11509 ( .A1(n12491), .A2(n9148), .ZN(n9108) );
  NAND2_X1 U11510 ( .A1(n8666), .A2(SI_28_), .ZN(n9107) );
  NAND2_X2 U11511 ( .A1(n9108), .A2(n9107), .ZN(n13118) );
  INV_X1 U11512 ( .A(n9110), .ZN(n9109) );
  INV_X1 U11513 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12571) );
  NAND2_X1 U11514 ( .A1(n9109), .A2(n12571), .ZN(n12860) );
  NAND2_X1 U11515 ( .A1(n9110), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U11516 ( .A1(n12860), .A2(n9111), .ZN(n12921) );
  INV_X1 U11517 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U11518 ( .A1(n9138), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U11519 ( .A1(n9151), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9112) );
  OAI211_X1 U11520 ( .C1(n9114), .C2(n7003), .A(n9113), .B(n9112), .ZN(n9115)
         );
  NAND2_X1 U11521 ( .A1(n13118), .A2(n12930), .ZN(n9202) );
  INV_X1 U11522 ( .A(n9202), .ZN(n9117) );
  OR2_X2 U11523 ( .A1(n13118), .A2(n12930), .ZN(n9204) );
  NOR2_X1 U11524 ( .A1(n12464), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U11525 ( .A1(n12464), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9120) );
  XNOR2_X1 U11526 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n9129) );
  XNOR2_X1 U11527 ( .A(n9131), .B(n9129), .ZN(n13247) );
  NAND2_X1 U11528 ( .A1(n13247), .A2(n9148), .ZN(n9122) );
  NAND2_X1 U11529 ( .A1(n8666), .A2(SI_29_), .ZN(n9121) );
  INV_X1 U11530 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U11531 ( .A1(n9151), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9125) );
  NAND2_X1 U11532 ( .A1(n9138), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9124) );
  OAI211_X1 U11533 ( .C1(n7003), .C2(n9126), .A(n9125), .B(n9124), .ZN(n9127)
         );
  INV_X1 U11534 ( .A(n9127), .ZN(n9128) );
  INV_X1 U11535 ( .A(n9129), .ZN(n9130) );
  NAND2_X1 U11536 ( .A1(n13886), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9133) );
  INV_X1 U11537 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14682) );
  NAND2_X1 U11538 ( .A1(n14682), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U11539 ( .A1(n9133), .A2(n9132), .ZN(n9144) );
  XNOR2_X1 U11540 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n9134) );
  XNOR2_X1 U11541 ( .A(n9135), .B(n9134), .ZN(n13237) );
  NAND2_X1 U11542 ( .A1(n13237), .A2(n9148), .ZN(n9137) );
  NAND2_X1 U11543 ( .A1(n8666), .A2(SI_31_), .ZN(n9136) );
  INV_X1 U11544 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13109) );
  NAND2_X1 U11545 ( .A1(n9138), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9141) );
  INV_X1 U11546 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12862) );
  OR2_X1 U11547 ( .A1(n9139), .A2(n12862), .ZN(n9140) );
  OAI211_X1 U11548 ( .C1(n13109), .C2(n7003), .A(n9141), .B(n9140), .ZN(n9142)
         );
  INV_X1 U11549 ( .A(n9142), .ZN(n9143) );
  NAND2_X1 U11550 ( .A1(n9145), .A2(n9144), .ZN(n9146) );
  NAND2_X1 U11551 ( .A1(n9147), .A2(n9146), .ZN(n13244) );
  NAND2_X1 U11552 ( .A1(n13244), .A2(n9148), .ZN(n9150) );
  NAND2_X1 U11553 ( .A1(n8666), .A2(SI_30_), .ZN(n9149) );
  INV_X1 U11554 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n9155) );
  NAND2_X1 U11555 ( .A1(n9138), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U11556 ( .A1(n9151), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9152) );
  OAI211_X1 U11557 ( .C1(n9155), .C2(n7003), .A(n9153), .B(n9152), .ZN(n9156)
         );
  INV_X1 U11558 ( .A(n9156), .ZN(n9157) );
  NAND2_X1 U11559 ( .A1(n9158), .A2(n9157), .ZN(n12907) );
  INV_X1 U11560 ( .A(n12907), .ZN(n9163) );
  NAND2_X1 U11561 ( .A1(n13111), .A2(n9163), .ZN(n9159) );
  NAND2_X1 U11562 ( .A1(n9160), .A2(n9159), .ZN(n9344) );
  INV_X1 U11563 ( .A(n9162), .ZN(n12859) );
  NAND2_X1 U11564 ( .A1(n12910), .A2(n12916), .ZN(n9340) );
  OAI21_X1 U11565 ( .B1(n13189), .B2(n12859), .A(n9340), .ZN(n9161) );
  NOR2_X1 U11566 ( .A1(n9344), .A2(n9161), .ZN(n9165) );
  NOR2_X1 U11567 ( .A1(n13111), .A2(n9163), .ZN(n9346) );
  NAND2_X1 U11568 ( .A1(n9175), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9171) );
  MUX2_X1 U11569 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9171), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9172) );
  NAND2_X1 U11570 ( .A1(n9173), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9174) );
  MUX2_X1 U11571 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9174), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9176) );
  NAND2_X1 U11572 ( .A1(n9176), .A2(n9175), .ZN(n11107) );
  INV_X1 U11573 ( .A(n11107), .ZN(n10815) );
  NAND2_X1 U11574 ( .A1(n10860), .A2(n10815), .ZN(n11578) );
  NAND2_X1 U11575 ( .A1(n11565), .A2(n10815), .ZN(n10862) );
  INV_X1 U11576 ( .A(n9346), .ZN(n9196) );
  NAND2_X1 U11577 ( .A1(n9331), .A2(n9332), .ZN(n12940) );
  AND2_X1 U11578 ( .A1(n13010), .A2(n12648), .ZN(n12887) );
  INV_X1 U11579 ( .A(n12887), .ZN(n9177) );
  OR2_X1 U11580 ( .A1(n13010), .A2(n12648), .ZN(n12888) );
  INV_X1 U11581 ( .A(n9178), .ZN(n9320) );
  NAND2_X1 U11582 ( .A1(n9283), .A2(n9179), .ZN(n14836) );
  INV_X1 U11583 ( .A(n14836), .ZN(n14831) );
  OR2_X1 U11584 ( .A1(n9278), .A2(n6741), .ZN(n14841) );
  NAND2_X1 U11585 ( .A1(n15397), .A2(n12131), .ZN(n12075) );
  OAI21_X1 U11586 ( .B1(n15397), .B2(n12131), .A(n12075), .ZN(n12152) );
  INV_X1 U11587 ( .A(n12152), .ZN(n9180) );
  NOR2_X1 U11588 ( .A1(n9180), .A2(n11570), .ZN(n9182) );
  NOR2_X1 U11589 ( .A1(n11571), .A2(n11595), .ZN(n9181) );
  AND4_X1 U11590 ( .A1(n9182), .A2(n9181), .A3(n11600), .A4(n11616), .ZN(n9185) );
  NOR2_X1 U11591 ( .A1(n15412), .A2(n11775), .ZN(n9183) );
  NAND2_X1 U11592 ( .A1(n9261), .A2(n9265), .ZN(n12326) );
  INV_X1 U11593 ( .A(n12326), .ZN(n12079) );
  AND2_X1 U11594 ( .A1(n15448), .A2(n10927), .ZN(n9215) );
  NOR2_X1 U11595 ( .A1(n15457), .A2(n9215), .ZN(n10809) );
  AND4_X1 U11596 ( .A1(n9183), .A2(n15396), .A3(n12079), .A4(n10809), .ZN(
        n9184) );
  NAND4_X1 U11597 ( .A1(n9185), .A2(n9184), .A3(n12334), .A4(n14861), .ZN(
        n9186) );
  NOR2_X1 U11598 ( .A1(n14841), .A2(n9186), .ZN(n9187) );
  NAND4_X1 U11599 ( .A1(n13087), .A2(n13097), .A3(n14831), .A4(n9187), .ZN(
        n9188) );
  NOR2_X1 U11600 ( .A1(n12878), .A2(n9188), .ZN(n9189) );
  NAND4_X1 U11601 ( .A1(n9297), .A2(n9189), .A3(n12881), .A4(n9303), .ZN(n9190) );
  OR4_X1 U11602 ( .A1(n13008), .A2(n12999), .A3(n13020), .A4(n9190), .ZN(n9191) );
  OR3_X1 U11603 ( .A1(n12966), .A2(n12891), .A3(n9191), .ZN(n9192) );
  NOR2_X1 U11604 ( .A1(n12940), .A2(n9192), .ZN(n9193) );
  AND3_X1 U11605 ( .A1(n12919), .A2(n9193), .A3(n12958), .ZN(n9195) );
  NAND4_X1 U11606 ( .A1(n9196), .A2(n12903), .A3(n9195), .A4(n9194), .ZN(n9197) );
  NOR3_X1 U11607 ( .A1(n9344), .A2(n9347), .A3(n9197), .ZN(n9198) );
  NAND2_X2 U11608 ( .A1(n13115), .A2(n10860), .ZN(n10820) );
  NAND2_X1 U11609 ( .A1(n9202), .A2(n9201), .ZN(n9203) );
  NAND2_X1 U11610 ( .A1(n9203), .A2(n11580), .ZN(n9205) );
  INV_X1 U11611 ( .A(n12940), .ZN(n12941) );
  XNOR2_X1 U11612 ( .A(n9206), .B(n10820), .ZN(n9207) );
  OAI21_X1 U11613 ( .B1(n12966), .B2(n6757), .A(n9207), .ZN(n9327) );
  INV_X1 U11614 ( .A(n13008), .ZN(n9312) );
  OR3_X1 U11615 ( .A1(n13019), .A2(n13031), .A3(n10820), .ZN(n9209) );
  NAND3_X1 U11616 ( .A1(n13019), .A2(n13031), .A3(n10820), .ZN(n9208) );
  AND2_X1 U11617 ( .A1(n9209), .A2(n9208), .ZN(n9311) );
  MUX2_X1 U11618 ( .A(n12881), .B(n12882), .S(n10820), .Z(n9210) );
  INV_X1 U11619 ( .A(n9210), .ZN(n9211) );
  OR2_X1 U11620 ( .A1(n13020), .A2(n9211), .ZN(n9308) );
  NAND2_X1 U11621 ( .A1(n9244), .A2(n9213), .ZN(n9214) );
  AOI21_X1 U11622 ( .B1(n11600), .B2(n7307), .A(n9214), .ZN(n9247) );
  INV_X1 U11623 ( .A(n9215), .ZN(n9216) );
  NAND2_X1 U11624 ( .A1(n9216), .A2(n13115), .ZN(n9219) );
  NAND2_X1 U11625 ( .A1(n9216), .A2(n10860), .ZN(n9217) );
  NAND3_X1 U11626 ( .A1(n10867), .A2(n10820), .A3(n9217), .ZN(n9218) );
  OAI21_X1 U11627 ( .B1(n11570), .B2(n9219), .A(n9218), .ZN(n9221) );
  NAND2_X1 U11628 ( .A1(n15457), .A2(n11565), .ZN(n9220) );
  NAND2_X1 U11629 ( .A1(n9221), .A2(n9220), .ZN(n9224) );
  MUX2_X1 U11630 ( .A(n9222), .B(n10867), .S(n11580), .Z(n9223) );
  NAND3_X1 U11631 ( .A1(n9224), .A2(n15429), .A3(n9223), .ZN(n9235) );
  NAND2_X1 U11632 ( .A1(n9230), .A2(n9225), .ZN(n9228) );
  NAND2_X1 U11633 ( .A1(n9231), .A2(n9226), .ZN(n9227) );
  MUX2_X1 U11634 ( .A(n9228), .B(n9227), .S(n11580), .Z(n9229) );
  INV_X1 U11635 ( .A(n9229), .ZN(n9234) );
  MUX2_X1 U11636 ( .A(n9231), .B(n9230), .S(n11580), .Z(n9232) );
  INV_X1 U11637 ( .A(n9232), .ZN(n9233) );
  NAND2_X1 U11638 ( .A1(n7759), .A2(n11600), .ZN(n9242) );
  INV_X1 U11639 ( .A(n9236), .ZN(n9240) );
  NAND2_X1 U11640 ( .A1(n9238), .A2(n9237), .ZN(n9239) );
  AOI21_X1 U11641 ( .B1(n11600), .B2(n9240), .A(n9239), .ZN(n9241) );
  OAI22_X1 U11642 ( .A1(n9243), .A2(n9242), .B1(n11580), .B2(n9241), .ZN(n9245) );
  NAND2_X1 U11643 ( .A1(n9245), .A2(n9244), .ZN(n9246) );
  MUX2_X1 U11644 ( .A(n9250), .B(n9249), .S(n11580), .Z(n9251) );
  NAND3_X1 U11645 ( .A1(n9252), .A2(n15396), .A3(n9251), .ZN(n9256) );
  MUX2_X1 U11646 ( .A(n9254), .B(n9253), .S(n10820), .Z(n9255) );
  NAND3_X1 U11647 ( .A1(n9256), .A2(n12152), .A3(n9255), .ZN(n9260) );
  NAND2_X1 U11648 ( .A1(n12113), .A2(n11580), .ZN(n9258) );
  NAND2_X1 U11649 ( .A1(n15397), .A2(n10820), .ZN(n9257) );
  MUX2_X1 U11650 ( .A(n9258), .B(n9257), .S(n12159), .Z(n9259) );
  NAND4_X1 U11651 ( .A1(n9260), .A2(n12334), .A3(n12079), .A4(n9259), .ZN(
        n9273) );
  INV_X1 U11652 ( .A(n9261), .ZN(n9262) );
  NAND2_X1 U11653 ( .A1(n12334), .A2(n9262), .ZN(n9264) );
  NAND3_X1 U11654 ( .A1(n9264), .A2(n9274), .A3(n9263), .ZN(n9270) );
  INV_X1 U11655 ( .A(n9265), .ZN(n9266) );
  NAND2_X1 U11656 ( .A1(n12334), .A2(n9266), .ZN(n9268) );
  NAND3_X1 U11657 ( .A1(n9268), .A2(n9267), .A3(n9275), .ZN(n9269) );
  MUX2_X1 U11658 ( .A(n9270), .B(n9269), .S(n11580), .Z(n9271) );
  INV_X1 U11659 ( .A(n9271), .ZN(n9272) );
  NAND2_X1 U11660 ( .A1(n9273), .A2(n9272), .ZN(n9277) );
  INV_X1 U11661 ( .A(n14841), .ZN(n14848) );
  MUX2_X1 U11662 ( .A(n9275), .B(n9274), .S(n11580), .Z(n9276) );
  NAND3_X1 U11663 ( .A1(n9277), .A2(n14848), .A3(n9276), .ZN(n9281) );
  MUX2_X1 U11664 ( .A(n9278), .B(n6741), .S(n11580), .Z(n9279) );
  NOR2_X1 U11665 ( .A1(n14836), .A2(n9279), .ZN(n9280) );
  NAND2_X1 U11666 ( .A1(n9281), .A2(n9280), .ZN(n9282) );
  NAND2_X1 U11667 ( .A1(n13097), .A2(n9284), .ZN(n9286) );
  NAND3_X1 U11668 ( .A1(n9286), .A2(n9293), .A3(n9285), .ZN(n9287) );
  NAND2_X1 U11669 ( .A1(n9287), .A2(n10820), .ZN(n9289) );
  INV_X1 U11670 ( .A(n9292), .ZN(n9288) );
  AOI21_X1 U11671 ( .B1(n9290), .B2(n9289), .A(n9288), .ZN(n9295) );
  AOI21_X1 U11672 ( .B1(n9292), .B2(n9291), .A(n10820), .ZN(n9294) );
  OAI22_X1 U11673 ( .A1(n9295), .A2(n9294), .B1(n10820), .B2(n9293), .ZN(n9299) );
  INV_X1 U11674 ( .A(n9296), .ZN(n9298) );
  NAND2_X1 U11675 ( .A1(n9297), .A2(n11580), .ZN(n9306) );
  AOI22_X1 U11676 ( .A1(n9299), .A2(n13066), .B1(n9298), .B2(n9306), .ZN(n9300) );
  INV_X1 U11677 ( .A(n9301), .ZN(n9302) );
  AND2_X1 U11678 ( .A1(n9303), .A2(n9302), .ZN(n9305) );
  NAND3_X1 U11679 ( .A1(n12881), .A2(n10820), .A3(n9303), .ZN(n9304) );
  OAI21_X1 U11680 ( .B1(n9306), .B2(n9305), .A(n9304), .ZN(n9307) );
  OR2_X1 U11681 ( .A1(n9308), .A2(n9307), .ZN(n9309) );
  NAND4_X1 U11682 ( .A1(n9312), .A2(n9311), .A3(n9310), .A4(n9309), .ZN(n9318)
         );
  INV_X1 U11683 ( .A(n9313), .ZN(n9314) );
  MUX2_X1 U11684 ( .A(n9315), .B(n9314), .S(n11580), .Z(n9316) );
  INV_X1 U11685 ( .A(n9316), .ZN(n9317) );
  NAND2_X1 U11686 ( .A1(n9318), .A2(n9317), .ZN(n9319) );
  NOR2_X1 U11687 ( .A1(n12999), .A2(n9319), .ZN(n9323) );
  MUX2_X1 U11688 ( .A(n9321), .B(n9320), .S(n11580), .Z(n9322) );
  NAND3_X1 U11689 ( .A1(n13139), .A2(n12997), .A3(n11580), .ZN(n9324) );
  NAND2_X1 U11690 ( .A1(n9325), .A2(n9324), .ZN(n9326) );
  OR3_X1 U11691 ( .A1(n12960), .A2(n12970), .A3(n10820), .ZN(n9329) );
  NAND3_X1 U11692 ( .A1(n12960), .A2(n12970), .A3(n10820), .ZN(n9328) );
  NAND4_X1 U11693 ( .A1(n12941), .A2(n9330), .A3(n9329), .A4(n9328), .ZN(n9334) );
  MUX2_X1 U11694 ( .A(n9332), .B(n9331), .S(n10820), .Z(n9333) );
  AND2_X1 U11695 ( .A1(n9334), .A2(n9333), .ZN(n9336) );
  OR3_X1 U11696 ( .A1(n12933), .A2(n11580), .A3(n12943), .ZN(n9335) );
  OAI21_X1 U11697 ( .B1(n9336), .B2(n12929), .A(n9335), .ZN(n9337) );
  NAND2_X1 U11698 ( .A1(n9342), .A2(n9341), .ZN(n9343) );
  INV_X1 U11699 ( .A(n9344), .ZN(n9345) );
  INV_X1 U11700 ( .A(n9347), .ZN(n9348) );
  NAND2_X1 U11701 ( .A1(n11577), .A2(n11107), .ZN(n15438) );
  OAI21_X1 U11702 ( .B1(n9349), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9351) );
  XNOR2_X1 U11703 ( .A(n9351), .B(n9350), .ZN(n10497) );
  OR2_X1 U11704 ( .A1(n10497), .A2(P3_U3151), .ZN(n11563) );
  NAND2_X1 U11705 ( .A1(n9354), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9355) );
  MUX2_X1 U11706 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9355), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9356) );
  OR2_X1 U11707 ( .A1(n9354), .A2(P3_IR_REG_25__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U11708 ( .A1(n9356), .A2(n9361), .ZN(n12014) );
  INV_X1 U11709 ( .A(n9357), .ZN(n9358) );
  NAND2_X1 U11710 ( .A1(n9358), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9359) );
  MUX2_X1 U11711 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9359), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9360) );
  NAND2_X1 U11712 ( .A1(n9360), .A2(n9354), .ZN(n11899) );
  NOR2_X1 U11713 ( .A1(n12014), .A2(n11899), .ZN(n9363) );
  NAND2_X1 U11714 ( .A1(n9361), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9362) );
  XNOR2_X1 U11715 ( .A(n9362), .B(P3_IR_REG_26__SCAN_IN), .ZN(n10604) );
  OR2_X1 U11716 ( .A1(n11583), .A2(n10820), .ZN(n10807) );
  NOR3_X1 U11717 ( .A1(n10918), .A2(n12840), .A3(n12857), .ZN(n9365) );
  OAI21_X1 U11718 ( .B1(n11563), .B2(n13115), .A(P3_B_REG_SCAN_IN), .ZN(n9364)
         );
  OR2_X1 U11719 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  OR2_X1 U11720 ( .A1(n9367), .A2(n10188), .ZN(n10192) );
  INV_X2 U11721 ( .A(n7798), .ZN(n13720) );
  NOR2_X1 U11722 ( .A1(n10428), .A2(n9379), .ZN(n10660) );
  AOI21_X1 U11723 ( .B1(n6697), .B2(n13720), .A(n10660), .ZN(n9370) );
  NAND2_X1 U11724 ( .A1(n13364), .A2(n12389), .ZN(n9372) );
  INV_X1 U11725 ( .A(n10740), .ZN(n9371) );
  NAND2_X1 U11726 ( .A1(n9372), .A2(n9371), .ZN(n9373) );
  NAND2_X1 U11727 ( .A1(n10741), .A2(n9373), .ZN(n9374) );
  XNOR2_X1 U11728 ( .A(n9379), .B(n10469), .ZN(n9375) );
  NAND2_X1 U11729 ( .A1(n13363), .A2(n12389), .ZN(n9376) );
  XNOR2_X1 U11730 ( .A(n9375), .B(n9376), .ZN(n10742) );
  NAND2_X1 U11731 ( .A1(n9374), .A2(n10742), .ZN(n10749) );
  INV_X1 U11732 ( .A(n9375), .ZN(n9377) );
  NAND2_X1 U11733 ( .A1(n9377), .A2(n9376), .ZN(n9378) );
  NAND2_X1 U11734 ( .A1(n10749), .A2(n9378), .ZN(n10114) );
  XNOR2_X1 U11735 ( .A(n10580), .B(n11089), .ZN(n9380) );
  AND2_X1 U11736 ( .A1(n8584), .A2(n13720), .ZN(n9381) );
  NAND2_X1 U11737 ( .A1(n9380), .A2(n9381), .ZN(n9384) );
  INV_X1 U11738 ( .A(n9380), .ZN(n10690) );
  INV_X1 U11739 ( .A(n9381), .ZN(n9382) );
  NAND2_X1 U11740 ( .A1(n10690), .A2(n9382), .ZN(n9383) );
  NAND2_X1 U11741 ( .A1(n9384), .A2(n9383), .ZN(n10113) );
  OR2_X1 U11742 ( .A1(n10114), .A2(n10113), .ZN(n10112) );
  XNOR2_X1 U11743 ( .A(n10899), .B(n11089), .ZN(n9386) );
  NAND2_X1 U11744 ( .A1(n13362), .A2(n12389), .ZN(n9387) );
  XNOR2_X1 U11745 ( .A(n9386), .B(n9387), .ZN(n10700) );
  AND2_X1 U11746 ( .A1(n10700), .A2(n9384), .ZN(n9385) );
  INV_X1 U11747 ( .A(n9386), .ZN(n10650) );
  XNOR2_X1 U11748 ( .A(n11084), .B(n11089), .ZN(n9388) );
  NAND2_X1 U11749 ( .A1(n13361), .A2(n12389), .ZN(n9389) );
  XNOR2_X1 U11750 ( .A(n9388), .B(n9389), .ZN(n10652) );
  INV_X1 U11751 ( .A(n9388), .ZN(n9390) );
  XNOR2_X1 U11752 ( .A(n11211), .B(n11089), .ZN(n9391) );
  AND2_X1 U11753 ( .A1(n13360), .A2(n13720), .ZN(n9392) );
  NAND2_X1 U11754 ( .A1(n9391), .A2(n9392), .ZN(n9396) );
  INV_X1 U11755 ( .A(n9391), .ZN(n11122) );
  INV_X1 U11756 ( .A(n9392), .ZN(n9393) );
  NAND2_X1 U11757 ( .A1(n11122), .A2(n9393), .ZN(n9394) );
  NAND2_X1 U11758 ( .A1(n9396), .A2(n9394), .ZN(n11035) );
  INV_X1 U11759 ( .A(n11035), .ZN(n9395) );
  XNOR2_X1 U11760 ( .A(n11375), .B(n11089), .ZN(n9397) );
  AND2_X1 U11761 ( .A1(n13359), .A2(n13720), .ZN(n9398) );
  NAND2_X1 U11762 ( .A1(n9397), .A2(n9398), .ZN(n9401) );
  INV_X1 U11763 ( .A(n9397), .ZN(n11393) );
  INV_X1 U11764 ( .A(n9398), .ZN(n9399) );
  NAND2_X1 U11765 ( .A1(n11393), .A2(n9399), .ZN(n9400) );
  AND2_X1 U11766 ( .A1(n9401), .A2(n9400), .ZN(n11119) );
  XNOR2_X1 U11767 ( .A(n11504), .B(n11089), .ZN(n11304) );
  NOR2_X1 U11768 ( .A1(n11503), .A2(n14928), .ZN(n9402) );
  XNOR2_X1 U11769 ( .A(n11304), .B(n9402), .ZN(n11404) );
  INV_X1 U11770 ( .A(n9402), .ZN(n9403) );
  XNOR2_X1 U11771 ( .A(n11677), .B(n11089), .ZN(n9405) );
  NAND2_X1 U11772 ( .A1(n13357), .A2(n12389), .ZN(n9406) );
  XNOR2_X1 U11773 ( .A(n9405), .B(n9406), .ZN(n11303) );
  NAND2_X1 U11774 ( .A1(n9404), .A2(n11303), .ZN(n11309) );
  INV_X1 U11775 ( .A(n9405), .ZN(n9407) );
  NAND2_X1 U11776 ( .A1(n9407), .A2(n9406), .ZN(n9408) );
  NAND2_X1 U11777 ( .A1(n11309), .A2(n9408), .ZN(n11856) );
  XNOR2_X1 U11778 ( .A(n15382), .B(n9464), .ZN(n9409) );
  NOR2_X1 U11779 ( .A1(n13354), .A2(n14928), .ZN(n9410) );
  NAND2_X1 U11780 ( .A1(n9409), .A2(n9410), .ZN(n9414) );
  INV_X1 U11781 ( .A(n9409), .ZN(n11811) );
  INV_X1 U11782 ( .A(n9410), .ZN(n9411) );
  NAND2_X1 U11783 ( .A1(n11811), .A2(n9411), .ZN(n9412) );
  NAND2_X1 U11784 ( .A1(n9414), .A2(n9412), .ZN(n11857) );
  XNOR2_X1 U11785 ( .A(n12064), .B(n11089), .ZN(n11867) );
  NAND2_X1 U11786 ( .A1(n13353), .A2(n12389), .ZN(n9416) );
  XNOR2_X1 U11787 ( .A(n11867), .B(n9416), .ZN(n11813) );
  AND2_X1 U11788 ( .A1(n11813), .A2(n9414), .ZN(n9415) );
  INV_X1 U11789 ( .A(n11867), .ZN(n9417) );
  XNOR2_X1 U11790 ( .A(n14945), .B(n11089), .ZN(n9420) );
  NOR2_X1 U11791 ( .A1(n11996), .A2(n14928), .ZN(n9418) );
  XNOR2_X1 U11792 ( .A(n9420), .B(n9418), .ZN(n11868) );
  INV_X1 U11793 ( .A(n9418), .ZN(n9419) );
  NAND2_X1 U11794 ( .A1(n9420), .A2(n9419), .ZN(n9421) );
  XNOR2_X1 U11795 ( .A(n12195), .B(n9464), .ZN(n12483) );
  NOR2_X1 U11796 ( .A1(n12477), .A2(n14928), .ZN(n9422) );
  NAND2_X1 U11797 ( .A1(n12483), .A2(n9422), .ZN(n9426) );
  INV_X1 U11798 ( .A(n12483), .ZN(n9424) );
  INV_X1 U11799 ( .A(n9422), .ZN(n9423) );
  NAND2_X1 U11800 ( .A1(n9424), .A2(n9423), .ZN(n9425) );
  NAND2_X1 U11801 ( .A1(n9426), .A2(n9425), .ZN(n12239) );
  XNOR2_X1 U11802 ( .A(n14921), .B(n9487), .ZN(n9427) );
  NAND2_X1 U11803 ( .A1(n13350), .A2(n13720), .ZN(n9428) );
  XNOR2_X1 U11804 ( .A(n9427), .B(n9428), .ZN(n12484) );
  INV_X1 U11805 ( .A(n9427), .ZN(n9429) );
  NAND2_X1 U11806 ( .A1(n9429), .A2(n9428), .ZN(n9430) );
  XNOR2_X1 U11807 ( .A(n12364), .B(n9487), .ZN(n9432) );
  AND2_X1 U11808 ( .A1(n13349), .A2(n13720), .ZN(n9431) );
  INV_X1 U11809 ( .A(n9432), .ZN(n9433) );
  INV_X1 U11810 ( .A(n14889), .ZN(n9435) );
  XNOR2_X1 U11811 ( .A(n12383), .B(n9487), .ZN(n9437) );
  NAND2_X1 U11812 ( .A1(n13348), .A2(n13720), .ZN(n9436) );
  XNOR2_X1 U11813 ( .A(n9437), .B(n9436), .ZN(n14888) );
  NAND2_X1 U11814 ( .A1(n9437), .A2(n9436), .ZN(n14898) );
  XNOR2_X1 U11815 ( .A(n13550), .B(n9487), .ZN(n9440) );
  NOR2_X1 U11816 ( .A1(n13549), .A2(n14928), .ZN(n9438) );
  XNOR2_X1 U11817 ( .A(n9440), .B(n9438), .ZN(n14897) );
  INV_X1 U11818 ( .A(n9438), .ZN(n9439) );
  NAND2_X1 U11819 ( .A1(n9440), .A2(n9439), .ZN(n9441) );
  XNOR2_X1 U11820 ( .A(n13744), .B(n9464), .ZN(n9444) );
  NOR2_X1 U11821 ( .A1(n13553), .A2(n14928), .ZN(n9443) );
  XNOR2_X1 U11822 ( .A(n9444), .B(n9443), .ZN(n13322) );
  INV_X1 U11823 ( .A(n13322), .ZN(n9442) );
  NAND2_X1 U11824 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  XNOR2_X1 U11825 ( .A(n13725), .B(n9487), .ZN(n9446) );
  NAND2_X1 U11826 ( .A1(n13517), .A2(n13720), .ZN(n9447) );
  NAND2_X1 U11827 ( .A1(n9446), .A2(n9447), .ZN(n13272) );
  INV_X1 U11828 ( .A(n9446), .ZN(n9449) );
  INV_X1 U11829 ( .A(n9447), .ZN(n9448) );
  NAND2_X1 U11830 ( .A1(n9449), .A2(n9448), .ZN(n13271) );
  INV_X1 U11831 ( .A(n13304), .ZN(n9456) );
  XNOR2_X1 U11832 ( .A(n13816), .B(n9487), .ZN(n9450) );
  INV_X1 U11833 ( .A(n13556), .ZN(n13347) );
  NAND2_X1 U11834 ( .A1(n13347), .A2(n13720), .ZN(n9451) );
  NAND2_X1 U11835 ( .A1(n9450), .A2(n9451), .ZN(n9457) );
  INV_X1 U11836 ( .A(n9450), .ZN(n9453) );
  INV_X1 U11837 ( .A(n9451), .ZN(n9452) );
  NAND2_X1 U11838 ( .A1(n9453), .A2(n9452), .ZN(n9454) );
  NAND2_X1 U11839 ( .A1(n9457), .A2(n9454), .ZN(n13305) );
  INV_X1 U11840 ( .A(n13305), .ZN(n9455) );
  XNOR2_X1 U11841 ( .A(n13699), .B(n9464), .ZN(n9459) );
  NAND2_X1 U11842 ( .A1(n13557), .A2(n13720), .ZN(n9458) );
  XNOR2_X1 U11843 ( .A(n9459), .B(n9458), .ZN(n13279) );
  XNOR2_X1 U11844 ( .A(n13802), .B(n9464), .ZN(n9460) );
  AND2_X1 U11845 ( .A1(n13559), .A2(n13720), .ZN(n13314) );
  INV_X1 U11846 ( .A(n9460), .ZN(n9461) );
  NAND2_X1 U11847 ( .A1(n9462), .A2(n9461), .ZN(n9463) );
  XNOR2_X1 U11848 ( .A(n13865), .B(n9464), .ZN(n9466) );
  NOR2_X1 U11849 ( .A1(n13561), .A2(n14928), .ZN(n9467) );
  AND2_X1 U11850 ( .A1(n9466), .A2(n9467), .ZN(n9465) );
  INV_X1 U11851 ( .A(n9466), .ZN(n13259) );
  INV_X1 U11852 ( .A(n9467), .ZN(n13261) );
  NAND2_X1 U11853 ( .A1(n13259), .A2(n13261), .ZN(n9468) );
  XNOR2_X1 U11854 ( .A(n13659), .B(n9487), .ZN(n9469) );
  NAND2_X1 U11855 ( .A1(n13564), .A2(n12389), .ZN(n9470) );
  XNOR2_X1 U11856 ( .A(n9469), .B(n9470), .ZN(n13295) );
  INV_X1 U11857 ( .A(n9469), .ZN(n9472) );
  INV_X1 U11858 ( .A(n9470), .ZN(n9471) );
  NAND2_X1 U11859 ( .A1(n9472), .A2(n9471), .ZN(n9473) );
  XNOR2_X1 U11860 ( .A(n13639), .B(n9487), .ZN(n9475) );
  NOR2_X1 U11861 ( .A1(n13567), .A2(n14928), .ZN(n9476) );
  XNOR2_X1 U11862 ( .A(n9475), .B(n9476), .ZN(n13286) );
  INV_X1 U11863 ( .A(n9475), .ZN(n9477) );
  NAND2_X1 U11864 ( .A1(n9477), .A2(n9476), .ZN(n9478) );
  XNOR2_X1 U11865 ( .A(n13619), .B(n9487), .ZN(n9479) );
  NAND2_X1 U11866 ( .A1(n13569), .A2(n13720), .ZN(n9480) );
  NAND2_X1 U11867 ( .A1(n9479), .A2(n9480), .ZN(n9484) );
  INV_X1 U11868 ( .A(n9479), .ZN(n9482) );
  INV_X1 U11869 ( .A(n9480), .ZN(n9481) );
  NAND2_X1 U11870 ( .A1(n9482), .A2(n9481), .ZN(n9483) );
  NAND2_X1 U11871 ( .A1(n9484), .A2(n9483), .ZN(n13333) );
  XNOR2_X1 U11872 ( .A(n13609), .B(n9487), .ZN(n9486) );
  NAND2_X1 U11873 ( .A1(n13537), .A2(n12389), .ZN(n9485) );
  NOR2_X1 U11874 ( .A1(n13545), .A2(n14928), .ZN(n9488) );
  XNOR2_X1 U11875 ( .A(n9488), .B(n9487), .ZN(n9489) );
  INV_X1 U11876 ( .A(P2_B_REG_SCAN_IN), .ZN(n12449) );
  XNOR2_X1 U11877 ( .A(n9493), .B(n12449), .ZN(n9490) );
  NAND2_X1 U11878 ( .A1(n9490), .A2(n13891), .ZN(n9492) );
  INV_X1 U11879 ( .A(n13889), .ZN(n9491) );
  INV_X1 U11880 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15366) );
  NAND2_X1 U11881 ( .A1(n15332), .A2(n15366), .ZN(n9495) );
  INV_X1 U11882 ( .A(n9493), .ZN(n12429) );
  NAND2_X1 U11883 ( .A1(n12429), .A2(n13889), .ZN(n9494) );
  NAND2_X1 U11884 ( .A1(n9495), .A2(n9494), .ZN(n15367) );
  INV_X1 U11885 ( .A(n15367), .ZN(n9506) );
  NOR4_X1 U11886 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9499) );
  NOR4_X1 U11887 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9498) );
  NOR4_X1 U11888 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9497) );
  NOR4_X1 U11889 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9496) );
  NAND4_X1 U11890 ( .A1(n9499), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n9505)
         );
  NOR2_X1 U11891 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9503) );
  NOR4_X1 U11892 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9502) );
  NOR4_X1 U11893 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9501) );
  NOR4_X1 U11894 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n9500) );
  NAND4_X1 U11895 ( .A1(n9503), .A2(n9502), .A3(n9501), .A4(n9500), .ZN(n9504)
         );
  OAI21_X1 U11896 ( .B1(n9505), .B2(n9504), .A(n15332), .ZN(n11076) );
  NAND2_X1 U11897 ( .A1(n9506), .A2(n11076), .ZN(n10195) );
  INV_X1 U11898 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15369) );
  NAND2_X1 U11899 ( .A1(n15332), .A2(n15369), .ZN(n9508) );
  NAND2_X1 U11900 ( .A1(n13889), .A2(n13891), .ZN(n9507) );
  NAND2_X1 U11901 ( .A1(n9508), .A2(n9507), .ZN(n11077) );
  OR2_X1 U11902 ( .A1(n9520), .A2(P2_U3088), .ZN(n15365) );
  OR2_X1 U11903 ( .A1(n11077), .A2(n15365), .ZN(n15368) );
  NOR2_X1 U11904 ( .A1(n10195), .A2(n15368), .ZN(n9518) );
  NAND2_X1 U11905 ( .A1(n9522), .A2(n11227), .ZN(n15381) );
  AND2_X1 U11906 ( .A1(n15381), .A2(n9519), .ZN(n9509) );
  NOR2_X1 U11907 ( .A1(n10192), .A2(n11695), .ZN(n11093) );
  NAND2_X1 U11908 ( .A1(n9518), .A2(n11093), .ZN(n9511) );
  NAND2_X1 U11909 ( .A1(n9510), .A2(n11901), .ZN(n10194) );
  NAND2_X1 U11910 ( .A1(n9511), .A2(n13737), .ZN(n14908) );
  AOI21_X1 U11911 ( .B1(n9512), .B2(n14903), .A(n14908), .ZN(n9528) );
  INV_X1 U11912 ( .A(n9512), .ZN(n9513) );
  OR2_X1 U11913 ( .A1(n9519), .A2(n8626), .ZN(n13544) );
  INV_X1 U11914 ( .A(n13544), .ZN(n13307) );
  NAND2_X1 U11915 ( .A1(n13537), .A2(n13307), .ZN(n9516) );
  OR2_X1 U11916 ( .A1(n9514), .A2(n13326), .ZN(n9515) );
  AND2_X1 U11917 ( .A1(n9516), .A2(n9515), .ZN(n13587) );
  NAND2_X1 U11918 ( .A1(n9518), .A2(n9517), .ZN(n13339) );
  OAI21_X1 U11919 ( .B1(n10195), .B2(n11077), .A(n10194), .ZN(n9523) );
  INV_X1 U11920 ( .A(n9519), .ZN(n9521) );
  AOI21_X1 U11921 ( .B1(n9522), .B2(n9521), .A(n9520), .ZN(n11078) );
  NAND2_X1 U11922 ( .A1(n9523), .A2(n11078), .ZN(n10427) );
  NAND2_X1 U11923 ( .A1(n10427), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14911) );
  INV_X1 U11924 ( .A(n14911), .ZN(n13337) );
  AOI22_X1 U11925 ( .A1(n13594), .A2(n13337), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9524) );
  OAI21_X1 U11926 ( .B1(n13587), .B2(n13339), .A(n9524), .ZN(n9525) );
  OAI211_X1 U11927 ( .C1(n9528), .C2(n13596), .A(n9527), .B(n9526), .ZN(
        P2_U3192) );
  INV_X2 U11928 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9689) );
  NAND4_X1 U11929 ( .A1(n9602), .A2(n9533), .A3(n9532), .A4(n9672), .ZN(n9534)
         );
  NAND4_X1 U11930 ( .A1(n9538), .A2(n9537), .A3(n9536), .A4(n9535), .ZN(n9539)
         );
  NOR2_X1 U11931 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9540) );
  NAND4_X1 U11932 ( .A1(n9540), .A2(n10086), .A3(n9562), .A4(n9569), .ZN(
        n10092) );
  INV_X1 U11933 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9541) );
  NAND3_X1 U11934 ( .A1(n9822), .A2(n10094), .A3(n9541), .ZN(n9542) );
  INV_X1 U11935 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9556) );
  INV_X1 U11936 ( .A(n9545), .ZN(n9544) );
  INV_X1 U11937 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U11938 ( .A1(n9544), .A2(n9546), .ZN(n14677) );
  INV_X1 U11939 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9548) );
  XNOR2_X2 U11940 ( .A(n9549), .B(n9548), .ZN(n14684) );
  AND2_X4 U11941 ( .A1(n14684), .A2(n12445), .ZN(n10013) );
  NAND2_X1 U11942 ( .A1(n10013), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9554) );
  INV_X1 U11944 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11456) );
  OR2_X1 U11945 ( .A1(n6689), .A2(n11456), .ZN(n9553) );
  NAND2_X4 U11946 ( .A1(n14684), .A2(n9550), .ZN(n10018) );
  INV_X1 U11947 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15019) );
  INV_X1 U11948 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n14195) );
  OR2_X1 U11949 ( .A1(n10020), .A2(n14195), .ZN(n9551) );
  INV_X1 U11950 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14198) );
  NOR2_X1 U11951 ( .A1(n10154), .A2(n10135), .ZN(n9555) );
  XNOR2_X1 U11952 ( .A(n9555), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14698) );
  XNOR2_X2 U11953 ( .A(n9557), .B(n9556), .ZN(n10107) );
  MUX2_X1 U11954 ( .A(n14198), .B(n14698), .S(n9910), .Z(n11480) );
  NAND2_X1 U11955 ( .A1(n14182), .A2(n11480), .ZN(n10051) );
  INV_X1 U11956 ( .A(n9564), .ZN(n9565) );
  NAND2_X1 U11957 ( .A1(n10093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U11958 ( .A1(n14696), .A2(n14511), .ZN(n10724) );
  INV_X1 U11959 ( .A(n14696), .ZN(n10035) );
  NAND2_X1 U11960 ( .A1(n10035), .A2(n14448), .ZN(n9571) );
  INV_X1 U11961 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11667) );
  OR2_X1 U11962 ( .A1(n6689), .A2(n11667), .ZN(n9575) );
  INV_X1 U11963 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9572) );
  INV_X1 U11964 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10285) );
  OR2_X1 U11965 ( .A1(n10020), .A2(n10285), .ZN(n9573) );
  INV_X1 U11966 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U11967 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9577) );
  MUX2_X1 U11968 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9577), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9578) );
  INV_X1 U11969 ( .A(n9578), .ZN(n9580) );
  MUX2_X1 U11970 ( .A(n11669), .B(n11488), .S(n9660), .Z(n9581) );
  OAI21_X1 U11971 ( .B1(n9582), .B2(n11473), .A(n9581), .ZN(n9584) );
  NAND2_X1 U11972 ( .A1(n9582), .A2(n10052), .ZN(n9583) );
  NAND2_X1 U11973 ( .A1(n10013), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9588) );
  INV_X1 U11974 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11526) );
  OR2_X1 U11975 ( .A1(n9886), .A2(n11526), .ZN(n9587) );
  INV_X1 U11976 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10280) );
  INV_X1 U11977 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10288) );
  OR2_X1 U11978 ( .A1(n10020), .A2(n10288), .ZN(n9585) );
  NOR2_X1 U11979 ( .A1(n9579), .A2(n14676), .ZN(n9589) );
  MUX2_X1 U11980 ( .A(n14676), .B(n9589), .S(P1_IR_REG_2__SCAN_IN), .Z(n9590)
         );
  NAND2_X1 U11981 ( .A1(n10177), .A2(n10289), .ZN(n9592) );
  OR2_X1 U11982 ( .A1(n9997), .A2(n10129), .ZN(n9591) );
  NAND2_X1 U11983 ( .A1(n14181), .A2(n11524), .ZN(n9594) );
  INV_X1 U11984 ( .A(n9594), .ZN(n9596) );
  INV_X1 U11985 ( .A(n11491), .ZN(n9595) );
  MUX2_X1 U11986 ( .A(n9596), .B(n9595), .S(n9660), .Z(n9607) );
  NAND2_X1 U11987 ( .A1(n10013), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9601) );
  OR2_X1 U11988 ( .A1(n6689), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9600) );
  INV_X1 U11989 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9597) );
  OR2_X1 U11990 ( .A1(n10018), .A2(n9597), .ZN(n9599) );
  INV_X1 U11991 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14214) );
  OR2_X1 U11992 ( .A1(n10020), .A2(n14214), .ZN(n9598) );
  NAND4_X1 U11993 ( .A1(n9601), .A2(n9600), .A3(n9599), .A4(n9598), .ZN(n14179) );
  NAND2_X1 U11994 ( .A1(n9603), .A2(n9602), .ZN(n9631) );
  INV_X1 U11995 ( .A(n9631), .ZN(n9604) );
  NOR2_X1 U11996 ( .A1(n9605), .A2(n9604), .ZN(n14218) );
  NAND2_X1 U11997 ( .A1(n14179), .A2(n15159), .ZN(n9610) );
  NOR2_X1 U11998 ( .A1(n9607), .A2(n15088), .ZN(n9608) );
  INV_X1 U11999 ( .A(n9610), .ZN(n9612) );
  INV_X1 U12000 ( .A(n11494), .ZN(n9611) );
  MUX2_X1 U12001 ( .A(n9612), .B(n9611), .S(n10011), .Z(n9613) );
  INV_X1 U12002 ( .A(n9613), .ZN(n9614) );
  NAND2_X1 U12003 ( .A1(n9615), .A2(n9614), .ZN(n9627) );
  INV_X1 U12004 ( .A(n9627), .ZN(n9630) );
  OR2_X1 U12005 ( .A1(n9878), .A2(n10155), .ZN(n9619) );
  OR2_X1 U12006 ( .A1(n9997), .A2(n10131), .ZN(n9618) );
  NAND2_X1 U12007 ( .A1(n9631), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9616) );
  XNOR2_X1 U12008 ( .A(n9616), .B(P1_IR_REG_4__SCAN_IN), .ZN(n15038) );
  NAND2_X1 U12009 ( .A1(n10177), .A2(n15038), .ZN(n9617) );
  NAND2_X1 U12010 ( .A1(n10012), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9624) );
  INV_X1 U12011 ( .A(n10013), .ZN(n10022) );
  INV_X1 U12012 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9620) );
  NAND2_X1 U12013 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9637) );
  OAI21_X1 U12014 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9637), .ZN(n11534) );
  OR2_X1 U12015 ( .A1(n6689), .A2(n11534), .ZN(n9622) );
  INV_X1 U12016 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10281) );
  OR2_X1 U12017 ( .A1(n10018), .A2(n10281), .ZN(n9621) );
  MUX2_X1 U12018 ( .A(n15167), .B(n14023), .S(n10011), .Z(n9626) );
  INV_X1 U12019 ( .A(n9626), .ZN(n9629) );
  INV_X1 U12020 ( .A(n14023), .ZN(n10054) );
  MUX2_X1 U12021 ( .A(n10054), .B(n6901), .S(n10011), .Z(n9625) );
  OR2_X1 U12022 ( .A1(n10157), .A2(n6690), .ZN(n9634) );
  NAND2_X1 U12023 ( .A1(n9655), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9632) );
  XNOR2_X1 U12024 ( .A(n9632), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U12025 ( .A1(n10177), .A2(n10293), .ZN(n9633) );
  OAI211_X1 U12026 ( .C1(n9997), .C2(n10130), .A(n9634), .B(n9633), .ZN(n11556) );
  NAND2_X1 U12027 ( .A1(n10013), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9642) );
  INV_X1 U12028 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11549) );
  OR2_X1 U12029 ( .A1(n10020), .A2(n11549), .ZN(n9641) );
  INV_X1 U12030 ( .A(n9637), .ZN(n9635) );
  NAND2_X1 U12031 ( .A1(n9635), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9649) );
  INV_X1 U12032 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U12033 ( .A1(n9637), .A2(n9636), .ZN(n9638) );
  NAND2_X1 U12034 ( .A1(n9649), .A2(n9638), .ZN(n11554) );
  OR2_X1 U12035 ( .A1(n6689), .A2(n11554), .ZN(n9640) );
  INV_X1 U12036 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10282) );
  NAND4_X1 U12037 ( .A1(n9642), .A2(n9641), .A3(n9640), .A4(n9639), .ZN(n14178) );
  MUX2_X1 U12038 ( .A(n11556), .B(n14178), .S(n10075), .Z(n9644) );
  MUX2_X1 U12039 ( .A(n14178), .B(n11556), .S(n9660), .Z(n9643) );
  NAND2_X1 U12040 ( .A1(n10012), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9654) );
  INV_X1 U12041 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9646) );
  OR2_X1 U12042 ( .A1(n10022), .A2(n9646), .ZN(n9653) );
  INV_X1 U12043 ( .A(n9649), .ZN(n9647) );
  NAND2_X1 U12044 ( .A1(n9647), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9666) );
  INV_X1 U12045 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U12046 ( .A1(n9649), .A2(n9648), .ZN(n9650) );
  NAND2_X1 U12047 ( .A1(n9666), .A2(n9650), .ZN(n11482) );
  OR2_X1 U12048 ( .A1(n6689), .A2(n11482), .ZN(n9652) );
  INV_X1 U12049 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10278) );
  OR2_X1 U12050 ( .A1(n10018), .A2(n10278), .ZN(n9651) );
  NAND4_X1 U12051 ( .A1(n9654), .A2(n9653), .A3(n9652), .A4(n9651), .ZN(n14177) );
  OR2_X1 U12052 ( .A1(n10160), .A2(n6690), .ZN(n9659) );
  INV_X1 U12053 ( .A(n9673), .ZN(n9656) );
  NAND2_X1 U12054 ( .A1(n9656), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9657) );
  XNOR2_X1 U12055 ( .A(n9657), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U12056 ( .A1(n10039), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10177), 
        .B2(n10358), .ZN(n9658) );
  NAND2_X1 U12057 ( .A1(n9659), .A2(n9658), .ZN(n11637) );
  MUX2_X1 U12058 ( .A(n14177), .B(n11637), .S(n9660), .Z(n9663) );
  MUX2_X1 U12059 ( .A(n11637), .B(n14177), .S(n10075), .Z(n9661) );
  INV_X1 U12060 ( .A(n9663), .ZN(n9664) );
  NAND2_X1 U12061 ( .A1(n10013), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9671) );
  INV_X1 U12062 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10364) );
  OR2_X1 U12063 ( .A1(n10020), .A2(n10364), .ZN(n9670) );
  NAND2_X1 U12064 ( .A1(n9666), .A2(n9665), .ZN(n9667) );
  NAND2_X1 U12065 ( .A1(n9683), .A2(n9667), .ZN(n15076) );
  OR2_X1 U12066 ( .A1(n6689), .A2(n15076), .ZN(n9669) );
  INV_X1 U12067 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10359) );
  OR2_X1 U12068 ( .A1(n10018), .A2(n10359), .ZN(n9668) );
  NAND4_X1 U12069 ( .A1(n9671), .A2(n9670), .A3(n9669), .A4(n9668), .ZN(n14176) );
  INV_X1 U12070 ( .A(n9690), .ZN(n9674) );
  NAND2_X1 U12071 ( .A1(n9674), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9675) );
  XNOR2_X1 U12072 ( .A(n9675), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U12073 ( .A1(n10039), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10177), 
        .B2(n10414), .ZN(n9676) );
  NAND2_X1 U12074 ( .A1(n9677), .A2(n9676), .ZN(n15193) );
  MUX2_X1 U12075 ( .A(n14176), .B(n15193), .S(n10011), .Z(n9680) );
  MUX2_X1 U12076 ( .A(n15193), .B(n14176), .S(n10011), .Z(n9678) );
  NAND2_X1 U12077 ( .A1(n10012), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9688) );
  INV_X1 U12078 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9681) );
  OR2_X1 U12079 ( .A1(n10022), .A2(n9681), .ZN(n9687) );
  INV_X1 U12080 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9682) );
  NAND2_X1 U12081 ( .A1(n9683), .A2(n9682), .ZN(n9684) );
  NAND2_X1 U12082 ( .A1(n9703), .A2(n9684), .ZN(n11642) );
  OR2_X1 U12083 ( .A1(n6689), .A2(n11642), .ZN(n9686) );
  INV_X1 U12084 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10415) );
  OR2_X1 U12085 ( .A1(n10018), .A2(n10415), .ZN(n9685) );
  NAND4_X1 U12086 ( .A1(n9688), .A2(n9687), .A3(n9686), .A4(n9685), .ZN(n14175) );
  INV_X1 U12087 ( .A(n9694), .ZN(n9691) );
  NAND2_X1 U12088 ( .A1(n9691), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9692) );
  MUX2_X1 U12089 ( .A(n9692), .B(P1_IR_REG_31__SCAN_IN), .S(n9693), .Z(n9695)
         );
  NAND2_X1 U12090 ( .A1(n9694), .A2(n9693), .ZN(n9720) );
  NAND2_X1 U12091 ( .A1(n9695), .A2(n9720), .ZN(n10441) );
  INV_X1 U12092 ( .A(n10441), .ZN(n10437) );
  AOI22_X1 U12093 ( .A1(n10039), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10177), 
        .B2(n10437), .ZN(n9696) );
  MUX2_X1 U12094 ( .A(n14175), .B(n11879), .S(n10075), .Z(n9700) );
  MUX2_X1 U12095 ( .A(n14175), .B(n11879), .S(n9858), .Z(n9698) );
  NAND2_X1 U12096 ( .A1(n9699), .A2(n9698), .ZN(n9702) );
  NAND2_X1 U12097 ( .A1(n10013), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9708) );
  INV_X1 U12098 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10435) );
  OR2_X1 U12099 ( .A1(n10018), .A2(n10435), .ZN(n9707) );
  INV_X1 U12100 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U12101 ( .A1(n9703), .A2(n10447), .ZN(n9704) );
  NAND2_X1 U12102 ( .A1(n9734), .A2(n9704), .ZN(n11918) );
  OR2_X1 U12103 ( .A1(n6689), .A2(n11918), .ZN(n9706) );
  INV_X1 U12104 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11826) );
  OR2_X1 U12105 ( .A1(n10020), .A2(n11826), .ZN(n9705) );
  NAND4_X1 U12106 ( .A1(n9708), .A2(n9707), .A3(n9706), .A4(n9705), .ZN(n14174) );
  OR2_X1 U12107 ( .A1(n10172), .A2(n6690), .ZN(n9711) );
  NAND2_X1 U12108 ( .A1(n9720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9709) );
  XNOR2_X1 U12109 ( .A(n9709), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U12110 ( .A1(n10039), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10177), 
        .B2(n10484), .ZN(n9710) );
  MUX2_X1 U12111 ( .A(n14174), .B(n11912), .S(n10011), .Z(n9713) );
  MUX2_X1 U12112 ( .A(n14174), .B(n11912), .S(n10075), .Z(n9712) );
  INV_X1 U12113 ( .A(n9713), .ZN(n9714) );
  NAND2_X1 U12114 ( .A1(n10013), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9719) );
  INV_X1 U12115 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9715) );
  OR2_X1 U12116 ( .A1(n10020), .A2(n9715), .ZN(n9718) );
  INV_X1 U12117 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9733) );
  XNOR2_X1 U12118 ( .A(n9734), .B(n9733), .ZN(n11750) );
  OR2_X1 U12119 ( .A1(n6689), .A2(n11750), .ZN(n9717) );
  INV_X1 U12120 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10480) );
  OR2_X1 U12121 ( .A1(n10018), .A2(n10480), .ZN(n9716) );
  NAND4_X1 U12122 ( .A1(n9719), .A2(n9718), .A3(n9717), .A4(n9716), .ZN(n14173) );
  NAND2_X1 U12123 ( .A1(n9742), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9721) );
  XNOR2_X1 U12124 ( .A(n9721), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U12125 ( .A1(n10039), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10177), 
        .B2(n10593), .ZN(n9722) );
  MUX2_X1 U12126 ( .A(n14173), .B(n11978), .S(n10075), .Z(n9727) );
  NAND2_X1 U12127 ( .A1(n9726), .A2(n9727), .ZN(n9725) );
  MUX2_X1 U12128 ( .A(n14173), .B(n11978), .S(n9858), .Z(n9724) );
  NAND2_X1 U12129 ( .A1(n9725), .A2(n9724), .ZN(n9731) );
  INV_X1 U12130 ( .A(n9727), .ZN(n9728) );
  NAND2_X1 U12131 ( .A1(n9729), .A2(n9728), .ZN(n9730) );
  NAND2_X1 U12132 ( .A1(n10013), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9741) );
  INV_X1 U12133 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9732) );
  OAI21_X1 U12134 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9737) );
  INV_X1 U12135 ( .A(n9734), .ZN(n9736) );
  AND2_X1 U12136 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n9735) );
  NAND2_X1 U12137 ( .A1(n9737), .A2(n9750), .ZN(n12228) );
  OR2_X1 U12138 ( .A1(n6689), .A2(n12228), .ZN(n9740) );
  INV_X1 U12139 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10594) );
  OR2_X1 U12140 ( .A1(n10018), .A2(n10594), .ZN(n9739) );
  INV_X1 U12141 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11846) );
  OR2_X1 U12142 ( .A1(n10020), .A2(n11846), .ZN(n9738) );
  NAND4_X1 U12143 ( .A1(n9741), .A2(n9740), .A3(n9739), .A4(n9738), .ZN(n14172) );
  NAND2_X1 U12144 ( .A1(n10234), .A2(n10038), .ZN(n9745) );
  OAI21_X1 U12145 ( .B1(n9742), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9743) );
  XNOR2_X1 U12146 ( .A(n9743), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U12147 ( .A1(n10039), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10937), 
        .B2(n10177), .ZN(n9744) );
  NAND2_X1 U12148 ( .A1(n9745), .A2(n9744), .ZN(n12230) );
  MUX2_X1 U12149 ( .A(n14172), .B(n12230), .S(n9858), .Z(n9747) );
  MUX2_X1 U12150 ( .A(n14172), .B(n12230), .S(n10075), .Z(n9746) );
  INV_X1 U12151 ( .A(n9747), .ZN(n9748) );
  NAND2_X1 U12152 ( .A1(n10013), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9756) );
  INV_X1 U12153 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12094) );
  OR2_X1 U12154 ( .A1(n10020), .A2(n12094), .ZN(n9755) );
  INV_X1 U12155 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U12156 ( .A1(n9750), .A2(n9749), .ZN(n9751) );
  NAND2_X1 U12157 ( .A1(n9767), .A2(n9751), .ZN(n12275) );
  OR2_X1 U12158 ( .A1(n6689), .A2(n12275), .ZN(n9754) );
  INV_X1 U12159 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9752) );
  OR2_X1 U12160 ( .A1(n10018), .A2(n9752), .ZN(n9753) );
  NAND4_X1 U12161 ( .A1(n9756), .A2(n9755), .A3(n9754), .A4(n9753), .ZN(n14171) );
  NAND2_X1 U12162 ( .A1(n10353), .A2(n10038), .ZN(n9760) );
  NAND2_X1 U12163 ( .A1(n9757), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9758) );
  XNOR2_X1 U12164 ( .A(n9758), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U12165 ( .A1(n10039), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10177), 
        .B2(n11257), .ZN(n9759) );
  MUX2_X1 U12166 ( .A(n14171), .B(n14819), .S(n10075), .Z(n9763) );
  MUX2_X1 U12167 ( .A(n14171), .B(n14819), .S(n10011), .Z(n9761) );
  INV_X1 U12168 ( .A(n9763), .ZN(n9764) );
  NAND2_X1 U12169 ( .A1(n10013), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9772) );
  INV_X1 U12170 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12055) );
  OR2_X1 U12171 ( .A1(n10020), .A2(n12055), .ZN(n9771) );
  INV_X1 U12172 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9766) );
  NAND2_X1 U12173 ( .A1(n9767), .A2(n9766), .ZN(n9768) );
  NAND2_X1 U12174 ( .A1(n9784), .A2(n9768), .ZN(n12320) );
  OR2_X1 U12175 ( .A1(n6689), .A2(n12320), .ZN(n9770) );
  INV_X1 U12176 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11248) );
  OR2_X1 U12177 ( .A1(n6688), .A2(n11248), .ZN(n9769) );
  NAND4_X1 U12178 ( .A1(n9772), .A2(n9771), .A3(n9770), .A4(n9769), .ZN(n14170) );
  NAND2_X1 U12179 ( .A1(n10455), .A2(n10038), .ZN(n9775) );
  OR2_X1 U12180 ( .A1(n9757), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n9779) );
  NAND2_X1 U12181 ( .A1(n9779), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9773) );
  XNOR2_X1 U12182 ( .A(n9773), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U12183 ( .A1(n10039), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10177), 
        .B2(n11339), .ZN(n9774) );
  MUX2_X1 U12184 ( .A(n14170), .B(n14976), .S(n10011), .Z(n9777) );
  MUX2_X1 U12185 ( .A(n14170), .B(n14976), .S(n10075), .Z(n9776) );
  INV_X1 U12186 ( .A(n9777), .ZN(n9778) );
  NAND2_X1 U12187 ( .A1(n10913), .A2(n10038), .ZN(n9782) );
  NOR2_X1 U12188 ( .A1(n9779), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n9790) );
  OR2_X1 U12189 ( .A1(n9790), .A2(n14676), .ZN(n9780) );
  XNOR2_X1 U12190 ( .A(n9780), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U12191 ( .A1(n10039), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n10177), 
        .B2(n12018), .ZN(n9781) );
  NAND2_X1 U12192 ( .A1(n10013), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9789) );
  INV_X1 U12193 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12256) );
  OR2_X1 U12194 ( .A1(n10020), .A2(n12256), .ZN(n9788) );
  INV_X1 U12195 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9783) );
  NAND2_X1 U12196 ( .A1(n9784), .A2(n9783), .ZN(n9785) );
  NAND2_X1 U12197 ( .A1(n9797), .A2(n9785), .ZN(n12411) );
  OR2_X1 U12198 ( .A1(n6689), .A2(n12411), .ZN(n9787) );
  INV_X1 U12199 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11336) );
  OR2_X1 U12200 ( .A1(n10018), .A2(n11336), .ZN(n9786) );
  XNOR2_X1 U12201 ( .A(n14292), .B(n14155), .ZN(n12251) );
  INV_X1 U12202 ( .A(n14155), .ZN(n14291) );
  NAND2_X1 U12203 ( .A1(n11102), .A2(n10038), .ZN(n9793) );
  INV_X1 U12204 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n15827) );
  NAND2_X1 U12205 ( .A1(n9790), .A2(n15827), .ZN(n9845) );
  NAND2_X1 U12206 ( .A1(n9845), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9791) );
  XNOR2_X1 U12207 ( .A(n9791), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U12208 ( .A1(n10039), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10177), 
        .B2(n12027), .ZN(n9792) );
  NAND2_X1 U12209 ( .A1(n10012), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9803) );
  INV_X1 U12210 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9794) );
  OR2_X1 U12211 ( .A1(n10022), .A2(n9794), .ZN(n9802) );
  INV_X1 U12212 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9796) );
  NAND2_X1 U12213 ( .A1(n9797), .A2(n9796), .ZN(n9798) );
  NAND2_X1 U12214 ( .A1(n9837), .A2(n9798), .ZN(n14955) );
  OR2_X1 U12215 ( .A1(n6689), .A2(n14955), .ZN(n9801) );
  INV_X1 U12216 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9799) );
  OR2_X1 U12217 ( .A1(n10018), .A2(n9799), .ZN(n9800) );
  NAND2_X1 U12218 ( .A1(n14963), .A2(n14294), .ZN(n10048) );
  OAI21_X1 U12219 ( .B1(n7088), .B2(n14291), .A(n10048), .ZN(n9805) );
  OR2_X1 U12220 ( .A1(n14292), .A2(n14155), .ZN(n14324) );
  NAND2_X1 U12221 ( .A1(n14326), .A2(n14324), .ZN(n9804) );
  MUX2_X1 U12222 ( .A(n9805), .B(n9804), .S(n10011), .Z(n9807) );
  MUX2_X1 U12223 ( .A(n10048), .B(n14326), .S(n10075), .Z(n9806) );
  NAND2_X1 U12224 ( .A1(n11310), .A2(n10038), .ZN(n9815) );
  INV_X1 U12225 ( .A(n9809), .ZN(n9810) );
  NAND2_X1 U12226 ( .A1(n9810), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9812) );
  MUX2_X1 U12227 ( .A(n9812), .B(P1_IR_REG_31__SCAN_IN), .S(n9811), .Z(n9813)
         );
  NAND2_X1 U12228 ( .A1(n9813), .A2(n9821), .ZN(n14246) );
  INV_X1 U12229 ( .A(n14246), .ZN(n14249) );
  AOI22_X1 U12230 ( .A1(n10039), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10177), 
        .B2(n14249), .ZN(n9814) );
  NAND2_X1 U12231 ( .A1(n10013), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9820) );
  INV_X1 U12232 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9836) );
  INV_X1 U12233 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n14091) );
  INV_X1 U12234 ( .A(n9827), .ZN(n9829) );
  NAND2_X1 U12235 ( .A1(n9839), .A2(n14091), .ZN(n9816) );
  NAND2_X1 U12236 ( .A1(n9829), .A2(n9816), .ZN(n14542) );
  OR2_X1 U12237 ( .A1(n14542), .A2(n6689), .ZN(n9819) );
  INV_X1 U12238 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14227) );
  OR2_X1 U12239 ( .A1(n10020), .A2(n14227), .ZN(n9818) );
  INV_X1 U12240 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14235) );
  OR2_X1 U12241 ( .A1(n10018), .A2(n14235), .ZN(n9817) );
  NAND2_X1 U12242 ( .A1(n14650), .A2(n14132), .ZN(n9861) );
  NAND2_X1 U12243 ( .A1(n9821), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9823) );
  MUX2_X1 U12244 ( .A(n9823), .B(P1_IR_REG_31__SCAN_IN), .S(n9822), .Z(n9824)
         );
  NAND2_X1 U12245 ( .A1(n9824), .A2(n10093), .ZN(n14257) );
  INV_X1 U12246 ( .A(n14257), .ZN(n14263) );
  AOI22_X1 U12247 ( .A1(n10039), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10177), 
        .B2(n14263), .ZN(n9825) );
  INV_X1 U12248 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14251) );
  NAND2_X1 U12249 ( .A1(n9827), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9853) );
  INV_X1 U12250 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U12251 ( .A1(n9829), .A2(n9828), .ZN(n9830) );
  NAND2_X1 U12252 ( .A1(n9853), .A2(n9830), .ZN(n14530) );
  OR2_X1 U12253 ( .A1(n14530), .A2(n6689), .ZN(n9835) );
  INV_X1 U12254 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14531) );
  OR2_X1 U12255 ( .A1(n10020), .A2(n14531), .ZN(n9833) );
  INV_X1 U12256 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9831) );
  OR2_X1 U12257 ( .A1(n10022), .A2(n9831), .ZN(n9832) );
  AND2_X1 U12258 ( .A1(n9833), .A2(n9832), .ZN(n9834) );
  OAI211_X1 U12259 ( .C1(n6688), .C2(n14251), .A(n9835), .B(n9834), .ZN(n14330) );
  NAND2_X1 U12260 ( .A1(n10013), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9844) );
  INV_X1 U12261 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12030) );
  OR2_X1 U12262 ( .A1(n10020), .A2(n12030), .ZN(n9843) );
  NAND2_X1 U12263 ( .A1(n9837), .A2(n9836), .ZN(n9838) );
  NAND2_X1 U12264 ( .A1(n9839), .A2(n9838), .ZN(n14077) );
  OR2_X1 U12265 ( .A1(n6689), .A2(n14077), .ZN(n9842) );
  INV_X1 U12266 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9840) );
  OR2_X1 U12267 ( .A1(n10018), .A2(n9840), .ZN(n9841) );
  NAND2_X1 U12268 ( .A1(n11194), .A2(n10038), .ZN(n9848) );
  OAI21_X1 U12269 ( .B1(n9845), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9846) );
  XNOR2_X1 U12270 ( .A(n9846), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14234) );
  AOI22_X1 U12271 ( .A1(n10039), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10177), 
        .B2(n14234), .ZN(n9847) );
  MUX2_X1 U12272 ( .A(n14298), .B(n14562), .S(n10011), .Z(n9867) );
  INV_X1 U12273 ( .A(n14298), .ZN(n14327) );
  MUX2_X1 U12274 ( .A(n14327), .B(n14656), .S(n10075), .Z(n9866) );
  NAND2_X1 U12275 ( .A1(n9867), .A2(n9866), .ZN(n9849) );
  AOI22_X1 U12276 ( .A1(n10039), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14448), 
        .B2(n10177), .ZN(n9851) );
  INV_X1 U12277 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U12278 ( .A1(n9853), .A2(n9852), .ZN(n9854) );
  NAND2_X1 U12279 ( .A1(n9874), .A2(n9854), .ZN(n14509) );
  OR2_X1 U12280 ( .A1(n14509), .A2(n6689), .ZN(n9857) );
  AOI22_X1 U12281 ( .A1(n10012), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10013), 
        .B2(P1_REG0_REG_19__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U12282 ( .A1(n6669), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9855) );
  AND2_X2 U12283 ( .A1(n9872), .A2(n14333), .ZN(n14507) );
  INV_X1 U12284 ( .A(n14329), .ZN(n9859) );
  OAI211_X1 U12285 ( .C1(n9859), .C2(n14330), .A(n14529), .B(n10075), .ZN(
        n9865) );
  INV_X1 U12286 ( .A(n14330), .ZN(n14302) );
  INV_X1 U12287 ( .A(n9861), .ZN(n9860) );
  OAI211_X1 U12288 ( .C1(n14302), .C2(n9860), .A(n14646), .B(n10011), .ZN(
        n9864) );
  OR3_X1 U12289 ( .A1(n14329), .A2(n14302), .A3(n10011), .ZN(n9863) );
  OR3_X1 U12290 ( .A1(n9861), .A2(n9660), .A3(n14330), .ZN(n9862) );
  AND4_X1 U12291 ( .A1(n9865), .A2(n9864), .A3(n9863), .A4(n9862), .ZN(n9871)
         );
  INV_X1 U12292 ( .A(n9866), .ZN(n9869) );
  INV_X1 U12293 ( .A(n9867), .ZN(n9868) );
  NAND4_X1 U12294 ( .A1(n14520), .A2(n10047), .A3(n9869), .A4(n9868), .ZN(
        n9870) );
  INV_X1 U12295 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U12296 ( .A1(n9874), .A2(n14111), .ZN(n9875) );
  NAND2_X1 U12297 ( .A1(n9884), .A2(n9875), .ZN(n14493) );
  AOI22_X1 U12298 ( .A1(n10012), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10013), 
        .B2(P1_REG0_REG_20__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U12299 ( .A1(n6669), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9876) );
  OAI211_X1 U12300 ( .C1(n14493), .C2(n6689), .A(n9877), .B(n9876), .ZN(n14334) );
  INV_X1 U12301 ( .A(n14334), .ZN(n14309) );
  OR2_X1 U12302 ( .A1(n9997), .A2(n11673), .ZN(n9879) );
  MUX2_X1 U12303 ( .A(n14309), .B(n14634), .S(n10011), .Z(n9882) );
  MUX2_X1 U12304 ( .A(n14334), .B(n14499), .S(n10075), .Z(n9881) );
  INV_X1 U12305 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14058) );
  NAND2_X1 U12306 ( .A1(n9884), .A2(n14058), .ZN(n9885) );
  AND2_X1 U12307 ( .A1(n9900), .A2(n9885), .ZN(n14483) );
  INV_X1 U12308 ( .A(n6689), .ZN(n10009) );
  NAND2_X1 U12309 ( .A1(n14483), .A2(n10009), .ZN(n9892) );
  INV_X1 U12310 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U12311 ( .A1(n10012), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9888) );
  NAND2_X1 U12312 ( .A1(n10013), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9887) );
  OAI211_X1 U12313 ( .C1(n9889), .C2(n6688), .A(n9888), .B(n9887), .ZN(n9890)
         );
  INV_X1 U12314 ( .A(n9890), .ZN(n9891) );
  NAND2_X1 U12315 ( .A1(n9892), .A2(n9891), .ZN(n14336) );
  NAND2_X1 U12316 ( .A1(n11900), .A2(n10038), .ZN(n9894) );
  OR2_X1 U12317 ( .A1(n9997), .A2(n11903), .ZN(n9893) );
  MUX2_X1 U12318 ( .A(n14336), .B(n14484), .S(n10075), .Z(n9897) );
  MUX2_X1 U12319 ( .A(n14336), .B(n14484), .S(n10011), .Z(n9895) );
  INV_X1 U12320 ( .A(n9897), .ZN(n9898) );
  INV_X1 U12321 ( .A(n9900), .ZN(n9899) );
  NAND2_X1 U12322 ( .A1(n9899), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9919) );
  INV_X1 U12323 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14122) );
  NAND2_X1 U12324 ( .A1(n9900), .A2(n14122), .ZN(n9901) );
  NAND2_X1 U12325 ( .A1(n9919), .A2(n9901), .ZN(n14462) );
  OR2_X1 U12326 ( .A1(n14462), .A2(n6689), .ZN(n9907) );
  INV_X1 U12327 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U12328 ( .A1(n10012), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9903) );
  NAND2_X1 U12329 ( .A1(n10013), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9902) );
  OAI211_X1 U12330 ( .C1(n9904), .C2(n10018), .A(n9903), .B(n9902), .ZN(n9905)
         );
  INV_X1 U12331 ( .A(n9905), .ZN(n9906) );
  NAND2_X1 U12332 ( .A1(n9907), .A2(n9906), .ZN(n14311) );
  XNOR2_X1 U12333 ( .A(n9909), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14697) );
  MUX2_X1 U12334 ( .A(n14311), .B(n14461), .S(n10011), .Z(n9914) );
  MUX2_X1 U12335 ( .A(n14311), .B(n14461), .S(n10075), .Z(n9911) );
  NAND2_X1 U12336 ( .A1(n9912), .A2(n9911), .ZN(n9918) );
  INV_X1 U12337 ( .A(n9913), .ZN(n9916) );
  INV_X1 U12338 ( .A(n9914), .ZN(n9915) );
  INV_X1 U12339 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14015) );
  NAND2_X1 U12340 ( .A1(n9919), .A2(n14015), .ZN(n9920) );
  AND2_X1 U12341 ( .A1(n9934), .A2(n9920), .ZN(n14451) );
  NAND2_X1 U12342 ( .A1(n14451), .A2(n10009), .ZN(n9926) );
  INV_X1 U12343 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U12344 ( .A1(n10013), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12345 ( .A1(n10012), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9921) );
  OAI211_X1 U12346 ( .C1(n10018), .C2(n9923), .A(n9922), .B(n9921), .ZN(n9924)
         );
  INV_X1 U12347 ( .A(n9924), .ZN(n9925) );
  NAND2_X1 U12348 ( .A1(n9926), .A2(n9925), .ZN(n14313) );
  NAND2_X1 U12349 ( .A1(n12146), .A2(n10038), .ZN(n9928) );
  INV_X1 U12350 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12144) );
  OR2_X1 U12351 ( .A1(n9997), .A2(n12144), .ZN(n9927) );
  MUX2_X1 U12352 ( .A(n14313), .B(n14452), .S(n10075), .Z(n9930) );
  MUX2_X1 U12353 ( .A(n14313), .B(n14452), .S(n10011), .Z(n9929) );
  INV_X1 U12354 ( .A(n9930), .ZN(n9931) );
  NAND2_X1 U12355 ( .A1(n10039), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9932) );
  INV_X1 U12356 ( .A(n9934), .ZN(n9933) );
  NAND2_X1 U12357 ( .A1(n9933), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9945) );
  INV_X1 U12358 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14102) );
  NAND2_X1 U12359 ( .A1(n9934), .A2(n14102), .ZN(n9935) );
  NAND2_X1 U12360 ( .A1(n9945), .A2(n9935), .ZN(n14100) );
  OR2_X1 U12361 ( .A1(n14100), .A2(n6689), .ZN(n9941) );
  INV_X1 U12362 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U12363 ( .A1(n10012), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U12364 ( .A1(n10013), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9936) );
  OAI211_X1 U12365 ( .C1(n9938), .C2(n10018), .A(n9937), .B(n9936), .ZN(n9939)
         );
  INV_X1 U12366 ( .A(n9939), .ZN(n9940) );
  NAND2_X1 U12367 ( .A1(n9941), .A2(n9940), .ZN(n14169) );
  MUX2_X1 U12368 ( .A(n14169), .B(n14437), .S(n9660), .Z(n9942) );
  INV_X1 U12369 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14068) );
  NAND2_X1 U12370 ( .A1(n9945), .A2(n14068), .ZN(n9946) );
  AND2_X1 U12371 ( .A1(n9961), .A2(n9946), .ZN(n14419) );
  NAND2_X1 U12372 ( .A1(n14419), .A2(n10009), .ZN(n9952) );
  INV_X1 U12373 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U12374 ( .A1(n10013), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12375 ( .A1(n10012), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9947) );
  OAI211_X1 U12376 ( .C1(n9949), .C2(n10018), .A(n9948), .B(n9947), .ZN(n9950)
         );
  INV_X1 U12377 ( .A(n9950), .ZN(n9951) );
  NAND2_X1 U12378 ( .A1(n9952), .A2(n9951), .ZN(n14321) );
  NAND2_X1 U12379 ( .A1(n13890), .A2(n10038), .ZN(n9954) );
  OR2_X1 U12380 ( .A1(n9997), .A2(n14692), .ZN(n9953) );
  MUX2_X1 U12381 ( .A(n14321), .B(n14420), .S(n10075), .Z(n9957) );
  MUX2_X1 U12382 ( .A(n14420), .B(n14321), .S(n10075), .Z(n9955) );
  NAND2_X1 U12383 ( .A1(n9956), .A2(n9955), .ZN(n9959) );
  INV_X1 U12384 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14146) );
  NAND2_X1 U12385 ( .A1(n9961), .A2(n14146), .ZN(n9962) );
  NAND2_X1 U12386 ( .A1(n9989), .A2(n9962), .ZN(n14403) );
  OR2_X1 U12387 ( .A1(n14403), .A2(n6689), .ZN(n9968) );
  INV_X1 U12388 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U12389 ( .A1(n10012), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U12390 ( .A1(n10013), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9963) );
  OAI211_X1 U12391 ( .C1(n9965), .C2(n10018), .A(n9964), .B(n9963), .ZN(n9966)
         );
  INV_X1 U12392 ( .A(n9966), .ZN(n9967) );
  NAND2_X1 U12393 ( .A1(n9968), .A2(n9967), .ZN(n14342) );
  NAND2_X1 U12394 ( .A1(n13887), .A2(n10038), .ZN(n9970) );
  INV_X1 U12395 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14687) );
  OR2_X1 U12396 ( .A1(n9997), .A2(n14687), .ZN(n9969) );
  MUX2_X1 U12397 ( .A(n14342), .B(n14596), .S(n10011), .Z(n9973) );
  MUX2_X1 U12398 ( .A(n14596), .B(n14342), .S(n9858), .Z(n9971) );
  XNOR2_X1 U12399 ( .A(n9989), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n14387) );
  NAND2_X1 U12400 ( .A1(n14387), .A2(n10009), .ZN(n9979) );
  INV_X1 U12401 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U12402 ( .A1(n10012), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U12403 ( .A1(n10013), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9974) );
  OAI211_X1 U12404 ( .C1(n9976), .C2(n10018), .A(n9975), .B(n9974), .ZN(n9977)
         );
  INV_X1 U12405 ( .A(n9977), .ZN(n9978) );
  NAND2_X1 U12406 ( .A1(n12457), .A2(n10038), .ZN(n9981) );
  OR2_X1 U12407 ( .A1(n9997), .A2(n14685), .ZN(n9980) );
  MUX2_X1 U12408 ( .A(n14344), .B(n14589), .S(n9660), .Z(n9983) );
  MUX2_X1 U12409 ( .A(n14344), .B(n14589), .S(n9858), .Z(n9982) );
  INV_X1 U12410 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9987) );
  INV_X1 U12411 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9986) );
  OAI21_X1 U12412 ( .B1(n9989), .B2(n9987), .A(n9986), .ZN(n9990) );
  NAND2_X1 U12413 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9988) );
  NAND2_X1 U12414 ( .A1(n14371), .A2(n10009), .ZN(n9996) );
  INV_X1 U12415 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U12416 ( .A1(n10012), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9992) );
  NAND2_X1 U12417 ( .A1(n10013), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9991) );
  OAI211_X1 U12418 ( .C1(n9993), .C2(n10018), .A(n9992), .B(n9991), .ZN(n9994)
         );
  INV_X1 U12419 ( .A(n9994), .ZN(n9995) );
  NAND2_X1 U12420 ( .A1(n12446), .A2(n10038), .ZN(n9999) );
  INV_X1 U12421 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12447) );
  OR2_X1 U12422 ( .A1(n9997), .A2(n12447), .ZN(n9998) );
  NAND2_X4 U12423 ( .A1(n9999), .A2(n9998), .ZN(n14583) );
  MUX2_X1 U12424 ( .A(n14346), .B(n14583), .S(n10011), .Z(n10000) );
  MUX2_X1 U12425 ( .A(n14583), .B(n14346), .S(n9858), .Z(n10002) );
  INV_X1 U12426 ( .A(n10000), .ZN(n10001) );
  NAND2_X1 U12427 ( .A1(n12443), .A2(n10038), .ZN(n10004) );
  NAND2_X1 U12428 ( .A1(n10039), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n10003) );
  INV_X1 U12429 ( .A(n14355), .ZN(n10010) );
  INV_X1 U12430 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U12431 ( .A1(n10012), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n10006) );
  NAND2_X1 U12432 ( .A1(n10013), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n10005) );
  OAI211_X1 U12433 ( .C1(n10007), .C2(n10018), .A(n10006), .B(n10005), .ZN(
        n10008) );
  AOI21_X1 U12434 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(n10043) );
  MUX2_X1 U12435 ( .A(n14361), .B(n10043), .S(n10011), .Z(n10030) );
  INV_X1 U12436 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U12437 ( .A1(n10012), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U12438 ( .A1(n10013), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n10014) );
  OAI211_X1 U12439 ( .C1(n10018), .C2(n10016), .A(n10015), .B(n10014), .ZN(
        n14283) );
  NAND2_X1 U12440 ( .A1(n10540), .A2(n10728), .ZN(n10090) );
  INV_X1 U12441 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10017) );
  OR2_X1 U12442 ( .A1(n10018), .A2(n10017), .ZN(n10025) );
  INV_X1 U12443 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10019) );
  OR2_X1 U12444 ( .A1(n10020), .A2(n10019), .ZN(n10024) );
  INV_X1 U12445 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10021) );
  OR2_X1 U12446 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  AND3_X1 U12447 ( .A1(n10025), .A2(n10024), .A3(n10023), .ZN(n14352) );
  INV_X1 U12448 ( .A(n14352), .ZN(n14167) );
  OAI21_X1 U12449 ( .B1(n14283), .B2(n10090), .A(n14167), .ZN(n10026) );
  MUX2_X1 U12450 ( .A(n10026), .B(n14573), .S(n9660), .Z(n10031) );
  AOI22_X1 U12451 ( .A1(n9660), .A2(n14283), .B1(n11905), .B2(n10027), .ZN(
        n10028) );
  OAI22_X1 U12452 ( .A1(n14573), .A2(n9660), .B1(n14352), .B2(n10028), .ZN(
        n10032) );
  INV_X1 U12453 ( .A(n10043), .ZN(n14168) );
  MUX2_X1 U12454 ( .A(n14576), .B(n14168), .S(n10075), .Z(n10029) );
  INV_X1 U12455 ( .A(n10031), .ZN(n10034) );
  INV_X1 U12456 ( .A(n10032), .ZN(n10033) );
  NAND2_X1 U12457 ( .A1(n14696), .A2(n10540), .ZN(n10552) );
  NAND2_X1 U12458 ( .A1(n10035), .A2(n11674), .ZN(n10036) );
  NAND2_X1 U12459 ( .A1(n10552), .A2(n10036), .ZN(n10037) );
  OR2_X1 U12460 ( .A1(n10725), .A2(n14511), .ZN(n11668) );
  NAND2_X1 U12461 ( .A1(n10037), .A2(n11668), .ZN(n10073) );
  INV_X1 U12462 ( .A(n10073), .ZN(n10042) );
  NAND2_X1 U12463 ( .A1(n13876), .A2(n10038), .ZN(n10041) );
  NAND2_X1 U12464 ( .A1(n10039), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10040) );
  INV_X1 U12465 ( .A(n14283), .ZN(n10074) );
  XNOR2_X1 U12466 ( .A(n14573), .B(n14167), .ZN(n10068) );
  INV_X1 U12467 ( .A(n14344), .ZN(n10044) );
  NAND2_X1 U12468 ( .A1(n14583), .A2(n14346), .ZN(n14319) );
  NAND2_X1 U12469 ( .A1(n14435), .A2(n14169), .ZN(n14340) );
  INV_X1 U12470 ( .A(n14169), .ZN(n14315) );
  NAND2_X1 U12471 ( .A1(n14437), .A2(n14315), .ZN(n10046) );
  NAND2_X1 U12472 ( .A1(n14340), .A2(n10046), .ZN(n14432) );
  INV_X1 U12473 ( .A(n14313), .ZN(n14339) );
  XNOR2_X1 U12474 ( .A(n14452), .B(n14339), .ZN(n14442) );
  INV_X1 U12475 ( .A(n14311), .ZN(n14337) );
  NAND2_X1 U12476 ( .A1(n14326), .A2(n10048), .ZN(n14961) );
  INV_X1 U12477 ( .A(n14170), .ZN(n12253) );
  XNOR2_X1 U12478 ( .A(n14976), .B(n12253), .ZN(n12246) );
  INV_X1 U12479 ( .A(n14171), .ZN(n12042) );
  XNOR2_X1 U12480 ( .A(n12230), .B(n14172), .ZN(n12036) );
  INV_X1 U12481 ( .A(n14173), .ZN(n10049) );
  NAND2_X1 U12482 ( .A1(n11978), .A2(n10049), .ZN(n10050) );
  INV_X1 U12483 ( .A(n14175), .ZN(n11734) );
  XNOR2_X1 U12484 ( .A(n11879), .B(n11734), .ZN(n11744) );
  AND2_X1 U12485 ( .A1(n10051), .A2(n7058), .ZN(n11464) );
  NAND4_X1 U12486 ( .A1(n11493), .A2(n11529), .A3(n11464), .A4(n11658), .ZN(
        n10055) );
  XNOR2_X1 U12487 ( .A(n10054), .B(n15167), .ZN(n11496) );
  NOR2_X1 U12488 ( .A1(n10055), .A2(n11496), .ZN(n10056) );
  XNOR2_X1 U12489 ( .A(n15193), .B(n14176), .ZN(n15071) );
  XNOR2_X1 U12490 ( .A(n14177), .B(n11637), .ZN(n11479) );
  XNOR2_X1 U12491 ( .A(n14178), .B(n11556), .ZN(n11542) );
  NAND4_X1 U12492 ( .A1(n10056), .A2(n15071), .A3(n11479), .A4(n11542), .ZN(
        n10057) );
  NOR2_X1 U12493 ( .A1(n11744), .A2(n10057), .ZN(n10058) );
  XNOR2_X1 U12494 ( .A(n11912), .B(n14174), .ZN(n11737) );
  NAND4_X1 U12495 ( .A1(n12036), .A2(n11747), .A3(n10058), .A4(n11737), .ZN(
        n10059) );
  OR3_X1 U12496 ( .A1(n12246), .A2(n12086), .A3(n10059), .ZN(n10060) );
  OR3_X1 U12497 ( .A1(n14961), .A2(n12251), .A3(n10060), .ZN(n10061) );
  NOR2_X1 U12498 ( .A1(n14546), .A2(n10061), .ZN(n10062) );
  XNOR2_X1 U12499 ( .A(n14656), .B(n14327), .ZN(n14563) );
  NAND3_X1 U12500 ( .A1(n14520), .A2(n10062), .A3(n14563), .ZN(n10063) );
  NOR2_X1 U12501 ( .A1(n14332), .A2(n10063), .ZN(n10064) );
  XNOR2_X1 U12502 ( .A(n14499), .B(n14334), .ZN(n14500) );
  XNOR2_X1 U12503 ( .A(n14484), .B(n14336), .ZN(n14477) );
  NAND4_X1 U12504 ( .A1(n14338), .A2(n10064), .A3(n14500), .A4(n14477), .ZN(
        n10065) );
  NOR3_X1 U12505 ( .A1(n14432), .A2(n14442), .A3(n10065), .ZN(n10066) );
  XNOR2_X1 U12506 ( .A(n14420), .B(n14321), .ZN(n14424) );
  XNOR2_X1 U12507 ( .A(n14596), .B(n14342), .ZN(n14317) );
  NAND4_X1 U12508 ( .A1(n14375), .A2(n10066), .A3(n14424), .A4(n14317), .ZN(
        n10067) );
  NOR4_X1 U12509 ( .A1(n10068), .A2(n14348), .A3(n14379), .A4(n10067), .ZN(
        n10069) );
  NAND2_X1 U12510 ( .A1(n10069), .A2(n6720), .ZN(n10070) );
  XOR2_X1 U12511 ( .A(n14448), .B(n10070), .Z(n10071) );
  NAND2_X1 U12512 ( .A1(n11905), .A2(n10728), .ZN(n10072) );
  NOR2_X1 U12513 ( .A1(n10071), .A2(n10072), .ZN(n10081) );
  NAND2_X1 U12514 ( .A1(n10073), .A2(n10072), .ZN(n10082) );
  NOR2_X1 U12515 ( .A1(n6720), .A2(n10082), .ZN(n10079) );
  NOR2_X1 U12516 ( .A1(n14284), .A2(n10074), .ZN(n10077) );
  AND2_X1 U12517 ( .A1(n14284), .A2(n10074), .ZN(n10076) );
  MUX2_X1 U12518 ( .A(n10077), .B(n10076), .S(n10075), .Z(n10083) );
  INV_X1 U12519 ( .A(n10083), .ZN(n10078) );
  MUX2_X1 U12520 ( .A(n10042), .B(n10079), .S(n10078), .Z(n10080) );
  OAI21_X1 U12521 ( .B1(n10085), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10087) );
  XNOR2_X1 U12522 ( .A(n10087), .B(n10086), .ZN(n10178) );
  INV_X1 U12523 ( .A(n10178), .ZN(n10088) );
  NAND2_X1 U12524 ( .A1(n10088), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12142) );
  NAND2_X1 U12525 ( .A1(n14696), .A2(n14448), .ZN(n10091) );
  INV_X1 U12526 ( .A(n10552), .ZN(n10179) );
  NAND2_X1 U12527 ( .A1(n15189), .A2(n10179), .ZN(n10553) );
  NAND2_X1 U12528 ( .A1(n10098), .A2(n10094), .ZN(n10101) );
  NAND2_X1 U12529 ( .A1(n10101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10095) );
  MUX2_X1 U12530 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10095), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n10097) );
  INV_X1 U12531 ( .A(n10098), .ZN(n10099) );
  NAND2_X1 U12532 ( .A1(n10099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U12533 ( .A1(n10096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10103) );
  MUX2_X1 U12534 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10103), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n10105) );
  NAND2_X1 U12535 ( .A1(n10105), .A2(n10104), .ZN(n14689) );
  NAND2_X1 U12536 ( .A1(n10553), .A2(n10546), .ZN(n11266) );
  NAND2_X1 U12537 ( .A1(n10178), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10244) );
  NOR2_X1 U12538 ( .A1(n11266), .A2(n10244), .ZN(n10735) );
  INV_X1 U12539 ( .A(n15020), .ZN(n14279) );
  INV_X1 U12540 ( .A(n10107), .ZN(n14197) );
  NAND3_X1 U12541 ( .A1(n10735), .A2(n14279), .A3(n14521), .ZN(n10108) );
  OAI211_X1 U12542 ( .C1(n14696), .C2(n12142), .A(n10108), .B(P1_B_REG_SCAN_IN), .ZN(n10109) );
  INV_X1 U12543 ( .A(n13356), .ZN(P2_U3947) );
  INV_X1 U12544 ( .A(n13235), .ZN(n10111) );
  INV_X1 U12545 ( .A(n11368), .ZN(P3_U3897) );
  INV_X2 U12546 ( .A(n14903), .ZN(n13342) );
  INV_X1 U12547 ( .A(n10112), .ZN(n10692) );
  AOI211_X1 U12548 ( .C1(n10114), .C2(n10113), .A(n13342), .B(n10692), .ZN(
        n10119) );
  MUX2_X1 U12549 ( .A(n13337), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n10118) );
  INV_X1 U12550 ( .A(n10580), .ZN(n11221) );
  INV_X1 U12551 ( .A(n14908), .ZN(n13330) );
  INV_X1 U12552 ( .A(n13362), .ZN(n10651) );
  INV_X1 U12553 ( .A(n13363), .ZN(n10115) );
  OAI22_X1 U12554 ( .A1(n10651), .A2(n13326), .B1(n10115), .B2(n13544), .ZN(
        n10472) );
  INV_X1 U12555 ( .A(n10472), .ZN(n10116) );
  OAI22_X1 U12556 ( .A1(n11221), .A2(n13330), .B1(n10116), .B2(n13339), .ZN(
        n10117) );
  OR3_X1 U12557 ( .A1(n10119), .A2(n10118), .A3(n10117), .ZN(P2_U3190) );
  MUX2_X1 U12558 ( .A(P2_RD_REG_SCAN_IN), .B(n7804), .S(P1_RD_REG_SCAN_IN), 
        .Z(n10120) );
  INV_X1 U12559 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15886) );
  NAND2_X1 U12560 ( .A1(n10120), .A2(n15886), .ZN(U29) );
  AND2_X1 U12561 ( .A1(n10154), .A2(P1_U3086), .ZN(n14679) );
  INV_X2 U12562 ( .A(n14679), .ZN(n14691) );
  AND2_X1 U12563 ( .A1(n10153), .A2(P1_U3086), .ZN(n12141) );
  INV_X2 U12564 ( .A(n12141), .ZN(n14694) );
  INV_X1 U12565 ( .A(n14188), .ZN(n10121) );
  OAI222_X1 U12566 ( .A1(n14691), .A2(n10122), .B1(n14694), .B2(n10181), .C1(
        P1_U3086), .C2(n10121), .ZN(P1_U3354) );
  AND2_X1 U12567 ( .A1(n10123), .A2(P3_U3151), .ZN(n11561) );
  NAND2_X1 U12568 ( .A1(n10154), .A2(P3_U3151), .ZN(n13251) );
  OAI222_X1 U12569 ( .A1(n6670), .A2(n10124), .B1(n13251), .B2(n15789), .C1(
        n11157), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12570 ( .A1(n6670), .A2(n10126), .B1(n13251), .B2(n10125), .C1(
        n10953), .C2(P3_U3151), .ZN(P3_U3288) );
  OAI222_X1 U12571 ( .A1(n6670), .A2(n10127), .B1(n13251), .B2(n15867), .C1(
        n7463), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12572 ( .A(n10289), .ZN(n14208) );
  INV_X1 U12573 ( .A(n10128), .ZN(n10166) );
  OAI222_X1 U12574 ( .A1(P1_U3086), .A2(n14208), .B1(n14694), .B2(n10166), 
        .C1(n10129), .C2(n14691), .ZN(P1_U3353) );
  INV_X1 U12575 ( .A(n10293), .ZN(n10389) );
  OAI222_X1 U12576 ( .A1(P1_U3086), .A2(n10389), .B1(n14694), .B2(n10157), 
        .C1(n10130), .C2(n14691), .ZN(P1_U3350) );
  INV_X1 U12577 ( .A(n15038), .ZN(n10292) );
  OAI222_X1 U12578 ( .A1(P1_U3086), .A2(n10292), .B1(n14694), .B2(n10155), 
        .C1(n10131), .C2(n14691), .ZN(P1_U3351) );
  INV_X1 U12579 ( .A(n10964), .ZN(n10793) );
  INV_X1 U12580 ( .A(n10132), .ZN(n10133) );
  OAI222_X1 U12581 ( .A1(n10793), .A2(P3_U3151), .B1(n6670), .B2(n10133), .C1(
        n15843), .C2(n13251), .ZN(P3_U3289) );
  INV_X1 U12582 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10507) );
  INV_X1 U12583 ( .A(n10134), .ZN(n10136) );
  OAI222_X1 U12584 ( .A1(n10507), .A2(P3_U3151), .B1(n6670), .B2(n10136), .C1(
        n10135), .C2(n13251), .ZN(P3_U3295) );
  INV_X1 U12585 ( .A(n14218), .ZN(n10139) );
  INV_X1 U12586 ( .A(n10137), .ZN(n10163) );
  OAI222_X1 U12587 ( .A1(P1_U3086), .A2(n10139), .B1(n14694), .B2(n10163), 
        .C1(n10138), .C2(n14691), .ZN(P1_U3352) );
  INV_X1 U12588 ( .A(SI_8_), .ZN(n15800) );
  OAI222_X1 U12589 ( .A1(P3_U3151), .A2(n11165), .B1(n13251), .B2(n15800), 
        .C1(n6670), .C2(n10140), .ZN(P3_U3287) );
  INV_X1 U12590 ( .A(n10358), .ZN(n10363) );
  OAI222_X1 U12591 ( .A1(P1_U3086), .A2(n10363), .B1(n14694), .B2(n10160), 
        .C1(n10141), .C2(n14691), .ZN(P1_U3349) );
  NOR2_X1 U12592 ( .A1(n15328), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U12593 ( .A(n13251), .ZN(n13240) );
  INV_X1 U12594 ( .A(n13240), .ZN(n12166) );
  OAI222_X1 U12595 ( .A1(n6670), .A2(n10142), .B1(n12166), .B2(n7067), .C1(
        n10783), .C2(P3_U3151), .ZN(P3_U3292) );
  OAI222_X1 U12596 ( .A1(n6670), .A2(n10143), .B1(n12166), .B2(n15586), .C1(
        n10787), .C2(P3_U3151), .ZN(P3_U3291) );
  OAI222_X1 U12597 ( .A1(n6670), .A2(n10145), .B1(n12166), .B2(n10144), .C1(
        n10780), .C2(P3_U3151), .ZN(P3_U3293) );
  INV_X1 U12598 ( .A(n10508), .ZN(n10524) );
  INV_X1 U12599 ( .A(SI_1_), .ZN(n15612) );
  OAI222_X1 U12600 ( .A1(P3_U3151), .A2(n10524), .B1(n12166), .B2(n15612), 
        .C1(n6670), .C2(n10146), .ZN(P3_U3294) );
  OAI222_X1 U12601 ( .A1(n6670), .A2(n10147), .B1(n12166), .B2(n15823), .C1(
        n11727), .C2(P3_U3151), .ZN(P3_U3285) );
  OAI222_X1 U12602 ( .A1(n6670), .A2(n10149), .B1(n12166), .B2(n10148), .C1(
        n11957), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12603 ( .A(n10414), .ZN(n10371) );
  OAI222_X1 U12604 ( .A1(P1_U3086), .A2(n10371), .B1(n14694), .B2(n10174), 
        .C1(n10150), .C2(n14691), .ZN(P1_U3348) );
  OAI222_X1 U12605 ( .A1(n6670), .A2(n10151), .B1(n12183), .B2(P3_U3151), .C1(
        n15814), .C2(n13251), .ZN(P3_U3283) );
  OAI222_X1 U12606 ( .A1(P1_U3086), .A2(n10441), .B1(n14694), .B2(n10168), 
        .C1(n10152), .C2(n14691), .ZN(P1_U3347) );
  NAND2_X1 U12607 ( .A1(n10154), .A2(P2_U3088), .ZN(n13892) );
  INV_X1 U12608 ( .A(n13892), .ZN(n12145) );
  INV_X1 U12609 ( .A(n12145), .ZN(n13883) );
  OAI222_X1 U12610 ( .A1(n13894), .A2(n10247), .B1(n13883), .B2(n10155), .C1(
        n15249), .C2(P2_U3088), .ZN(P2_U3323) );
  INV_X1 U12611 ( .A(n13399), .ZN(n10156) );
  OAI222_X1 U12612 ( .A1(n13894), .A2(n10158), .B1(n13883), .B2(n10157), .C1(
        n10156), .C2(P2_U3088), .ZN(P2_U3322) );
  INV_X1 U12613 ( .A(n13410), .ZN(n10159) );
  OAI222_X1 U12614 ( .A1(n13894), .A2(n10161), .B1(n13883), .B2(n10160), .C1(
        n10159), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U12615 ( .A(n13386), .ZN(n10162) );
  OAI222_X1 U12616 ( .A1(n13894), .A2(n10164), .B1(n13883), .B2(n10163), .C1(
        n10162), .C2(P2_U3088), .ZN(P2_U3324) );
  INV_X1 U12617 ( .A(n15239), .ZN(n10165) );
  OAI222_X1 U12618 ( .A1(n13894), .A2(n10167), .B1(n13883), .B2(n10166), .C1(
        n10165), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U12619 ( .A(n13438), .ZN(n10315) );
  OAI222_X1 U12620 ( .A1(n13894), .A2(n10169), .B1(n13883), .B2(n10168), .C1(
        n10315), .C2(P2_U3088), .ZN(P2_U3319) );
  OAI222_X1 U12621 ( .A1(n13894), .A2(n10170), .B1(n13883), .B2(n10172), .C1(
        n10339), .C2(P2_U3088), .ZN(P2_U3318) );
  INV_X1 U12622 ( .A(n10484), .ZN(n10449) );
  OAI222_X1 U12623 ( .A1(P1_U3086), .A2(n10449), .B1(n14694), .B2(n10172), 
        .C1(n10171), .C2(n14691), .ZN(P1_U3346) );
  INV_X1 U12624 ( .A(n13424), .ZN(n10173) );
  OAI222_X1 U12625 ( .A1(n13894), .A2(n10175), .B1(n13892), .B2(n10174), .C1(
        n10173), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U12626 ( .A(n10546), .ZN(n10176) );
  OR2_X1 U12627 ( .A1(n11453), .A2(n10089), .ZN(n10277) );
  AOI21_X1 U12628 ( .B1(n10179), .B2(n10178), .A(n10177), .ZN(n10276) );
  INV_X1 U12629 ( .A(n10276), .ZN(n10180) );
  AND2_X1 U12630 ( .A1(n10277), .A2(n10180), .ZN(n15027) );
  NOR2_X1 U12631 ( .A1(n15027), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U12632 ( .A1(P2_U3088), .A2(n13368), .B1(n13894), .B2(n10232), 
        .C1(n13883), .C2(n10181), .ZN(P2_U3326) );
  OAI222_X1 U12633 ( .A1(n6670), .A2(n10183), .B1(n12166), .B2(n10182), .C1(
        n12714), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12634 ( .A(n10593), .ZN(n10490) );
  OAI222_X1 U12635 ( .A1(P1_U3086), .A2(n10490), .B1(n14694), .B2(n10185), 
        .C1(n10184), .C2(n14691), .ZN(P1_U3345) );
  INV_X1 U12636 ( .A(n10564), .ZN(n10348) );
  OAI222_X1 U12637 ( .A1(n13894), .A2(n10186), .B1(n13883), .B2(n10185), .C1(
        n10348), .C2(P2_U3088), .ZN(P2_U3317) );
  INV_X1 U12638 ( .A(n11933), .ZN(n13652) );
  NAND2_X1 U12639 ( .A1(n10188), .A2(n10187), .ZN(n10189) );
  INV_X1 U12640 ( .A(n11230), .ZN(n10430) );
  OAI21_X1 U12641 ( .B1(n13652), .B2(n14915), .A(n10430), .ZN(n10191) );
  INV_X1 U12642 ( .A(n13326), .ZN(n13336) );
  NAND2_X1 U12643 ( .A1(n13364), .A2(n13336), .ZN(n10433) );
  NAND2_X1 U12644 ( .A1(n10191), .A2(n10433), .ZN(n11233) );
  OAI22_X1 U12645 ( .A1(n11230), .A2(n15377), .B1(n10192), .B2(n7919), .ZN(
        n10193) );
  NOR2_X1 U12646 ( .A1(n11233), .A2(n10193), .ZN(n10253) );
  NAND4_X1 U12647 ( .A1(n11078), .A2(P2_STATE_REG_SCAN_IN), .A3(n10194), .A4(
        n11077), .ZN(n10249) );
  NAND2_X1 U12648 ( .A1(n15389), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10196) );
  OAI21_X1 U12649 ( .B1(n10253), .B2(n15389), .A(n10196), .ZN(P2_U3499) );
  XNOR2_X1 U12650 ( .A(n11899), .B(P3_B_REG_SCAN_IN), .ZN(n10197) );
  NAND2_X1 U12651 ( .A1(n10197), .A2(n12014), .ZN(n10198) );
  NOR2_X1 U12652 ( .A1(n13235), .A2(n10618), .ZN(n10201) );
  INV_X1 U12653 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10199) );
  NOR2_X1 U12654 ( .A1(n10230), .A2(n10199), .ZN(P3_U3244) );
  INV_X1 U12655 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U12656 ( .A1(n10230), .A2(n10200), .ZN(P3_U3243) );
  CLKBUF_X1 U12657 ( .A(n10201), .Z(n10230) );
  INV_X1 U12658 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10202) );
  NOR2_X1 U12659 ( .A1(n10230), .A2(n10202), .ZN(P3_U3261) );
  INV_X1 U12660 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10203) );
  NOR2_X1 U12661 ( .A1(n10230), .A2(n10203), .ZN(P3_U3242) );
  INV_X1 U12662 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10204) );
  NOR2_X1 U12663 ( .A1(n10201), .A2(n10204), .ZN(P3_U3260) );
  INV_X1 U12664 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10205) );
  NOR2_X1 U12665 ( .A1(n10201), .A2(n10205), .ZN(P3_U3245) );
  INV_X1 U12666 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10206) );
  NOR2_X1 U12667 ( .A1(n10201), .A2(n10206), .ZN(P3_U3239) );
  INV_X1 U12668 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10207) );
  NOR2_X1 U12669 ( .A1(n10201), .A2(n10207), .ZN(P3_U3238) );
  INV_X1 U12670 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U12671 ( .A1(n10201), .A2(n10208), .ZN(P3_U3235) );
  INV_X1 U12672 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10209) );
  NOR2_X1 U12673 ( .A1(n10230), .A2(n10209), .ZN(P3_U3263) );
  INV_X1 U12674 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U12675 ( .A1(n10201), .A2(n10210), .ZN(P3_U3262) );
  INV_X1 U12676 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U12677 ( .A1(n10201), .A2(n10211), .ZN(P3_U3241) );
  INV_X1 U12678 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U12679 ( .A1(n10201), .A2(n10212), .ZN(P3_U3237) );
  INV_X1 U12680 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U12681 ( .A1(n10201), .A2(n10213), .ZN(P3_U3236) );
  INV_X1 U12682 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U12683 ( .A1(n10201), .A2(n10214), .ZN(P3_U3234) );
  INV_X1 U12684 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U12685 ( .A1(n10201), .A2(n10215), .ZN(P3_U3240) );
  INV_X1 U12686 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10216) );
  NOR2_X1 U12687 ( .A1(n10230), .A2(n10216), .ZN(P3_U3258) );
  INV_X1 U12688 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U12689 ( .A1(n10230), .A2(n10217), .ZN(P3_U3257) );
  INV_X1 U12690 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U12691 ( .A1(n10230), .A2(n10218), .ZN(P3_U3256) );
  INV_X1 U12692 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U12693 ( .A1(n10230), .A2(n10219), .ZN(P3_U3255) );
  INV_X1 U12694 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U12695 ( .A1(n10230), .A2(n10220), .ZN(P3_U3254) );
  INV_X1 U12696 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U12697 ( .A1(n10230), .A2(n10221), .ZN(P3_U3253) );
  INV_X1 U12698 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U12699 ( .A1(n10230), .A2(n10222), .ZN(P3_U3252) );
  INV_X1 U12700 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U12701 ( .A1(n10230), .A2(n10223), .ZN(P3_U3247) );
  INV_X1 U12702 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U12703 ( .A1(n10230), .A2(n10224), .ZN(P3_U3246) );
  INV_X1 U12704 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U12705 ( .A1(n10230), .A2(n10225), .ZN(P3_U3249) );
  INV_X1 U12706 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U12707 ( .A1(n10230), .A2(n10226), .ZN(P3_U3248) );
  INV_X1 U12708 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10227) );
  NOR2_X1 U12709 ( .A1(n10230), .A2(n10227), .ZN(P3_U3250) );
  INV_X1 U12710 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10228) );
  NOR2_X1 U12711 ( .A1(n10230), .A2(n10228), .ZN(P3_U3259) );
  INV_X1 U12712 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10229) );
  NOR2_X1 U12713 ( .A1(n10230), .A2(n10229), .ZN(P3_U3251) );
  OAI222_X1 U12714 ( .A1(n6670), .A2(n10231), .B1(n13251), .B2(n15873), .C1(
        n12729), .C2(P3_U3151), .ZN(P3_U3281) );
  MUX2_X1 U12715 ( .A(n10232), .B(n11488), .S(P1_U4016), .Z(n10233) );
  INV_X1 U12716 ( .A(n10233), .ZN(P1_U3561) );
  INV_X1 U12717 ( .A(n10937), .ZN(n10933) );
  INV_X1 U12718 ( .A(n10234), .ZN(n10236) );
  OAI222_X1 U12719 ( .A1(n10933), .A2(P1_U3086), .B1(n14694), .B2(n10236), 
        .C1(n10235), .C2(n14691), .ZN(P1_U3344) );
  INV_X1 U12720 ( .A(n10831), .ZN(n10562) );
  OAI222_X1 U12721 ( .A1(n13894), .A2(n10237), .B1(n13883), .B2(n10236), .C1(
        P2_U3088), .C2(n10562), .ZN(P2_U3316) );
  INV_X1 U12722 ( .A(P1_B_REG_SCAN_IN), .ZN(n10239) );
  NOR2_X1 U12723 ( .A1(n14690), .A2(n10239), .ZN(n10238) );
  MUX2_X1 U12724 ( .A(n10239), .B(n10238), .S(n12426), .Z(n10240) );
  INV_X1 U12725 ( .A(n10240), .ZN(n10241) );
  INV_X1 U12726 ( .A(n14689), .ZN(n10242) );
  NAND2_X1 U12727 ( .A1(n10241), .A2(n10242), .ZN(n10539) );
  AND2_X2 U12728 ( .A1(n10539), .A2(n11453), .ZN(n15139) );
  OR2_X1 U12729 ( .A1(n14690), .A2(n10242), .ZN(n10525) );
  OAI22_X1 U12730 ( .A1(n15139), .A2(P1_D_REG_1__SCAN_IN), .B1(n10244), .B2(
        n10525), .ZN(n10243) );
  INV_X1 U12731 ( .A(n10243), .ZN(P1_U3446) );
  NAND2_X1 U12732 ( .A1(n12426), .A2(n14689), .ZN(n10527) );
  OAI22_X1 U12733 ( .A1(n15139), .A2(P1_D_REG_0__SCAN_IN), .B1(n10244), .B2(
        n10527), .ZN(n10245) );
  INV_X1 U12734 ( .A(n10245), .ZN(P1_U3445) );
  MUX2_X1 U12735 ( .A(n10914), .B(n14155), .S(P1_U4016), .Z(n10246) );
  INV_X1 U12736 ( .A(n10246), .ZN(P1_U3574) );
  MUX2_X1 U12737 ( .A(n10247), .B(n14023), .S(P1_U4016), .Z(n10248) );
  INV_X1 U12738 ( .A(n10248), .ZN(P1_U3564) );
  NAND2_X1 U12739 ( .A1(n11076), .A2(n15367), .ZN(n10250) );
  INV_X2 U12740 ( .A(n15386), .ZN(n15387) );
  INV_X1 U12741 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10251) );
  OR2_X1 U12742 ( .A1(n15387), .A2(n10251), .ZN(n10252) );
  OAI21_X1 U12743 ( .B1(n10253), .B2(n15386), .A(n10252), .ZN(P2_U3430) );
  MUX2_X1 U12744 ( .A(n11105), .B(n14294), .S(P1_U4016), .Z(n10254) );
  INV_X1 U12745 ( .A(n10254), .ZN(P1_U3575) );
  OAI222_X1 U12746 ( .A1(n6670), .A2(n10255), .B1(n13251), .B2(n15875), .C1(
        n12775), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12747 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U12748 ( .A1(n14833), .A2(n11422), .ZN(n10256) );
  OAI21_X1 U12749 ( .B1(n11422), .B2(n10257), .A(n10256), .ZN(P3_U3506) );
  INV_X1 U12750 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10264) );
  XOR2_X1 U12751 ( .A(n6697), .B(n10400), .Z(n11184) );
  NAND2_X1 U12752 ( .A1(n15377), .A2(n11933), .ZN(n14941) );
  INV_X1 U12753 ( .A(n10258), .ZN(n10399) );
  XNOR2_X1 U12754 ( .A(n10400), .B(n10399), .ZN(n11182) );
  NAND2_X1 U12755 ( .A1(n8582), .A2(n13307), .ZN(n10260) );
  NAND2_X1 U12756 ( .A1(n13363), .A2(n13336), .ZN(n10259) );
  NAND2_X1 U12757 ( .A1(n10260), .A2(n10259), .ZN(n10658) );
  INV_X1 U12758 ( .A(n8585), .ZN(n10659) );
  OR2_X1 U12759 ( .A1(n8585), .A2(n10428), .ZN(n10398) );
  OAI211_X1 U12760 ( .C1(n10659), .C2(n7919), .A(n14928), .B(n10398), .ZN(
        n11180) );
  OAI21_X1 U12761 ( .B1(n10659), .B2(n15381), .A(n11180), .ZN(n10261) );
  AOI211_X1 U12762 ( .C1(n11182), .C2(n14915), .A(n10658), .B(n10261), .ZN(
        n10262) );
  OAI21_X1 U12763 ( .B1(n11184), .B2(n13842), .A(n10262), .ZN(n10394) );
  NAND2_X1 U12764 ( .A1(n10394), .A2(n15387), .ZN(n10263) );
  OAI21_X1 U12765 ( .B1(n15387), .B2(n10264), .A(n10263), .ZN(P2_U3433) );
  INV_X2 U12766 ( .A(n11368), .ZN(n11422) );
  INV_X1 U12767 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n10267) );
  NAND2_X1 U12768 ( .A1(n10265), .A2(n11422), .ZN(n10266) );
  OAI21_X1 U12769 ( .B1(n11422), .B2(n10267), .A(n10266), .ZN(P3_U3496) );
  INV_X1 U12770 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n15889) );
  NAND2_X1 U12771 ( .A1(n12656), .A2(n11422), .ZN(n10268) );
  OAI21_X1 U12772 ( .B1(P3_U3897), .B2(n15889), .A(n10268), .ZN(P3_U3508) );
  INV_X1 U12773 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n15810) );
  NAND2_X1 U12774 ( .A1(n15397), .A2(n11422), .ZN(n10269) );
  OAI21_X1 U12775 ( .B1(P3_U3897), .B2(n15810), .A(n10269), .ZN(P3_U3500) );
  INV_X1 U12776 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n15610) );
  NAND2_X1 U12777 ( .A1(n15399), .A2(n11422), .ZN(n10270) );
  OAI21_X1 U12778 ( .B1(n11422), .B2(n15610), .A(n10270), .ZN(P3_U3498) );
  INV_X1 U12779 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n15850) );
  NAND2_X1 U12780 ( .A1(n11575), .A2(n11422), .ZN(n10271) );
  OAI21_X1 U12781 ( .B1(n11422), .B2(n15850), .A(n10271), .ZN(P3_U3494) );
  INV_X1 U12782 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n15834) );
  NAND2_X1 U12783 ( .A1(n14843), .A2(n11422), .ZN(n10272) );
  OAI21_X1 U12784 ( .B1(P3_U3897), .B2(n15834), .A(n10272), .ZN(P3_U3505) );
  INV_X1 U12785 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U12786 ( .A1(n14857), .A2(n11422), .ZN(n10273) );
  OAI21_X1 U12787 ( .B1(P3_U3897), .B2(n10274), .A(n10273), .ZN(P3_U3502) );
  INV_X1 U12788 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n15880) );
  NAND2_X1 U12789 ( .A1(n15448), .A2(n11422), .ZN(n10275) );
  OAI21_X1 U12790 ( .B1(P3_U3897), .B2(n15880), .A(n10275), .ZN(P3_U3491) );
  NAND2_X1 U12791 ( .A1(n10277), .A2(n10276), .ZN(n15030) );
  MUX2_X1 U12792 ( .A(n10278), .B(P1_REG1_REG_6__SCAN_IN), .S(n10358), .Z(
        n10284) );
  MUX2_X1 U12793 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9572), .S(n14188), .Z(
        n14185) );
  AND2_X1 U12794 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14184) );
  NAND2_X1 U12795 ( .A1(n14185), .A2(n14184), .ZN(n14183) );
  NAND2_X1 U12796 ( .A1(n14188), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U12797 ( .A1(n14183), .A2(n10279), .ZN(n14201) );
  XNOR2_X1 U12798 ( .A(n10289), .B(n10280), .ZN(n14202) );
  NAND2_X1 U12799 ( .A1(n14201), .A2(n14202), .ZN(n14200) );
  MUX2_X1 U12800 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9597), .S(n14218), .Z(
        n14213) );
  NAND2_X1 U12801 ( .A1(n14212), .A2(n14213), .ZN(n15033) );
  NAND2_X1 U12802 ( .A1(n14218), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n15031) );
  MUX2_X1 U12803 ( .A(n10281), .B(P1_REG1_REG_4__SCAN_IN), .S(n15038), .Z(
        n15032) );
  AOI21_X1 U12804 ( .B1(n15033), .B2(n15031), .A(n15032), .ZN(n15035) );
  MUX2_X1 U12805 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10282), .S(n10293), .Z(
        n10377) );
  OR2_X1 U12806 ( .A1(n15030), .A2(n14279), .ZN(n15036) );
  AOI211_X1 U12807 ( .C1(n10284), .C2(n10283), .A(n10357), .B(n15036), .ZN(
        n10298) );
  OR3_X1 U12808 ( .A1(n15030), .A2(n15020), .A3(n10107), .ZN(n15055) );
  MUX2_X1 U12809 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10285), .S(n14188), .Z(
        n14187) );
  AND2_X1 U12810 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10286) );
  NAND2_X1 U12811 ( .A1(n14187), .A2(n10286), .ZN(n14186) );
  NAND2_X1 U12812 ( .A1(n14188), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10287) );
  NAND2_X1 U12813 ( .A1(n14186), .A2(n10287), .ZN(n14203) );
  XNOR2_X1 U12814 ( .A(n10289), .B(n10288), .ZN(n14204) );
  AOI22_X1 U12815 ( .A1(n14203), .A2(n14204), .B1(n10289), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n14215) );
  MUX2_X1 U12816 ( .A(n14214), .B(P1_REG2_REG_3__SCAN_IN), .S(n14218), .Z(
        n10290) );
  OR2_X1 U12817 ( .A1(n14215), .A2(n10290), .ZN(n15043) );
  NAND2_X1 U12818 ( .A1(n14218), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n15042) );
  INV_X1 U12819 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10291) );
  MUX2_X1 U12820 ( .A(n10291), .B(P1_REG2_REG_4__SCAN_IN), .S(n15038), .Z(
        n15041) );
  AOI21_X1 U12821 ( .B1(n15043), .B2(n15042), .A(n15041), .ZN(n15040) );
  NOR2_X1 U12822 ( .A1(n10292), .A2(n10291), .ZN(n10381) );
  MUX2_X1 U12823 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11549), .S(n10293), .Z(
        n10380) );
  OAI21_X1 U12824 ( .B1(n15040), .B2(n10381), .A(n10380), .ZN(n10379) );
  NAND2_X1 U12825 ( .A1(n10293), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10295) );
  INV_X1 U12826 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10362) );
  MUX2_X1 U12827 ( .A(n10362), .B(P1_REG2_REG_6__SCAN_IN), .S(n10358), .Z(
        n10294) );
  AOI21_X1 U12828 ( .B1(n10379), .B2(n10295), .A(n10294), .ZN(n10367) );
  AND3_X1 U12829 ( .A1(n10379), .A2(n10295), .A3(n10294), .ZN(n10296) );
  NOR3_X1 U12830 ( .A1(n15055), .A2(n10367), .A3(n10296), .ZN(n10297) );
  NOR2_X1 U12831 ( .A1(n10298), .A2(n10297), .ZN(n10301) );
  NOR2_X1 U12832 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9648), .ZN(n10299) );
  AOI21_X1 U12833 ( .B1(n15027), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10299), .ZN(
        n10300) );
  OAI211_X1 U12834 ( .C1(n10363), .C2(n15064), .A(n10301), .B(n10300), .ZN(
        P1_U3249) );
  INV_X1 U12835 ( .A(n12778), .ZN(n12793) );
  OAI222_X1 U12836 ( .A1(n6670), .A2(n10302), .B1(n13251), .B2(n15595), .C1(
        n12793), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12837 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10303) );
  MUX2_X1 U12838 ( .A(n10303), .B(P2_REG1_REG_10__SCAN_IN), .S(n10564), .Z(
        n10319) );
  INV_X1 U12839 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10314) );
  MUX2_X1 U12840 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7961), .S(n13386), .Z(
        n13380) );
  MUX2_X1 U12841 ( .A(n7893), .B(P2_REG1_REG_1__SCAN_IN), .S(n13368), .Z(
        n13367) );
  AND2_X1 U12842 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13366) );
  NAND2_X1 U12843 ( .A1(n13367), .A2(n13366), .ZN(n13365) );
  INV_X1 U12844 ( .A(n13368), .ZN(n13373) );
  NAND2_X1 U12845 ( .A1(n13373), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U12846 ( .A1(n13365), .A2(n10304), .ZN(n15235) );
  XNOR2_X1 U12847 ( .A(n15239), .B(n10305), .ZN(n15236) );
  NAND2_X1 U12848 ( .A1(n15235), .A2(n15236), .ZN(n15234) );
  NAND2_X1 U12849 ( .A1(n15239), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10306) );
  NAND2_X1 U12850 ( .A1(n15234), .A2(n10306), .ZN(n13379) );
  NAND2_X1 U12851 ( .A1(n13380), .A2(n13379), .ZN(n13378) );
  NAND2_X1 U12852 ( .A1(n13386), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U12853 ( .A1(n13378), .A2(n10307), .ZN(n15247) );
  INV_X1 U12854 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10590) );
  MUX2_X1 U12855 ( .A(n10590), .B(P2_REG1_REG_4__SCAN_IN), .S(n15249), .Z(
        n15248) );
  NAND2_X1 U12856 ( .A1(n15247), .A2(n15248), .ZN(n15246) );
  OR2_X1 U12857 ( .A1(n15249), .A2(n10590), .ZN(n10308) );
  NAND2_X1 U12858 ( .A1(n15246), .A2(n10308), .ZN(n13392) );
  INV_X1 U12859 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10912) );
  MUX2_X1 U12860 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10912), .S(n13399), .Z(
        n13393) );
  NAND2_X1 U12861 ( .A1(n13392), .A2(n13393), .ZN(n13391) );
  NAND2_X1 U12862 ( .A1(n13399), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10309) );
  NAND2_X1 U12863 ( .A1(n13391), .A2(n10309), .ZN(n13408) );
  INV_X1 U12864 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10310) );
  MUX2_X1 U12865 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10310), .S(n13410), .Z(
        n13409) );
  NAND2_X1 U12866 ( .A1(n13408), .A2(n13409), .ZN(n13407) );
  NAND2_X1 U12867 ( .A1(n13410), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10311) );
  NAND2_X1 U12868 ( .A1(n13407), .A2(n10311), .ZN(n13422) );
  INV_X1 U12869 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10312) );
  MUX2_X1 U12870 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10312), .S(n13424), .Z(
        n13423) );
  NAND2_X1 U12871 ( .A1(n13422), .A2(n13423), .ZN(n13421) );
  NAND2_X1 U12872 ( .A1(n13424), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10313) );
  NAND2_X1 U12873 ( .A1(n13421), .A2(n10313), .ZN(n13436) );
  MUX2_X1 U12874 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10314), .S(n13438), .Z(
        n13437) );
  NAND2_X1 U12875 ( .A1(n13436), .A2(n13437), .ZN(n13435) );
  OAI21_X1 U12876 ( .B1(n10315), .B2(n10314), .A(n13435), .ZN(n15268) );
  INV_X1 U12877 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10316) );
  MUX2_X1 U12878 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10316), .S(n10339), .Z(
        n15267) );
  OAI21_X1 U12879 ( .B1(n15259), .B2(P2_REG1_REG_9__SCAN_IN), .A(n15265), .ZN(
        n10318) );
  OR2_X1 U12880 ( .A1(n10317), .A2(P2_U3088), .ZN(n10321) );
  NOR2_X1 U12881 ( .A1(n10321), .A2(n8626), .ZN(n10342) );
  NAND2_X1 U12882 ( .A1(n10342), .A2(n12458), .ZN(n15319) );
  NOR2_X1 U12883 ( .A1(n10318), .A2(n10319), .ZN(n10563) );
  AOI211_X1 U12884 ( .C1(n10319), .C2(n10318), .A(n15319), .B(n10563), .ZN(
        n10350) );
  NOR2_X2 U12885 ( .A1(n10321), .A2(n10320), .ZN(n15310) );
  INV_X1 U12886 ( .A(n15310), .ZN(n15325) );
  MUX2_X1 U12887 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11515), .S(n10339), .Z(
        n15263) );
  INV_X1 U12888 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11220) );
  MUX2_X1 U12889 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11220), .S(n13386), .Z(
        n10327) );
  INV_X1 U12890 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11176) );
  MUX2_X1 U12891 ( .A(n11176), .B(P2_REG2_REG_1__SCAN_IN), .S(n13368), .Z(
        n10323) );
  AND2_X1 U12892 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10322) );
  NAND2_X1 U12893 ( .A1(n10323), .A2(n10322), .ZN(n13372) );
  NAND2_X1 U12894 ( .A1(n13373), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10324) );
  NAND2_X1 U12895 ( .A1(n13372), .A2(n10324), .ZN(n15242) );
  INV_X1 U12896 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10325) );
  MUX2_X1 U12897 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10325), .S(n15239), .Z(
        n15241) );
  NAND2_X1 U12898 ( .A1(n15242), .A2(n15241), .ZN(n15240) );
  NAND2_X1 U12899 ( .A1(n15239), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13382) );
  NAND2_X1 U12900 ( .A1(n15240), .A2(n13382), .ZN(n10326) );
  NAND2_X1 U12901 ( .A1(n10327), .A2(n10326), .ZN(n13385) );
  NAND2_X1 U12902 ( .A1(n13386), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10328) );
  NAND2_X1 U12903 ( .A1(n13385), .A2(n10328), .ZN(n15255) );
  MUX2_X1 U12904 ( .A(n11199), .B(P2_REG2_REG_4__SCAN_IN), .S(n15249), .Z(
        n15254) );
  NAND2_X1 U12905 ( .A1(n15255), .A2(n15254), .ZN(n15253) );
  OR2_X1 U12906 ( .A1(n15249), .A2(n11199), .ZN(n13397) );
  NAND2_X1 U12907 ( .A1(n15253), .A2(n13397), .ZN(n10331) );
  MUX2_X1 U12908 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10329), .S(n13399), .Z(
        n10330) );
  NAND2_X1 U12909 ( .A1(n10331), .A2(n10330), .ZN(n13413) );
  NAND2_X1 U12910 ( .A1(n13399), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13412) );
  NAND2_X1 U12911 ( .A1(n13413), .A2(n13412), .ZN(n10333) );
  MUX2_X1 U12912 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11210), .S(n13410), .Z(
        n10332) );
  NAND2_X1 U12913 ( .A1(n10333), .A2(n10332), .ZN(n13427) );
  NAND2_X1 U12914 ( .A1(n13410), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13426) );
  NAND2_X1 U12915 ( .A1(n13427), .A2(n13426), .ZN(n10335) );
  MUX2_X1 U12916 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11097), .S(n13424), .Z(
        n10334) );
  NAND2_X1 U12917 ( .A1(n10335), .A2(n10334), .ZN(n13441) );
  NAND2_X1 U12918 ( .A1(n13424), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13440) );
  NAND2_X1 U12919 ( .A1(n13441), .A2(n13440), .ZN(n10337) );
  MUX2_X1 U12920 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11383), .S(n13438), .Z(
        n10336) );
  NAND2_X1 U12921 ( .A1(n10337), .A2(n10336), .ZN(n13443) );
  NAND2_X1 U12922 ( .A1(n13438), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10338) );
  NAND2_X1 U12923 ( .A1(n13443), .A2(n10338), .ZN(n15262) );
  OR2_X1 U12924 ( .A1(n15263), .A2(n15262), .ZN(n15260) );
  NAND2_X1 U12925 ( .A1(n10339), .A2(n11515), .ZN(n10340) );
  AND2_X1 U12926 ( .A1(n15260), .A2(n10340), .ZN(n10344) );
  MUX2_X1 U12927 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n11687), .S(n10564), .Z(
        n10343) );
  NAND2_X1 U12928 ( .A1(n10344), .A2(n10343), .ZN(n10557) );
  OAI211_X1 U12929 ( .C1(n10344), .C2(n10343), .A(n10557), .B(n15306), .ZN(
        n10347) );
  NAND2_X1 U12930 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11852)
         );
  INV_X1 U12931 ( .A(n11852), .ZN(n10345) );
  AOI21_X1 U12932 ( .B1(n15328), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10345), 
        .ZN(n10346) );
  OAI211_X1 U12933 ( .C1(n15325), .C2(n10348), .A(n10347), .B(n10346), .ZN(
        n10349) );
  OR2_X1 U12934 ( .A1(n10350), .A2(n10349), .ZN(P2_U3224) );
  INV_X1 U12935 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n10352) );
  INV_X1 U12936 ( .A(n13062), .ZN(n13094) );
  NAND2_X1 U12937 ( .A1(n13094), .A2(n11422), .ZN(n10351) );
  OAI21_X1 U12938 ( .B1(P3_U3897), .B2(n10352), .A(n10351), .ZN(P3_U3507) );
  INV_X1 U12939 ( .A(n11257), .ZN(n10941) );
  INV_X1 U12940 ( .A(n10353), .ZN(n10355) );
  OAI222_X1 U12941 ( .A1(P1_U3086), .A2(n10941), .B1(n14694), .B2(n10355), 
        .C1(n10354), .C2(n14691), .ZN(P1_U3343) );
  OAI222_X1 U12942 ( .A1(n13894), .A2(n10356), .B1(n13883), .B2(n10355), .C1(
        n11135), .C2(P2_U3088), .ZN(P2_U3315) );
  MUX2_X1 U12943 ( .A(n10359), .B(P1_REG1_REG_7__SCAN_IN), .S(n10414), .Z(
        n10360) );
  NOR2_X1 U12944 ( .A1(n10361), .A2(n10360), .ZN(n10413) );
  AOI211_X1 U12945 ( .C1(n10361), .C2(n10360), .A(n15036), .B(n10413), .ZN(
        n10374) );
  NOR2_X1 U12946 ( .A1(n10363), .A2(n10362), .ZN(n10366) );
  MUX2_X1 U12947 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10364), .S(n10414), .Z(
        n10365) );
  OAI21_X1 U12948 ( .B1(n10367), .B2(n10366), .A(n10365), .ZN(n10411) );
  INV_X1 U12949 ( .A(n10411), .ZN(n10369) );
  NOR3_X1 U12950 ( .A1(n10367), .A2(n10366), .A3(n10365), .ZN(n10368) );
  NOR3_X1 U12951 ( .A1(n15055), .A2(n10369), .A3(n10368), .ZN(n10373) );
  NAND2_X1 U12952 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11710) );
  NAND2_X1 U12953 ( .A1(n15027), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10370) );
  OAI211_X1 U12954 ( .C1(n15064), .C2(n10371), .A(n11710), .B(n10370), .ZN(
        n10372) );
  OR3_X1 U12955 ( .A1(n10374), .A2(n10373), .A3(n10372), .ZN(P1_U3250) );
  INV_X1 U12956 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n15832) );
  NAND2_X1 U12957 ( .A1(n11598), .A2(n11422), .ZN(n10375) );
  OAI21_X1 U12958 ( .B1(n11422), .B2(n15832), .A(n10375), .ZN(P3_U3495) );
  OAI21_X1 U12959 ( .B1(n10378), .B2(n10377), .A(n10376), .ZN(n10385) );
  INV_X1 U12960 ( .A(n10379), .ZN(n10383) );
  NOR3_X1 U12961 ( .A1(n15040), .A2(n10381), .A3(n10380), .ZN(n10382) );
  NOR3_X1 U12962 ( .A1(n15055), .A2(n10383), .A3(n10382), .ZN(n10384) );
  AOI21_X1 U12963 ( .B1(n15059), .B2(n10385), .A(n10384), .ZN(n10388) );
  NAND2_X1 U12964 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11362) );
  INV_X1 U12965 ( .A(n11362), .ZN(n10386) );
  AOI21_X1 U12966 ( .B1(n15027), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10386), .ZN(
        n10387) );
  OAI211_X1 U12967 ( .C1(n10389), .C2(n15064), .A(n10388), .B(n10387), .ZN(
        P1_U3248) );
  INV_X1 U12968 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U12969 ( .A1(n12110), .A2(n11422), .ZN(n10390) );
  OAI21_X1 U12970 ( .B1(P3_U3897), .B2(n10391), .A(n10390), .ZN(P3_U3499) );
  INV_X1 U12971 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n15583) );
  NAND2_X1 U12972 ( .A1(n14856), .A2(n11422), .ZN(n10392) );
  OAI21_X1 U12973 ( .B1(n11422), .B2(n15583), .A(n10392), .ZN(P3_U3504) );
  INV_X1 U12974 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n15833) );
  NAND2_X1 U12975 ( .A1(n12342), .A2(n11422), .ZN(n10393) );
  OAI21_X1 U12976 ( .B1(n11422), .B2(n15833), .A(n10393), .ZN(P3_U3501) );
  INV_X2 U12977 ( .A(n15389), .ZN(n15391) );
  NAND2_X1 U12978 ( .A1(n10394), .A2(n15391), .ZN(n10395) );
  OAI21_X1 U12979 ( .B1(n15391), .B2(n7893), .A(n10395), .ZN(P2_U3500) );
  INV_X1 U12980 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n15647) );
  NAND2_X1 U12981 ( .A1(n12104), .A2(n11422), .ZN(n10396) );
  OAI21_X1 U12982 ( .B1(n11422), .B2(n15647), .A(n10396), .ZN(P3_U3497) );
  OR2_X1 U12983 ( .A1(n13364), .A2(n8585), .ZN(n10397) );
  XNOR2_X1 U12984 ( .A(n10462), .B(n10467), .ZN(n11467) );
  INV_X1 U12985 ( .A(n15381), .ZN(n15373) );
  AOI211_X1 U12986 ( .C1(n10469), .C2(n10398), .A(n13720), .B(n10465), .ZN(
        n11470) );
  AOI21_X1 U12987 ( .B1(n15373), .B2(n10469), .A(n11470), .ZN(n10404) );
  NAND2_X1 U12988 ( .A1(n10400), .A2(n10399), .ZN(n10402) );
  OR2_X1 U12989 ( .A1(n13364), .A2(n10659), .ZN(n10401) );
  NAND2_X1 U12990 ( .A1(n10402), .A2(n10401), .ZN(n10468) );
  XNOR2_X1 U12991 ( .A(n10468), .B(n10467), .ZN(n10403) );
  INV_X1 U12992 ( .A(n8584), .ZN(n10689) );
  OAI22_X1 U12993 ( .A1(n10689), .A2(n13326), .B1(n7172), .B2(n13544), .ZN(
        n10738) );
  AOI21_X1 U12994 ( .B1(n10403), .B2(n14915), .A(n10738), .ZN(n11472) );
  OAI211_X1 U12995 ( .C1(n13842), .C2(n11467), .A(n10404), .B(n11472), .ZN(
        n10406) );
  NAND2_X1 U12996 ( .A1(n10406), .A2(n15387), .ZN(n10405) );
  OAI21_X1 U12997 ( .B1(n15387), .B2(n7928), .A(n10405), .ZN(P2_U3436) );
  NAND2_X1 U12998 ( .A1(n10406), .A2(n15391), .ZN(n10407) );
  OAI21_X1 U12999 ( .B1(n15391), .B2(n10305), .A(n10407), .ZN(P2_U3501) );
  INV_X1 U13000 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n15866) );
  NAND2_X1 U13001 ( .A1(n10999), .A2(n11422), .ZN(n10408) );
  OAI21_X1 U13002 ( .B1(P3_U3897), .B2(n15866), .A(n10408), .ZN(P3_U3492) );
  NAND2_X1 U13003 ( .A1(n10414), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10410) );
  INV_X1 U13004 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10440) );
  MUX2_X1 U13005 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10440), .S(n10441), .Z(
        n10409) );
  AOI21_X1 U13006 ( .B1(n10411), .B2(n10410), .A(n10409), .ZN(n10444) );
  NAND3_X1 U13007 ( .A1(n10411), .A2(n10410), .A3(n10409), .ZN(n10412) );
  NAND2_X1 U13008 ( .A1(n15046), .A2(n10412), .ZN(n10422) );
  MUX2_X1 U13009 ( .A(n10415), .B(P1_REG1_REG_8__SCAN_IN), .S(n10441), .Z(
        n10416) );
  OAI21_X1 U13010 ( .B1(n10417), .B2(n10416), .A(n10436), .ZN(n10418) );
  NAND2_X1 U13011 ( .A1(n10418), .A2(n15059), .ZN(n10421) );
  AND2_X1 U13012 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11890) );
  NOR2_X1 U13013 ( .A1(n15064), .A2(n10441), .ZN(n10419) );
  AOI211_X1 U13014 ( .C1(n15027), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11890), .B(
        n10419), .ZN(n10420) );
  OAI211_X1 U13015 ( .C1(n10444), .C2(n10422), .A(n10421), .B(n10420), .ZN(
        P1_U3251) );
  INV_X1 U13016 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n10425) );
  NAND2_X1 U13017 ( .A1(n10423), .A2(n11422), .ZN(n10424) );
  OAI21_X1 U13018 ( .B1(P3_U3897), .B2(n10425), .A(n10424), .ZN(P3_U3493) );
  INV_X1 U13019 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n15892) );
  INV_X1 U13020 ( .A(n13061), .ZN(n12880) );
  NAND2_X1 U13021 ( .A1(n12880), .A2(n11422), .ZN(n10426) );
  OAI21_X1 U13022 ( .B1(P3_U3897), .B2(n15892), .A(n10426), .ZN(P3_U3509) );
  OAI21_X1 U13023 ( .B1(n13342), .B2(n12389), .A(n13330), .ZN(n10429) );
  OR2_X1 U13024 ( .A1(n10427), .A2(P2_U3088), .ZN(n10747) );
  AOI22_X1 U13025 ( .A1(n10429), .A2(n10428), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n10747), .ZN(n10432) );
  NOR2_X1 U13026 ( .A1(n13342), .A2(n14928), .ZN(n13313) );
  NAND2_X1 U13027 ( .A1(n13313), .A2(n10430), .ZN(n10431) );
  OAI211_X1 U13028 ( .C1(n13339), .C2(n10433), .A(n10432), .B(n10431), .ZN(
        P2_U3204) );
  INV_X1 U13029 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n15636) );
  NAND2_X1 U13030 ( .A1(n14844), .A2(n11422), .ZN(n10434) );
  OAI21_X1 U13031 ( .B1(n11422), .B2(n15636), .A(n10434), .ZN(P3_U3503) );
  MUX2_X1 U13032 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10435), .S(n10484), .Z(
        n10439) );
  OAI21_X1 U13033 ( .B1(n10439), .B2(n10438), .A(n10481), .ZN(n10452) );
  NOR2_X1 U13034 ( .A1(n10441), .A2(n10440), .ZN(n10443) );
  MUX2_X1 U13035 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11826), .S(n10484), .Z(
        n10442) );
  OAI21_X1 U13036 ( .B1(n10444), .B2(n10443), .A(n10442), .ZN(n10487) );
  INV_X1 U13037 ( .A(n10487), .ZN(n10446) );
  NOR3_X1 U13038 ( .A1(n10444), .A2(n10443), .A3(n10442), .ZN(n10445) );
  NOR3_X1 U13039 ( .A1(n10446), .A2(n10445), .A3(n15055), .ZN(n10451) );
  NOR2_X1 U13040 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10447), .ZN(n11920) );
  AOI21_X1 U13041 ( .B1(n15027), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n11920), .ZN(
        n10448) );
  OAI21_X1 U13042 ( .B1(n15064), .B2(n10449), .A(n10448), .ZN(n10450) );
  AOI211_X1 U13043 ( .C1(n10452), .C2(n15059), .A(n10451), .B(n10450), .ZN(
        n10453) );
  INV_X1 U13044 ( .A(n10453), .ZN(P1_U3252) );
  INV_X1 U13045 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n15584) );
  INV_X1 U13046 ( .A(n13051), .ZN(n12883) );
  NAND2_X1 U13047 ( .A1(n12883), .A2(n11422), .ZN(n10454) );
  OAI21_X1 U13048 ( .B1(P3_U3897), .B2(n15584), .A(n10454), .ZN(P3_U3510) );
  INV_X1 U13049 ( .A(n10455), .ZN(n10458) );
  OAI222_X1 U13050 ( .A1(P2_U3088), .A2(n11148), .B1(n13883), .B2(n10458), 
        .C1(n10456), .C2(n13894), .ZN(P2_U3314) );
  INV_X1 U13051 ( .A(n11339), .ZN(n11261) );
  OAI222_X1 U13052 ( .A1(P1_U3086), .A2(n11261), .B1(n14694), .B2(n10458), 
        .C1(n10457), .C2(n14691), .ZN(P1_U3342) );
  OAI222_X1 U13053 ( .A1(n6670), .A2(n10460), .B1(n13251), .B2(n10459), .C1(
        n12824), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13054 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10476) );
  INV_X1 U13055 ( .A(n10467), .ZN(n10461) );
  OR2_X1 U13056 ( .A1(n13363), .A2(n10469), .ZN(n10463) );
  NAND2_X1 U13057 ( .A1(n10464), .A2(n10463), .ZN(n10573) );
  XNOR2_X1 U13058 ( .A(n10573), .B(n10578), .ZN(n11226) );
  INV_X1 U13059 ( .A(n10465), .ZN(n10466) );
  AND2_X1 U13060 ( .A1(n10465), .A2(n11221), .ZN(n10576) );
  AOI211_X1 U13061 ( .C1(n10580), .C2(n10466), .A(n13720), .B(n10576), .ZN(
        n11223) );
  AOI21_X1 U13062 ( .B1(n15373), .B2(n10580), .A(n11223), .ZN(n10474) );
  NAND2_X1 U13063 ( .A1(n10468), .A2(n10467), .ZN(n10471) );
  INV_X1 U13064 ( .A(n10469), .ZN(n11466) );
  OR2_X1 U13065 ( .A1(n13363), .A2(n11466), .ZN(n10470) );
  NAND2_X1 U13066 ( .A1(n10471), .A2(n10470), .ZN(n10579) );
  XNOR2_X1 U13067 ( .A(n10579), .B(n10578), .ZN(n10473) );
  AOI21_X1 U13068 ( .B1(n10473), .B2(n14915), .A(n10472), .ZN(n11219) );
  OAI211_X1 U13069 ( .C1(n13842), .C2(n11226), .A(n10474), .B(n11219), .ZN(
        n10477) );
  NAND2_X1 U13070 ( .A1(n10477), .A2(n15387), .ZN(n10475) );
  OAI21_X1 U13071 ( .B1(n15387), .B2(n10476), .A(n10475), .ZN(P2_U3439) );
  NAND2_X1 U13072 ( .A1(n10477), .A2(n15391), .ZN(n10478) );
  OAI21_X1 U13073 ( .B1(n15391), .B2(n7961), .A(n10478), .ZN(P2_U3502) );
  INV_X1 U13074 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n15664) );
  INV_X1 U13075 ( .A(n13031), .ZN(n12885) );
  NAND2_X1 U13076 ( .A1(n12885), .A2(n11422), .ZN(n10479) );
  OAI21_X1 U13077 ( .B1(P3_U3897), .B2(n15664), .A(n10479), .ZN(P3_U3511) );
  MUX2_X1 U13078 ( .A(n10480), .B(P1_REG1_REG_10__SCAN_IN), .S(n10593), .Z(
        n10483) );
  OAI21_X1 U13079 ( .B1(n10484), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10481), .ZN(
        n10482) );
  NOR2_X1 U13080 ( .A1(n10482), .A2(n10483), .ZN(n10592) );
  AOI211_X1 U13081 ( .C1(n10483), .C2(n10482), .A(n15036), .B(n10592), .ZN(
        n10493) );
  NAND2_X1 U13082 ( .A1(n10484), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10486) );
  MUX2_X1 U13083 ( .A(n9715), .B(P1_REG2_REG_10__SCAN_IN), .S(n10593), .Z(
        n10485) );
  AOI21_X1 U13084 ( .B1(n10487), .B2(n10486), .A(n10485), .ZN(n10591) );
  AND3_X1 U13085 ( .A1(n10487), .A2(n10486), .A3(n10485), .ZN(n10488) );
  NOR3_X1 U13086 ( .A1(n10591), .A2(n10488), .A3(n15055), .ZN(n10492) );
  AND2_X1 U13087 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11979) );
  AOI21_X1 U13088 ( .B1(n15027), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11979), 
        .ZN(n10489) );
  OAI21_X1 U13089 ( .B1(n15064), .B2(n10490), .A(n10489), .ZN(n10491) );
  OR3_X1 U13090 ( .A1(n10493), .A2(n10492), .A3(n10491), .ZN(P1_U3253) );
  INV_X1 U13091 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n15796) );
  NAND2_X1 U13092 ( .A1(n12648), .A2(n11422), .ZN(n10494) );
  OAI21_X1 U13093 ( .B1(n11422), .B2(n15796), .A(n10494), .ZN(P3_U3512) );
  INV_X1 U13094 ( .A(n12838), .ZN(n12826) );
  OAI222_X1 U13095 ( .A1(n6670), .A2(n10496), .B1(n13251), .B2(n10495), .C1(
        n12826), .C2(P3_U3151), .ZN(P3_U3277) );
  NAND2_X1 U13096 ( .A1(n11580), .A2(n10497), .ZN(n10498) );
  NAND2_X1 U13097 ( .A1(n10639), .A2(n10498), .ZN(n10506) );
  NAND2_X1 U13098 ( .A1(n10920), .A2(n11563), .ZN(n10505) );
  INV_X1 U13099 ( .A(n10505), .ZN(n10499) );
  NOR2_X1 U13100 ( .A1(n10506), .A2(n10499), .ZN(n10513) );
  INV_X1 U13101 ( .A(n10513), .ZN(n10500) );
  INV_X1 U13102 ( .A(n12857), .ZN(n10511) );
  MUX2_X1 U13103 ( .A(n10500), .B(n11368), .S(n10511), .Z(n12851) );
  NAND2_X1 U13104 ( .A1(n10513), .A2(n12814), .ZN(n12855) );
  INV_X1 U13105 ( .A(n12855), .ZN(n11030) );
  NAND2_X1 U13106 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10507), .ZN(n11050) );
  INV_X1 U13107 ( .A(n11050), .ZN(n10503) );
  NAND2_X1 U13108 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10503), .ZN(n10502) );
  OAI21_X1 U13109 ( .B1(n10508), .B2(n10503), .A(n10502), .ZN(n10504) );
  NAND2_X1 U13110 ( .A1(n10504), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10676) );
  OAI21_X1 U13111 ( .B1(n10504), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10676), .ZN(
        n10517) );
  OAI22_X1 U13112 ( .A1(n12813), .A2(n15864), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15459), .ZN(n10516) );
  NAND2_X1 U13113 ( .A1(n10507), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11045) );
  NAND2_X1 U13114 ( .A1(n10508), .A2(n11045), .ZN(n10509) );
  NAND2_X1 U13115 ( .A1(n8678), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10679) );
  NAND2_X1 U13116 ( .A1(n10509), .A2(n10679), .ZN(n10510) );
  OR2_X1 U13117 ( .A1(n10510), .A2(n8662), .ZN(n10680) );
  NAND2_X1 U13118 ( .A1(n10510), .A2(n8662), .ZN(n10514) );
  NAND2_X1 U13119 ( .A1(n10511), .A2(n12840), .ZN(n10640) );
  INV_X1 U13120 ( .A(n10640), .ZN(n10512) );
  NAND2_X1 U13121 ( .A1(n10513), .A2(n10512), .ZN(n12847) );
  AOI21_X1 U13122 ( .B1(n10680), .B2(n10514), .A(n12847), .ZN(n10515) );
  AOI211_X1 U13123 ( .C1(n11030), .C2(n10517), .A(n10516), .B(n10515), .ZN(
        n10523) );
  INV_X1 U13124 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10985) );
  MUX2_X1 U13125 ( .A(n10985), .B(n10519), .S(n12814), .Z(n11051) );
  AND2_X1 U13126 ( .A1(n11051), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11056) );
  OAI21_X1 U13127 ( .B1(n10520), .B2(n11056), .A(n10673), .ZN(n10521) );
  AND2_X1 U13128 ( .A1(P3_U3897), .A2(n12857), .ZN(n12853) );
  NAND2_X1 U13129 ( .A1(n10521), .A2(n12853), .ZN(n10522) );
  OAI211_X1 U13130 ( .C1(n12851), .C2(n10524), .A(n10523), .B(n10522), .ZN(
        P3_U3183) );
  OR2_X1 U13131 ( .A1(n10539), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10526) );
  AND2_X1 U13132 ( .A1(n10526), .A2(n10525), .ZN(n11452) );
  OR2_X1 U13133 ( .A1(n10539), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10528) );
  AND2_X1 U13134 ( .A1(n10528), .A2(n10527), .ZN(n11449) );
  NOR4_X1 U13135 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10537) );
  NOR4_X1 U13136 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n10536) );
  INV_X1 U13137 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15138) );
  INV_X1 U13138 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15137) );
  INV_X1 U13139 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15136) );
  INV_X1 U13140 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15135) );
  NAND4_X1 U13141 ( .A1(n15138), .A2(n15137), .A3(n15136), .A4(n15135), .ZN(
        n10534) );
  NOR4_X1 U13142 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10532) );
  NOR4_X1 U13143 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n10531) );
  NOR4_X1 U13144 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10530) );
  NOR4_X1 U13145 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10529) );
  NAND4_X1 U13146 ( .A1(n10532), .A2(n10531), .A3(n10530), .A4(n10529), .ZN(
        n10533) );
  NOR4_X1 U13147 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n10534), .A4(n10533), .ZN(n10535) );
  AND3_X1 U13148 ( .A1(n10537), .A2(n10536), .A3(n10535), .ZN(n10538) );
  OR2_X1 U13149 ( .A1(n10539), .A2(n10538), .ZN(n10734) );
  NAND3_X1 U13150 ( .A1(n11452), .A2(n11449), .A3(n10734), .ZN(n10541) );
  NAND2_X2 U13151 ( .A1(n10732), .A2(n11674), .ZN(n15205) );
  NAND2_X1 U13152 ( .A1(n10541), .A2(n10733), .ZN(n11268) );
  AND2_X1 U13153 ( .A1(n11268), .A2(n11453), .ZN(n14062) );
  NAND2_X1 U13154 ( .A1(n10732), .A2(n10728), .ZN(n11459) );
  INV_X1 U13155 ( .A(n14163), .ZN(n14150) );
  INV_X1 U13156 ( .A(n10541), .ZN(n10551) );
  NAND2_X1 U13157 ( .A1(n11453), .A2(n10552), .ZN(n10542) );
  NOR2_X1 U13158 ( .A1(n15192), .A2(n10542), .ZN(n10543) );
  NAND2_X2 U13159 ( .A1(n10546), .A2(n10544), .ZN(n13941) );
  OAI22_X1 U13160 ( .A1(n11480), .A2(n13941), .B1(n10546), .B2(n14198), .ZN(
        n10545) );
  NAND2_X1 U13161 ( .A1(n14182), .A2(n6666), .ZN(n10549) );
  OAI22_X1 U13162 ( .A1(n11480), .A2(n13942), .B1(n10546), .B2(n15019), .ZN(
        n10547) );
  INV_X1 U13163 ( .A(n10547), .ZN(n10548) );
  NAND2_X1 U13164 ( .A1(n10549), .A2(n10548), .ZN(n10703) );
  OAI21_X1 U13165 ( .B1(n10550), .B2(n10703), .A(n10705), .ZN(n14193) );
  NAND2_X1 U13166 ( .A1(n10551), .A2(n10735), .ZN(n14133) );
  OR2_X1 U13167 ( .A1(n10552), .A2(n14197), .ZN(n14156) );
  OR2_X1 U13168 ( .A1(n11488), .A2(n14156), .ZN(n11457) );
  INV_X1 U13169 ( .A(n11457), .ZN(n10731) );
  AOI22_X1 U13170 ( .A1(n14142), .A2(n14193), .B1(n14159), .B2(n10731), .ZN(
        n10555) );
  NAND2_X1 U13171 ( .A1(n14062), .A2(n10553), .ZN(n10804) );
  NAND2_X1 U13172 ( .A1(n10804), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10554) );
  OAI211_X1 U13173 ( .C1(n14150), .C2(n11480), .A(n10555), .B(n10554), .ZN(
        P1_U3232) );
  NAND2_X1 U13174 ( .A1(n10564), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10556) );
  AND2_X1 U13175 ( .A1(n10557), .A2(n10556), .ZN(n10559) );
  MUX2_X1 U13176 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11767), .S(n10831), .Z(
        n10558) );
  NAND2_X1 U13177 ( .A1(n10559), .A2(n10558), .ZN(n10836) );
  OAI21_X1 U13178 ( .B1(n10559), .B2(n10558), .A(n10836), .ZN(n10570) );
  NAND2_X1 U13179 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11806)
         );
  INV_X1 U13180 ( .A(n11806), .ZN(n10560) );
  AOI21_X1 U13181 ( .B1(n15328), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10560), 
        .ZN(n10561) );
  OAI21_X1 U13182 ( .B1(n15325), .B2(n10562), .A(n10561), .ZN(n10569) );
  INV_X1 U13183 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10565) );
  MUX2_X1 U13184 ( .A(n10565), .B(P2_REG1_REG_11__SCAN_IN), .S(n10831), .Z(
        n10566) );
  NOR2_X1 U13185 ( .A1(n10567), .A2(n10566), .ZN(n10827) );
  AOI211_X1 U13186 ( .C1(n10567), .C2(n10566), .A(n15319), .B(n10827), .ZN(
        n10568) );
  AOI211_X1 U13187 ( .C1(n15306), .C2(n10570), .A(n10569), .B(n10568), .ZN(
        n10571) );
  INV_X1 U13188 ( .A(n10571), .ZN(P2_U3225) );
  INV_X1 U13189 ( .A(n10578), .ZN(n10572) );
  NAND2_X1 U13190 ( .A1(n10573), .A2(n10572), .ZN(n10575) );
  OR2_X1 U13191 ( .A1(n10580), .A2(n8584), .ZN(n10574) );
  NAND2_X1 U13192 ( .A1(n10575), .A2(n10574), .ZN(n10898) );
  XNOR2_X1 U13193 ( .A(n10898), .B(n10901), .ZN(n11206) );
  INV_X1 U13194 ( .A(n10576), .ZN(n10577) );
  INV_X1 U13195 ( .A(n10899), .ZN(n11201) );
  AOI211_X1 U13196 ( .C1(n10899), .C2(n10577), .A(n13720), .B(n10905), .ZN(
        n11203) );
  AOI21_X1 U13197 ( .B1(n15373), .B2(n10899), .A(n11203), .ZN(n10586) );
  NAND2_X1 U13198 ( .A1(n10579), .A2(n10578), .ZN(n10582) );
  NAND2_X1 U13199 ( .A1(n10689), .A2(n10580), .ZN(n10581) );
  NAND2_X1 U13200 ( .A1(n10582), .A2(n10581), .ZN(n10902) );
  XNOR2_X1 U13201 ( .A(n10902), .B(n10901), .ZN(n10585) );
  NAND2_X1 U13202 ( .A1(n8584), .A2(n13307), .ZN(n10584) );
  NAND2_X1 U13203 ( .A1(n13361), .A2(n13336), .ZN(n10583) );
  NAND2_X1 U13204 ( .A1(n10584), .A2(n10583), .ZN(n10694) );
  AOI21_X1 U13205 ( .B1(n10585), .B2(n14915), .A(n10694), .ZN(n11198) );
  OAI211_X1 U13206 ( .C1(n13842), .C2(n11206), .A(n10586), .B(n11198), .ZN(
        n10588) );
  NAND2_X1 U13207 ( .A1(n10588), .A2(n15387), .ZN(n10587) );
  OAI21_X1 U13208 ( .B1(n15387), .B2(n7978), .A(n10587), .ZN(P2_U3442) );
  NAND2_X1 U13209 ( .A1(n10588), .A2(n15391), .ZN(n10589) );
  OAI21_X1 U13210 ( .B1(n15391), .B2(n10590), .A(n10589), .ZN(P2_U3503) );
  AOI21_X1 U13211 ( .B1(n10593), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10591), 
        .ZN(n10931) );
  MUX2_X1 U13212 ( .A(n11846), .B(P1_REG2_REG_11__SCAN_IN), .S(n10937), .Z(
        n10930) );
  XNOR2_X1 U13213 ( .A(n10931), .B(n10930), .ZN(n10602) );
  MUX2_X1 U13214 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10594), .S(n10937), .Z(
        n10595) );
  OAI21_X1 U13215 ( .B1(n10596), .B2(n10595), .A(n10936), .ZN(n10597) );
  NAND2_X1 U13216 ( .A1(n10597), .A2(n15059), .ZN(n10601) );
  NAND2_X1 U13217 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12227)
         );
  INV_X1 U13218 ( .A(n12227), .ZN(n10599) );
  NOR2_X1 U13219 ( .A1(n15064), .A2(n10933), .ZN(n10598) );
  AOI211_X1 U13220 ( .C1(n15027), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10599), 
        .B(n10598), .ZN(n10600) );
  OAI211_X1 U13221 ( .C1(n15055), .C2(n10602), .A(n10601), .B(n10600), .ZN(
        P1_U3254) );
  INV_X1 U13222 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10603) );
  NAND2_X1 U13223 ( .A1(n10618), .A2(n10603), .ZN(n10606) );
  INV_X1 U13224 ( .A(n10604), .ZN(n12167) );
  NAND2_X1 U13225 ( .A1(n12167), .A2(n12014), .ZN(n10605) );
  INV_X1 U13226 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U13227 ( .A1(n10618), .A2(n10607), .ZN(n10609) );
  NAND2_X1 U13228 ( .A1(n12167), .A2(n11899), .ZN(n10608) );
  NOR2_X1 U13229 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n10613) );
  NOR4_X1 U13230 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n10612) );
  NOR4_X1 U13231 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n10611) );
  NOR4_X1 U13232 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n10610) );
  NAND4_X1 U13233 ( .A1(n10613), .A2(n10612), .A3(n10611), .A4(n10610), .ZN(
        n10620) );
  NOR4_X1 U13234 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n10617) );
  NOR4_X1 U13235 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n10616) );
  NOR4_X1 U13236 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n10615) );
  NOR4_X1 U13237 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n10614) );
  NAND4_X1 U13238 ( .A1(n10617), .A2(n10616), .A3(n10615), .A4(n10614), .ZN(
        n10619) );
  OAI21_X1 U13239 ( .B1(n10620), .B2(n10619), .A(n10618), .ZN(n10811) );
  AND3_X1 U13240 ( .A1(n13234), .A2(n13236), .A3(n10811), .ZN(n10921) );
  NAND2_X1 U13241 ( .A1(n12850), .A2(n11565), .ZN(n10623) );
  NAND2_X1 U13242 ( .A1(n11565), .A2(n11107), .ZN(n10621) );
  XNOR2_X1 U13243 ( .A(n13115), .B(n10621), .ZN(n10622) );
  NAND2_X1 U13244 ( .A1(n10623), .A2(n10622), .ZN(n11585) );
  INV_X1 U13245 ( .A(n11585), .ZN(n10624) );
  NOR2_X1 U13246 ( .A1(n10921), .A2(n10624), .ZN(n10630) );
  INV_X1 U13247 ( .A(n13236), .ZN(n10625) );
  INV_X1 U13248 ( .A(n13234), .ZN(n10976) );
  AND3_X1 U13249 ( .A1(n10625), .A2(n10976), .A3(n10811), .ZN(n10924) );
  NOR2_X1 U13250 ( .A1(n10862), .A2(n10819), .ZN(n10626) );
  NAND2_X1 U13251 ( .A1(n11577), .A2(n10626), .ZN(n10919) );
  INV_X1 U13252 ( .A(n10627), .ZN(n10628) );
  NAND2_X1 U13253 ( .A1(n11583), .A2(n11580), .ZN(n10975) );
  OAI211_X1 U13254 ( .C1(n10924), .C2(n10919), .A(n10628), .B(n10975), .ZN(
        n10629) );
  OAI21_X1 U13255 ( .B1(n10630), .B2(n10629), .A(P3_STATE_REG_SCAN_IN), .ZN(
        n10633) );
  INV_X1 U13256 ( .A(n10918), .ZN(n10631) );
  INV_X1 U13257 ( .A(n10924), .ZN(n10638) );
  NAND2_X1 U13258 ( .A1(n10631), .A2(n10638), .ZN(n10632) );
  NAND2_X1 U13259 ( .A1(n10633), .A2(n10632), .ZN(n11058) );
  NOR2_X1 U13260 ( .A1(n11058), .A2(n13235), .ZN(n11002) );
  INV_X1 U13261 ( .A(n10809), .ZN(n10644) );
  NAND3_X1 U13262 ( .A1(n10921), .A2(n15512), .A3(n11585), .ZN(n10636) );
  INV_X1 U13263 ( .A(n10919), .ZN(n10634) );
  NAND2_X1 U13264 ( .A1(n10924), .A2(n10634), .ZN(n10635) );
  NAND2_X1 U13265 ( .A1(n10636), .A2(n10635), .ZN(n10637) );
  INV_X1 U13266 ( .A(n10920), .ZN(n10923) );
  NAND2_X1 U13267 ( .A1(n10637), .A2(n10923), .ZN(n12672) );
  NOR2_X1 U13268 ( .A1(n10638), .A2(n10918), .ZN(n10875) );
  NAND2_X1 U13269 ( .A1(n10640), .A2(n10639), .ZN(n10874) );
  NAND2_X1 U13270 ( .A1(n10875), .A2(n10874), .ZN(n12668) );
  INV_X1 U13271 ( .A(n10921), .ZN(n10641) );
  NAND2_X1 U13272 ( .A1(n10641), .A2(n15438), .ZN(n10642) );
  NOR2_X1 U13273 ( .A1(n10920), .A2(n15512), .ZN(n10983) );
  INV_X1 U13274 ( .A(n12670), .ZN(n12684) );
  OAI22_X1 U13275 ( .A1(n15426), .A2(n12668), .B1(n12684), .B2(n10927), .ZN(
        n10643) );
  AOI21_X1 U13276 ( .B1(n10644), .B2(n7432), .A(n10643), .ZN(n10645) );
  OAI21_X1 U13277 ( .B1(n11002), .B2(n11046), .A(n10645), .ZN(P3_U3172) );
  NAND2_X1 U13278 ( .A1(n13362), .A2(n13307), .ZN(n10647) );
  NAND2_X1 U13279 ( .A1(n13360), .A2(n13336), .ZN(n10646) );
  AND2_X1 U13280 ( .A1(n10647), .A2(n10646), .ZN(n11237) );
  NAND2_X1 U13281 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13394) );
  OAI21_X1 U13282 ( .B1(n13339), .B2(n11237), .A(n13394), .ZN(n10649) );
  NOR2_X1 U13283 ( .A1(n14911), .A2(n11239), .ZN(n10648) );
  AOI211_X1 U13284 ( .C1(n11084), .C2(n14908), .A(n10649), .B(n10648), .ZN(
        n10656) );
  INV_X1 U13285 ( .A(n13313), .ZN(n11810) );
  OAI22_X1 U13286 ( .A1(n11810), .A2(n10651), .B1(n10650), .B2(n13342), .ZN(
        n10654) );
  INV_X1 U13287 ( .A(n10652), .ZN(n10653) );
  NAND3_X1 U13288 ( .A1(n10654), .A2(n10693), .A3(n10653), .ZN(n10655) );
  OAI211_X1 U13289 ( .C1(n10657), .C2(n13342), .A(n10656), .B(n10655), .ZN(
        P2_U3199) );
  INV_X1 U13290 ( .A(n10658), .ZN(n11177) );
  OAI22_X1 U13291 ( .A1(n13330), .A2(n10659), .B1(n11177), .B2(n13339), .ZN(
        n10664) );
  AOI22_X1 U13292 ( .A1(n13313), .A2(n6697), .B1(n10660), .B2(n14903), .ZN(
        n10662) );
  NOR2_X1 U13293 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  AOI211_X1 U13294 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(n10747), .A(n10664), .B(
        n10663), .ZN(n10665) );
  OAI21_X1 U13295 ( .B1(n10741), .B2(n13342), .A(n10665), .ZN(P2_U3194) );
  MUX2_X1 U13296 ( .A(n10667), .B(n10666), .S(n12814), .Z(n10669) );
  INV_X1 U13297 ( .A(n10780), .ZN(n10668) );
  NAND2_X1 U13298 ( .A1(n10669), .A2(n10668), .ZN(n10758) );
  INV_X1 U13299 ( .A(n10669), .ZN(n10670) );
  NAND2_X1 U13300 ( .A1(n10670), .A2(n10780), .ZN(n10671) );
  NAND2_X1 U13301 ( .A1(n10758), .A2(n10671), .ZN(n10672) );
  AND3_X1 U13302 ( .A1(n10673), .A2(n7040), .A3(n10672), .ZN(n10674) );
  OAI21_X1 U13303 ( .B1(n10854), .B2(n10674), .A(n12853), .ZN(n10688) );
  MUX2_X1 U13304 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10666), .S(n10780), .Z(
        n10678) );
  OR2_X1 U13305 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11050), .ZN(n10675) );
  NAND2_X1 U13306 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  NAND2_X1 U13307 ( .A1(n10678), .A2(n10677), .ZN(n10782) );
  OAI21_X1 U13308 ( .B1(n10678), .B2(n10677), .A(n10782), .ZN(n10686) );
  OAI22_X1 U13309 ( .A1(n12813), .A2(n15894), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8670), .ZN(n10685) );
  INV_X1 U13310 ( .A(n12847), .ZN(n12702) );
  NAND2_X1 U13311 ( .A1(n10680), .A2(n10679), .ZN(n10681) );
  OAI21_X1 U13312 ( .B1(n10682), .B2(n10681), .A(n10751), .ZN(n10683) );
  AND2_X1 U13313 ( .A1(n12702), .A2(n10683), .ZN(n10684) );
  AOI211_X1 U13314 ( .C1(n11030), .C2(n10686), .A(n10685), .B(n10684), .ZN(
        n10687) );
  OAI211_X1 U13315 ( .C1(n12851), .C2(n10780), .A(n10688), .B(n10687), .ZN(
        P3_U3184) );
  NOR3_X1 U13316 ( .A1(n11810), .A2(n10690), .A3(n10689), .ZN(n10691) );
  AOI21_X1 U13317 ( .B1(n14903), .B2(n10692), .A(n10691), .ZN(n10701) );
  INV_X1 U13318 ( .A(n10693), .ZN(n10698) );
  AOI22_X1 U13319 ( .A1(n14905), .A2(n10694), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10696) );
  NAND2_X1 U13320 ( .A1(n14908), .A2(n10899), .ZN(n10695) );
  OAI211_X1 U13321 ( .C1(n14911), .C2(n11200), .A(n10696), .B(n10695), .ZN(
        n10697) );
  AOI21_X1 U13322 ( .B1(n10698), .B2(n14903), .A(n10697), .ZN(n10699) );
  OAI21_X1 U13323 ( .B1(n10701), .B2(n10700), .A(n10699), .ZN(P2_U3202) );
  OAI222_X1 U13324 ( .A1(n6670), .A2(n10702), .B1(n12850), .B2(P3_U3151), .C1(
        n15895), .C2(n13251), .ZN(P3_U3276) );
  OR2_X1 U13325 ( .A1(n10703), .A2(n13985), .ZN(n10704) );
  NAND2_X1 U13326 ( .A1(n10705), .A2(n10704), .ZN(n10800) );
  XNOR2_X1 U13327 ( .A(n10706), .B(n13985), .ZN(n10710) );
  NAND2_X1 U13328 ( .A1(n15142), .A2(n6666), .ZN(n10707) );
  XNOR2_X1 U13329 ( .A(n10710), .B(n10708), .ZN(n10799) );
  NAND2_X1 U13330 ( .A1(n10800), .A2(n10799), .ZN(n10712) );
  INV_X1 U13331 ( .A(n10708), .ZN(n10709) );
  NAND2_X1 U13332 ( .A1(n10710), .A2(n10709), .ZN(n10711) );
  NAND2_X1 U13333 ( .A1(n14181), .A2(n6666), .ZN(n10714) );
  NAND2_X1 U13334 ( .A1(n7010), .A2(n14042), .ZN(n10713) );
  NAND2_X1 U13335 ( .A1(n10714), .A2(n10713), .ZN(n10715) );
  XNOR2_X1 U13336 ( .A(n10715), .B(n13985), .ZN(n11275) );
  NAND2_X1 U13337 ( .A1(n14181), .A2(n14045), .ZN(n10717) );
  NAND2_X1 U13338 ( .A1(n7010), .A2(n6666), .ZN(n10716) );
  NAND2_X1 U13339 ( .A1(n10717), .A2(n10716), .ZN(n11273) );
  XNOR2_X1 U13340 ( .A(n11273), .B(n11275), .ZN(n11271) );
  XNOR2_X1 U13341 ( .A(n11272), .B(n11271), .ZN(n10718) );
  NAND2_X1 U13342 ( .A1(n10718), .A2(n14142), .ZN(n10722) );
  OR2_X1 U13343 ( .A1(n11488), .A2(n14357), .ZN(n10720) );
  NAND2_X1 U13344 ( .A1(n14179), .A2(n14281), .ZN(n10719) );
  NAND2_X1 U13345 ( .A1(n10720), .A2(n10719), .ZN(n15150) );
  AOI22_X1 U13346 ( .A1(n10804), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14159), 
        .B2(n15150), .ZN(n10721) );
  OAI211_X1 U13347 ( .C1(n11524), .C2(n14150), .A(n10722), .B(n10721), .ZN(
        P1_U3237) );
  INV_X1 U13348 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n15890) );
  NAND2_X1 U13349 ( .A1(n12985), .A2(n11422), .ZN(n10723) );
  OAI21_X1 U13350 ( .B1(n11422), .B2(n15890), .A(n10723), .ZN(P3_U3513) );
  INV_X1 U13351 ( .A(n11480), .ZN(n11486) );
  INV_X1 U13352 ( .A(n15189), .ZN(n15089) );
  NOR2_X1 U13353 ( .A1(n10725), .A2(n10724), .ZN(n10726) );
  OR2_X1 U13354 ( .A1(n13985), .A2(n10726), .ZN(n11455) );
  INV_X1 U13355 ( .A(n11455), .ZN(n10727) );
  NAND2_X1 U13356 ( .A1(n10727), .A2(n14511), .ZN(n15187) );
  OR2_X1 U13357 ( .A1(n10728), .A2(n14511), .ZN(n10729) );
  OR2_X1 U13358 ( .A1(n14696), .A2(n10729), .ZN(n15197) );
  AOI21_X1 U13359 ( .B1(n15089), .B2(n15176), .A(n11464), .ZN(n10730) );
  AOI211_X1 U13360 ( .C1(n10732), .C2(n11486), .A(n10731), .B(n10730), .ZN(
        n15141) );
  INV_X1 U13361 ( .A(n10733), .ZN(n11454) );
  AND2_X1 U13362 ( .A1(n10735), .A2(n10734), .ZN(n11450) );
  AND2_X1 U13363 ( .A1(n11450), .A2(n11449), .ZN(n10736) );
  AND2_X2 U13364 ( .A1(n12303), .A2(n10736), .ZN(n15233) );
  NAND2_X1 U13365 ( .A1(n15231), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10737) );
  OAI21_X1 U13366 ( .B1(n15141), .B2(n15231), .A(n10737), .ZN(P1_U3528) );
  INV_X1 U13367 ( .A(n10738), .ZN(n10739) );
  OAI22_X1 U13368 ( .A1(n11466), .A2(n13330), .B1(n10739), .B2(n13339), .ZN(
        n10746) );
  AOI22_X1 U13369 ( .A1(n13313), .A2(n13364), .B1(n14903), .B2(n10740), .ZN(
        n10744) );
  INV_X1 U13370 ( .A(n10741), .ZN(n10743) );
  NOR3_X1 U13371 ( .A1(n10744), .A2(n10743), .A3(n10742), .ZN(n10745) );
  AOI211_X1 U13372 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n10747), .A(n10746), .B(
        n10745), .ZN(n10748) );
  OAI21_X1 U13373 ( .B1(n10749), .B2(n13342), .A(n10748), .ZN(P2_U3209) );
  NAND2_X1 U13374 ( .A1(n10780), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U13375 ( .A1(n10752), .A2(n10783), .ZN(n12699) );
  MUX2_X1 U13376 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10765), .S(n10787), .Z(
        n12701) );
  INV_X1 U13377 ( .A(n12701), .ZN(n10753) );
  AOI21_X1 U13378 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10787), .A(n12704), .ZN(
        n10754) );
  MUX2_X1 U13379 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n10963), .S(n10964), .Z(
        n10756) );
  INV_X1 U13380 ( .A(n10966), .ZN(n10755) );
  AOI21_X1 U13381 ( .B1(n10757), .B2(n10756), .A(n10755), .ZN(n10798) );
  INV_X1 U13382 ( .A(n10758), .ZN(n10853) );
  MUX2_X1 U13383 ( .A(n10760), .B(n10759), .S(n12814), .Z(n10761) );
  INV_X1 U13384 ( .A(n10783), .ZN(n10851) );
  NAND2_X1 U13385 ( .A1(n10761), .A2(n10851), .ZN(n12686) );
  INV_X1 U13386 ( .A(n10761), .ZN(n10762) );
  NAND2_X1 U13387 ( .A1(n10762), .A2(n10783), .ZN(n10763) );
  AND2_X1 U13388 ( .A1(n12686), .A2(n10763), .ZN(n10852) );
  MUX2_X1 U13389 ( .A(n10765), .B(n10764), .S(n12814), .Z(n10766) );
  INV_X1 U13390 ( .A(n10787), .ZN(n12698) );
  NAND2_X1 U13391 ( .A1(n10766), .A2(n12698), .ZN(n10769) );
  INV_X1 U13392 ( .A(n10766), .ZN(n10767) );
  NAND2_X1 U13393 ( .A1(n10767), .A2(n10787), .ZN(n10768) );
  NAND2_X1 U13394 ( .A1(n10769), .A2(n10768), .ZN(n12685) );
  INV_X1 U13395 ( .A(n10769), .ZN(n10882) );
  MUX2_X1 U13396 ( .A(n11607), .B(n10770), .S(n12814), .Z(n10771) );
  NAND2_X1 U13397 ( .A1(n10771), .A2(n10894), .ZN(n10778) );
  INV_X1 U13398 ( .A(n10771), .ZN(n10772) );
  NAND2_X1 U13399 ( .A1(n10772), .A2(n7463), .ZN(n10773) );
  AND2_X1 U13400 ( .A1(n10778), .A2(n10773), .ZN(n10881) );
  MUX2_X1 U13401 ( .A(n10963), .B(n10946), .S(n12814), .Z(n10774) );
  NAND2_X1 U13402 ( .A1(n10774), .A2(n10964), .ZN(n10950) );
  INV_X1 U13403 ( .A(n10774), .ZN(n10775) );
  NAND2_X1 U13404 ( .A1(n10775), .A2(n10793), .ZN(n10776) );
  NAND2_X1 U13405 ( .A1(n10950), .A2(n10776), .ZN(n10777) );
  AND3_X1 U13406 ( .A1(n10880), .A2(n10778), .A3(n10777), .ZN(n10779) );
  OAI21_X1 U13407 ( .B1(n10958), .B2(n10779), .A(n12853), .ZN(n10797) );
  MUX2_X1 U13408 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10946), .S(n10964), .Z(
        n10790) );
  NAND2_X1 U13409 ( .A1(n10780), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U13410 ( .A1(n10784), .A2(n10783), .ZN(n12691) );
  NAND2_X1 U13411 ( .A1(n10785), .A2(n12691), .ZN(n10845) );
  NOR2_X1 U13412 ( .A1(n10845), .A2(n10759), .ZN(n10844) );
  INV_X1 U13413 ( .A(n12691), .ZN(n10786) );
  MUX2_X1 U13414 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10764), .S(n10787), .Z(
        n12690) );
  OAI21_X1 U13415 ( .B1(n10844), .B2(n10786), .A(n12690), .ZN(n12695) );
  NOR2_X1 U13416 ( .A1(n10894), .A2(n10788), .ZN(n10789) );
  OAI21_X1 U13417 ( .B1(n7282), .B2(n7283), .A(n10948), .ZN(n10795) );
  INV_X1 U13418 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10791) );
  NOR2_X1 U13419 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10791), .ZN(n11788) );
  AOI21_X1 U13420 ( .B1(n15392), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11788), .ZN(
        n10792) );
  OAI21_X1 U13421 ( .B1(n12851), .B2(n10793), .A(n10792), .ZN(n10794) );
  AOI21_X1 U13422 ( .B1(n10795), .B2(n11030), .A(n10794), .ZN(n10796) );
  OAI211_X1 U13423 ( .C1(n10798), .C2(n12847), .A(n10797), .B(n10796), .ZN(
        P3_U3188) );
  XOR2_X1 U13424 ( .A(n10799), .B(n10800), .Z(n10806) );
  NOR2_X1 U13425 ( .A1(n14133), .A2(n14357), .ZN(n14136) );
  INV_X1 U13426 ( .A(n14136), .ZN(n10801) );
  INV_X1 U13427 ( .A(n14182), .ZN(n11662) );
  NAND2_X1 U13428 ( .A1(n14159), .A2(n14281), .ZN(n11982) );
  OAI22_X1 U13429 ( .A1(n10801), .A2(n11662), .B1(n7011), .B2(n11982), .ZN(
        n10803) );
  NOR2_X1 U13430 ( .A1(n14150), .A2(n11669), .ZN(n10802) );
  AOI211_X1 U13431 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n10804), .A(n10803), .B(
        n10802), .ZN(n10805) );
  OAI21_X1 U13432 ( .B1(n14165), .B2(n10806), .A(n10805), .ZN(P1_U3222) );
  INV_X1 U13433 ( .A(n10807), .ZN(n10808) );
  NOR3_X1 U13434 ( .A1(n10809), .A2(n10808), .A3(n15495), .ZN(n10810) );
  AOI21_X1 U13435 ( .B1(n15398), .B2(n10999), .A(n10810), .ZN(n10984) );
  XNOR2_X1 U13436 ( .A(n13236), .B(n13234), .ZN(n10813) );
  NAND2_X1 U13437 ( .A1(n10923), .A2(n10811), .ZN(n10812) );
  NOR2_X1 U13438 ( .A1(n10813), .A2(n10812), .ZN(n10982) );
  NAND2_X1 U13439 ( .A1(n12850), .A2(n13115), .ZN(n10814) );
  OAI21_X1 U13440 ( .B1(n10815), .B2(n15512), .A(n10814), .ZN(n10816) );
  NAND2_X1 U13441 ( .A1(n10816), .A2(n11583), .ZN(n10817) );
  NAND2_X1 U13442 ( .A1(n10817), .A2(n10820), .ZN(n10818) );
  NAND2_X1 U13443 ( .A1(n10818), .A2(n10976), .ZN(n10823) );
  OR3_X1 U13444 ( .A1(n11577), .A2(n11107), .A3(n10819), .ZN(n11586) );
  NAND2_X1 U13445 ( .A1(n11586), .A2(n10820), .ZN(n10977) );
  NAND2_X1 U13446 ( .A1(n10975), .A2(n10977), .ZN(n10821) );
  NAND2_X1 U13447 ( .A1(n10821), .A2(n13234), .ZN(n10822) );
  NAND2_X1 U13448 ( .A1(n15532), .A2(n15495), .ZN(n13168) );
  OAI22_X1 U13449 ( .A1(n13168), .A2(n10927), .B1(n15532), .B2(n10519), .ZN(
        n10825) );
  INV_X1 U13450 ( .A(n10825), .ZN(n10826) );
  OAI21_X1 U13451 ( .B1(n10984), .B2(n15530), .A(n10826), .ZN(P3_U3459) );
  MUX2_X1 U13452 ( .A(n10828), .B(P2_REG1_REG_12__SCAN_IN), .S(n11135), .Z(
        n10829) );
  NAND2_X1 U13453 ( .A1(n10830), .A2(n10829), .ZN(n11131) );
  OAI21_X1 U13454 ( .B1(n10830), .B2(n10829), .A(n11131), .ZN(n10841) );
  INV_X1 U13455 ( .A(n15319), .ZN(n15299) );
  OR2_X1 U13456 ( .A1(n10831), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10834) );
  NAND2_X1 U13457 ( .A1(n10836), .A2(n10834), .ZN(n10832) );
  MUX2_X1 U13458 ( .A(n11935), .B(P2_REG2_REG_12__SCAN_IN), .S(n11135), .Z(
        n10833) );
  NAND2_X1 U13459 ( .A1(n10832), .A2(n10833), .ZN(n11137) );
  INV_X1 U13460 ( .A(n10833), .ZN(n10835) );
  NAND3_X1 U13461 ( .A1(n10836), .A2(n10835), .A3(n10834), .ZN(n10837) );
  INV_X1 U13462 ( .A(n15306), .ZN(n15330) );
  AOI21_X1 U13463 ( .B1(n11137), .B2(n10837), .A(n15330), .ZN(n10840) );
  NAND2_X1 U13464 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11864)
         );
  NAND2_X1 U13465 ( .A1(n15328), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n10838) );
  OAI211_X1 U13466 ( .C1(n15325), .C2(n11135), .A(n11864), .B(n10838), .ZN(
        n10839) );
  AOI211_X1 U13467 ( .C1(n10841), .C2(n15299), .A(n10840), .B(n10839), .ZN(
        n10842) );
  INV_X1 U13468 ( .A(n10842), .ZN(P2_U3226) );
  AOI21_X1 U13469 ( .B1(n10760), .B2(n10843), .A(n6719), .ZN(n10849) );
  INV_X1 U13470 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15581) );
  NOR2_X1 U13471 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15581), .ZN(n11067) );
  INV_X1 U13472 ( .A(n10844), .ZN(n12693) );
  NAND2_X1 U13473 ( .A1(n10845), .A2(n10759), .ZN(n10846) );
  AOI21_X1 U13474 ( .B1(n12693), .B2(n10846), .A(n12855), .ZN(n10847) );
  AOI211_X1 U13475 ( .C1(n15392), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n11067), .B(
        n10847), .ZN(n10848) );
  OAI21_X1 U13476 ( .B1(n10849), .B2(n12847), .A(n10848), .ZN(n10850) );
  AOI21_X1 U13477 ( .B1(n10851), .B2(n12822), .A(n10850), .ZN(n10858) );
  INV_X1 U13478 ( .A(n12687), .ZN(n10856) );
  NOR3_X1 U13479 ( .A1(n10854), .A2(n10853), .A3(n10852), .ZN(n10855) );
  OAI21_X1 U13480 ( .B1(n10856), .B2(n10855), .A(n12853), .ZN(n10857) );
  NAND2_X1 U13481 ( .A1(n10858), .A2(n10857), .ZN(P3_U3185) );
  OAI21_X1 U13482 ( .B1(n10876), .B2(n15426), .A(n15428), .ZN(n10859) );
  INV_X1 U13483 ( .A(n10859), .ZN(n10866) );
  NAND2_X1 U13484 ( .A1(n10860), .A2(n11107), .ZN(n10861) );
  AND2_X1 U13485 ( .A1(n11583), .A2(n10861), .ZN(n10865) );
  INV_X1 U13486 ( .A(n10862), .ZN(n10863) );
  NAND2_X1 U13487 ( .A1(n13236), .A2(n10863), .ZN(n10864) );
  MUX2_X1 U13488 ( .A(n10867), .B(n10866), .S(n12532), .Z(n10872) );
  NAND2_X1 U13489 ( .A1(n15445), .A2(n12532), .ZN(n10868) );
  INV_X1 U13490 ( .A(n15457), .ZN(n10870) );
  OAI211_X1 U13491 ( .C1(n10872), .C2(n15445), .A(n10994), .B(n10871), .ZN(
        n10873) );
  NAND2_X1 U13492 ( .A1(n10873), .A2(n7432), .ZN(n10879) );
  INV_X1 U13493 ( .A(n10874), .ZN(n11581) );
  NAND2_X1 U13494 ( .A1(n10875), .A2(n11581), .ZN(n12677) );
  OAI22_X1 U13495 ( .A1(n15451), .A2(n12668), .B1(n12684), .B2(n10876), .ZN(
        n10877) );
  AOI21_X1 U13496 ( .B1(n12657), .B2(n15448), .A(n10877), .ZN(n10878) );
  OAI211_X1 U13497 ( .C1(n11002), .C2(n15459), .A(n10879), .B(n10878), .ZN(
        P3_U3162) );
  INV_X1 U13498 ( .A(n10880), .ZN(n10884) );
  NOR3_X1 U13499 ( .A1(n12689), .A2(n10882), .A3(n10881), .ZN(n10883) );
  OAI21_X1 U13500 ( .B1(n10884), .B2(n10883), .A(n12853), .ZN(n10896) );
  AOI21_X1 U13501 ( .B1(n10770), .B2(n10886), .A(n10885), .ZN(n10892) );
  NOR2_X1 U13502 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8720), .ZN(n12611) );
  AOI21_X1 U13503 ( .B1(n11607), .B2(n10888), .A(n10887), .ZN(n10889) );
  NOR2_X1 U13504 ( .A1(n10889), .A2(n12847), .ZN(n10890) );
  AOI211_X1 U13505 ( .C1(n15392), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n12611), .B(
        n10890), .ZN(n10891) );
  OAI21_X1 U13506 ( .B1(n10892), .B2(n12855), .A(n10891), .ZN(n10893) );
  AOI21_X1 U13507 ( .B1(n10894), .B2(n12822), .A(n10893), .ZN(n10895) );
  NAND2_X1 U13508 ( .A1(n10896), .A2(n10895), .ZN(P3_U3187) );
  INV_X1 U13509 ( .A(n10901), .ZN(n10897) );
  OR2_X1 U13510 ( .A1(n13362), .A2(n10899), .ZN(n10900) );
  XNOR2_X1 U13511 ( .A(n11083), .B(n11070), .ZN(n11246) );
  NAND2_X1 U13512 ( .A1(n10902), .A2(n10901), .ZN(n10904) );
  OR2_X1 U13513 ( .A1(n13362), .A2(n11201), .ZN(n10903) );
  NAND2_X1 U13514 ( .A1(n10904), .A2(n10903), .ZN(n11071) );
  XNOR2_X1 U13515 ( .A(n11071), .B(n11070), .ZN(n11236) );
  OR2_X1 U13516 ( .A1(n10905), .A2(n11240), .ZN(n10906) );
  AND3_X1 U13517 ( .A1(n11110), .A2(n10906), .A3(n14928), .ZN(n11243) );
  OAI21_X1 U13518 ( .B1(n11240), .B2(n15381), .A(n11237), .ZN(n10907) );
  AOI211_X1 U13519 ( .C1(n11236), .C2(n14915), .A(n11243), .B(n10907), .ZN(
        n10908) );
  OAI21_X1 U13520 ( .B1(n13842), .B2(n11246), .A(n10908), .ZN(n10910) );
  NAND2_X1 U13521 ( .A1(n10910), .A2(n15387), .ZN(n10909) );
  OAI21_X1 U13522 ( .B1(n15387), .B2(n8004), .A(n10909), .ZN(P2_U3445) );
  NAND2_X1 U13523 ( .A1(n10910), .A2(n15391), .ZN(n10911) );
  OAI21_X1 U13524 ( .B1(n15391), .B2(n10912), .A(n10911), .ZN(P2_U3504) );
  INV_X1 U13525 ( .A(n15284), .ZN(n10915) );
  INV_X1 U13526 ( .A(n10913), .ZN(n10917) );
  OAI222_X1 U13527 ( .A1(P2_U3088), .A2(n10915), .B1(n13883), .B2(n10917), 
        .C1(n10914), .C2(n13894), .ZN(P2_U3313) );
  INV_X1 U13528 ( .A(n12018), .ZN(n12026) );
  OAI222_X1 U13529 ( .A1(P1_U3086), .A2(n12026), .B1(n14694), .B2(n10917), 
        .C1(n10916), .C2(n14691), .ZN(P1_U3341) );
  OAI21_X1 U13530 ( .B1(n10920), .B2(n10919), .A(n10918), .ZN(n10922) );
  NAND2_X1 U13531 ( .A1(n10922), .A2(n10921), .ZN(n10926) );
  NAND3_X1 U13532 ( .A1(n10924), .A2(n10923), .A3(n11585), .ZN(n10925) );
  AND2_X2 U13533 ( .A1(n10926), .A2(n10925), .ZN(n15517) );
  INV_X2 U13534 ( .A(n15517), .ZN(n15519) );
  OAI22_X1 U13535 ( .A1(n10927), .A2(n13229), .B1(n15519), .B2(n8649), .ZN(
        n10928) );
  INV_X1 U13536 ( .A(n10928), .ZN(n10929) );
  OAI21_X1 U13537 ( .B1(n10984), .B2(n15517), .A(n10929), .ZN(P3_U3390) );
  AOI22_X1 U13538 ( .A1(n11257), .A2(n12094), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10941), .ZN(n10935) );
  OR2_X1 U13539 ( .A1(n10931), .A2(n10930), .ZN(n10932) );
  OAI21_X1 U13540 ( .B1(n10933), .B2(n11846), .A(n10932), .ZN(n10934) );
  NOR2_X1 U13541 ( .A1(n10935), .A2(n10934), .ZN(n11258) );
  AOI21_X1 U13542 ( .B1(n10935), .B2(n10934), .A(n11258), .ZN(n10945) );
  AOI22_X1 U13543 ( .A1(n11257), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9752), 
        .B2(n10941), .ZN(n10939) );
  OAI21_X1 U13544 ( .B1(n10939), .B2(n10938), .A(n11247), .ZN(n10943) );
  AND2_X1 U13545 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n12277) );
  AOI21_X1 U13546 ( .B1(n15027), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n12277), 
        .ZN(n10940) );
  OAI21_X1 U13547 ( .B1(n10941), .B2(n15064), .A(n10940), .ZN(n10942) );
  AOI21_X1 U13548 ( .B1(n10943), .B2(n15059), .A(n10942), .ZN(n10944) );
  OAI21_X1 U13549 ( .B1(n10945), .B2(n15055), .A(n10944), .ZN(P1_U3255) );
  INV_X1 U13550 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15526) );
  OR2_X1 U13551 ( .A1(n10964), .A2(n10946), .ZN(n10947) );
  AOI21_X1 U13552 ( .B1(n15526), .B2(n10949), .A(n11020), .ZN(n10973) );
  INV_X1 U13553 ( .A(n10950), .ZN(n10957) );
  MUX2_X1 U13554 ( .A(n10951), .B(n15526), .S(n12814), .Z(n10952) );
  NAND2_X1 U13555 ( .A1(n10952), .A2(n11019), .ZN(n11015) );
  INV_X1 U13556 ( .A(n10952), .ZN(n10954) );
  NAND2_X1 U13557 ( .A1(n10954), .A2(n10953), .ZN(n10955) );
  AND2_X1 U13558 ( .A1(n11015), .A2(n10955), .ZN(n10956) );
  INV_X1 U13559 ( .A(n11016), .ZN(n10960) );
  NOR3_X1 U13560 ( .A1(n10958), .A2(n10957), .A3(n10956), .ZN(n10959) );
  OAI21_X1 U13561 ( .B1(n10960), .B2(n10959), .A(n12853), .ZN(n10972) );
  INV_X1 U13562 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10962) );
  INV_X1 U13563 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15587) );
  NOR2_X1 U13564 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15587), .ZN(n12496) );
  INV_X1 U13565 ( .A(n12496), .ZN(n10961) );
  OAI21_X1 U13566 ( .B1(n12813), .B2(n10962), .A(n10961), .ZN(n10970) );
  OR2_X1 U13567 ( .A1(n10964), .A2(n10963), .ZN(n10965) );
  AOI21_X1 U13568 ( .B1(n10951), .B2(n10967), .A(n11004), .ZN(n10968) );
  NOR2_X1 U13569 ( .A1(n10968), .A2(n12847), .ZN(n10969) );
  AOI211_X1 U13570 ( .C1(n12822), .C2(n11019), .A(n10970), .B(n10969), .ZN(
        n10971) );
  OAI211_X1 U13571 ( .C1(n10973), .C2(n12855), .A(n10972), .B(n10971), .ZN(
        P3_U3189) );
  INV_X1 U13572 ( .A(n10977), .ZN(n10974) );
  NAND2_X1 U13573 ( .A1(n10974), .A2(n10976), .ZN(n10980) );
  NAND2_X1 U13574 ( .A1(n10976), .A2(n10975), .ZN(n10978) );
  NAND2_X1 U13575 ( .A1(n10978), .A2(n10977), .ZN(n10979) );
  AND2_X1 U13576 ( .A1(n10980), .A2(n10979), .ZN(n10981) );
  NAND2_X1 U13577 ( .A1(n10982), .A2(n10981), .ZN(n10986) );
  NAND2_X2 U13578 ( .A1(n10986), .A2(n15458), .ZN(n15463) );
  MUX2_X1 U13579 ( .A(n10985), .B(n10984), .S(n15463), .Z(n10989) );
  OR2_X1 U13580 ( .A1(n10986), .A2(n15455), .ZN(n11774) );
  NAND2_X1 U13581 ( .A1(n15419), .A2(n15495), .ZN(n13104) );
  AOI22_X1 U13582 ( .A1(n13085), .A2(n10987), .B1(n15442), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U13583 ( .A1(n10989), .A2(n10988), .ZN(P3_U3233) );
  INV_X1 U13584 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n15809) );
  INV_X1 U13585 ( .A(n12997), .ZN(n12892) );
  NAND2_X1 U13586 ( .A1(n12892), .A2(n11422), .ZN(n10990) );
  OAI21_X1 U13587 ( .B1(n11422), .B2(n15809), .A(n10990), .ZN(P3_U3514) );
  XNOR2_X1 U13588 ( .A(n10991), .B(n12532), .ZN(n11059) );
  XNOR2_X1 U13589 ( .A(n11059), .B(n15451), .ZN(n10996) );
  NAND2_X1 U13590 ( .A1(n15426), .A2(n10992), .ZN(n10993) );
  NAND2_X1 U13591 ( .A1(n10994), .A2(n10993), .ZN(n10995) );
  NAND2_X1 U13592 ( .A1(n10995), .A2(n10996), .ZN(n11063) );
  OAI21_X1 U13593 ( .B1(n10996), .B2(n10995), .A(n11063), .ZN(n10997) );
  NAND2_X1 U13594 ( .A1(n10997), .A2(n7432), .ZN(n11001) );
  OAI22_X1 U13595 ( .A1(n15424), .A2(n12668), .B1(n12684), .B2(n15437), .ZN(
        n10998) );
  AOI21_X1 U13596 ( .B1(n12657), .B2(n10999), .A(n10998), .ZN(n11000) );
  OAI211_X1 U13597 ( .C1(n11002), .C2(n8670), .A(n11001), .B(n11000), .ZN(
        P3_U3177) );
  NOR2_X1 U13598 ( .A1(n11019), .A2(n11003), .ZN(n11005) );
  MUX2_X1 U13599 ( .A(n11009), .B(P3_REG2_REG_8__SCAN_IN), .S(n11165), .Z(
        n11007) );
  INV_X1 U13600 ( .A(n11167), .ZN(n11006) );
  AOI21_X1 U13601 ( .B1(n11008), .B2(n11007), .A(n11006), .ZN(n11034) );
  MUX2_X1 U13602 ( .A(n11009), .B(n11022), .S(n12814), .Z(n11011) );
  NAND2_X1 U13603 ( .A1(n11011), .A2(n11010), .ZN(n11154) );
  INV_X1 U13604 ( .A(n11011), .ZN(n11012) );
  NAND2_X1 U13605 ( .A1(n11012), .A2(n11165), .ZN(n11013) );
  NAND2_X1 U13606 ( .A1(n11154), .A2(n11013), .ZN(n11014) );
  AND3_X1 U13607 ( .A1(n11016), .A2(n11015), .A3(n11014), .ZN(n11017) );
  OAI21_X1 U13608 ( .B1(n11162), .B2(n11017), .A(n12853), .ZN(n11033) );
  NOR2_X1 U13609 ( .A1(n11019), .A2(n11018), .ZN(n11021) );
  INV_X1 U13610 ( .A(n11024), .ZN(n11026) );
  MUX2_X1 U13611 ( .A(n11022), .B(P3_REG1_REG_8__SCAN_IN), .S(n11165), .Z(
        n11023) );
  INV_X1 U13612 ( .A(n11023), .ZN(n11025) );
  OR2_X2 U13613 ( .A1(n11024), .A2(n11023), .ZN(n11152) );
  OAI21_X1 U13614 ( .B1(n11026), .B2(n11025), .A(n11152), .ZN(n11031) );
  NOR2_X1 U13615 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11027), .ZN(n12579) );
  AOI21_X1 U13616 ( .B1(n15392), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12579), .ZN(
        n11028) );
  OAI21_X1 U13617 ( .B1(n12851), .B2(n11165), .A(n11028), .ZN(n11029) );
  AOI21_X1 U13618 ( .B1(n11031), .B2(n11030), .A(n11029), .ZN(n11032) );
  OAI211_X1 U13619 ( .C1(n11034), .C2(n12847), .A(n11033), .B(n11032), .ZN(
        P3_U3190) );
  AOI21_X1 U13620 ( .B1(n11036), .B2(n11035), .A(n13342), .ZN(n11037) );
  NAND2_X1 U13621 ( .A1(n11037), .A2(n7108), .ZN(n11042) );
  NAND2_X1 U13622 ( .A1(n13361), .A2(n13307), .ZN(n11039) );
  NAND2_X1 U13623 ( .A1(n13359), .A2(n13336), .ZN(n11038) );
  AND2_X1 U13624 ( .A1(n11039), .A2(n11038), .ZN(n11114) );
  INV_X1 U13625 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n13404) );
  OAI22_X1 U13626 ( .A1(n13339), .A2(n11114), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13404), .ZN(n11040) );
  AOI21_X1 U13627 ( .B1(n11211), .B2(n14908), .A(n11040), .ZN(n11041) );
  OAI211_X1 U13628 ( .C1(n14911), .C2(n11212), .A(n11042), .B(n11041), .ZN(
        P2_U3211) );
  INV_X1 U13629 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n11044) );
  NAND2_X1 U13630 ( .A1(n12986), .A2(n11422), .ZN(n11043) );
  OAI21_X1 U13631 ( .B1(n11422), .B2(n11044), .A(n11043), .ZN(P3_U3515) );
  INV_X1 U13632 ( .A(n12853), .ZN(n12819) );
  NAND3_X1 U13633 ( .A1(n12855), .A2(n12847), .A3(n12819), .ZN(n11055) );
  OR2_X1 U13634 ( .A1(n12847), .A2(n11045), .ZN(n11049) );
  NOR2_X1 U13635 ( .A1(n11046), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11047) );
  AOI21_X1 U13636 ( .B1(n15392), .B2(P3_ADDR_REG_0__SCAN_IN), .A(n11047), .ZN(
        n11048) );
  OAI211_X1 U13637 ( .C1(n12855), .C2(n11050), .A(n11049), .B(n11048), .ZN(
        n11054) );
  NOR2_X1 U13638 ( .A1(n12819), .A2(n11051), .ZN(n11052) );
  MUX2_X1 U13639 ( .A(n11052), .B(n12822), .S(P3_IR_REG_0__SCAN_IN), .Z(n11053) );
  AOI211_X1 U13640 ( .C1(n11056), .C2(n11055), .A(n11054), .B(n11053), .ZN(
        n11057) );
  INV_X1 U13641 ( .A(n11057), .ZN(P3_U3182) );
  INV_X1 U13642 ( .A(n12666), .ZN(n12678) );
  INV_X1 U13643 ( .A(n11059), .ZN(n11060) );
  NAND2_X1 U13644 ( .A1(n11060), .A2(n15451), .ZN(n11061) );
  AND2_X1 U13645 ( .A1(n11063), .A2(n11061), .ZN(n11065) );
  XNOR2_X1 U13646 ( .A(n11574), .B(n12532), .ZN(n11314) );
  XNOR2_X1 U13647 ( .A(n11314), .B(n15424), .ZN(n11064) );
  AND2_X1 U13648 ( .A1(n11064), .A2(n11061), .ZN(n11062) );
  NAND2_X1 U13649 ( .A1(n11063), .A2(n11062), .ZN(n11316) );
  OAI211_X1 U13650 ( .C1(n11065), .C2(n11064), .A(n7432), .B(n11316), .ZN(
        n11069) );
  OAI22_X1 U13651 ( .A1(n15408), .A2(n12668), .B1(n15451), .B2(n12677), .ZN(
        n11066) );
  AOI211_X1 U13652 ( .C1(n12670), .C2(n11574), .A(n11067), .B(n11066), .ZN(
        n11068) );
  OAI211_X1 U13653 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12678), .A(n11069), .B(
        n11068), .ZN(P3_U3158) );
  INV_X1 U13654 ( .A(n13361), .ZN(n11072) );
  NAND2_X1 U13655 ( .A1(n11072), .A2(n11084), .ZN(n11073) );
  INV_X1 U13656 ( .A(n13360), .ZN(n11121) );
  NAND2_X1 U13657 ( .A1(n11211), .A2(n11121), .ZN(n11075) );
  INV_X1 U13658 ( .A(n11087), .ZN(n11369) );
  XNOR2_X1 U13659 ( .A(n11374), .B(n11369), .ZN(n11187) );
  AND2_X1 U13660 ( .A1(n11076), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11080) );
  INV_X1 U13661 ( .A(n11077), .ZN(n11079) );
  NAND4_X1 U13662 ( .A1(n11080), .A2(n11079), .A3(n11078), .A4(n15367), .ZN(
        n11081) );
  NAND2_X1 U13663 ( .A1(n13741), .A2(n14915), .ZN(n13688) );
  NOR2_X1 U13664 ( .A1(n13361), .A2(n11084), .ZN(n11082) );
  NAND2_X1 U13665 ( .A1(n11109), .A2(n7339), .ZN(n11086) );
  NAND2_X1 U13666 ( .A1(n11211), .A2(n13360), .ZN(n11085) );
  NAND2_X1 U13667 ( .A1(n11086), .A2(n11085), .ZN(n11370) );
  XNOR2_X1 U13668 ( .A(n11370), .B(n11087), .ZN(n11189) );
  NAND2_X1 U13669 ( .A1(n11933), .A2(n12465), .ZN(n11088) );
  NAND2_X1 U13670 ( .A1(n11089), .A2(n11088), .ZN(n11090) );
  NAND2_X1 U13671 ( .A1(n11111), .A2(n11375), .ZN(n11091) );
  NAND2_X1 U13672 ( .A1(n11091), .A2(n14928), .ZN(n11092) );
  OR2_X1 U13673 ( .A1(n11092), .A2(n11384), .ZN(n11185) );
  NAND2_X1 U13674 ( .A1(n13741), .A2(n12465), .ZN(n13713) );
  NAND2_X1 U13675 ( .A1(n13741), .A2(n11093), .ZN(n13743) );
  INV_X1 U13676 ( .A(n13737), .ZN(n14918) );
  INV_X1 U13677 ( .A(n11125), .ZN(n11094) );
  AOI22_X1 U13678 ( .A1(n14920), .A2(n11375), .B1(n14918), .B2(n11094), .ZN(
        n11099) );
  OR2_X1 U13679 ( .A1(n11503), .A2(n13326), .ZN(n11096) );
  NAND2_X1 U13680 ( .A1(n13360), .A2(n13307), .ZN(n11095) );
  AND2_X1 U13681 ( .A1(n11096), .A2(n11095), .ZN(n11186) );
  MUX2_X1 U13682 ( .A(n11186), .B(n11097), .S(n14935), .Z(n11098) );
  OAI211_X1 U13683 ( .C1(n11185), .C2(n13713), .A(n11099), .B(n11098), .ZN(
        n11100) );
  AOI21_X1 U13684 ( .B1(n11189), .B2(n14932), .A(n11100), .ZN(n11101) );
  OAI21_X1 U13685 ( .B1(n11187), .B2(n13688), .A(n11101), .ZN(P2_U3258) );
  INV_X1 U13686 ( .A(n12027), .ZN(n15063) );
  INV_X1 U13687 ( .A(n11102), .ZN(n11104) );
  OAI222_X1 U13688 ( .A1(P1_U3086), .A2(n15063), .B1(n14694), .B2(n11104), 
        .C1(n11103), .C2(n14691), .ZN(P1_U3340) );
  INV_X1 U13689 ( .A(n15293), .ZN(n13461) );
  OAI222_X1 U13690 ( .A1(n13894), .A2(n11105), .B1(n13892), .B2(n11104), .C1(
        n13461), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI222_X1 U13691 ( .A1(P3_U3151), .A2(n11107), .B1(n12166), .B2(n15844), 
        .C1(n6670), .C2(n11106), .ZN(P3_U3275) );
  XNOR2_X1 U13692 ( .A(n11109), .B(n11108), .ZN(n11207) );
  AOI21_X1 U13693 ( .B1(n11110), .B2(n11211), .A(n13720), .ZN(n11112) );
  AND2_X1 U13694 ( .A1(n11112), .A2(n11111), .ZN(n11215) );
  XNOR2_X1 U13695 ( .A(n11113), .B(n7339), .ZN(n11115) );
  OAI21_X1 U13696 ( .B1(n11115), .B2(n13806), .A(n11114), .ZN(n11208) );
  AOI211_X1 U13697 ( .C1(n14941), .C2(n11207), .A(n11215), .B(n11208), .ZN(
        n11118) );
  NOR2_X1 U13698 ( .A1(n15386), .A2(n15381), .ZN(n13873) );
  AOI22_X1 U13699 ( .A1(n13873), .A2(n11211), .B1(n15386), .B2(
        P2_REG0_REG_6__SCAN_IN), .ZN(n11116) );
  OAI21_X1 U13700 ( .B1(n11118), .B2(n15386), .A(n11116), .ZN(P2_U3448) );
  AOI22_X1 U13701 ( .A1(n13837), .A2(n11211), .B1(n15389), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11117) );
  OAI21_X1 U13702 ( .B1(n11118), .B2(n15389), .A(n11117), .ZN(P2_U3505) );
  AOI21_X1 U13703 ( .B1(n7108), .B2(n7571), .A(n13342), .ZN(n11124) );
  NOR3_X1 U13704 ( .A1(n11810), .A2(n11122), .A3(n11121), .ZN(n11123) );
  OAI21_X1 U13705 ( .B1(n11124), .B2(n11123), .A(n11391), .ZN(n11129) );
  NAND2_X1 U13706 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13418) );
  OAI21_X1 U13707 ( .B1(n11186), .B2(n13339), .A(n13418), .ZN(n11127) );
  NOR2_X1 U13708 ( .A1(n14911), .A2(n11125), .ZN(n11126) );
  AOI211_X1 U13709 ( .C1(n11375), .C2(n14908), .A(n11127), .B(n11126), .ZN(
        n11128) );
  NAND2_X1 U13710 ( .A1(n11129), .A2(n11128), .ZN(P2_U3185) );
  NOR2_X1 U13711 ( .A1(n11148), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11130) );
  AOI21_X1 U13712 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n11148), .A(n11130), 
        .ZN(n11134) );
  OAI21_X1 U13713 ( .B1(n11132), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11131), 
        .ZN(n11133) );
  NOR2_X1 U13714 ( .A1(n11133), .A2(n11134), .ZN(n13447) );
  AOI211_X1 U13715 ( .C1(n11134), .C2(n11133), .A(n15319), .B(n13447), .ZN(
        n11150) );
  NAND2_X1 U13716 ( .A1(n11135), .A2(n11935), .ZN(n11136) );
  NAND2_X1 U13717 ( .A1(n11137), .A2(n11136), .ZN(n11142) );
  NAND2_X1 U13718 ( .A1(n11148), .A2(n11139), .ZN(n11138) );
  OAI21_X1 U13719 ( .B1(n11148), .B2(n11139), .A(n11138), .ZN(n11140) );
  NAND2_X1 U13720 ( .A1(n11148), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11141) );
  OAI211_X1 U13721 ( .C1(P2_REG2_REG_13__SCAN_IN), .C2(n11148), .A(n11142), 
        .B(n11141), .ZN(n11143) );
  NAND3_X1 U13722 ( .A1(n13458), .A2(n11143), .A3(n15306), .ZN(n11147) );
  INV_X1 U13723 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11144) );
  NOR2_X1 U13724 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11144), .ZN(n11145) );
  AOI21_X1 U13725 ( .B1(n15328), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n11145), 
        .ZN(n11146) );
  OAI211_X1 U13726 ( .C1(n15325), .C2(n11148), .A(n11147), .B(n11146), .ZN(
        n11149) );
  OR2_X1 U13727 ( .A1(n11150), .A2(n11149), .ZN(P2_U3227) );
  NAND2_X1 U13728 ( .A1(n11165), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11151) );
  AOI21_X1 U13729 ( .B1(n11155), .B2(n11153), .A(n11439), .ZN(n11175) );
  INV_X1 U13730 ( .A(n11154), .ZN(n11161) );
  MUX2_X1 U13731 ( .A(n12158), .B(n11155), .S(n12814), .Z(n11156) );
  NAND2_X1 U13732 ( .A1(n11156), .A2(n11438), .ZN(n11427) );
  INV_X1 U13733 ( .A(n11156), .ZN(n11158) );
  NAND2_X1 U13734 ( .A1(n11158), .A2(n11157), .ZN(n11159) );
  AND2_X1 U13735 ( .A1(n11427), .A2(n11159), .ZN(n11160) );
  INV_X1 U13736 ( .A(n11428), .ZN(n11164) );
  NOR3_X1 U13737 ( .A1(n11162), .A2(n11161), .A3(n11160), .ZN(n11163) );
  OAI21_X1 U13738 ( .B1(n11164), .B2(n11163), .A(n12853), .ZN(n11174) );
  NAND2_X1 U13739 ( .A1(n11165), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11166) );
  AOI21_X1 U13740 ( .B1(n12158), .B2(n11168), .A(n11431), .ZN(n11171) );
  NOR2_X1 U13741 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8790), .ZN(n12130) );
  AOI21_X1 U13742 ( .B1(n15392), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12130), .ZN(
        n11170) );
  NAND2_X1 U13743 ( .A1(n12822), .A2(n11438), .ZN(n11169) );
  OAI211_X1 U13744 ( .C1(n11171), .C2(n12847), .A(n11170), .B(n11169), .ZN(
        n11172) );
  INV_X1 U13745 ( .A(n11172), .ZN(n11173) );
  OAI211_X1 U13746 ( .C1(n11175), .C2(n12855), .A(n11174), .B(n11173), .ZN(
        P3_U3191) );
  INV_X1 U13747 ( .A(n14932), .ZN(n13751) );
  INV_X1 U13748 ( .A(n13688), .ZN(n13748) );
  AOI22_X1 U13749 ( .A1(n14920), .A2(n8585), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n14918), .ZN(n11179) );
  MUX2_X1 U13750 ( .A(n11177), .B(n11176), .S(n14935), .Z(n11178) );
  OAI211_X1 U13751 ( .C1(n11180), .C2(n13713), .A(n11179), .B(n11178), .ZN(
        n11181) );
  AOI21_X1 U13752 ( .B1(n13748), .B2(n11182), .A(n11181), .ZN(n11183) );
  OAI21_X1 U13753 ( .B1(n13751), .B2(n11184), .A(n11183), .ZN(P2_U3264) );
  OAI211_X1 U13754 ( .C1(n11187), .C2(n13806), .A(n11186), .B(n11185), .ZN(
        n11188) );
  AOI21_X1 U13755 ( .B1(n14941), .B2(n11189), .A(n11188), .ZN(n11192) );
  AOI22_X1 U13756 ( .A1(n13837), .A2(n11375), .B1(n15389), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11190) );
  OAI21_X1 U13757 ( .B1(n11192), .B2(n15389), .A(n11190), .ZN(P2_U3506) );
  AOI22_X1 U13758 ( .A1(n13873), .A2(n11375), .B1(n15386), .B2(
        P2_REG0_REG_7__SCAN_IN), .ZN(n11191) );
  OAI21_X1 U13759 ( .B1(n11192), .B2(n15386), .A(n11191), .ZN(P2_U3451) );
  INV_X1 U13760 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n15641) );
  NAND2_X1 U13761 ( .A1(n12897), .A2(n11422), .ZN(n11193) );
  OAI21_X1 U13762 ( .B1(n11422), .B2(n15641), .A(n11193), .ZN(P3_U3516) );
  INV_X1 U13763 ( .A(n14234), .ZN(n14230) );
  INV_X1 U13764 ( .A(n11194), .ZN(n11197) );
  OAI222_X1 U13765 ( .A1(P1_U3086), .A2(n14230), .B1(n14694), .B2(n11197), 
        .C1(n11195), .C2(n14691), .ZN(P1_U3339) );
  INV_X1 U13766 ( .A(n13481), .ZN(n13475) );
  OAI222_X1 U13767 ( .A1(P2_U3088), .A2(n13475), .B1(n13892), .B2(n11197), 
        .C1(n11196), .C2(n13894), .ZN(P2_U3311) );
  MUX2_X1 U13768 ( .A(n11199), .B(n11198), .S(n13741), .Z(n11205) );
  OAI22_X1 U13769 ( .A1(n13743), .A2(n11201), .B1(n11200), .B2(n13737), .ZN(
        n11202) );
  AOI21_X1 U13770 ( .B1(n11203), .B2(n14931), .A(n11202), .ZN(n11204) );
  OAI211_X1 U13771 ( .C1(n13751), .C2(n11206), .A(n11205), .B(n11204), .ZN(
        P2_U3261) );
  INV_X1 U13772 ( .A(n11207), .ZN(n11218) );
  INV_X1 U13773 ( .A(n11208), .ZN(n11209) );
  MUX2_X1 U13774 ( .A(n11210), .B(n11209), .S(n13741), .Z(n11217) );
  INV_X1 U13775 ( .A(n11211), .ZN(n11213) );
  OAI22_X1 U13776 ( .A1(n13743), .A2(n11213), .B1(n13737), .B2(n11212), .ZN(
        n11214) );
  AOI21_X1 U13777 ( .B1(n11215), .B2(n14931), .A(n11214), .ZN(n11216) );
  OAI211_X1 U13778 ( .C1(n13751), .C2(n11218), .A(n11217), .B(n11216), .ZN(
        P2_U3259) );
  MUX2_X1 U13779 ( .A(n11220), .B(n11219), .S(n13741), .Z(n11225) );
  OAI22_X1 U13780 ( .A1(n13743), .A2(n11221), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13737), .ZN(n11222) );
  AOI21_X1 U13781 ( .B1(n11223), .B2(n14931), .A(n11222), .ZN(n11224) );
  OAI211_X1 U13782 ( .C1(n13751), .C2(n11226), .A(n11225), .B(n11224), .ZN(
        P2_U3262) );
  AOI21_X1 U13783 ( .B1(n14931), .B2(n11227), .A(n14920), .ZN(n11235) );
  INV_X1 U13784 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n13370) );
  OAI22_X1 U13785 ( .A1(n13741), .A2(n13370), .B1(n12473), .B2(n13737), .ZN(
        n11232) );
  NAND2_X1 U13786 ( .A1(n6686), .A2(n11228), .ZN(n11229) );
  NOR2_X1 U13787 ( .A1(n14919), .A2(n11229), .ZN(n13661) );
  INV_X1 U13788 ( .A(n13661), .ZN(n11942) );
  NOR2_X1 U13789 ( .A1(n11942), .A2(n11230), .ZN(n11231) );
  AOI211_X1 U13790 ( .C1(n13741), .C2(n11233), .A(n11232), .B(n11231), .ZN(
        n11234) );
  OAI21_X1 U13791 ( .B1(n11235), .B2(n7919), .A(n11234), .ZN(P2_U3265) );
  NAND2_X1 U13792 ( .A1(n11236), .A2(n13748), .ZN(n11245) );
  INV_X1 U13793 ( .A(n11237), .ZN(n11238) );
  MUX2_X1 U13794 ( .A(n11238), .B(P2_REG2_REG_5__SCAN_IN), .S(n14935), .Z(
        n11242) );
  OAI22_X1 U13795 ( .A1(n13743), .A2(n11240), .B1(n13737), .B2(n11239), .ZN(
        n11241) );
  AOI211_X1 U13796 ( .C1(n11243), .C2(n14931), .A(n11242), .B(n11241), .ZN(
        n11244) );
  OAI211_X1 U13797 ( .C1(n11246), .C2(n13751), .A(n11245), .B(n11244), .ZN(
        P2_U3260) );
  OAI21_X1 U13798 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n11257), .A(n11247), 
        .ZN(n11252) );
  OR2_X1 U13799 ( .A1(n11339), .A2(n11248), .ZN(n11250) );
  NAND2_X1 U13800 ( .A1(n11339), .A2(n11248), .ZN(n11249) );
  AND2_X1 U13801 ( .A1(n11250), .A2(n11249), .ZN(n11251) );
  AOI211_X1 U13802 ( .C1(n11252), .C2(n11251), .A(n11338), .B(n15036), .ZN(
        n11256) );
  NAND2_X1 U13803 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n12319)
         );
  INV_X1 U13804 ( .A(n12319), .ZN(n11253) );
  AOI21_X1 U13805 ( .B1(n15027), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11253), 
        .ZN(n11254) );
  OAI21_X1 U13806 ( .B1(n15064), .B2(n11261), .A(n11254), .ZN(n11255) );
  NOR2_X1 U13807 ( .A1(n11256), .A2(n11255), .ZN(n11265) );
  NOR2_X1 U13808 ( .A1(n11257), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11259) );
  NOR2_X1 U13809 ( .A1(n11259), .A2(n11258), .ZN(n11263) );
  NAND2_X1 U13810 ( .A1(n11339), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11332) );
  INV_X1 U13811 ( .A(n11332), .ZN(n11260) );
  AOI21_X1 U13812 ( .B1(n12055), .B2(n11261), .A(n11260), .ZN(n11262) );
  NAND2_X1 U13813 ( .A1(n11262), .A2(n11263), .ZN(n11331) );
  OAI211_X1 U13814 ( .C1(n11263), .C2(n11262), .A(n15046), .B(n11331), .ZN(
        n11264) );
  NAND2_X1 U13815 ( .A1(n11265), .A2(n11264), .ZN(P1_U3256) );
  INV_X1 U13816 ( .A(n11266), .ZN(n11267) );
  NAND2_X1 U13817 ( .A1(n11268), .A2(n11267), .ZN(n11269) );
  NAND2_X1 U13818 ( .A1(n11269), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11270) );
  NAND2_X1 U13819 ( .A1(n11270), .A2(n12142), .ZN(n14124) );
  INV_X1 U13820 ( .A(n11273), .ZN(n11274) );
  NAND2_X1 U13821 ( .A1(n14026), .A2(n14042), .ZN(n11278) );
  NAND2_X1 U13822 ( .A1(n14179), .A2(n6666), .ZN(n11277) );
  NAND2_X1 U13823 ( .A1(n11278), .A2(n11277), .ZN(n11279) );
  XNOR2_X1 U13824 ( .A(n11279), .B(n14043), .ZN(n11282) );
  NAND2_X1 U13825 ( .A1(n14179), .A2(n14045), .ZN(n11280) );
  NAND2_X1 U13826 ( .A1(n11282), .A2(n11281), .ZN(n11283) );
  OR2_X1 U13827 ( .A1(n14023), .A2(n13940), .ZN(n11285) );
  NAND2_X1 U13828 ( .A1(n6901), .A2(n6666), .ZN(n11284) );
  AND2_X1 U13829 ( .A1(n11285), .A2(n11284), .ZN(n11348) );
  OAI22_X1 U13830 ( .A1(n14023), .A2(n13941), .B1(n15167), .B2(n13942), .ZN(
        n11286) );
  XNOR2_X1 U13831 ( .A(n11286), .B(n14043), .ZN(n11287) );
  OAI211_X1 U13832 ( .C1(n11288), .C2(n11287), .A(n11352), .B(n14142), .ZN(
        n11294) );
  NAND2_X1 U13833 ( .A1(n14179), .A2(n14521), .ZN(n11290) );
  NAND2_X1 U13834 ( .A1(n14178), .A2(n14281), .ZN(n11289) );
  AND2_X1 U13835 ( .A1(n11290), .A2(n11289), .ZN(n15165) );
  INV_X1 U13836 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n11291) );
  OAI22_X1 U13837 ( .A1(n14133), .A2(n15165), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11291), .ZN(n11292) );
  AOI21_X1 U13838 ( .B1(n14163), .B2(n6901), .A(n11292), .ZN(n11293) );
  OAI211_X1 U13839 ( .C1(n14161), .C2(n11534), .A(n11294), .B(n11293), .ZN(
        P1_U3230) );
  OAI222_X1 U13840 ( .A1(P3_U3151), .A2(n11565), .B1(n12166), .B2(n11296), 
        .C1(n6670), .C2(n11295), .ZN(P3_U3274) );
  INV_X1 U13841 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n11298) );
  NAND2_X1 U13842 ( .A1(n12898), .A2(n11422), .ZN(n11297) );
  OAI21_X1 U13843 ( .B1(n11422), .B2(n11298), .A(n11297), .ZN(P3_U3517) );
  OR2_X1 U13844 ( .A1(n11503), .A2(n13544), .ZN(n11300) );
  OR2_X1 U13845 ( .A1(n13354), .A2(n13326), .ZN(n11299) );
  NAND2_X1 U13846 ( .A1(n11300), .A2(n11299), .ZN(n11509) );
  NAND2_X1 U13847 ( .A1(n14905), .A2(n11509), .ZN(n11301) );
  NAND2_X1 U13848 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n15272) );
  OAI211_X1 U13849 ( .C1(n14911), .C2(n11514), .A(n11301), .B(n15272), .ZN(
        n11302) );
  AOI21_X1 U13850 ( .B1(n11677), .B2(n14908), .A(n11302), .ZN(n11308) );
  INV_X1 U13851 ( .A(n11303), .ZN(n11306) );
  OAI22_X1 U13852 ( .A1(n11304), .A2(n13342), .B1(n11810), .B2(n11503), .ZN(
        n11305) );
  NAND3_X1 U13853 ( .A1(n11400), .A2(n11306), .A3(n11305), .ZN(n11307) );
  OAI211_X1 U13854 ( .C1(n11309), .C2(n13342), .A(n11308), .B(n11307), .ZN(
        P2_U3203) );
  INV_X1 U13855 ( .A(n11310), .ZN(n11312) );
  OAI222_X1 U13856 ( .A1(P1_U3086), .A2(n14246), .B1(n14694), .B2(n11312), 
        .C1(n11311), .C2(n14691), .ZN(P1_U3338) );
  INV_X1 U13857 ( .A(n15309), .ZN(n13472) );
  OAI222_X1 U13858 ( .A1(n13894), .A2(n11313), .B1(n13892), .B2(n11312), .C1(
        n13472), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U13859 ( .A1(n11575), .A2(n11314), .ZN(n11315) );
  NAND2_X1 U13860 ( .A1(n11316), .A2(n11315), .ZN(n11322) );
  XNOR2_X1 U13861 ( .A(n11597), .B(n12532), .ZN(n11317) );
  NAND2_X1 U13862 ( .A1(n11598), .A2(n11317), .ZN(n11319) );
  INV_X1 U13863 ( .A(n11317), .ZN(n11318) );
  NAND2_X1 U13864 ( .A1(n11318), .A2(n15408), .ZN(n11792) );
  NAND2_X1 U13865 ( .A1(n11319), .A2(n11792), .ZN(n11321) );
  INV_X1 U13866 ( .A(n11793), .ZN(n11320) );
  AOI21_X1 U13867 ( .B1(n11322), .B2(n11321), .A(n11320), .ZN(n11327) );
  INV_X1 U13868 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15598) );
  NOR2_X1 U13869 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15598), .ZN(n12697) );
  OAI22_X1 U13870 ( .A1(n11795), .A2(n12668), .B1(n15424), .B2(n12677), .ZN(
        n11323) );
  AOI211_X1 U13871 ( .C1(n12670), .C2(n11597), .A(n12697), .B(n11323), .ZN(
        n11326) );
  INV_X1 U13872 ( .A(n11569), .ZN(n11324) );
  NAND2_X1 U13873 ( .A1(n12666), .A2(n11324), .ZN(n11325) );
  OAI211_X1 U13874 ( .C1(n11327), .C2(n12672), .A(n11326), .B(n11325), .ZN(
        P3_U3170) );
  INV_X1 U13875 ( .A(n11328), .ZN(n11330) );
  OAI22_X1 U13876 ( .A1(n13115), .A2(P3_U3151), .B1(SI_22_), .B2(n12166), .ZN(
        n11329) );
  AOI21_X1 U13877 ( .B1(n11330), .B2(n11561), .A(n11329), .ZN(P3_U3273) );
  NAND2_X1 U13878 ( .A1(n11332), .A2(n11331), .ZN(n11335) );
  NOR2_X1 U13879 ( .A1(n12026), .A2(n12256), .ZN(n11333) );
  AOI21_X1 U13880 ( .B1(n12256), .B2(n12026), .A(n11333), .ZN(n11334) );
  NAND2_X1 U13881 ( .A1(n11334), .A2(n11335), .ZN(n12025) );
  OAI211_X1 U13882 ( .C1(n11335), .C2(n11334), .A(n15046), .B(n12025), .ZN(
        n11347) );
  NOR2_X1 U13883 ( .A1(n12026), .A2(n11336), .ZN(n11337) );
  AOI21_X1 U13884 ( .B1(n11336), .B2(n12026), .A(n11337), .ZN(n11341) );
  OAI21_X1 U13885 ( .B1(n11341), .B2(n11340), .A(n12017), .ZN(n11345) );
  NAND2_X1 U13886 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n12410)
         );
  INV_X1 U13887 ( .A(n12410), .ZN(n11342) );
  AOI21_X1 U13888 ( .B1(n15027), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n11342), 
        .ZN(n11343) );
  OAI21_X1 U13889 ( .B1(n15064), .B2(n12026), .A(n11343), .ZN(n11344) );
  AOI21_X1 U13890 ( .B1(n15059), .B2(n11345), .A(n11344), .ZN(n11346) );
  NAND2_X1 U13891 ( .A1(n11347), .A2(n11346), .ZN(P1_U3257) );
  INV_X1 U13892 ( .A(n11348), .ZN(n11349) );
  NAND2_X1 U13893 ( .A1(n11350), .A2(n11349), .ZN(n11351) );
  NAND2_X1 U13894 ( .A1(n14178), .A2(n6666), .ZN(n11354) );
  NAND2_X1 U13895 ( .A1(n11556), .A2(n14042), .ZN(n11353) );
  NAND2_X1 U13896 ( .A1(n11354), .A2(n11353), .ZN(n11355) );
  XNOR2_X1 U13897 ( .A(n11355), .B(n14043), .ZN(n11407) );
  NAND2_X1 U13898 ( .A1(n14178), .A2(n14045), .ZN(n11357) );
  NAND2_X1 U13899 ( .A1(n11556), .A2(n6666), .ZN(n11356) );
  NAND2_X1 U13900 ( .A1(n11357), .A2(n11356), .ZN(n11408) );
  XNOR2_X1 U13901 ( .A(n11407), .B(n11408), .ZN(n11358) );
  XNOR2_X1 U13902 ( .A(n11409), .B(n11358), .ZN(n11359) );
  NAND2_X1 U13903 ( .A1(n11359), .A2(n14142), .ZN(n11366) );
  OR2_X1 U13904 ( .A1(n14023), .A2(n14357), .ZN(n11361) );
  NAND2_X1 U13905 ( .A1(n14177), .A2(n14281), .ZN(n11360) );
  AND2_X1 U13906 ( .A1(n11361), .A2(n11360), .ZN(n11547) );
  AND2_X1 U13907 ( .A1(n15192), .A2(n11556), .ZN(n15172) );
  NAND2_X1 U13908 ( .A1(n14062), .A2(n15172), .ZN(n11363) );
  OAI211_X1 U13909 ( .C1(n11547), .C2(n14133), .A(n11363), .B(n11362), .ZN(
        n11364) );
  INV_X1 U13910 ( .A(n11364), .ZN(n11365) );
  OAI211_X1 U13911 ( .C1(n14161), .C2(n11554), .A(n11366), .B(n11365), .ZN(
        P1_U3227) );
  NAND2_X1 U13912 ( .A1(n11368), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11367) );
  OAI21_X1 U13913 ( .B1(n12916), .B2(n11368), .A(n11367), .ZN(P3_U3520) );
  NAND2_X1 U13914 ( .A1(n11375), .A2(n13359), .ZN(n11371) );
  XNOR2_X1 U13915 ( .A(n11502), .B(n11378), .ZN(n11382) );
  INV_X1 U13916 ( .A(n11382), .ZN(n15376) );
  NAND2_X1 U13917 ( .A1(n13359), .A2(n13307), .ZN(n11373) );
  NAND2_X1 U13918 ( .A1(n13357), .A2(n13336), .ZN(n11372) );
  NAND2_X1 U13919 ( .A1(n11373), .A2(n11372), .ZN(n11396) );
  INV_X1 U13920 ( .A(n13359), .ZN(n11392) );
  OR2_X1 U13921 ( .A1(n11375), .A2(n11392), .ZN(n11376) );
  NAND2_X1 U13922 ( .A1(n11377), .A2(n11376), .ZN(n11379) );
  NAND2_X1 U13923 ( .A1(n11379), .A2(n11501), .ZN(n11380) );
  AOI21_X1 U13924 ( .B1(n11506), .B2(n11380), .A(n13806), .ZN(n11381) );
  AOI211_X1 U13925 ( .C1(n11382), .C2(n13652), .A(n11396), .B(n11381), .ZN(
        n15375) );
  MUX2_X1 U13926 ( .A(n11383), .B(n15375), .S(n13741), .Z(n11388) );
  INV_X1 U13927 ( .A(n11384), .ZN(n11385) );
  AOI211_X1 U13928 ( .C1(n15372), .C2(n11385), .A(n13720), .B(n11512), .ZN(
        n15371) );
  OAI22_X1 U13929 ( .A1(n11504), .A2(n13743), .B1(n11399), .B2(n13737), .ZN(
        n11386) );
  AOI21_X1 U13930 ( .B1(n15371), .B2(n14931), .A(n11386), .ZN(n11387) );
  OAI211_X1 U13931 ( .C1(n15376), .C2(n11942), .A(n11388), .B(n11387), .ZN(
        P2_U3257) );
  INV_X1 U13932 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n11390) );
  INV_X1 U13933 ( .A(n12943), .ZN(n12901) );
  NAND2_X1 U13934 ( .A1(n12901), .A2(n11422), .ZN(n11389) );
  OAI21_X1 U13935 ( .B1(P3_U3897), .B2(n11390), .A(n11389), .ZN(P3_U3518) );
  INV_X1 U13936 ( .A(n11391), .ZN(n11395) );
  NOR3_X1 U13937 ( .A1(n11810), .A2(n11393), .A3(n11392), .ZN(n11394) );
  AOI21_X1 U13938 ( .B1(n11395), .B2(n14903), .A(n11394), .ZN(n11405) );
  NAND2_X1 U13939 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n13432) );
  INV_X1 U13940 ( .A(n11396), .ZN(n11397) );
  OR2_X1 U13941 ( .A1(n13339), .A2(n11397), .ZN(n11398) );
  OAI211_X1 U13942 ( .C1(n14911), .C2(n11399), .A(n13432), .B(n11398), .ZN(
        n11402) );
  NOR2_X1 U13943 ( .A1(n11400), .A2(n13342), .ZN(n11401) );
  AOI211_X1 U13944 ( .C1(n15372), .C2(n14908), .A(n11402), .B(n11401), .ZN(
        n11403) );
  OAI21_X1 U13945 ( .B1(n11405), .B2(n11404), .A(n11403), .ZN(P2_U3193) );
  INV_X1 U13946 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n15608) );
  NAND2_X1 U13947 ( .A1(n12907), .A2(n11422), .ZN(n11406) );
  OAI21_X1 U13948 ( .B1(P3_U3897), .B2(n15608), .A(n11406), .ZN(P3_U3521) );
  NAND2_X1 U13949 ( .A1(n14177), .A2(n6666), .ZN(n11411) );
  NAND2_X1 U13950 ( .A1(n11637), .A2(n14042), .ZN(n11410) );
  NAND2_X1 U13951 ( .A1(n11411), .A2(n11410), .ZN(n11412) );
  XNOR2_X1 U13952 ( .A(n11412), .B(n13985), .ZN(n11704) );
  NAND2_X1 U13953 ( .A1(n14177), .A2(n14045), .ZN(n11414) );
  NAND2_X1 U13954 ( .A1(n11637), .A2(n6666), .ZN(n11413) );
  NAND2_X1 U13955 ( .A1(n11414), .A2(n11413), .ZN(n11705) );
  XNOR2_X1 U13956 ( .A(n11704), .B(n11705), .ZN(n11702) );
  XNOR2_X1 U13957 ( .A(n11703), .B(n11702), .ZN(n11420) );
  NAND2_X1 U13958 ( .A1(n14178), .A2(n14521), .ZN(n11416) );
  NAND2_X1 U13959 ( .A1(n14176), .A2(n14281), .ZN(n11415) );
  AND2_X1 U13960 ( .A1(n11416), .A2(n11415), .ZN(n15181) );
  OAI22_X1 U13961 ( .A1(n14133), .A2(n15181), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9648), .ZN(n11418) );
  NOR2_X1 U13962 ( .A1(n14161), .A2(n11482), .ZN(n11417) );
  AOI211_X1 U13963 ( .C1(n14163), .C2(n11637), .A(n11418), .B(n11417), .ZN(
        n11419) );
  OAI21_X1 U13964 ( .B1(n11420), .B2(n14165), .A(n11419), .ZN(P1_U3239) );
  INV_X1 U13965 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n15879) );
  INV_X1 U13966 ( .A(n12930), .ZN(n12908) );
  NAND2_X1 U13967 ( .A1(n12908), .A2(n11422), .ZN(n11421) );
  OAI21_X1 U13968 ( .B1(n11422), .B2(n15879), .A(n11421), .ZN(P3_U3519) );
  MUX2_X1 U13969 ( .A(n12077), .B(n11440), .S(n12814), .Z(n11423) );
  INV_X1 U13970 ( .A(n11727), .ZN(n11446) );
  NAND2_X1 U13971 ( .A1(n11423), .A2(n11446), .ZN(n11718) );
  INV_X1 U13972 ( .A(n11423), .ZN(n11424) );
  NAND2_X1 U13973 ( .A1(n11424), .A2(n11727), .ZN(n11425) );
  NAND2_X1 U13974 ( .A1(n11718), .A2(n11425), .ZN(n11426) );
  AND3_X1 U13975 ( .A1(n11428), .A2(n11427), .A3(n11426), .ZN(n11429) );
  OAI21_X1 U13976 ( .B1(n11720), .B2(n11429), .A(n12853), .ZN(n11448) );
  NOR2_X1 U13977 ( .A1(n11438), .A2(n11430), .ZN(n11432) );
  MUX2_X1 U13978 ( .A(n12077), .B(P3_REG2_REG_10__SCAN_IN), .S(n11727), .Z(
        n11433) );
  NOR2_X1 U13979 ( .A1(n11434), .A2(n11433), .ZN(n11726) );
  AOI21_X1 U13980 ( .B1(n11434), .B2(n11433), .A(n11726), .ZN(n11436) );
  INV_X1 U13981 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15849) );
  NOR2_X1 U13982 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15849), .ZN(n12120) );
  AOI21_X1 U13983 ( .B1(n15392), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12120), 
        .ZN(n11435) );
  OAI21_X1 U13984 ( .B1(n12847), .B2(n11436), .A(n11435), .ZN(n11445) );
  MUX2_X1 U13985 ( .A(n11440), .B(P3_REG1_REG_10__SCAN_IN), .S(n11727), .Z(
        n11441) );
  NAND2_X1 U13986 ( .A1(n11442), .A2(n11441), .ZN(n11443) );
  AOI21_X1 U13987 ( .B1(n11715), .B2(n11443), .A(n12855), .ZN(n11444) );
  AOI211_X1 U13988 ( .C1(n12822), .C2(n11446), .A(n11445), .B(n11444), .ZN(
        n11447) );
  NAND2_X1 U13989 ( .A1(n11448), .A2(n11447), .ZN(P3_U3192) );
  INV_X1 U13990 ( .A(n11449), .ZN(n11451) );
  AND2_X1 U13991 ( .A1(n11451), .A2(n11450), .ZN(n12304) );
  NAND2_X1 U13992 ( .A1(n12304), .A2(n11452), .ZN(n14353) );
  INV_X2 U13993 ( .A(n14532), .ZN(n15108) );
  NOR2_X1 U13994 ( .A1(n15108), .A2(n15089), .ZN(n14516) );
  NOR2_X1 U13995 ( .A1(n14516), .A2(n14967), .ZN(n11463) );
  OAI22_X1 U13996 ( .A1(n15108), .A2(n11457), .B1(n11456), .B2(n15094), .ZN(
        n11461) );
  INV_X1 U13997 ( .A(n14353), .ZN(n11458) );
  NAND2_X1 U13998 ( .A1(n11458), .A2(n14511), .ZN(n14496) );
  OR2_X1 U13999 ( .A1(n14496), .A2(n15205), .ZN(n14350) );
  AOI21_X1 U14000 ( .B1(n14350), .B2(n15098), .A(n11480), .ZN(n11460) );
  AOI211_X1 U14001 ( .C1(n15108), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11461), .B(
        n11460), .ZN(n11462) );
  OAI21_X1 U14002 ( .B1(n11464), .B2(n11463), .A(n11462), .ZN(P1_U3293) );
  AOI22_X1 U14003 ( .A1(n14919), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14918), .ZN(n11465) );
  OAI21_X1 U14004 ( .B1(n13743), .B2(n11466), .A(n11465), .ZN(n11469) );
  NOR2_X1 U14005 ( .A1(n11467), .A2(n13751), .ZN(n11468) );
  AOI211_X1 U14006 ( .C1(n11470), .C2(n14931), .A(n11469), .B(n11468), .ZN(
        n11471) );
  OAI21_X1 U14007 ( .B1(n14919), .B2(n11472), .A(n11471), .ZN(P2_U3263) );
  AND2_X1 U14008 ( .A1(n14182), .A2(n11486), .ZN(n11657) );
  OR2_X1 U14009 ( .A1(n7010), .A2(n14181), .ZN(n11474) );
  NAND2_X1 U14010 ( .A1(n15086), .A2(n15088), .ZN(n11476) );
  OR2_X1 U14011 ( .A1(n14026), .A2(n14179), .ZN(n11475) );
  NAND2_X1 U14012 ( .A1(n11476), .A2(n11475), .ZN(n11533) );
  NAND2_X1 U14013 ( .A1(n14023), .A2(n15167), .ZN(n11477) );
  OR2_X1 U14014 ( .A1(n14178), .A2(n11556), .ZN(n11478) );
  INV_X1 U14015 ( .A(n11479), .ZN(n11635) );
  XNOR2_X1 U14016 ( .A(n11636), .B(n11635), .ZN(n15184) );
  INV_X1 U14017 ( .A(n15184), .ZN(n15186) );
  AND2_X1 U14018 ( .A1(n11669), .A2(n11480), .ZN(n11525) );
  NAND2_X1 U14019 ( .A1(n11525), .A2(n11524), .ZN(n15100) );
  OAI211_X1 U14020 ( .C1(n7285), .C2(n7284), .A(n15143), .B(n15082), .ZN(
        n15182) );
  INV_X1 U14021 ( .A(n15182), .ZN(n11485) );
  INV_X1 U14022 ( .A(n14496), .ZN(n15104) );
  INV_X1 U14023 ( .A(n15181), .ZN(n11481) );
  MUX2_X1 U14024 ( .A(n11481), .B(P1_REG2_REG_6__SCAN_IN), .S(n15108), .Z(
        n11484) );
  OAI22_X1 U14025 ( .A1(n15098), .A2(n7284), .B1(n11482), .B2(n15094), .ZN(
        n11483) );
  AOI211_X1 U14026 ( .C1(n11485), .C2(n15104), .A(n11484), .B(n11483), .ZN(
        n11500) );
  NAND2_X1 U14027 ( .A1(n11661), .A2(n15144), .ZN(n11660) );
  NAND2_X1 U14028 ( .A1(n11660), .A2(n11487), .ZN(n11490) );
  NAND2_X1 U14029 ( .A1(n11488), .A2(n15142), .ZN(n11489) );
  NAND2_X1 U14030 ( .A1(n11490), .A2(n11489), .ZN(n11530) );
  NAND2_X1 U14031 ( .A1(n11530), .A2(n11529), .ZN(n11492) );
  NAND2_X1 U14032 ( .A1(n11492), .A2(n11491), .ZN(n15087) );
  NAND2_X1 U14033 ( .A1(n15087), .A2(n11493), .ZN(n11495) );
  INV_X1 U14034 ( .A(n11496), .ZN(n11538) );
  NAND2_X1 U14035 ( .A1(n14023), .A2(n6901), .ZN(n11497) );
  INV_X1 U14036 ( .A(n11556), .ZN(n11552) );
  NOR2_X1 U14037 ( .A1(n14178), .A2(n11552), .ZN(n11498) );
  XNOR2_X1 U14038 ( .A(n11628), .B(n11635), .ZN(n15190) );
  NAND2_X1 U14039 ( .A1(n15190), .A2(n14516), .ZN(n11499) );
  OAI211_X1 U14040 ( .C1(n15186), .C2(n14564), .A(n11500), .B(n11499), .ZN(
        P1_U3287) );
  XNOR2_X1 U14041 ( .A(n11676), .B(n11675), .ZN(n11648) );
  INV_X1 U14042 ( .A(n11675), .ZN(n11508) );
  OAI21_X1 U14043 ( .B1(n11508), .B2(n11507), .A(n11681), .ZN(n11510) );
  AOI21_X1 U14044 ( .B1(n11510), .B2(n14915), .A(n11509), .ZN(n11511) );
  OAI21_X1 U14045 ( .B1(n11933), .B2(n11648), .A(n11511), .ZN(n11649) );
  NAND2_X1 U14046 ( .A1(n11649), .A2(n13741), .ZN(n11519) );
  INV_X1 U14047 ( .A(n11512), .ZN(n11513) );
  NAND2_X1 U14048 ( .A1(n11512), .A2(n11653), .ZN(n11688) );
  INV_X1 U14049 ( .A(n11688), .ZN(n11689) );
  AOI211_X1 U14050 ( .C1(n11677), .C2(n11513), .A(n13720), .B(n11689), .ZN(
        n11650) );
  NOR2_X1 U14051 ( .A1(n11653), .A2(n13743), .ZN(n11517) );
  OAI22_X1 U14052 ( .A1(n13741), .A2(n11515), .B1(n11514), .B2(n13737), .ZN(
        n11516) );
  AOI211_X1 U14053 ( .C1(n11650), .C2(n14931), .A(n11517), .B(n11516), .ZN(
        n11518) );
  OAI211_X1 U14054 ( .C1(n11648), .C2(n11942), .A(n11519), .B(n11518), .ZN(
        P2_U3256) );
  INV_X1 U14055 ( .A(n11520), .ZN(n15324) );
  OAI222_X1 U14056 ( .A1(P2_U3088), .A2(n15324), .B1(n13892), .B2(n11523), 
        .C1(n11521), .C2(n13894), .ZN(P2_U3309) );
  OAI222_X1 U14057 ( .A1(P1_U3086), .A2(n14257), .B1(n14694), .B2(n11523), 
        .C1(n11522), .C2(n14691), .ZN(P1_U3337) );
  OAI211_X1 U14058 ( .C1(n11525), .C2(n11524), .A(n15143), .B(n15100), .ZN(
        n15151) );
  OAI22_X1 U14059 ( .A1(n14496), .A2(n15151), .B1(n11526), .B2(n15094), .ZN(
        n11528) );
  MUX2_X1 U14060 ( .A(n15150), .B(P1_REG2_REG_2__SCAN_IN), .S(n15108), .Z(
        n11527) );
  AOI211_X1 U14061 ( .C1(n14958), .C2(n7010), .A(n11528), .B(n11527), .ZN(
        n11532) );
  XNOR2_X1 U14062 ( .A(n11529), .B(n11530), .ZN(n15156) );
  NAND2_X1 U14063 ( .A1(n14516), .A2(n15156), .ZN(n11531) );
  OAI211_X1 U14064 ( .C1(n14564), .C2(n15153), .A(n11532), .B(n11531), .ZN(
        P1_U3291) );
  XNOR2_X1 U14065 ( .A(n11533), .B(n11538), .ZN(n15168) );
  OAI211_X1 U14066 ( .C1(n15101), .C2(n15167), .A(n11550), .B(n15143), .ZN(
        n15166) );
  OAI22_X1 U14067 ( .A1(n14496), .A2(n15166), .B1(n11534), .B2(n15094), .ZN(
        n11537) );
  INV_X1 U14068 ( .A(n15165), .ZN(n11535) );
  MUX2_X1 U14069 ( .A(n11535), .B(P1_REG2_REG_4__SCAN_IN), .S(n15108), .Z(
        n11536) );
  AOI211_X1 U14070 ( .C1(n14958), .C2(n6901), .A(n11537), .B(n11536), .ZN(
        n11541) );
  XNOR2_X1 U14071 ( .A(n11539), .B(n11538), .ZN(n15171) );
  NAND2_X1 U14072 ( .A1(n15171), .A2(n14516), .ZN(n11540) );
  OAI211_X1 U14073 ( .C1(n15168), .C2(n14564), .A(n11541), .B(n11540), .ZN(
        P1_U3289) );
  XNOR2_X1 U14074 ( .A(n11543), .B(n11542), .ZN(n15177) );
  XNOR2_X1 U14075 ( .A(n11545), .B(n11544), .ZN(n11546) );
  NOR2_X1 U14076 ( .A1(n11546), .A2(n15089), .ZN(n15178) );
  INV_X1 U14077 ( .A(n11547), .ZN(n15173) );
  NOR2_X1 U14078 ( .A1(n15178), .A2(n15173), .ZN(n11548) );
  MUX2_X1 U14079 ( .A(n11549), .B(n11548), .S(n14532), .Z(n11558) );
  INV_X1 U14080 ( .A(n11550), .ZN(n11553) );
  OAI211_X1 U14081 ( .C1(n11553), .C2(n11552), .A(n15143), .B(n11551), .ZN(
        n15174) );
  OAI22_X1 U14082 ( .A1(n15174), .A2(n14496), .B1(n11554), .B2(n15094), .ZN(
        n11555) );
  AOI21_X1 U14083 ( .B1(n14958), .B2(n11556), .A(n11555), .ZN(n11557) );
  OAI211_X1 U14084 ( .C1(n14564), .C2(n15177), .A(n11558), .B(n11557), .ZN(
        P1_U3288) );
  INV_X1 U14085 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U14086 ( .A1(n12859), .A2(n11422), .ZN(n11559) );
  OAI21_X1 U14087 ( .B1(P3_U3897), .B2(n11560), .A(n11559), .ZN(P3_U3522) );
  NAND2_X1 U14088 ( .A1(n11562), .A2(n11561), .ZN(n11564) );
  OAI211_X1 U14089 ( .C1(n15662), .C2(n12166), .A(n11564), .B(n11563), .ZN(
        P3_U3272) );
  NOR2_X1 U14090 ( .A1(n15438), .A2(n11565), .ZN(n15439) );
  NAND2_X1 U14091 ( .A1(n15463), .A2(n15439), .ZN(n12992) );
  INV_X1 U14092 ( .A(n12992), .ZN(n12978) );
  OR2_X1 U14093 ( .A1(n11566), .A2(n7759), .ZN(n11567) );
  NAND2_X1 U14094 ( .A1(n11568), .A2(n11567), .ZN(n15482) );
  NAND2_X1 U14095 ( .A1(n11597), .A2(n15495), .ZN(n15479) );
  OAI22_X1 U14096 ( .A1(n11774), .A2(n15479), .B1(n11569), .B2(n15458), .ZN(
        n11592) );
  NAND2_X1 U14097 ( .A1(n15427), .A2(n15428), .ZN(n11572) );
  NAND2_X1 U14098 ( .A1(n15451), .A2(n15437), .ZN(n15410) );
  NAND2_X1 U14099 ( .A1(n11575), .A2(n11574), .ZN(n11576) );
  XNOR2_X1 U14100 ( .A(n11596), .B(n11595), .ZN(n11590) );
  NAND2_X1 U14101 ( .A1(n11577), .A2(n13115), .ZN(n11579) );
  OAI22_X1 U14102 ( .A1(n11795), .A2(n15450), .B1(n15424), .B2(n15425), .ZN(
        n11582) );
  INV_X1 U14103 ( .A(n11582), .ZN(n11589) );
  INV_X1 U14104 ( .A(n11583), .ZN(n11584) );
  NAND3_X1 U14105 ( .A1(n11585), .A2(n11584), .A3(n15512), .ZN(n11587) );
  NAND2_X1 U14106 ( .A1(n15482), .A2(n15435), .ZN(n11588) );
  OAI211_X1 U14107 ( .C1(n11590), .C2(n15430), .A(n11589), .B(n11588), .ZN(
        n15480) );
  MUX2_X1 U14108 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15480), .S(n15463), .Z(
        n11591) );
  AOI211_X1 U14109 ( .C1(n12978), .C2(n15482), .A(n11592), .B(n11591), .ZN(
        n11593) );
  INV_X1 U14110 ( .A(n11593), .ZN(P3_U3229) );
  XNOR2_X1 U14111 ( .A(n11594), .B(n11600), .ZN(n15485) );
  INV_X1 U14112 ( .A(n15485), .ZN(n11611) );
  NAND2_X1 U14113 ( .A1(n15485), .A2(n15435), .ZN(n11606) );
  NAND2_X1 U14114 ( .A1(n11598), .A2(n11597), .ZN(n11599) );
  NAND2_X1 U14115 ( .A1(n11601), .A2(n11600), .ZN(n11602) );
  NAND2_X1 U14116 ( .A1(n11777), .A2(n11602), .ZN(n11604) );
  OAI22_X1 U14117 ( .A1(n15408), .A2(n15425), .B1(n12613), .B2(n15450), .ZN(
        n11603) );
  AOI21_X1 U14118 ( .B1(n11604), .B2(n15453), .A(n11603), .ZN(n11605) );
  AND2_X1 U14119 ( .A1(n11606), .A2(n11605), .ZN(n15487) );
  MUX2_X1 U14120 ( .A(n11607), .B(n15487), .S(n15463), .Z(n11610) );
  AND2_X1 U14121 ( .A1(n12612), .A2(n15495), .ZN(n15484) );
  INV_X1 U14122 ( .A(n11608), .ZN(n12615) );
  AOI22_X1 U14123 ( .A1(n15419), .A2(n15484), .B1(n15442), .B2(n12615), .ZN(
        n11609) );
  OAI211_X1 U14124 ( .C1(n11611), .C2(n12992), .A(n11610), .B(n11609), .ZN(
        P3_U3228) );
  XNOR2_X1 U14125 ( .A(n11612), .B(n11616), .ZN(n15497) );
  NAND2_X1 U14126 ( .A1(n15497), .A2(n15435), .ZN(n11620) );
  NAND2_X1 U14127 ( .A1(n11795), .A2(n11613), .ZN(n11776) );
  AND2_X1 U14128 ( .A1(n11775), .A2(n11776), .ZN(n11614) );
  NAND2_X1 U14129 ( .A1(n12104), .A2(n11791), .ZN(n11615) );
  XNOR2_X1 U14130 ( .A(n12071), .B(n11616), .ZN(n11618) );
  OAI22_X1 U14131 ( .A1(n12497), .A2(n15450), .B1(n12613), .B2(n15425), .ZN(
        n11617) );
  AOI21_X1 U14132 ( .B1(n11618), .B2(n15453), .A(n11617), .ZN(n11619) );
  AND2_X1 U14133 ( .A1(n11620), .A2(n11619), .ZN(n15499) );
  INV_X2 U14134 ( .A(n15463), .ZN(n15465) );
  NOR2_X1 U14135 ( .A1(n13104), .A2(n11621), .ZN(n11623) );
  OAI22_X1 U14136 ( .A1(n15463), .A2(n10951), .B1(n12499), .B2(n15458), .ZN(
        n11622) );
  AOI211_X1 U14137 ( .C1(n15497), .C2(n12978), .A(n11623), .B(n11622), .ZN(
        n11624) );
  OAI21_X1 U14138 ( .B1(n15499), .B2(n15465), .A(n11624), .ZN(P3_U3226) );
  AND2_X1 U14139 ( .A1(n7284), .A2(n14177), .ZN(n11627) );
  INV_X1 U14140 ( .A(n14177), .ZN(n11625) );
  NAND2_X1 U14141 ( .A1(n11625), .A2(n11637), .ZN(n11626) );
  INV_X1 U14142 ( .A(n14176), .ZN(n11629) );
  AND2_X1 U14143 ( .A1(n15193), .A2(n11629), .ZN(n11630) );
  OAI22_X1 U14144 ( .A1(n15070), .A2(n11630), .B1(n11629), .B2(n15193), .ZN(
        n11733) );
  XNOR2_X1 U14145 ( .A(n11733), .B(n6667), .ZN(n11634) );
  NAND2_X1 U14146 ( .A1(n14176), .A2(n14521), .ZN(n11632) );
  NAND2_X1 U14147 ( .A1(n14174), .A2(n14281), .ZN(n11631) );
  NAND2_X1 U14148 ( .A1(n11632), .A2(n11631), .ZN(n11891) );
  INV_X1 U14149 ( .A(n11891), .ZN(n11633) );
  OAI21_X1 U14150 ( .B1(n11634), .B2(n15089), .A(n11633), .ZN(n15202) );
  INV_X1 U14151 ( .A(n15202), .ZN(n11647) );
  NAND2_X1 U14152 ( .A1(n11636), .A2(n11635), .ZN(n11639) );
  OR2_X1 U14153 ( .A1(n14177), .A2(n11637), .ZN(n11638) );
  INV_X1 U14154 ( .A(n15071), .ZN(n11640) );
  OR2_X1 U14155 ( .A1(n15193), .A2(n14176), .ZN(n11641) );
  XNOR2_X1 U14156 ( .A(n11745), .B(n11744), .ZN(n15204) );
  INV_X1 U14157 ( .A(n11879), .ZN(n15201) );
  OAI211_X1 U14158 ( .C1(n15081), .C2(n15201), .A(n11827), .B(n15143), .ZN(
        n15200) );
  INV_X1 U14159 ( .A(n11642), .ZN(n11894) );
  INV_X1 U14160 ( .A(n15094), .ZN(n14956) );
  AOI22_X1 U14161 ( .A1(n15108), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n11894), 
        .B2(n14956), .ZN(n11644) );
  NAND2_X1 U14162 ( .A1(n14958), .A2(n11879), .ZN(n11643) );
  OAI211_X1 U14163 ( .C1(n15200), .C2(n14496), .A(n11644), .B(n11643), .ZN(
        n11645) );
  AOI21_X1 U14164 ( .B1(n15204), .B2(n14967), .A(n11645), .ZN(n11646) );
  OAI21_X1 U14165 ( .B1(n11647), .B2(n15096), .A(n11646), .ZN(P1_U3285) );
  INV_X1 U14166 ( .A(n11648), .ZN(n11651) );
  AOI211_X1 U14167 ( .C1(n11651), .C2(n9510), .A(n11650), .B(n11649), .ZN(
        n11656) );
  AOI22_X1 U14168 ( .A1(n11677), .A2(n13837), .B1(n15389), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11652) );
  OAI21_X1 U14169 ( .B1(n11656), .B2(n15389), .A(n11652), .ZN(P2_U3508) );
  INV_X1 U14170 ( .A(n13873), .ZN(n13864) );
  OAI22_X1 U14171 ( .A1(n11653), .A2(n13864), .B1(n15387), .B2(n8103), .ZN(
        n11654) );
  INV_X1 U14172 ( .A(n11654), .ZN(n11655) );
  OAI21_X1 U14173 ( .B1(n11656), .B2(n15386), .A(n11655), .ZN(P2_U3457) );
  XOR2_X1 U14174 ( .A(n11657), .B(n11658), .Z(n15147) );
  OAI22_X1 U14175 ( .A1(n15147), .A2(n15187), .B1(n7011), .B2(n14156), .ZN(
        n11666) );
  INV_X1 U14176 ( .A(n11658), .ZN(n11659) );
  OAI21_X1 U14177 ( .B1(n11659), .B2(n11662), .A(n15189), .ZN(n11664) );
  OAI211_X1 U14178 ( .C1(n11661), .C2(n15144), .A(n11660), .B(n15189), .ZN(
        n11663) );
  AOI22_X1 U14179 ( .A1(n11664), .A2(n14357), .B1(n11663), .B2(n11662), .ZN(
        n11665) );
  NOR2_X1 U14180 ( .A1(n11666), .A2(n11665), .ZN(n15146) );
  INV_X1 U14181 ( .A(n14350), .ZN(n14550) );
  OAI22_X1 U14182 ( .A1(n14532), .A2(n10285), .B1(n11667), .B2(n15094), .ZN(
        n11671) );
  NOR2_X1 U14183 ( .A1(n15096), .A2(n11668), .ZN(n15105) );
  INV_X1 U14184 ( .A(n15105), .ZN(n12101) );
  OAI22_X1 U14185 ( .A1(n12101), .A2(n15147), .B1(n11669), .B2(n15098), .ZN(
        n11670) );
  AOI211_X1 U14186 ( .C1(n14550), .C2(n15144), .A(n11671), .B(n11670), .ZN(
        n11672) );
  OAI21_X1 U14187 ( .B1(n15108), .B2(n15146), .A(n11672), .ZN(P1_U3292) );
  OAI222_X1 U14188 ( .A1(P1_U3086), .A2(n11674), .B1(n14694), .B2(n11694), 
        .C1(n11673), .C2(n14691), .ZN(P1_U3335) );
  NAND2_X1 U14189 ( .A1(n11676), .A2(n11675), .ZN(n11679) );
  NAND2_X1 U14190 ( .A1(n11677), .A2(n13357), .ZN(n11678) );
  NAND2_X1 U14191 ( .A1(n11679), .A2(n11678), .ZN(n11757) );
  XNOR2_X1 U14192 ( .A(n11757), .B(n11756), .ZN(n15379) );
  OAI21_X1 U14193 ( .B1(n11683), .B2(n11682), .A(n11763), .ZN(n11685) );
  OAI22_X1 U14194 ( .A1(n11926), .A2(n13326), .B1(n11684), .B2(n13544), .ZN(
        n11851) );
  AOI21_X1 U14195 ( .B1(n11685), .B2(n14915), .A(n11851), .ZN(n11686) );
  OAI21_X1 U14196 ( .B1(n11933), .B2(n15379), .A(n11686), .ZN(n15383) );
  NAND2_X1 U14197 ( .A1(n15383), .A2(n13741), .ZN(n11693) );
  OAI22_X1 U14198 ( .A1(n13741), .A2(n11687), .B1(n11854), .B2(n13737), .ZN(
        n11691) );
  OAI211_X1 U14199 ( .C1(n11689), .C2(n15382), .A(n14928), .B(n11766), .ZN(
        n15380) );
  NOR2_X1 U14200 ( .A1(n15380), .A2(n13713), .ZN(n11690) );
  AOI211_X1 U14201 ( .C1(n14920), .C2(n11860), .A(n11691), .B(n11690), .ZN(
        n11692) );
  OAI211_X1 U14202 ( .C1(n15379), .C2(n11942), .A(n11693), .B(n11692), .ZN(
        P2_U3255) );
  OAI222_X1 U14203 ( .A1(n13894), .A2(n11696), .B1(P2_U3088), .B2(n11695), 
        .C1(n13883), .C2(n11694), .ZN(P2_U3307) );
  INV_X1 U14204 ( .A(n11697), .ZN(n12466) );
  OAI222_X1 U14205 ( .A1(n14511), .A2(P1_U3086), .B1(n14694), .B2(n12466), 
        .C1(n11698), .C2(n14691), .ZN(P1_U3336) );
  NAND2_X1 U14206 ( .A1(n15193), .A2(n14042), .ZN(n11700) );
  NAND2_X1 U14207 ( .A1(n14176), .A2(n6666), .ZN(n11699) );
  NAND2_X1 U14208 ( .A1(n11700), .A2(n11699), .ZN(n11701) );
  XNOR2_X1 U14209 ( .A(n11701), .B(n14043), .ZN(n11882) );
  AOI22_X1 U14210 ( .A1(n15193), .A2(n6666), .B1(n14045), .B2(n14176), .ZN(
        n11883) );
  XNOR2_X1 U14211 ( .A(n11882), .B(n11883), .ZN(n11880) );
  INV_X1 U14212 ( .A(n11704), .ZN(n11706) );
  XOR2_X1 U14213 ( .A(n11881), .B(n11880), .Z(n11707) );
  NAND2_X1 U14214 ( .A1(n11707), .A2(n14142), .ZN(n11713) );
  NAND2_X1 U14215 ( .A1(n14177), .A2(n14521), .ZN(n11709) );
  NAND2_X1 U14216 ( .A1(n14175), .A2(n14281), .ZN(n11708) );
  AND2_X1 U14217 ( .A1(n11709), .A2(n11708), .ZN(n15073) );
  OAI21_X1 U14218 ( .B1(n14133), .B2(n15073), .A(n11710), .ZN(n11711) );
  AOI21_X1 U14219 ( .B1(n14163), .B2(n15193), .A(n11711), .ZN(n11712) );
  OAI211_X1 U14220 ( .C1(n14161), .C2(n15076), .A(n11713), .B(n11712), .ZN(
        P1_U3213) );
  NAND2_X1 U14221 ( .A1(n11727), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11714) );
  AOI21_X1 U14222 ( .B1(n8828), .B2(n11716), .A(n11944), .ZN(n11732) );
  INV_X1 U14223 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14724) );
  INV_X1 U14224 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15797) );
  NOR2_X1 U14225 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15797), .ZN(n12348) );
  INV_X1 U14226 ( .A(n12348), .ZN(n11717) );
  OAI21_X1 U14227 ( .B1(n12813), .B2(n14724), .A(n11717), .ZN(n11725) );
  INV_X1 U14228 ( .A(n11718), .ZN(n11719) );
  MUX2_X1 U14229 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12814), .Z(n11958) );
  XNOR2_X1 U14230 ( .A(n11958), .B(n11957), .ZN(n11721) );
  AOI21_X1 U14231 ( .B1(n11722), .B2(n11721), .A(n11960), .ZN(n11723) );
  NOR2_X1 U14232 ( .A1(n11723), .A2(n12819), .ZN(n11724) );
  AOI211_X1 U14233 ( .C1(n12822), .C2(n11951), .A(n11725), .B(n11724), .ZN(
        n11731) );
  XNOR2_X1 U14234 ( .A(n11951), .B(n11950), .ZN(n11728) );
  AOI21_X1 U14235 ( .B1(n12336), .B2(n11728), .A(n11952), .ZN(n11729) );
  OR2_X1 U14236 ( .A1(n11729), .A2(n12847), .ZN(n11730) );
  OAI211_X1 U14237 ( .C1(n11732), .C2(n12855), .A(n11731), .B(n11730), .ZN(
        P3_U3193) );
  NAND2_X1 U14238 ( .A1(n11733), .A2(n6667), .ZN(n11736) );
  OR2_X1 U14239 ( .A1(n11879), .A2(n11734), .ZN(n11735) );
  INV_X1 U14240 ( .A(n14174), .ZN(n11741) );
  NAND2_X1 U14241 ( .A1(n11912), .A2(n11741), .ZN(n11740) );
  AND2_X1 U14242 ( .A1(n11747), .A2(n11740), .ZN(n11738) );
  NAND2_X1 U14243 ( .A1(n11835), .A2(n15189), .ZN(n11743) );
  AOI21_X1 U14244 ( .B1(n11739), .B2(n11740), .A(n11747), .ZN(n11742) );
  OAI22_X1 U14245 ( .A1(n11743), .A2(n11742), .B1(n11741), .B2(n14357), .ZN(
        n15215) );
  INV_X1 U14246 ( .A(n15215), .ZN(n11755) );
  OR2_X1 U14247 ( .A1(n11912), .A2(n14174), .ZN(n11746) );
  INV_X1 U14248 ( .A(n11747), .ZN(n11839) );
  XNOR2_X1 U14249 ( .A(n11840), .B(n11839), .ZN(n15217) );
  INV_X1 U14250 ( .A(n11978), .ZN(n15214) );
  XNOR2_X1 U14251 ( .A(n11843), .B(n15214), .ZN(n11749) );
  AND2_X1 U14252 ( .A1(n14172), .A2(n14281), .ZN(n11748) );
  AOI21_X1 U14253 ( .B1(n11749), .B2(n15143), .A(n11748), .ZN(n15212) );
  INV_X1 U14254 ( .A(n11750), .ZN(n11985) );
  AOI22_X1 U14255 ( .A1(n15108), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11985), 
        .B2(n14956), .ZN(n11752) );
  NAND2_X1 U14256 ( .A1(n14958), .A2(n11978), .ZN(n11751) );
  OAI211_X1 U14257 ( .C1(n15212), .C2(n14496), .A(n11752), .B(n11751), .ZN(
        n11753) );
  AOI21_X1 U14258 ( .B1(n15217), .B2(n14967), .A(n11753), .ZN(n11754) );
  OAI21_X1 U14259 ( .B1(n11755), .B2(n15096), .A(n11754), .ZN(P1_U3283) );
  OR2_X1 U14260 ( .A1(n15382), .A2(n13354), .ZN(n11758) );
  XNOR2_X1 U14261 ( .A(n11925), .B(n11761), .ZN(n12063) );
  OR2_X1 U14262 ( .A1(n13354), .A2(n13544), .ZN(n11760) );
  OR2_X1 U14263 ( .A1(n11996), .A2(n13326), .ZN(n11759) );
  NAND2_X1 U14264 ( .A1(n11760), .A2(n11759), .ZN(n11805) );
  NAND3_X1 U14265 ( .A1(n11763), .A2(n7341), .A3(n11762), .ZN(n11764) );
  AOI21_X1 U14266 ( .B1(n11928), .B2(n11764), .A(n13806), .ZN(n11765) );
  AOI211_X1 U14267 ( .C1(n13652), .C2(n12063), .A(n11805), .B(n11765), .ZN(
        n12060) );
  AOI211_X1 U14268 ( .C1(n12064), .C2(n11766), .A(n13720), .B(n11937), .ZN(
        n12062) );
  NOR2_X1 U14269 ( .A1(n12066), .A2(n13743), .ZN(n11769) );
  OAI22_X1 U14270 ( .A1(n13741), .A2(n11767), .B1(n11808), .B2(n13737), .ZN(
        n11768) );
  AOI211_X1 U14271 ( .C1(n12062), .C2(n14931), .A(n11769), .B(n11768), .ZN(
        n11771) );
  NAND2_X1 U14272 ( .A1(n12063), .A2(n13661), .ZN(n11770) );
  OAI211_X1 U14273 ( .C1(n12060), .C2(n14919), .A(n11771), .B(n11770), .ZN(
        P2_U3254) );
  XNOR2_X1 U14274 ( .A(n11773), .B(n11772), .ZN(n15490) );
  NAND2_X1 U14275 ( .A1(n11791), .A2(n15495), .ZN(n15489) );
  OAI22_X1 U14276 ( .A1(n11774), .A2(n15489), .B1(n11787), .B2(n15458), .ZN(
        n11785) );
  AOI21_X1 U14277 ( .B1(n11777), .B2(n11776), .A(n11775), .ZN(n11783) );
  NAND2_X1 U14278 ( .A1(n11778), .A2(n15453), .ZN(n11782) );
  NAND2_X1 U14279 ( .A1(n15490), .A2(n15435), .ZN(n11781) );
  OAI22_X1 U14280 ( .A1(n12107), .A2(n15450), .B1(n11795), .B2(n15425), .ZN(
        n11779) );
  INV_X1 U14281 ( .A(n11779), .ZN(n11780) );
  OAI211_X1 U14282 ( .C1(n11783), .C2(n11782), .A(n11781), .B(n11780), .ZN(
        n15493) );
  MUX2_X1 U14283 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n15493), .S(n15463), .Z(
        n11784) );
  AOI211_X1 U14284 ( .C1(n15490), .C2(n12978), .A(n11785), .B(n11784), .ZN(
        n11786) );
  INV_X1 U14285 ( .A(n11786), .ZN(P3_U3227) );
  INV_X1 U14286 ( .A(n11787), .ZN(n11803) );
  OR2_X1 U14287 ( .A1(n12107), .A2(n12668), .ZN(n11790) );
  AOI21_X1 U14288 ( .B1(n12670), .B2(n11791), .A(n11788), .ZN(n11789) );
  OAI211_X1 U14289 ( .C1(n11795), .C2(n12677), .A(n11790), .B(n11789), .ZN(
        n11802) );
  XNOR2_X1 U14290 ( .A(n12613), .B(n12102), .ZN(n11800) );
  NAND2_X1 U14291 ( .A1(n11793), .A2(n11792), .ZN(n12608) );
  XNOR2_X1 U14292 ( .A(n12612), .B(n12532), .ZN(n11794) );
  XNOR2_X1 U14293 ( .A(n11794), .B(n11795), .ZN(n12609) );
  INV_X1 U14294 ( .A(n11794), .ZN(n11796) );
  NAND2_X1 U14295 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  INV_X1 U14296 ( .A(n12106), .ZN(n11798) );
  AOI211_X1 U14297 ( .C1(n11800), .C2(n11799), .A(n12672), .B(n11798), .ZN(
        n11801) );
  AOI211_X1 U14298 ( .C1(n11803), .C2(n12666), .A(n11802), .B(n11801), .ZN(
        n11804) );
  INV_X1 U14299 ( .A(n11804), .ZN(P3_U3179) );
  NAND2_X1 U14300 ( .A1(n14905), .A2(n11805), .ZN(n11807) );
  OAI211_X1 U14301 ( .C1(n14911), .C2(n11808), .A(n11807), .B(n11806), .ZN(
        n11816) );
  INV_X1 U14302 ( .A(n11809), .ZN(n11855) );
  NOR3_X1 U14303 ( .A1(n11811), .A2(n13354), .A3(n11810), .ZN(n11812) );
  AOI21_X1 U14304 ( .B1(n11855), .B2(n14903), .A(n11812), .ZN(n11814) );
  NOR2_X1 U14305 ( .A1(n11814), .A2(n11813), .ZN(n11815) );
  AOI211_X1 U14306 ( .C1(n12064), .C2(n14908), .A(n11816), .B(n11815), .ZN(
        n11817) );
  OAI21_X1 U14307 ( .B1(n11866), .B2(n13342), .A(n11817), .ZN(P2_U3208) );
  XNOR2_X1 U14308 ( .A(n11818), .B(n11821), .ZN(n15209) );
  INV_X1 U14309 ( .A(n15209), .ZN(n11833) );
  INV_X1 U14310 ( .A(n11739), .ZN(n11819) );
  AOI21_X1 U14311 ( .B1(n11821), .B2(n11820), .A(n11819), .ZN(n11825) );
  INV_X1 U14312 ( .A(n15187), .ZN(n15093) );
  NAND2_X1 U14313 ( .A1(n14175), .A2(n14521), .ZN(n11823) );
  NAND2_X1 U14314 ( .A1(n14173), .A2(n14281), .ZN(n11822) );
  NAND2_X1 U14315 ( .A1(n11823), .A2(n11822), .ZN(n11921) );
  AOI21_X1 U14316 ( .B1(n15209), .B2(n15093), .A(n11921), .ZN(n11824) );
  OAI21_X1 U14317 ( .B1(n11825), .B2(n15089), .A(n11824), .ZN(n15207) );
  NAND2_X1 U14318 ( .A1(n15207), .A2(n14532), .ZN(n11832) );
  OAI22_X1 U14319 ( .A1(n14532), .A2(n11826), .B1(n11918), .B2(n15094), .ZN(
        n11830) );
  NAND2_X1 U14320 ( .A1(n11827), .A2(n11912), .ZN(n11828) );
  NAND2_X1 U14321 ( .A1(n11843), .A2(n11828), .ZN(n15206) );
  NOR2_X1 U14322 ( .A1(n15206), .A2(n14350), .ZN(n11829) );
  AOI211_X1 U14323 ( .C1(n14958), .C2(n11912), .A(n11830), .B(n11829), .ZN(
        n11831) );
  OAI211_X1 U14324 ( .C1(n11833), .C2(n12101), .A(n11832), .B(n11831), .ZN(
        P1_U3284) );
  INV_X1 U14325 ( .A(n12036), .ZN(n12048) );
  XNOR2_X1 U14326 ( .A(n12037), .B(n12048), .ZN(n11838) );
  NAND2_X1 U14327 ( .A1(n14173), .A2(n14521), .ZN(n11837) );
  NAND2_X1 U14328 ( .A1(n14171), .A2(n14281), .ZN(n11836) );
  NAND2_X1 U14329 ( .A1(n11837), .A2(n11836), .ZN(n12225) );
  AOI21_X1 U14330 ( .B1(n11838), .B2(n15189), .A(n12225), .ZN(n14988) );
  NAND2_X1 U14331 ( .A1(n11840), .A2(n11839), .ZN(n11842) );
  OR2_X1 U14332 ( .A1(n11978), .A2(n14173), .ZN(n11841) );
  NAND2_X1 U14333 ( .A1(n11842), .A2(n11841), .ZN(n12049) );
  XNOR2_X1 U14334 ( .A(n12049), .B(n12048), .ZN(n14986) );
  INV_X1 U14335 ( .A(n12230), .ZN(n14984) );
  OAI21_X1 U14336 ( .B1(n11844), .B2(n14984), .A(n15143), .ZN(n11845) );
  OR2_X1 U14337 ( .A1(n11845), .A2(n12096), .ZN(n14983) );
  OAI22_X1 U14338 ( .A1(n14532), .A2(n11846), .B1(n12228), .B2(n15094), .ZN(
        n11847) );
  AOI21_X1 U14339 ( .B1(n12230), .B2(n14958), .A(n11847), .ZN(n11848) );
  OAI21_X1 U14340 ( .B1(n14983), .B2(n14496), .A(n11848), .ZN(n11849) );
  AOI21_X1 U14341 ( .B1(n14986), .B2(n14967), .A(n11849), .ZN(n11850) );
  OAI21_X1 U14342 ( .B1(n14988), .B2(n15108), .A(n11850), .ZN(P1_U3282) );
  NAND2_X1 U14343 ( .A1(n14905), .A2(n11851), .ZN(n11853) );
  OAI211_X1 U14344 ( .C1(n14911), .C2(n11854), .A(n11853), .B(n11852), .ZN(
        n11859) );
  AOI211_X1 U14345 ( .C1(n11857), .C2(n11856), .A(n13342), .B(n11855), .ZN(
        n11858) );
  AOI211_X1 U14346 ( .C1(n11860), .C2(n14908), .A(n11859), .B(n11858), .ZN(
        n11861) );
  INV_X1 U14347 ( .A(n11861), .ZN(P2_U3189) );
  OR2_X1 U14348 ( .A1(n12477), .A2(n13326), .ZN(n11863) );
  NAND2_X1 U14349 ( .A1(n13353), .A2(n13307), .ZN(n11862) );
  NAND2_X1 U14350 ( .A1(n11863), .A2(n11862), .ZN(n11930) );
  NAND2_X1 U14351 ( .A1(n14905), .A2(n11930), .ZN(n11865) );
  OAI211_X1 U14352 ( .C1(n14911), .C2(n11934), .A(n11865), .B(n11864), .ZN(
        n11872) );
  INV_X1 U14353 ( .A(n11866), .ZN(n11870) );
  AOI22_X1 U14354 ( .A1(n11867), .A2(n14903), .B1(n13313), .B2(n13353), .ZN(
        n11869) );
  NOR3_X1 U14355 ( .A1(n11870), .A2(n11869), .A3(n11868), .ZN(n11871) );
  AOI211_X1 U14356 ( .C1(n7230), .C2(n14908), .A(n11872), .B(n11871), .ZN(
        n11873) );
  OAI21_X1 U14357 ( .B1(n11874), .B2(n13342), .A(n11873), .ZN(P2_U3196) );
  NAND2_X1 U14358 ( .A1(n11879), .A2(n14042), .ZN(n11876) );
  NAND2_X1 U14359 ( .A1(n14175), .A2(n6666), .ZN(n11875) );
  NAND2_X1 U14360 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  XNOR2_X1 U14361 ( .A(n11877), .B(n13985), .ZN(n11907) );
  AND2_X1 U14362 ( .A1(n14175), .A2(n14045), .ZN(n11878) );
  AOI21_X1 U14363 ( .B1(n11879), .B2(n6666), .A(n11878), .ZN(n11906) );
  XNOR2_X1 U14364 ( .A(n11907), .B(n11906), .ZN(n11889) );
  INV_X1 U14365 ( .A(n11882), .ZN(n11884) );
  OR2_X1 U14366 ( .A1(n11884), .A2(n11883), .ZN(n11885) );
  INV_X1 U14367 ( .A(n11915), .ZN(n11887) );
  AOI21_X1 U14368 ( .B1(n11889), .B2(n11888), .A(n11887), .ZN(n11896) );
  AOI21_X1 U14369 ( .B1(n14159), .B2(n11891), .A(n11890), .ZN(n11892) );
  OAI21_X1 U14370 ( .B1(n14150), .B2(n15201), .A(n11892), .ZN(n11893) );
  AOI21_X1 U14371 ( .B1(n11894), .B2(n14124), .A(n11893), .ZN(n11895) );
  OAI21_X1 U14372 ( .B1(n11896), .B2(n14165), .A(n11895), .ZN(P1_U3221) );
  INV_X1 U14373 ( .A(n11897), .ZN(n11898) );
  OAI222_X1 U14374 ( .A1(P3_U3151), .A2(n11899), .B1(n6670), .B2(n11898), .C1(
        n15613), .C2(n13251), .ZN(P3_U3271) );
  INV_X1 U14375 ( .A(n11900), .ZN(n11904) );
  OAI222_X1 U14376 ( .A1(n13894), .A2(n11902), .B1(n13892), .B2(n11904), .C1(
        n11901), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U14377 ( .A1(n11905), .A2(P1_U3086), .B1(n14694), .B2(n11904), 
        .C1(n11903), .C2(n14691), .ZN(P1_U3334) );
  NAND2_X1 U14378 ( .A1(n11907), .A2(n11906), .ZN(n11913) );
  AND2_X1 U14379 ( .A1(n11915), .A2(n11913), .ZN(n11917) );
  NAND2_X1 U14380 ( .A1(n11912), .A2(n14042), .ZN(n11909) );
  NAND2_X1 U14381 ( .A1(n14174), .A2(n6666), .ZN(n11908) );
  NAND2_X1 U14382 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  XNOR2_X1 U14383 ( .A(n11910), .B(n14043), .ZN(n11972) );
  AND2_X1 U14384 ( .A1(n14174), .A2(n14045), .ZN(n11911) );
  AOI21_X1 U14385 ( .B1(n11912), .B2(n6666), .A(n11911), .ZN(n11970) );
  XNOR2_X1 U14386 ( .A(n11972), .B(n11970), .ZN(n11916) );
  AND2_X1 U14387 ( .A1(n11916), .A2(n11913), .ZN(n11914) );
  OAI211_X1 U14388 ( .C1(n11917), .C2(n11916), .A(n14142), .B(n11973), .ZN(
        n11923) );
  NOR2_X1 U14389 ( .A1(n14161), .A2(n11918), .ZN(n11919) );
  AOI211_X1 U14390 ( .C1(n14159), .C2(n11921), .A(n11920), .B(n11919), .ZN(
        n11922) );
  OAI211_X1 U14391 ( .C1(n7087), .C2(n14150), .A(n11923), .B(n11922), .ZN(
        P1_U3231) );
  AND2_X1 U14392 ( .A1(n12064), .A2(n13353), .ZN(n11924) );
  XNOR2_X1 U14393 ( .A(n11989), .B(n11929), .ZN(n14943) );
  NAND2_X1 U14394 ( .A1(n12064), .A2(n11926), .ZN(n11927) );
  NAND2_X1 U14395 ( .A1(n11928), .A2(n11927), .ZN(n11992) );
  XNOR2_X1 U14396 ( .A(n11992), .B(n11929), .ZN(n11931) );
  AOI21_X1 U14397 ( .B1(n11931), .B2(n14915), .A(n11930), .ZN(n11932) );
  OAI21_X1 U14398 ( .B1(n11933), .B2(n14943), .A(n11932), .ZN(n14946) );
  NAND2_X1 U14399 ( .A1(n14946), .A2(n13741), .ZN(n11941) );
  OAI22_X1 U14400 ( .A1(n13741), .A2(n11935), .B1(n11934), .B2(n13737), .ZN(
        n11939) );
  INV_X1 U14401 ( .A(n11995), .ZN(n11936) );
  OAI211_X1 U14402 ( .C1(n14945), .C2(n11937), .A(n11936), .B(n14928), .ZN(
        n14944) );
  NOR2_X1 U14403 ( .A1(n14944), .A2(n13713), .ZN(n11938) );
  AOI211_X1 U14404 ( .C1(n14920), .C2(n7230), .A(n11939), .B(n11938), .ZN(
        n11940) );
  OAI211_X1 U14405 ( .C1(n14943), .C2(n11942), .A(n11941), .B(n11940), .ZN(
        P2_U3253) );
  NOR2_X1 U14406 ( .A1(n11951), .A2(n11943), .ZN(n11945) );
  MUX2_X1 U14407 ( .A(n11946), .B(P3_REG1_REG_12__SCAN_IN), .S(n12183), .Z(
        n11948) );
  INV_X1 U14408 ( .A(n12169), .ZN(n11947) );
  AOI21_X1 U14409 ( .B1(n11949), .B2(n11948), .A(n11947), .ZN(n11966) );
  NOR2_X1 U14410 ( .A1(n11951), .A2(n11950), .ZN(n11953) );
  INV_X1 U14411 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11954) );
  MUX2_X1 U14412 ( .A(n11954), .B(P3_REG2_REG_12__SCAN_IN), .S(n12183), .Z(
        n12182) );
  INV_X1 U14413 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11955) );
  NOR2_X1 U14414 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11955), .ZN(n12417) );
  AOI21_X1 U14415 ( .B1(n15392), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12417), 
        .ZN(n11956) );
  OAI21_X1 U14416 ( .B1(n12847), .B2(n7795), .A(n11956), .ZN(n11964) );
  MUX2_X1 U14417 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12814), .Z(n12172) );
  XNOR2_X1 U14418 ( .A(n12172), .B(n12183), .ZN(n11962) );
  NOR2_X1 U14419 ( .A1(n11958), .A2(n11957), .ZN(n11959) );
  OR2_X1 U14420 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  AOI211_X1 U14421 ( .C1(n11962), .C2(n11961), .A(n12819), .B(n12177), .ZN(
        n11963) );
  AOI211_X1 U14422 ( .C1(n12822), .C2(n12173), .A(n11964), .B(n11963), .ZN(
        n11965) );
  OAI21_X1 U14423 ( .B1(n11966), .B2(n12855), .A(n11965), .ZN(P3_U3194) );
  OAI222_X1 U14424 ( .A1(n13894), .A2(n11969), .B1(P2_U3088), .B2(n11968), 
        .C1(n13892), .C2(n11967), .ZN(P2_U3305) );
  INV_X1 U14425 ( .A(n11970), .ZN(n11971) );
  NAND2_X1 U14426 ( .A1(n11978), .A2(n14042), .ZN(n11975) );
  NAND2_X1 U14427 ( .A1(n14173), .A2(n6666), .ZN(n11974) );
  NAND2_X1 U14428 ( .A1(n11975), .A2(n11974), .ZN(n11976) );
  XNOR2_X1 U14429 ( .A(n11976), .B(n14043), .ZN(n12217) );
  AND2_X1 U14430 ( .A1(n14173), .A2(n14045), .ZN(n11977) );
  AOI21_X1 U14431 ( .B1(n11978), .B2(n6666), .A(n11977), .ZN(n12215) );
  XNOR2_X1 U14432 ( .A(n12217), .B(n12215), .ZN(n12213) );
  XNOR2_X1 U14433 ( .A(n12214), .B(n12213), .ZN(n11987) );
  INV_X1 U14434 ( .A(n14172), .ZN(n12038) );
  NAND2_X1 U14435 ( .A1(n14136), .A2(n14174), .ZN(n11981) );
  INV_X1 U14436 ( .A(n11979), .ZN(n11980) );
  OAI211_X1 U14437 ( .C1(n11982), .C2(n12038), .A(n11981), .B(n11980), .ZN(
        n11984) );
  NOR2_X1 U14438 ( .A1(n15214), .A2(n14150), .ZN(n11983) );
  AOI211_X1 U14439 ( .C1(n11985), .C2(n14124), .A(n11984), .B(n11983), .ZN(
        n11986) );
  OAI21_X1 U14440 ( .B1(n11987), .B2(n14165), .A(n11986), .ZN(P1_U3217) );
  AND2_X1 U14441 ( .A1(n14945), .A2(n11996), .ZN(n11988) );
  OR2_X1 U14442 ( .A1(n14945), .A2(n11996), .ZN(n11990) );
  XNOR2_X1 U14443 ( .A(n12191), .B(n11994), .ZN(n12006) );
  NAND2_X1 U14444 ( .A1(n14945), .A2(n13352), .ZN(n11991) );
  OR2_X1 U14445 ( .A1(n14945), .A2(n13352), .ZN(n11993) );
  XOR2_X1 U14446 ( .A(n11994), .B(n12194), .Z(n12008) );
  NAND2_X1 U14447 ( .A1(n12008), .A2(n13748), .ZN(n12004) );
  OAI211_X1 U14448 ( .C1(n11995), .C2(n12195), .A(n14928), .B(n14926), .ZN(
        n12005) );
  INV_X1 U14449 ( .A(n12005), .ZN(n12002) );
  OR2_X1 U14450 ( .A1(n11996), .A2(n13544), .ZN(n11998) );
  NAND2_X1 U14451 ( .A1(n13350), .A2(n13336), .ZN(n11997) );
  AND2_X1 U14452 ( .A1(n11998), .A2(n11997), .ZN(n12233) );
  OAI22_X1 U14453 ( .A1(n12233), .A2(n14919), .B1(n12236), .B2(n13737), .ZN(
        n11999) );
  AOI21_X1 U14454 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n14919), .A(n11999), 
        .ZN(n12000) );
  OAI21_X1 U14455 ( .B1(n12195), .B2(n13743), .A(n12000), .ZN(n12001) );
  AOI21_X1 U14456 ( .B1(n12002), .B2(n14931), .A(n12001), .ZN(n12003) );
  OAI211_X1 U14457 ( .C1(n12006), .C2(n13751), .A(n12004), .B(n12003), .ZN(
        P2_U3252) );
  OAI211_X1 U14458 ( .C1(n12006), .C2(n13842), .A(n12233), .B(n12005), .ZN(
        n12007) );
  AOI21_X1 U14459 ( .B1(n12008), .B2(n14915), .A(n12007), .ZN(n12012) );
  AOI22_X1 U14460 ( .A1(n12242), .A2(n13837), .B1(n15389), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n12009) );
  OAI21_X1 U14461 ( .B1(n12012), .B2(n15389), .A(n12009), .ZN(P2_U3512) );
  OAI22_X1 U14462 ( .A1(n12195), .A2(n13864), .B1(n15387), .B2(n8181), .ZN(
        n12010) );
  INV_X1 U14463 ( .A(n12010), .ZN(n12011) );
  OAI21_X1 U14464 ( .B1(n12012), .B2(n15386), .A(n12011), .ZN(P2_U3469) );
  INV_X1 U14465 ( .A(n12013), .ZN(n12015) );
  INV_X1 U14466 ( .A(SI_25_), .ZN(n15846) );
  OAI222_X1 U14467 ( .A1(n6670), .A2(n12015), .B1(P3_U3151), .B2(n12014), .C1(
        n15846), .C2(n13251), .ZN(P3_U3270) );
  INV_X1 U14468 ( .A(n15064), .ZN(n15039) );
  INV_X1 U14469 ( .A(n15027), .ZN(n15068) );
  INV_X1 U14470 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n12016) );
  NAND2_X1 U14471 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14078)
         );
  OAI21_X1 U14472 ( .B1(n15068), .B2(n12016), .A(n14078), .ZN(n12024) );
  NAND2_X1 U14473 ( .A1(n15063), .A2(n12019), .ZN(n12020) );
  XNOR2_X1 U14474 ( .A(n14234), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12021) );
  AOI211_X1 U14475 ( .C1(n12022), .C2(n12021), .A(n14233), .B(n15036), .ZN(
        n12023) );
  AOI211_X1 U14476 ( .C1(n15039), .C2(n14234), .A(n12024), .B(n12023), .ZN(
        n12035) );
  OAI21_X1 U14477 ( .B1(n12256), .B2(n12026), .A(n12025), .ZN(n12028) );
  NOR2_X1 U14478 ( .A1(n12027), .A2(n12028), .ZN(n12029) );
  XNOR2_X1 U14479 ( .A(n12028), .B(n12027), .ZN(n15054) );
  NOR2_X1 U14480 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15054), .ZN(n15053) );
  NOR2_X1 U14481 ( .A1(n12029), .A2(n15053), .ZN(n12033) );
  NOR2_X1 U14482 ( .A1(n14230), .A2(n12030), .ZN(n12031) );
  AOI21_X1 U14483 ( .B1(n12030), .B2(n14230), .A(n12031), .ZN(n12032) );
  NAND2_X1 U14484 ( .A1(n12032), .A2(n12033), .ZN(n14229) );
  OAI211_X1 U14485 ( .C1(n12033), .C2(n12032), .A(n15046), .B(n14229), .ZN(
        n12034) );
  NAND2_X1 U14486 ( .A1(n12035), .A2(n12034), .ZN(P1_U3259) );
  OR2_X1 U14487 ( .A1(n12230), .A2(n12038), .ZN(n12039) );
  NAND2_X1 U14488 ( .A1(n12040), .A2(n12039), .ZN(n12085) );
  INV_X1 U14489 ( .A(n12086), .ZN(n12041) );
  NAND2_X1 U14490 ( .A1(n12085), .A2(n12041), .ZN(n12044) );
  OR2_X1 U14491 ( .A1(n14819), .A2(n12042), .ZN(n12043) );
  XNOR2_X1 U14492 ( .A(n12248), .B(n12246), .ZN(n12047) );
  OR2_X1 U14493 ( .A1(n14155), .A2(n14156), .ZN(n12046) );
  NAND2_X1 U14494 ( .A1(n14171), .A2(n14521), .ZN(n12045) );
  NAND2_X1 U14495 ( .A1(n12046), .A2(n12045), .ZN(n12317) );
  AOI21_X1 U14496 ( .B1(n12047), .B2(n15189), .A(n12317), .ZN(n14982) );
  NAND2_X1 U14497 ( .A1(n12049), .A2(n12048), .ZN(n12051) );
  OR2_X1 U14498 ( .A1(n12230), .A2(n14172), .ZN(n12050) );
  NAND2_X1 U14499 ( .A1(n12051), .A2(n12050), .ZN(n12084) );
  NAND2_X1 U14500 ( .A1(n12084), .A2(n12086), .ZN(n12053) );
  OR2_X1 U14501 ( .A1(n14819), .A2(n14171), .ZN(n12052) );
  XNOR2_X1 U14502 ( .A(n12244), .B(n12246), .ZN(n14980) );
  INV_X1 U14503 ( .A(n14819), .ZN(n12281) );
  NAND2_X1 U14504 ( .A1(n12096), .A2(n12281), .ZN(n12095) );
  AOI21_X1 U14505 ( .B1(n12095), .B2(n14976), .A(n15205), .ZN(n12054) );
  NAND2_X1 U14506 ( .A1(n12054), .A2(n12255), .ZN(n14977) );
  OAI22_X1 U14507 ( .A1(n14532), .A2(n12055), .B1(n12320), .B2(n15094), .ZN(
        n12056) );
  AOI21_X1 U14508 ( .B1(n14976), .B2(n14958), .A(n12056), .ZN(n12057) );
  OAI21_X1 U14509 ( .B1(n14977), .B2(n14496), .A(n12057), .ZN(n12058) );
  AOI21_X1 U14510 ( .B1(n14980), .B2(n14967), .A(n12058), .ZN(n12059) );
  OAI21_X1 U14511 ( .B1(n14982), .B2(n15108), .A(n12059), .ZN(P1_U3280) );
  INV_X1 U14512 ( .A(n12060), .ZN(n12061) );
  AOI22_X1 U14513 ( .A1(n12064), .A2(n13837), .B1(n15389), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n12065) );
  OAI21_X1 U14514 ( .B1(n12069), .B2(n15389), .A(n12065), .ZN(P2_U3510) );
  OAI22_X1 U14515 ( .A1(n12066), .A2(n13864), .B1(n15387), .B2(n8126), .ZN(
        n12067) );
  INV_X1 U14516 ( .A(n12067), .ZN(n12068) );
  OAI21_X1 U14517 ( .B1(n12069), .B2(n15386), .A(n12068), .ZN(P2_U3463) );
  NAND2_X1 U14518 ( .A1(n15399), .A2(n15496), .ZN(n12072) );
  NOR2_X1 U14519 ( .A1(n12110), .A2(n12580), .ZN(n12153) );
  NOR2_X1 U14520 ( .A1(n12152), .A2(n12153), .ZN(n12074) );
  XNOR2_X1 U14521 ( .A(n12327), .B(n12079), .ZN(n12076) );
  AOI222_X1 U14522 ( .A1(n15453), .A2(n12076), .B1(n14857), .B2(n15398), .C1(
        n15397), .C2(n15447), .ZN(n15511) );
  OAI22_X1 U14523 ( .A1(n15463), .A2(n12077), .B1(n12121), .B2(n15458), .ZN(
        n12078) );
  AOI21_X1 U14524 ( .B1(n13085), .B2(n12328), .A(n12078), .ZN(n12083) );
  XNOR2_X1 U14525 ( .A(n12080), .B(n12079), .ZN(n15516) );
  NAND2_X1 U14526 ( .A1(n15463), .A2(n15435), .ZN(n12081) );
  NAND2_X1 U14527 ( .A1(n15516), .A2(n14864), .ZN(n12082) );
  OAI211_X1 U14528 ( .C1(n15511), .C2(n15465), .A(n12083), .B(n12082), .ZN(
        P3_U3223) );
  XNOR2_X1 U14529 ( .A(n12084), .B(n12086), .ZN(n12088) );
  INV_X1 U14530 ( .A(n12088), .ZN(n14822) );
  XNOR2_X1 U14531 ( .A(n12085), .B(n12086), .ZN(n12087) );
  NAND2_X1 U14532 ( .A1(n12087), .A2(n15189), .ZN(n12093) );
  NAND2_X1 U14533 ( .A1(n12088), .A2(n15093), .ZN(n12092) );
  NAND2_X1 U14534 ( .A1(n14172), .A2(n14521), .ZN(n12090) );
  NAND2_X1 U14535 ( .A1(n14170), .A2(n14281), .ZN(n12089) );
  NAND2_X1 U14536 ( .A1(n12090), .A2(n12089), .ZN(n12278) );
  INV_X1 U14537 ( .A(n12278), .ZN(n12091) );
  NAND3_X1 U14538 ( .A1(n12093), .A2(n12092), .A3(n12091), .ZN(n14824) );
  NAND2_X1 U14539 ( .A1(n14824), .A2(n14532), .ZN(n12100) );
  OAI22_X1 U14540 ( .A1(n14532), .A2(n12094), .B1(n12275), .B2(n15094), .ZN(
        n12098) );
  OAI211_X1 U14541 ( .C1(n12096), .C2(n12281), .A(n15143), .B(n12095), .ZN(
        n14821) );
  NOR2_X1 U14542 ( .A1(n14821), .A2(n14496), .ZN(n12097) );
  AOI211_X1 U14543 ( .C1(n14958), .C2(n14819), .A(n12098), .B(n12097), .ZN(
        n12099) );
  OAI211_X1 U14544 ( .C1(n14822), .C2(n12101), .A(n12100), .B(n12099), .ZN(
        P1_U3281) );
  INV_X1 U14545 ( .A(n12102), .ZN(n12103) );
  NAND2_X1 U14546 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  XNOR2_X1 U14547 ( .A(n15496), .B(n12532), .ZN(n12108) );
  XNOR2_X1 U14548 ( .A(n12108), .B(n12107), .ZN(n12494) );
  XNOR2_X1 U14549 ( .A(n12580), .B(n12532), .ZN(n12109) );
  XNOR2_X1 U14550 ( .A(n12497), .B(n12109), .ZN(n12577) );
  NAND2_X1 U14551 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  NAND2_X1 U14552 ( .A1(n12112), .A2(n12111), .ZN(n12135) );
  XNOR2_X1 U14553 ( .A(n12114), .B(n12113), .ZN(n12134) );
  XNOR2_X1 U14554 ( .A(n12328), .B(n12532), .ZN(n12341) );
  XNOR2_X1 U14555 ( .A(n12341), .B(n12353), .ZN(n12116) );
  NAND2_X1 U14556 ( .A1(n12114), .A2(n12113), .ZN(n12117) );
  AND2_X1 U14557 ( .A1(n12116), .A2(n12117), .ZN(n12115) );
  NAND2_X1 U14558 ( .A1(n12137), .A2(n12115), .ZN(n12344) );
  INV_X1 U14559 ( .A(n12344), .ZN(n12119) );
  AOI21_X1 U14560 ( .B1(n12137), .B2(n12117), .A(n12116), .ZN(n12118) );
  NOR3_X1 U14561 ( .A1(n12119), .A2(n12118), .A3(n12672), .ZN(n12128) );
  INV_X1 U14562 ( .A(n12668), .ZN(n12681) );
  AOI21_X1 U14563 ( .B1(n14857), .B2(n12681), .A(n12120), .ZN(n12126) );
  INV_X1 U14564 ( .A(n12121), .ZN(n12122) );
  NAND2_X1 U14565 ( .A1(n12666), .A2(n12122), .ZN(n12125) );
  NAND2_X1 U14566 ( .A1(n12670), .A2(n12328), .ZN(n12124) );
  NAND2_X1 U14567 ( .A1(n12657), .A2(n15397), .ZN(n12123) );
  NAND4_X1 U14568 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n12123), .ZN(
        n12127) );
  OR2_X1 U14569 ( .A1(n12128), .A2(n12127), .ZN(P3_U3157) );
  INV_X1 U14570 ( .A(n12129), .ZN(n12160) );
  OR2_X1 U14571 ( .A1(n12497), .A2(n12677), .ZN(n12133) );
  AOI21_X1 U14572 ( .B1(n12670), .B2(n12131), .A(n12130), .ZN(n12132) );
  OAI211_X1 U14573 ( .C1(n12353), .C2(n12668), .A(n12133), .B(n12132), .ZN(
        n12139) );
  NAND2_X1 U14574 ( .A1(n12135), .A2(n12134), .ZN(n12136) );
  AOI21_X1 U14575 ( .B1(n12137), .B2(n12136), .A(n12672), .ZN(n12138) );
  AOI211_X1 U14576 ( .C1(n12160), .C2(n12666), .A(n12139), .B(n12138), .ZN(
        n12140) );
  INV_X1 U14577 ( .A(n12140), .ZN(P3_U3171) );
  NAND2_X1 U14578 ( .A1(n12146), .A2(n12141), .ZN(n12143) );
  OAI211_X1 U14579 ( .C1(n12144), .C2(n14691), .A(n12143), .B(n12142), .ZN(
        P1_U3332) );
  NAND2_X1 U14580 ( .A1(n12146), .A2(n12145), .ZN(n12148) );
  OAI211_X1 U14581 ( .C1(n12149), .C2(n13894), .A(n12148), .B(n12147), .ZN(
        P2_U3304) );
  XNOR2_X1 U14582 ( .A(n12150), .B(n12152), .ZN(n15508) );
  INV_X1 U14583 ( .A(n15508), .ZN(n12163) );
  OAI22_X1 U14584 ( .A1(n12497), .A2(n15425), .B1(n12353), .B2(n15450), .ZN(
        n12157) );
  INV_X1 U14585 ( .A(n12151), .ZN(n15394) );
  OAI21_X1 U14586 ( .B1(n15394), .B2(n12153), .A(n12152), .ZN(n12155) );
  AND3_X1 U14587 ( .A1(n12154), .A2(n15453), .A3(n12155), .ZN(n12156) );
  AOI211_X1 U14588 ( .C1(n15435), .C2(n15508), .A(n12157), .B(n12156), .ZN(
        n15505) );
  MUX2_X1 U14589 ( .A(n12158), .B(n15505), .S(n15463), .Z(n12162) );
  NOR2_X1 U14590 ( .A1(n12159), .A2(n15512), .ZN(n15507) );
  AOI22_X1 U14591 ( .A1(n15507), .A2(n15419), .B1(n15442), .B2(n12160), .ZN(
        n12161) );
  OAI211_X1 U14592 ( .C1(n12163), .C2(n12992), .A(n12162), .B(n12161), .ZN(
        P3_U3224) );
  INV_X1 U14593 ( .A(SI_26_), .ZN(n15877) );
  INV_X1 U14594 ( .A(n12164), .ZN(n12165) );
  OAI222_X1 U14595 ( .A1(n12167), .A2(P3_U3151), .B1(n12166), .B2(n15877), 
        .C1(n6670), .C2(n12165), .ZN(P3_U3269) );
  NAND2_X1 U14596 ( .A1(n12183), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12168) );
  AOI21_X1 U14597 ( .B1(n8877), .B2(n12170), .A(n12710), .ZN(n12189) );
  INV_X1 U14598 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14727) );
  AND2_X1 U14599 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12438) );
  INV_X1 U14600 ( .A(n12438), .ZN(n12171) );
  OAI21_X1 U14601 ( .B1(n12813), .B2(n14727), .A(n12171), .ZN(n12181) );
  INV_X1 U14602 ( .A(n12172), .ZN(n12174) );
  NOR2_X1 U14603 ( .A1(n12174), .A2(n12173), .ZN(n12176) );
  MUX2_X1 U14604 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12814), .Z(n12715) );
  XNOR2_X1 U14605 ( .A(n12715), .B(n12714), .ZN(n12175) );
  INV_X1 U14606 ( .A(n12720), .ZN(n12179) );
  OAI21_X1 U14607 ( .B1(n12177), .B2(n12176), .A(n12175), .ZN(n12178) );
  AOI21_X1 U14608 ( .B1(n12179), .B2(n12178), .A(n12819), .ZN(n12180) );
  AOI211_X1 U14609 ( .C1(n12822), .C2(n7101), .A(n12181), .B(n12180), .ZN(
        n12188) );
  NAND2_X1 U14610 ( .A1(n12183), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12184) );
  AOI21_X1 U14611 ( .B1(n8876), .B2(n12185), .A(n12722), .ZN(n12186) );
  OR2_X1 U14612 ( .A1(n12186), .A2(n12847), .ZN(n12187) );
  OAI211_X1 U14613 ( .C1(n12189), .C2(n12855), .A(n12188), .B(n12187), .ZN(
        P3_U3195) );
  NOR2_X1 U14614 ( .A1(n12195), .A2(n12477), .ZN(n12190) );
  INV_X1 U14615 ( .A(n12477), .ZN(n13351) );
  INV_X1 U14616 ( .A(n14912), .ZN(n14925) );
  NAND2_X1 U14617 ( .A1(n14921), .A2(n13350), .ZN(n12192) );
  NAND2_X1 U14618 ( .A1(n14922), .A2(n12192), .ZN(n12358) );
  XNOR2_X1 U14619 ( .A(n12358), .B(n12200), .ZN(n12283) );
  NOR2_X1 U14620 ( .A1(n12195), .A2(n13351), .ZN(n12193) );
  NAND2_X1 U14621 ( .A1(n12195), .A2(n13351), .ZN(n12196) );
  NAND2_X1 U14622 ( .A1(n14921), .A2(n12198), .ZN(n12199) );
  INV_X1 U14623 ( .A(n12200), .ZN(n12362) );
  XNOR2_X1 U14624 ( .A(n12363), .B(n12362), .ZN(n12285) );
  NAND2_X1 U14625 ( .A1(n12285), .A2(n13748), .ZN(n12208) );
  AND2_X1 U14626 ( .A1(n13350), .A2(n13307), .ZN(n12201) );
  AOI21_X1 U14627 ( .B1(n13348), .B2(n13336), .A(n12201), .ZN(n12293) );
  INV_X1 U14628 ( .A(n12292), .ZN(n12202) );
  AOI22_X1 U14629 ( .A1(n14919), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12202), 
        .B2(n14918), .ZN(n12203) );
  OAI21_X1 U14630 ( .B1(n12293), .B2(n14935), .A(n12203), .ZN(n12206) );
  AND2_X1 U14631 ( .A1(n12364), .A2(n14927), .ZN(n12204) );
  OR3_X1 U14632 ( .A1(n12371), .A2(n12204), .A3(n12389), .ZN(n12282) );
  NOR2_X1 U14633 ( .A1(n12282), .A2(n13713), .ZN(n12205) );
  AOI211_X1 U14634 ( .C1(n14920), .C2(n12364), .A(n12206), .B(n12205), .ZN(
        n12207) );
  OAI211_X1 U14635 ( .C1(n12283), .C2(n13751), .A(n12208), .B(n12207), .ZN(
        P2_U3250) );
  NAND2_X1 U14636 ( .A1(n12230), .A2(n14042), .ZN(n12210) );
  NAND2_X1 U14637 ( .A1(n14172), .A2(n6666), .ZN(n12209) );
  NAND2_X1 U14638 ( .A1(n12210), .A2(n12209), .ZN(n12211) );
  XNOR2_X1 U14639 ( .A(n12211), .B(n13985), .ZN(n12265) );
  AND2_X1 U14640 ( .A1(n14172), .A2(n14045), .ZN(n12212) );
  AOI21_X1 U14641 ( .B1(n12230), .B2(n6666), .A(n12212), .ZN(n12264) );
  XNOR2_X1 U14642 ( .A(n12265), .B(n12264), .ZN(n12224) );
  NAND2_X1 U14643 ( .A1(n12214), .A2(n12213), .ZN(n12219) );
  INV_X1 U14644 ( .A(n12215), .ZN(n12216) );
  NAND2_X1 U14645 ( .A1(n12217), .A2(n12216), .ZN(n12218) );
  INV_X1 U14646 ( .A(n12272), .ZN(n12222) );
  AOI21_X1 U14647 ( .B1(n12224), .B2(n12223), .A(n12222), .ZN(n12232) );
  NAND2_X1 U14648 ( .A1(n14159), .A2(n12225), .ZN(n12226) );
  OAI211_X1 U14649 ( .C1(n14161), .C2(n12228), .A(n12227), .B(n12226), .ZN(
        n12229) );
  AOI21_X1 U14650 ( .B1(n12230), .B2(n14163), .A(n12229), .ZN(n12231) );
  OAI21_X1 U14651 ( .B1(n12232), .B2(n14165), .A(n12231), .ZN(P1_U3236) );
  INV_X1 U14652 ( .A(n12233), .ZN(n12234) );
  AOI22_X1 U14653 ( .A1(n12234), .A2(n14905), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12235) );
  OAI21_X1 U14654 ( .B1(n12236), .B2(n14911), .A(n12235), .ZN(n12241) );
  INV_X1 U14655 ( .A(n12237), .ZN(n12482) );
  AOI211_X1 U14656 ( .C1(n12239), .C2(n12238), .A(n13342), .B(n12482), .ZN(
        n12240) );
  AOI211_X1 U14657 ( .C1(n12242), .C2(n14908), .A(n12241), .B(n12240), .ZN(
        n12243) );
  INV_X1 U14658 ( .A(n12243), .ZN(P2_U3206) );
  OR2_X1 U14659 ( .A1(n14976), .A2(n14170), .ZN(n12245) );
  XNOR2_X1 U14660 ( .A(n14290), .B(n14322), .ZN(n12301) );
  INV_X1 U14661 ( .A(n12246), .ZN(n12247) );
  NAND2_X1 U14662 ( .A1(n12248), .A2(n12247), .ZN(n12250) );
  OR2_X1 U14663 ( .A1(n14976), .A2(n12253), .ZN(n12249) );
  NAND2_X1 U14664 ( .A1(n12250), .A2(n12249), .ZN(n14323) );
  XNOR2_X1 U14665 ( .A(n14323), .B(n12251), .ZN(n12252) );
  NAND2_X1 U14666 ( .A1(n12252), .A2(n15189), .ZN(n12299) );
  INV_X1 U14667 ( .A(n12299), .ZN(n12254) );
  OAI22_X1 U14668 ( .A1(n12253), .A2(n14357), .B1(n14294), .B2(n14156), .ZN(
        n12408) );
  OAI21_X1 U14669 ( .B1(n12254), .B2(n12408), .A(n14532), .ZN(n12260) );
  INV_X1 U14670 ( .A(n14275), .ZN(n14965) );
  AOI211_X1 U14671 ( .C1(n14292), .C2(n12255), .A(n15205), .B(n14965), .ZN(
        n12298) );
  NOR2_X1 U14672 ( .A1(n7088), .A2(n15098), .ZN(n12258) );
  OAI22_X1 U14673 ( .A1(n14532), .A2(n12256), .B1(n12411), .B2(n15094), .ZN(
        n12257) );
  AOI211_X1 U14674 ( .C1(n12298), .C2(n15104), .A(n12258), .B(n12257), .ZN(
        n12259) );
  OAI211_X1 U14675 ( .C1(n12301), .C2(n14564), .A(n12260), .B(n12259), .ZN(
        P1_U3279) );
  INV_X1 U14676 ( .A(n12261), .ZN(n12263) );
  OAI222_X1 U14677 ( .A1(n12814), .A2(P3_U3151), .B1(n6670), .B2(n12263), .C1(
        n12262), .C2(n13251), .ZN(P3_U3268) );
  NAND2_X1 U14678 ( .A1(n12265), .A2(n12264), .ZN(n12270) );
  AND2_X1 U14679 ( .A1(n12272), .A2(n12270), .ZN(n12274) );
  NAND2_X1 U14680 ( .A1(n14819), .A2(n14042), .ZN(n12267) );
  NAND2_X1 U14681 ( .A1(n14171), .A2(n6666), .ZN(n12266) );
  NAND2_X1 U14682 ( .A1(n12267), .A2(n12266), .ZN(n12268) );
  XNOR2_X1 U14683 ( .A(n12268), .B(n14043), .ZN(n12310) );
  AND2_X1 U14684 ( .A1(n14171), .A2(n14045), .ZN(n12269) );
  AOI21_X1 U14685 ( .B1(n14819), .B2(n6666), .A(n12269), .ZN(n12308) );
  XNOR2_X1 U14686 ( .A(n12310), .B(n12308), .ZN(n12273) );
  AND2_X1 U14687 ( .A1(n12273), .A2(n12270), .ZN(n12271) );
  NAND2_X1 U14688 ( .A1(n12272), .A2(n12271), .ZN(n12312) );
  OAI211_X1 U14689 ( .C1(n12274), .C2(n12273), .A(n14142), .B(n12312), .ZN(
        n12280) );
  NOR2_X1 U14690 ( .A1(n14161), .A2(n12275), .ZN(n12276) );
  AOI211_X1 U14691 ( .C1(n14159), .C2(n12278), .A(n12277), .B(n12276), .ZN(
        n12279) );
  OAI211_X1 U14692 ( .C1(n12281), .C2(n14150), .A(n12280), .B(n12279), .ZN(
        P1_U3224) );
  OAI211_X1 U14693 ( .C1(n12283), .C2(n13842), .A(n12293), .B(n12282), .ZN(
        n12284) );
  AOI21_X1 U14694 ( .B1(n14915), .B2(n12285), .A(n12284), .ZN(n12290) );
  AOI22_X1 U14695 ( .A1(n12364), .A2(n13837), .B1(n15389), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n12286) );
  OAI21_X1 U14696 ( .B1(n12290), .B2(n15389), .A(n12286), .ZN(P2_U3514) );
  INV_X1 U14697 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n12287) );
  OAI22_X1 U14698 ( .A1(n7703), .A2(n13864), .B1(n15387), .B2(n12287), .ZN(
        n12288) );
  INV_X1 U14699 ( .A(n12288), .ZN(n12289) );
  OAI21_X1 U14700 ( .B1(n12290), .B2(n15386), .A(n12289), .ZN(P2_U3475) );
  AOI22_X1 U14701 ( .A1(n12291), .A2(n14903), .B1(n13313), .B2(n13349), .ZN(
        n12297) );
  NOR2_X1 U14702 ( .A1(n14911), .A2(n12292), .ZN(n12295) );
  INV_X1 U14703 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n15288) );
  OAI22_X1 U14704 ( .A1(n12293), .A2(n13339), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15288), .ZN(n12294) );
  AOI211_X1 U14705 ( .C1(n12364), .C2(n14908), .A(n12295), .B(n12294), .ZN(
        n12296) );
  OAI21_X1 U14706 ( .B1(n12297), .B2(n6818), .A(n12296), .ZN(P2_U3213) );
  AOI211_X1 U14707 ( .C1(n14292), .C2(n15192), .A(n12408), .B(n12298), .ZN(
        n12300) );
  OAI211_X1 U14708 ( .C1(n15176), .C2(n12301), .A(n12300), .B(n12299), .ZN(
        n12305) );
  NAND2_X1 U14709 ( .A1(n12305), .A2(n15233), .ZN(n12302) );
  OAI21_X1 U14710 ( .B1(n15233), .B2(n11336), .A(n12302), .ZN(P1_U3542) );
  AND2_X2 U14711 ( .A1(n12304), .A2(n12303), .ZN(n15221) );
  INV_X1 U14712 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U14713 ( .A1(n12305), .A2(n15221), .ZN(n12306) );
  OAI21_X1 U14714 ( .B1(n15221), .B2(n12307), .A(n12306), .ZN(P1_U3501) );
  INV_X1 U14715 ( .A(n12308), .ZN(n12309) );
  NAND2_X1 U14716 ( .A1(n12310), .A2(n12309), .ZN(n12311) );
  NAND2_X1 U14717 ( .A1(n14976), .A2(n14042), .ZN(n12314) );
  NAND2_X1 U14718 ( .A1(n14170), .A2(n6666), .ZN(n12313) );
  NAND2_X1 U14719 ( .A1(n12314), .A2(n12313), .ZN(n12315) );
  XNOR2_X1 U14720 ( .A(n12315), .B(n14043), .ZN(n12405) );
  AND2_X1 U14721 ( .A1(n14170), .A2(n14045), .ZN(n12316) );
  AOI21_X1 U14722 ( .B1(n14976), .B2(n6666), .A(n12316), .ZN(n12403) );
  XNOR2_X1 U14723 ( .A(n12405), .B(n12403), .ZN(n12401) );
  XNOR2_X1 U14724 ( .A(n12402), .B(n12401), .ZN(n12323) );
  NAND2_X1 U14725 ( .A1(n14159), .A2(n12317), .ZN(n12318) );
  OAI211_X1 U14726 ( .C1(n14161), .C2(n12320), .A(n12319), .B(n12318), .ZN(
        n12321) );
  AOI21_X1 U14727 ( .B1(n14976), .B2(n14163), .A(n12321), .ZN(n12322) );
  OAI21_X1 U14728 ( .B1(n12323), .B2(n14165), .A(n12322), .ZN(P1_U3234) );
  OAI21_X1 U14729 ( .B1(n12325), .B2(n12334), .A(n12324), .ZN(n14881) );
  INV_X1 U14730 ( .A(n14881), .ZN(n12340) );
  NAND2_X1 U14731 ( .A1(n12327), .A2(n12326), .ZN(n12330) );
  NAND2_X1 U14732 ( .A1(n12342), .A2(n12328), .ZN(n12329) );
  INV_X1 U14733 ( .A(n12333), .ZN(n12332) );
  AOI21_X1 U14734 ( .B1(n12334), .B2(n12333), .A(n6980), .ZN(n12335) );
  OAI222_X1 U14735 ( .A1(n15450), .A2(n12870), .B1(n15425), .B2(n12353), .C1(
        n15430), .C2(n12335), .ZN(n14879) );
  NAND2_X1 U14736 ( .A1(n14879), .A2(n15463), .ZN(n12339) );
  AND2_X1 U14737 ( .A1(n12355), .A2(n15495), .ZN(n14880) );
  OAI22_X1 U14738 ( .A1(n15463), .A2(n12336), .B1(n12349), .B2(n15458), .ZN(
        n12337) );
  AOI21_X1 U14739 ( .B1(n15419), .B2(n14880), .A(n12337), .ZN(n12338) );
  OAI211_X1 U14740 ( .C1(n15460), .C2(n12340), .A(n12339), .B(n12338), .ZN(
        P3_U3222) );
  NAND2_X1 U14741 ( .A1(n12342), .A2(n12341), .ZN(n12343) );
  INV_X1 U14742 ( .A(n12345), .ZN(n12346) );
  AOI21_X1 U14743 ( .B1(n14857), .B2(n12347), .A(n6816), .ZN(n12357) );
  AOI21_X1 U14744 ( .B1(n14844), .B2(n12681), .A(n12348), .ZN(n12352) );
  INV_X1 U14745 ( .A(n12349), .ZN(n12350) );
  NAND2_X1 U14746 ( .A1(n12666), .A2(n12350), .ZN(n12351) );
  OAI211_X1 U14747 ( .C1(n12353), .C2(n12677), .A(n12352), .B(n12351), .ZN(
        n12354) );
  AOI21_X1 U14748 ( .B1(n12355), .B2(n12670), .A(n12354), .ZN(n12356) );
  OAI21_X1 U14749 ( .B1(n12357), .B2(n12672), .A(n12356), .ZN(P3_U3176) );
  NAND2_X1 U14750 ( .A1(n12360), .A2(n12367), .ZN(n12361) );
  NAND2_X1 U14751 ( .A1(n12384), .A2(n12361), .ZN(n13843) );
  NAND2_X1 U14752 ( .A1(n12363), .A2(n12362), .ZN(n12366) );
  NAND2_X1 U14753 ( .A1(n12364), .A2(n12368), .ZN(n12365) );
  XNOR2_X1 U14754 ( .A(n12377), .B(n12367), .ZN(n12369) );
  OAI22_X1 U14755 ( .A1(n13549), .A2(n13326), .B1(n12368), .B2(n13544), .ZN(
        n14892) );
  AOI21_X1 U14756 ( .B1(n12369), .B2(n14915), .A(n14892), .ZN(n13841) );
  OAI21_X1 U14757 ( .B1(n14896), .B2(n13737), .A(n13841), .ZN(n12370) );
  NAND2_X1 U14758 ( .A1(n12370), .A2(n13741), .ZN(n12375) );
  INV_X1 U14759 ( .A(n12371), .ZN(n12372) );
  AOI211_X1 U14760 ( .C1(n14893), .C2(n12372), .A(n13720), .B(n12388), .ZN(
        n13839) );
  INV_X1 U14761 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13463) );
  OAI22_X1 U14762 ( .A1(n12383), .A2(n13743), .B1(n13463), .B2(n13741), .ZN(
        n12373) );
  AOI21_X1 U14763 ( .B1(n13839), .B2(n14931), .A(n12373), .ZN(n12374) );
  OAI211_X1 U14764 ( .C1(n13843), .C2(n13751), .A(n12375), .B(n12374), .ZN(
        P2_U3249) );
  NOR2_X1 U14765 ( .A1(n12383), .A2(n13348), .ZN(n12376) );
  NAND2_X1 U14766 ( .A1(n12383), .A2(n13348), .ZN(n12378) );
  INV_X1 U14767 ( .A(n13509), .ZN(n12385) );
  XNOR2_X1 U14768 ( .A(n13510), .B(n12385), .ZN(n12381) );
  OR2_X1 U14769 ( .A1(n13553), .A2(n13326), .ZN(n12380) );
  NAND2_X1 U14770 ( .A1(n13348), .A2(n13307), .ZN(n12379) );
  NAND2_X1 U14771 ( .A1(n12380), .A2(n12379), .ZN(n14906) );
  AOI21_X1 U14772 ( .B1(n12381), .B2(n14915), .A(n14906), .ZN(n13834) );
  OR2_X1 U14773 ( .A1(n12386), .A2(n12385), .ZN(n12387) );
  NAND2_X1 U14774 ( .A1(n13552), .A2(n12387), .ZN(n13835) );
  INV_X1 U14775 ( .A(n13835), .ZN(n12395) );
  NOR2_X1 U14776 ( .A1(n13550), .A2(n12388), .ZN(n12390) );
  OR3_X1 U14777 ( .A1(n12390), .A2(n13734), .A3(n12389), .ZN(n13833) );
  NAND2_X1 U14778 ( .A1(n14919), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12391) );
  OAI21_X1 U14779 ( .B1(n13737), .B2(n14910), .A(n12391), .ZN(n12392) );
  AOI21_X1 U14780 ( .B1(n14907), .B2(n14920), .A(n12392), .ZN(n12393) );
  OAI21_X1 U14781 ( .B1(n13833), .B2(n13713), .A(n12393), .ZN(n12394) );
  AOI21_X1 U14782 ( .B1(n12395), .B2(n14932), .A(n12394), .ZN(n12396) );
  OAI21_X1 U14783 ( .B1(n14935), .B2(n13834), .A(n12396), .ZN(P2_U3248) );
  NAND2_X1 U14784 ( .A1(n14292), .A2(n14042), .ZN(n12398) );
  OR2_X1 U14785 ( .A1(n14155), .A2(n13941), .ZN(n12397) );
  NAND2_X1 U14786 ( .A1(n12398), .A2(n12397), .ZN(n12399) );
  XNOR2_X1 U14787 ( .A(n12399), .B(n13985), .ZN(n13910) );
  NOR2_X1 U14788 ( .A1(n14155), .A2(n13940), .ZN(n12400) );
  AOI21_X1 U14789 ( .B1(n14292), .B2(n6666), .A(n12400), .ZN(n13909) );
  XNOR2_X1 U14790 ( .A(n13910), .B(n13909), .ZN(n13908) );
  NAND2_X1 U14791 ( .A1(n12402), .A2(n12401), .ZN(n12407) );
  INV_X1 U14792 ( .A(n12403), .ZN(n12404) );
  NAND2_X1 U14793 ( .A1(n12405), .A2(n12404), .ZN(n12406) );
  XOR2_X1 U14794 ( .A(n13907), .B(n13908), .Z(n12414) );
  NAND2_X1 U14795 ( .A1(n14159), .A2(n12408), .ZN(n12409) );
  OAI211_X1 U14796 ( .C1(n14161), .C2(n12411), .A(n12410), .B(n12409), .ZN(
        n12412) );
  AOI21_X1 U14797 ( .B1(n14292), .B2(n14163), .A(n12412), .ZN(n12413) );
  OAI21_X1 U14798 ( .B1(n12414), .B2(n14165), .A(n12413), .ZN(P1_U3215) );
  XNOR2_X1 U14799 ( .A(n12432), .B(n14844), .ZN(n12415) );
  XNOR2_X1 U14800 ( .A(n12431), .B(n12415), .ZN(n12423) );
  NOR2_X1 U14801 ( .A1(n12871), .A2(n12668), .ZN(n12416) );
  AOI211_X1 U14802 ( .C1(n12657), .C2(n14857), .A(n12417), .B(n12416), .ZN(
        n12418) );
  OAI21_X1 U14803 ( .B1(n12419), .B2(n12678), .A(n12418), .ZN(n12420) );
  AOI21_X1 U14804 ( .B1(n12670), .B2(n12421), .A(n12420), .ZN(n12422) );
  OAI21_X1 U14805 ( .B1(n12423), .B2(n12672), .A(n12422), .ZN(P3_U3164) );
  INV_X1 U14806 ( .A(n12424), .ZN(n12428) );
  OAI222_X1 U14807 ( .A1(P1_U3086), .A2(n12426), .B1(n14694), .B2(n12428), 
        .C1(n12425), .C2(n14691), .ZN(P1_U3331) );
  OAI222_X1 U14808 ( .A1(n12429), .A2(P2_U3088), .B1(n13892), .B2(n12428), 
        .C1(n12427), .C2(n13894), .ZN(P2_U3303) );
  NAND2_X1 U14809 ( .A1(n12432), .A2(n14844), .ZN(n12430) );
  NAND2_X1 U14810 ( .A1(n12431), .A2(n12430), .ZN(n12435) );
  INV_X1 U14811 ( .A(n12432), .ZN(n12433) );
  NAND2_X1 U14812 ( .A1(n12433), .A2(n12870), .ZN(n12434) );
  XNOR2_X1 U14813 ( .A(n12505), .B(n12871), .ZN(n12436) );
  XNOR2_X1 U14814 ( .A(n12507), .B(n12436), .ZN(n12442) );
  NOR2_X1 U14815 ( .A1(n12870), .A2(n12677), .ZN(n12437) );
  AOI211_X1 U14816 ( .C1(n12681), .C2(n14843), .A(n12438), .B(n12437), .ZN(
        n12439) );
  OAI21_X1 U14817 ( .B1(n14847), .B2(n12678), .A(n12439), .ZN(n12440) );
  AOI21_X1 U14818 ( .B1(n14850), .B2(n12670), .A(n12440), .ZN(n12441) );
  OAI21_X1 U14819 ( .B1(n12442), .B2(n12672), .A(n12441), .ZN(P3_U3174) );
  INV_X1 U14820 ( .A(n12443), .ZN(n12462) );
  INV_X1 U14821 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12444) );
  OAI222_X1 U14822 ( .A1(P1_U3086), .A2(n12445), .B1(n14694), .B2(n12462), 
        .C1(n12444), .C2(n14691), .ZN(P1_U3326) );
  INV_X1 U14823 ( .A(n12446), .ZN(n12463) );
  OAI222_X1 U14824 ( .A1(n10107), .A2(P1_U3086), .B1(n14694), .B2(n12463), 
        .C1(n12447), .C2(n14691), .ZN(P1_U3327) );
  NAND2_X1 U14825 ( .A1(n13719), .A2(n13816), .ZN(n13707) );
  OR2_X1 U14826 ( .A1(n13707), .A2(n13699), .ZN(n13694) );
  AND2_X2 U14827 ( .A1(n13619), .A2(n13641), .ZN(n13621) );
  NAND2_X1 U14828 ( .A1(n13580), .A2(n13593), .ZN(n13577) );
  NAND2_X1 U14829 ( .A1(n12448), .A2(n13504), .ZN(n13499) );
  OAI211_X1 U14830 ( .C1(n12448), .C2(n13504), .A(n14928), .B(n13499), .ZN(
        n13508) );
  NOR2_X1 U14831 ( .A1(n12458), .A2(n12449), .ZN(n12450) );
  OR2_X1 U14832 ( .A1(n13326), .A2(n12450), .ZN(n13542) );
  INV_X1 U14833 ( .A(n13542), .ZN(n12451) );
  AND2_X1 U14834 ( .A1(n13344), .A2(n12451), .ZN(n13752) );
  INV_X1 U14835 ( .A(n13752), .ZN(n13501) );
  AND2_X1 U14836 ( .A1(n13508), .A2(n13501), .ZN(n12454) );
  MUX2_X1 U14837 ( .A(n12454), .B(n12452), .S(n15386), .Z(n12453) );
  OAI21_X1 U14838 ( .B1(n13504), .B2(n13864), .A(n12453), .ZN(P2_U3497) );
  MUX2_X1 U14839 ( .A(n12455), .B(n12454), .S(n15391), .Z(n12456) );
  OAI21_X1 U14840 ( .B1(n13504), .B2(n7353), .A(n12456), .ZN(P2_U3529) );
  INV_X1 U14841 ( .A(n12457), .ZN(n14686) );
  OAI222_X1 U14842 ( .A1(n13894), .A2(n12459), .B1(n13892), .B2(n14686), .C1(
        P2_U3088), .C2(n12458), .ZN(P2_U3300) );
  OAI222_X1 U14843 ( .A1(n13892), .A2(n12462), .B1(P2_U3088), .B2(n12461), 
        .C1(n12460), .C2(n13894), .ZN(P2_U3298) );
  OAI222_X1 U14844 ( .A1(n13894), .A2(n12464), .B1(n13892), .B2(n12463), .C1(
        n8626), .C2(P2_U3088), .ZN(P2_U3299) );
  OAI222_X1 U14845 ( .A1(n13894), .A2(n12467), .B1(n13892), .B2(n12466), .C1(
        n12465), .C2(P2_U3088), .ZN(P2_U3308) );
  NAND2_X1 U14846 ( .A1(n15306), .A2(n13370), .ZN(n12468) );
  OAI211_X1 U14847 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15319), .A(n12468), .B(
        n15325), .ZN(n12472) );
  OAI22_X1 U14848 ( .A1(n15330), .A2(n13370), .B1(n12469), .B2(n15319), .ZN(
        n12471) );
  MUX2_X1 U14849 ( .A(n12472), .B(n12471), .S(n12470), .Z(n12476) );
  INV_X1 U14850 ( .A(n15328), .ZN(n15298) );
  INV_X1 U14851 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n12474) );
  OAI22_X1 U14852 ( .A1(n15298), .A2(n12474), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12473), .ZN(n12475) );
  OR2_X1 U14853 ( .A1(n12476), .A2(n12475), .ZN(P2_U3214) );
  OR2_X1 U14854 ( .A1(n12477), .A2(n13544), .ZN(n12479) );
  NAND2_X1 U14855 ( .A1(n13349), .A2(n13336), .ZN(n12478) );
  NAND2_X1 U14856 ( .A1(n12479), .A2(n12478), .ZN(n14914) );
  AOI22_X1 U14857 ( .A1(n14905), .A2(n14914), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12480) );
  OAI21_X1 U14858 ( .B1(n12481), .B2(n14911), .A(n12480), .ZN(n12488) );
  NAND2_X1 U14859 ( .A1(n12482), .A2(n14903), .ZN(n12486) );
  NAND3_X1 U14860 ( .A1(n12483), .A2(n13313), .A3(n13351), .ZN(n12485) );
  AOI21_X1 U14861 ( .B1(n12486), .B2(n12485), .A(n12484), .ZN(n12487) );
  AOI211_X1 U14862 ( .C1(n14921), .C2(n14908), .A(n12488), .B(n12487), .ZN(
        n12489) );
  OAI21_X1 U14863 ( .B1(n12490), .B2(n13342), .A(n12489), .ZN(P2_U3187) );
  INV_X1 U14864 ( .A(n12491), .ZN(n12492) );
  OAI222_X1 U14865 ( .A1(n6670), .A2(n12492), .B1(n12857), .B2(P3_U3151), .C1(
        n15799), .C2(n13251), .ZN(P3_U3267) );
  XOR2_X1 U14866 ( .A(n12494), .B(n12493), .Z(n12495) );
  NAND2_X1 U14867 ( .A1(n12495), .A2(n7432), .ZN(n12504) );
  AOI21_X1 U14868 ( .B1(n12670), .B2(n15496), .A(n12496), .ZN(n12503) );
  OAI22_X1 U14869 ( .A1(n12497), .A2(n12668), .B1(n12613), .B2(n12677), .ZN(
        n12498) );
  INV_X1 U14870 ( .A(n12498), .ZN(n12502) );
  INV_X1 U14871 ( .A(n12499), .ZN(n12500) );
  NAND2_X1 U14872 ( .A1(n12666), .A2(n12500), .ZN(n12501) );
  NAND4_X1 U14873 ( .A1(n12504), .A2(n12503), .A3(n12502), .A4(n12501), .ZN(
        P3_U3153) );
  XNOR2_X1 U14874 ( .A(n12933), .B(n12532), .ZN(n12566) );
  XNOR2_X1 U14875 ( .A(n12566), .B(n12943), .ZN(n12568) );
  INV_X1 U14876 ( .A(n12631), .ZN(n12529) );
  AOI21_X1 U14877 ( .B1(n12551), .B2(n12997), .A(n12630), .ZN(n12528) );
  XNOR2_X1 U14878 ( .A(n12889), .B(n12532), .ZN(n12547) );
  AND2_X1 U14879 ( .A1(n12505), .A2(n12871), .ZN(n12506) );
  AND2_X1 U14880 ( .A1(n12539), .A2(n14843), .ZN(n12508) );
  INV_X1 U14881 ( .A(n12539), .ZN(n12509) );
  INV_X1 U14882 ( .A(n14843), .ZN(n12872) );
  NAND2_X1 U14883 ( .A1(n12509), .A2(n12872), .ZN(n12510) );
  INV_X1 U14884 ( .A(n14833), .ZN(n13078) );
  XNOR2_X1 U14885 ( .A(n12511), .B(n13078), .ZN(n12675) );
  NAND2_X1 U14886 ( .A1(n12511), .A2(n14833), .ZN(n12512) );
  XNOR2_X1 U14887 ( .A(n13174), .B(n12532), .ZN(n12599) );
  INV_X1 U14888 ( .A(n12656), .ZN(n13077) );
  XNOR2_X1 U14889 ( .A(n12513), .B(n13077), .ZN(n12621) );
  XNOR2_X1 U14890 ( .A(n12514), .B(n12880), .ZN(n12654) );
  NAND2_X1 U14891 ( .A1(n12655), .A2(n12654), .ZN(n12517) );
  INV_X1 U14892 ( .A(n12514), .ZN(n12515) );
  NAND2_X1 U14893 ( .A1(n12515), .A2(n12880), .ZN(n12516) );
  NAND2_X1 U14894 ( .A1(n12517), .A2(n12516), .ZN(n12559) );
  NAND2_X1 U14895 ( .A1(n12518), .A2(n13051), .ZN(n12557) );
  NAND2_X1 U14896 ( .A1(n12559), .A2(n12557), .ZN(n12520) );
  INV_X1 U14897 ( .A(n12518), .ZN(n12519) );
  NAND2_X1 U14898 ( .A1(n12519), .A2(n12883), .ZN(n12558) );
  NAND2_X1 U14899 ( .A1(n12520), .A2(n12558), .ZN(n12641) );
  XNOR2_X1 U14900 ( .A(n12521), .B(n12885), .ZN(n12640) );
  INV_X1 U14901 ( .A(n12521), .ZN(n12522) );
  NAND2_X1 U14902 ( .A1(n12522), .A2(n12885), .ZN(n12523) );
  XNOR2_X1 U14903 ( .A(n12524), .B(n13018), .ZN(n12586) );
  INV_X1 U14904 ( .A(n12551), .ZN(n12628) );
  AOI22_X1 U14905 ( .A1(n12628), .A2(n12892), .B1(n12547), .B2(n12985), .ZN(
        n12525) );
  NAND3_X1 U14906 ( .A1(n12551), .A2(n12630), .A3(n12997), .ZN(n12526) );
  OAI211_X1 U14907 ( .C1(n12529), .C2(n12528), .A(n12527), .B(n12526), .ZN(
        n12592) );
  XNOR2_X1 U14908 ( .A(n12960), .B(n12532), .ZN(n12530) );
  XNOR2_X1 U14909 ( .A(n12530), .B(n12970), .ZN(n12593) );
  INV_X1 U14910 ( .A(n12530), .ZN(n12531) );
  AOI22_X1 U14911 ( .A1(n12592), .A2(n12593), .B1(n12970), .B2(n12531), .ZN(
        n12663) );
  XNOR2_X1 U14912 ( .A(n13125), .B(n12532), .ZN(n12533) );
  XNOR2_X1 U14913 ( .A(n12533), .B(n12898), .ZN(n12664) );
  XOR2_X1 U14914 ( .A(n12568), .B(n12569), .Z(n12538) );
  AOI22_X1 U14915 ( .A1(n12934), .A2(n12666), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12535) );
  NAND2_X1 U14916 ( .A1(n12898), .A2(n12657), .ZN(n12534) );
  OAI211_X1 U14917 ( .C1(n12930), .C2(n12668), .A(n12535), .B(n12534), .ZN(
        n12536) );
  AOI21_X1 U14918 ( .B1(n12933), .B2(n12670), .A(n12536), .ZN(n12537) );
  OAI21_X1 U14919 ( .B1(n12538), .B2(n12672), .A(n12537), .ZN(P3_U3154) );
  XNOR2_X1 U14920 ( .A(n12539), .B(n12872), .ZN(n12540) );
  XNOR2_X1 U14921 ( .A(n12541), .B(n12540), .ZN(n12546) );
  INV_X1 U14922 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15600) );
  NOR2_X1 U14923 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15600), .ZN(n12727) );
  AOI21_X1 U14924 ( .B1(n12681), .B2(n14833), .A(n12727), .ZN(n12542) );
  OAI21_X1 U14925 ( .B1(n12871), .B2(n12677), .A(n12542), .ZN(n12544) );
  NOR2_X1 U14926 ( .A1(n14838), .A2(n12684), .ZN(n12543) );
  AOI211_X1 U14927 ( .C1(n14835), .C2(n12666), .A(n12544), .B(n12543), .ZN(
        n12545) );
  OAI21_X1 U14928 ( .B1(n12546), .B2(n12672), .A(n12545), .ZN(P3_U3155) );
  XNOR2_X1 U14929 ( .A(n12549), .B(n12547), .ZN(n12647) );
  INV_X1 U14930 ( .A(n12547), .ZN(n12548) );
  AND2_X1 U14931 ( .A1(n12549), .A2(n12548), .ZN(n12550) );
  AOI21_X1 U14932 ( .B1(n12647), .B2(n13007), .A(n12550), .ZN(n12627) );
  XOR2_X1 U14933 ( .A(n12551), .B(n12627), .Z(n12629) );
  XNOR2_X1 U14934 ( .A(n12629), .B(n12997), .ZN(n12556) );
  AOI22_X1 U14935 ( .A1(n12985), .A2(n12657), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12553) );
  NAND2_X1 U14936 ( .A1(n12989), .A2(n12666), .ZN(n12552) );
  OAI211_X1 U14937 ( .C1(n12630), .C2(n12668), .A(n12553), .B(n12552), .ZN(
        n12554) );
  AOI21_X1 U14938 ( .B1(n13139), .B2(n12670), .A(n12554), .ZN(n12555) );
  OAI21_X1 U14939 ( .B1(n12556), .B2(n12672), .A(n12555), .ZN(P3_U3156) );
  NAND2_X1 U14940 ( .A1(n12558), .A2(n12557), .ZN(n12560) );
  XOR2_X1 U14941 ( .A(n12560), .B(n12559), .Z(n12565) );
  NAND2_X1 U14942 ( .A1(n12880), .A2(n12657), .ZN(n12561) );
  NAND2_X1 U14943 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12849)
         );
  OAI211_X1 U14944 ( .C1(n13031), .C2(n12668), .A(n12561), .B(n12849), .ZN(
        n12562) );
  AOI21_X1 U14945 ( .B1(n13035), .B2(n12666), .A(n12562), .ZN(n12564) );
  NAND2_X1 U14946 ( .A1(n13157), .A2(n12670), .ZN(n12563) );
  OAI211_X1 U14947 ( .C1(n12565), .C2(n12672), .A(n12564), .B(n12563), .ZN(
        P3_U3159) );
  INV_X1 U14948 ( .A(n12566), .ZN(n12567) );
  INV_X1 U14949 ( .A(n12921), .ZN(n12572) );
  OAI22_X1 U14950 ( .A1(n12572), .A2(n12678), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12571), .ZN(n12574) );
  OAI22_X1 U14951 ( .A1(n12916), .A2(n12668), .B1(n12943), .B2(n12677), .ZN(
        n12573) );
  AOI211_X1 U14952 ( .C1(n13118), .C2(n12670), .A(n12574), .B(n12573), .ZN(
        n12575) );
  XOR2_X1 U14953 ( .A(n12577), .B(n12576), .Z(n12578) );
  NAND2_X1 U14954 ( .A1(n12578), .A2(n7432), .ZN(n12584) );
  AOI21_X1 U14955 ( .B1(n12670), .B2(n12580), .A(n12579), .ZN(n12583) );
  AOI22_X1 U14956 ( .A1(n15399), .A2(n12657), .B1(n12681), .B2(n15397), .ZN(
        n12582) );
  NAND2_X1 U14957 ( .A1(n12666), .A2(n15404), .ZN(n12581) );
  NAND4_X1 U14958 ( .A1(n12584), .A2(n12583), .A3(n12582), .A4(n12581), .ZN(
        P3_U3161) );
  AOI21_X1 U14959 ( .B1(n12586), .B2(n12585), .A(n6752), .ZN(n12591) );
  AOI22_X1 U14960 ( .A1(n12885), .A2(n12657), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12588) );
  NAND2_X1 U14961 ( .A1(n12666), .A2(n13011), .ZN(n12587) );
  OAI211_X1 U14962 ( .C1(n13007), .C2(n12668), .A(n12588), .B(n12587), .ZN(
        n12589) );
  AOI21_X1 U14963 ( .B1(n13010), .B2(n12670), .A(n12589), .ZN(n12590) );
  OAI21_X1 U14964 ( .B1(n12591), .B2(n12672), .A(n12590), .ZN(P3_U3163) );
  XOR2_X1 U14965 ( .A(n12593), .B(n12592), .Z(n12598) );
  AOI22_X1 U14966 ( .A1(n12986), .A2(n12657), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12595) );
  NAND2_X1 U14967 ( .A1(n12961), .A2(n12666), .ZN(n12594) );
  OAI211_X1 U14968 ( .C1(n12956), .C2(n12668), .A(n12595), .B(n12594), .ZN(
        n12596) );
  AOI21_X1 U14969 ( .B1(n12960), .B2(n12670), .A(n12596), .ZN(n12597) );
  OAI21_X1 U14970 ( .B1(n12598), .B2(n12672), .A(n12597), .ZN(P3_U3165) );
  XNOR2_X1 U14971 ( .A(n12599), .B(n13062), .ZN(n12600) );
  XNOR2_X1 U14972 ( .A(n12601), .B(n12600), .ZN(n12606) );
  NAND2_X1 U14973 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12772)
         );
  OAI21_X1 U14974 ( .B1(n13077), .B2(n12668), .A(n12772), .ZN(n12602) );
  AOI21_X1 U14975 ( .B1(n12657), .B2(n14833), .A(n12602), .ZN(n12603) );
  OAI21_X1 U14976 ( .B1(n13082), .B2(n12678), .A(n12603), .ZN(n12604) );
  AOI21_X1 U14977 ( .B1(n13174), .B2(n12670), .A(n12604), .ZN(n12605) );
  OAI21_X1 U14978 ( .B1(n12606), .B2(n12672), .A(n12605), .ZN(P3_U3166) );
  OAI21_X1 U14979 ( .B1(n12609), .B2(n12608), .A(n12607), .ZN(n12610) );
  NAND2_X1 U14980 ( .A1(n12610), .A2(n7432), .ZN(n12619) );
  AOI21_X1 U14981 ( .B1(n12670), .B2(n12612), .A(n12611), .ZN(n12618) );
  OAI22_X1 U14982 ( .A1(n15408), .A2(n12677), .B1(n12613), .B2(n12668), .ZN(
        n12614) );
  INV_X1 U14983 ( .A(n12614), .ZN(n12617) );
  NAND2_X1 U14984 ( .A1(n12666), .A2(n12615), .ZN(n12616) );
  NAND4_X1 U14985 ( .A1(n12619), .A2(n12618), .A3(n12617), .A4(n12616), .ZN(
        P3_U3167) );
  XOR2_X1 U14986 ( .A(n12621), .B(n12620), .Z(n12622) );
  NAND2_X1 U14987 ( .A1(n12622), .A2(n7432), .ZN(n12626) );
  NAND2_X1 U14988 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12798)
         );
  OAI21_X1 U14989 ( .B1(n13061), .B2(n12668), .A(n12798), .ZN(n12624) );
  NOR2_X1 U14990 ( .A1(n12678), .A2(n13070), .ZN(n12623) );
  AOI211_X1 U14991 ( .C1(n12657), .C2(n13094), .A(n12624), .B(n12623), .ZN(
        n12625) );
  OAI211_X1 U14992 ( .C1(n12684), .C2(n13171), .A(n12626), .B(n12625), .ZN(
        P3_U3168) );
  OAI22_X1 U14993 ( .A1(n12629), .A2(n12892), .B1(n12628), .B2(n12627), .ZN(
        n12633) );
  XNOR2_X1 U14994 ( .A(n12631), .B(n12630), .ZN(n12632) );
  XNOR2_X1 U14995 ( .A(n12633), .B(n12632), .ZN(n12638) );
  OAI22_X1 U14996 ( .A1(n12997), .A2(n12677), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15847), .ZN(n12635) );
  NOR2_X1 U14997 ( .A1(n12970), .A2(n12668), .ZN(n12634) );
  AOI211_X1 U14998 ( .C1(n12975), .C2(n12666), .A(n12635), .B(n12634), .ZN(
        n12637) );
  NAND2_X1 U14999 ( .A1(n12974), .A2(n12670), .ZN(n12636) );
  OAI211_X1 U15000 ( .C1(n12638), .C2(n12672), .A(n12637), .B(n12636), .ZN(
        P3_U3169) );
  OAI211_X1 U15001 ( .C1(n12641), .C2(n12640), .A(n12639), .B(n7432), .ZN(
        n12646) );
  AOI22_X1 U15002 ( .A1(n12648), .A2(n12681), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12643) );
  NAND2_X1 U15003 ( .A1(n12666), .A2(n13024), .ZN(n12642) );
  OAI211_X1 U15004 ( .C1(n13051), .C2(n12677), .A(n12643), .B(n12642), .ZN(
        n12644) );
  AOI21_X1 U15005 ( .B1(n13019), .B2(n12670), .A(n12644), .ZN(n12645) );
  NAND2_X1 U15006 ( .A1(n12646), .A2(n12645), .ZN(P3_U3173) );
  XNOR2_X1 U15007 ( .A(n12647), .B(n12985), .ZN(n12653) );
  AOI22_X1 U15008 ( .A1(n12648), .A2(n12657), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12650) );
  NAND2_X1 U15009 ( .A1(n13000), .A2(n12666), .ZN(n12649) );
  OAI211_X1 U15010 ( .C1(n12997), .C2(n12668), .A(n12650), .B(n12649), .ZN(
        n12651) );
  AOI21_X1 U15011 ( .B1(n12889), .B2(n12670), .A(n12651), .ZN(n12652) );
  OAI21_X1 U15012 ( .B1(n12653), .B2(n12672), .A(n12652), .ZN(P3_U3175) );
  XNOR2_X1 U15013 ( .A(n12655), .B(n12654), .ZN(n12662) );
  NAND2_X1 U15014 ( .A1(n12657), .A2(n12656), .ZN(n12658) );
  NAND2_X1 U15015 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12812)
         );
  OAI211_X1 U15016 ( .C1(n13051), .C2(n12668), .A(n12658), .B(n12812), .ZN(
        n12659) );
  AOI21_X1 U15017 ( .B1(n13052), .B2(n12666), .A(n12659), .ZN(n12661) );
  NAND2_X1 U15018 ( .A1(n13163), .A2(n12670), .ZN(n12660) );
  OAI211_X1 U15019 ( .C1(n12662), .C2(n12672), .A(n12661), .B(n12660), .ZN(
        P3_U3178) );
  XOR2_X1 U15020 ( .A(n12664), .B(n12663), .Z(n12673) );
  OAI22_X1 U15021 ( .A1(n12970), .A2(n12677), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15812), .ZN(n12665) );
  AOI21_X1 U15022 ( .B1(n12947), .B2(n12666), .A(n12665), .ZN(n12667) );
  OAI21_X1 U15023 ( .B1(n12943), .B2(n12668), .A(n12667), .ZN(n12669) );
  AOI21_X1 U15024 ( .B1(n13125), .B2(n12670), .A(n12669), .ZN(n12671) );
  OAI21_X1 U15025 ( .B1(n12673), .B2(n12672), .A(n12671), .ZN(P3_U3180) );
  OAI211_X1 U15026 ( .C1(n12676), .C2(n12675), .A(n12674), .B(n7432), .ZN(
        n12683) );
  NAND2_X1 U15027 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12740)
         );
  OAI21_X1 U15028 ( .B1(n12872), .B2(n12677), .A(n12740), .ZN(n12680) );
  NOR2_X1 U15029 ( .A1(n12678), .A2(n13101), .ZN(n12679) );
  AOI211_X1 U15030 ( .C1(n12681), .C2(n13094), .A(n12680), .B(n12679), .ZN(
        n12682) );
  OAI211_X1 U15031 ( .C1(n12684), .C2(n13178), .A(n12683), .B(n12682), .ZN(
        P3_U3181) );
  AND3_X1 U15032 ( .A1(n12687), .A2(n12686), .A3(n12685), .ZN(n12688) );
  OAI21_X1 U15033 ( .B1(n12689), .B2(n12688), .A(n12853), .ZN(n12708) );
  INV_X1 U15034 ( .A(n12690), .ZN(n12692) );
  NAND3_X1 U15035 ( .A1(n12693), .A2(n12692), .A3(n12691), .ZN(n12694) );
  AOI21_X1 U15036 ( .B1(n12695), .B2(n12694), .A(n12855), .ZN(n12696) );
  AOI211_X1 U15037 ( .C1(n15392), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n12697), .B(
        n12696), .ZN(n12707) );
  NAND2_X1 U15038 ( .A1(n12822), .A2(n12698), .ZN(n12706) );
  INV_X1 U15039 ( .A(n12699), .ZN(n12700) );
  NOR3_X1 U15040 ( .A1(n6719), .A2(n12701), .A3(n12700), .ZN(n12703) );
  OAI21_X1 U15041 ( .B1(n12704), .B2(n12703), .A(n12702), .ZN(n12705) );
  NAND4_X1 U15042 ( .A1(n12708), .A2(n12707), .A3(n12706), .A4(n12705), .ZN(
        P3_U3186) );
  NOR2_X1 U15043 ( .A1(n7101), .A2(n12709), .ZN(n12711) );
  NAND2_X1 U15044 ( .A1(n12729), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12741) );
  OR2_X1 U15045 ( .A1(n12729), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12712) );
  NAND2_X1 U15046 ( .A1(n12741), .A2(n12712), .ZN(n12717) );
  AOI21_X1 U15047 ( .B1(n12713), .B2(n12717), .A(n12736), .ZN(n12735) );
  NOR2_X1 U15048 ( .A1(n12715), .A2(n12714), .ZN(n12719) );
  NAND2_X1 U15049 ( .A1(n12729), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12753) );
  OR2_X1 U15050 ( .A1(n12729), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12716) );
  NAND2_X1 U15051 ( .A1(n12753), .A2(n12716), .ZN(n12724) );
  MUX2_X1 U15052 ( .A(n12724), .B(n12717), .S(n12814), .Z(n12718) );
  NOR2_X1 U15053 ( .A1(n12745), .A2(n12819), .ZN(n12733) );
  OAI21_X1 U15054 ( .B1(n12720), .B2(n12719), .A(n12718), .ZN(n12732) );
  NOR2_X1 U15055 ( .A1(n7101), .A2(n12721), .ZN(n12723) );
  AOI21_X1 U15056 ( .B1(n12725), .B2(n12724), .A(n12751), .ZN(n12726) );
  NOR2_X1 U15057 ( .A1(n12726), .A2(n12847), .ZN(n12731) );
  AOI21_X1 U15058 ( .B1(n15392), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12727), 
        .ZN(n12728) );
  OAI21_X1 U15059 ( .B1(n12851), .B2(n12729), .A(n12728), .ZN(n12730) );
  AOI211_X1 U15060 ( .C1(n12733), .C2(n12732), .A(n12731), .B(n12730), .ZN(
        n12734) );
  OAI21_X1 U15061 ( .B1(n12735), .B2(n12855), .A(n12734), .ZN(P3_U3196) );
  NAND2_X1 U15062 ( .A1(n12741), .A2(n12737), .ZN(n12760) );
  AOI21_X1 U15063 ( .B1(n12739), .B2(n12738), .A(n12761), .ZN(n12759) );
  INV_X1 U15064 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14743) );
  OAI21_X1 U15065 ( .B1(n12813), .B2(n14743), .A(n12740), .ZN(n12750) );
  INV_X1 U15066 ( .A(n12753), .ZN(n12743) );
  INV_X1 U15067 ( .A(n12741), .ZN(n12742) );
  MUX2_X1 U15068 ( .A(n12743), .B(n12742), .S(n12814), .Z(n12744) );
  MUX2_X1 U15069 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12814), .Z(n12746) );
  NOR2_X1 U15070 ( .A1(n12747), .A2(n12746), .ZN(n12766) );
  AOI21_X1 U15071 ( .B1(n12747), .B2(n12746), .A(n12766), .ZN(n12748) );
  NOR2_X1 U15072 ( .A1(n12748), .A2(n12819), .ZN(n12749) );
  AOI211_X1 U15073 ( .C1(n12822), .C2(n7038), .A(n12750), .B(n12749), .ZN(
        n12758) );
  NAND2_X1 U15074 ( .A1(n12753), .A2(n12752), .ZN(n12774) );
  XNOR2_X1 U15075 ( .A(n12775), .B(n12774), .ZN(n12754) );
  AOI21_X1 U15076 ( .B1(n12755), .B2(n12754), .A(n12776), .ZN(n12756) );
  OR2_X1 U15077 ( .A1(n12756), .A2(n12847), .ZN(n12757) );
  OAI211_X1 U15078 ( .C1(n12759), .C2(n12855), .A(n12758), .B(n12757), .ZN(
        P3_U3197) );
  XNOR2_X1 U15079 ( .A(n12778), .B(n12768), .ZN(n12765) );
  AND2_X1 U15080 ( .A1(n12775), .A2(n12760), .ZN(n12762) );
  INV_X1 U15081 ( .A(n12790), .ZN(n12763) );
  AOI21_X1 U15082 ( .B1(n12765), .B2(n12764), .A(n12763), .ZN(n12788) );
  MUX2_X1 U15083 ( .A(n13083), .B(n12768), .S(n12814), .Z(n12769) );
  NOR2_X1 U15084 ( .A1(n12769), .A2(n12778), .ZN(n12801) );
  INV_X1 U15085 ( .A(n12801), .ZN(n12770) );
  NAND2_X1 U15086 ( .A1(n12769), .A2(n12778), .ZN(n12800) );
  NAND2_X1 U15087 ( .A1(n12770), .A2(n12800), .ZN(n12771) );
  XNOR2_X1 U15088 ( .A(n12802), .B(n12771), .ZN(n12786) );
  INV_X1 U15089 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14794) );
  NAND2_X1 U15090 ( .A1(n12822), .A2(n12778), .ZN(n12773) );
  OAI211_X1 U15091 ( .C1(n14794), .C2(n12813), .A(n12773), .B(n12772), .ZN(
        n12785) );
  AND2_X1 U15092 ( .A1(n12775), .A2(n12774), .ZN(n12777) );
  NAND2_X1 U15093 ( .A1(n12793), .A2(n13083), .ZN(n12780) );
  NAND2_X1 U15094 ( .A1(n12778), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12779) );
  AND2_X1 U15095 ( .A1(n12780), .A2(n12779), .ZN(n12781) );
  NAND2_X1 U15096 ( .A1(n12782), .A2(n12781), .ZN(n12783) );
  AOI21_X1 U15097 ( .B1(n12795), .B2(n12783), .A(n12847), .ZN(n12784) );
  AOI211_X1 U15098 ( .C1(n12786), .C2(n12853), .A(n12785), .B(n12784), .ZN(
        n12787) );
  OAI21_X1 U15099 ( .B1(n12788), .B2(n12855), .A(n12787), .ZN(P3_U3198) );
  NAND2_X1 U15100 ( .A1(n12793), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12789) );
  AOI21_X1 U15101 ( .B1(n12792), .B2(n12791), .A(n12809), .ZN(n12808) );
  NAND2_X1 U15102 ( .A1(n12793), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12794) );
  INV_X1 U15103 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14738) );
  OR2_X1 U15104 ( .A1(n12813), .A2(n14738), .ZN(n12797) );
  OAI211_X1 U15105 ( .C1(n12847), .C2(n12799), .A(n12798), .B(n12797), .ZN(
        n12806) );
  MUX2_X1 U15106 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12814), .Z(n12816) );
  XNOR2_X1 U15107 ( .A(n12816), .B(n12824), .ZN(n12804) );
  AOI211_X1 U15108 ( .C1(n12804), .C2(n12803), .A(n12819), .B(n12815), .ZN(
        n12805) );
  NAND2_X1 U15109 ( .A1(n12826), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12833) );
  OAI21_X1 U15110 ( .B1(n12826), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12833), 
        .ZN(n12811) );
  AOI21_X1 U15111 ( .B1(n6806), .B2(n12811), .A(n12835), .ZN(n12832) );
  INV_X1 U15112 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15536) );
  OAI21_X1 U15113 ( .B1(n12813), .B2(n15536), .A(n12812), .ZN(n12821) );
  MUX2_X1 U15114 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12814), .Z(n12818) );
  XNOR2_X1 U15115 ( .A(n12839), .B(n12838), .ZN(n12817) );
  NOR2_X1 U15116 ( .A1(n12817), .A2(n12818), .ZN(n12837) );
  AOI211_X1 U15117 ( .C1(n12822), .C2(n12838), .A(n12821), .B(n12820), .ZN(
        n12831) );
  NAND2_X1 U15118 ( .A1(n12826), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12844) );
  OAI21_X1 U15119 ( .B1(n12826), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12844), 
        .ZN(n12827) );
  AOI21_X1 U15120 ( .B1(n12828), .B2(n12827), .A(n12845), .ZN(n12829) );
  OR2_X1 U15121 ( .A1(n12829), .A2(n12847), .ZN(n12830) );
  OAI211_X1 U15122 ( .C1(n12832), .C2(n12855), .A(n12831), .B(n12830), .ZN(
        P3_U3200) );
  XNOR2_X1 U15123 ( .A(n12850), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12841) );
  INV_X1 U15124 ( .A(n12833), .ZN(n12834) );
  XOR2_X1 U15125 ( .A(n12841), .B(n12836), .Z(n12856) );
  XNOR2_X1 U15126 ( .A(n12850), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12846) );
  MUX2_X1 U15127 ( .A(n12841), .B(n12846), .S(n12840), .Z(n12842) );
  XNOR2_X1 U15128 ( .A(n12843), .B(n12842), .ZN(n12854) );
  NAND2_X1 U15129 ( .A1(n15392), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12848) );
  OAI211_X1 U15130 ( .C1(n12851), .C2(n12850), .A(n12849), .B(n12848), .ZN(
        n12852) );
  NAND2_X1 U15131 ( .A1(n13183), .A2(n13085), .ZN(n12861) );
  INV_X1 U15132 ( .A(P3_B_REG_SCAN_IN), .ZN(n15825) );
  NOR2_X1 U15133 ( .A1(n12857), .A2(n15825), .ZN(n12858) );
  NOR2_X1 U15134 ( .A1(n15450), .A2(n12858), .ZN(n12906) );
  NOR2_X1 U15135 ( .A1(n12860), .A2(n15458), .ZN(n12912) );
  AOI21_X1 U15136 ( .B1(n13184), .B2(n15463), .A(n12912), .ZN(n12864) );
  OAI211_X1 U15137 ( .C1(n15463), .C2(n12862), .A(n12861), .B(n12864), .ZN(
        P3_U3202) );
  NAND2_X1 U15138 ( .A1(n15465), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12863) );
  OAI211_X1 U15139 ( .C1(n13189), .C2(n13104), .A(n12864), .B(n12863), .ZN(
        P3_U3203) );
  NAND2_X1 U15140 ( .A1(n12867), .A2(n12866), .ZN(n12868) );
  OR2_X1 U15141 ( .A1(n14838), .A2(n12872), .ZN(n12873) );
  NAND2_X1 U15142 ( .A1(n13178), .A2(n13078), .ZN(n12875) );
  NAND2_X1 U15143 ( .A1(n13174), .A2(n13094), .ZN(n12877) );
  OR2_X1 U15144 ( .A1(n13171), .A2(n13077), .ZN(n12879) );
  NAND2_X1 U15145 ( .A1(n12882), .A2(n12881), .ZN(n13041) );
  NAND2_X1 U15146 ( .A1(n13157), .A2(n12883), .ZN(n12884) );
  NAND2_X1 U15147 ( .A1(n13019), .A2(n12885), .ZN(n12886) );
  NOR2_X1 U15148 ( .A1(n12889), .A2(n12985), .ZN(n12890) );
  INV_X1 U15149 ( .A(n12889), .ZN(n13213) );
  NAND2_X1 U15150 ( .A1(n13139), .A2(n12892), .ZN(n12893) );
  AND2_X1 U15151 ( .A1(n12974), .A2(n12986), .ZN(n12896) );
  OR2_X1 U15152 ( .A1(n12974), .A2(n12986), .ZN(n12895) );
  OR2_X1 U15153 ( .A1(n13125), .A2(n12898), .ZN(n12900) );
  AND2_X1 U15154 ( .A1(n13125), .A2(n12898), .ZN(n12899) );
  OR2_X1 U15155 ( .A1(n12933), .A2(n12901), .ZN(n12902) );
  XNOR2_X1 U15156 ( .A(n12904), .B(n12903), .ZN(n12905) );
  AOI22_X1 U15157 ( .A1(n12908), .A2(n15447), .B1(n12907), .B2(n12906), .ZN(
        n12909) );
  NAND2_X1 U15158 ( .A1(n13114), .A2(n15463), .ZN(n12914) );
  INV_X1 U15159 ( .A(n12910), .ZN(n13116) );
  NOR2_X1 U15160 ( .A1(n13116), .A2(n13104), .ZN(n12911) );
  AOI211_X1 U15161 ( .C1(n15465), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12912), 
        .B(n12911), .ZN(n12913) );
  OAI211_X1 U15162 ( .C1(n13117), .C2(n15460), .A(n12914), .B(n12913), .ZN(
        P3_U3204) );
  OAI22_X1 U15163 ( .A1(n12916), .A2(n15450), .B1(n12943), .B2(n15425), .ZN(
        n12917) );
  XNOR2_X1 U15164 ( .A(n12920), .B(n7775), .ZN(n13121) );
  AOI22_X1 U15165 ( .A1(n12921), .A2(n15442), .B1(n15465), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12923) );
  NAND2_X1 U15166 ( .A1(n13118), .A2(n13085), .ZN(n12922) );
  OAI211_X1 U15167 ( .C1(n13121), .C2(n15460), .A(n12923), .B(n12922), .ZN(
        n12924) );
  INV_X1 U15168 ( .A(n12924), .ZN(n12925) );
  OAI21_X1 U15169 ( .B1(n13120), .B2(n15465), .A(n12925), .ZN(P3_U3205) );
  OAI21_X1 U15170 ( .B1(n12929), .B2(n12928), .A(n12927), .ZN(n12932) );
  OAI22_X1 U15171 ( .A1(n12930), .A2(n15450), .B1(n12956), .B2(n15425), .ZN(
        n12931) );
  INV_X1 U15172 ( .A(n13123), .ZN(n12938) );
  INV_X1 U15173 ( .A(n12933), .ZN(n13193) );
  AOI22_X1 U15174 ( .A1(n12934), .A2(n15442), .B1(n15465), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12935) );
  OAI21_X1 U15175 ( .B1(n13193), .B2(n13104), .A(n12935), .ZN(n12936) );
  AOI21_X1 U15176 ( .B1(n6665), .B2(n12978), .A(n12936), .ZN(n12937) );
  OAI21_X1 U15177 ( .B1(n12938), .B2(n15465), .A(n12937), .ZN(P3_U3206) );
  XNOR2_X1 U15178 ( .A(n12940), .B(n12939), .ZN(n13126) );
  XNOR2_X1 U15179 ( .A(n12942), .B(n12941), .ZN(n12945) );
  OAI22_X1 U15180 ( .A1(n12943), .A2(n15450), .B1(n12970), .B2(n15425), .ZN(
        n12944) );
  AOI21_X1 U15181 ( .B1(n12945), .B2(n15453), .A(n12944), .ZN(n12946) );
  OAI21_X1 U15182 ( .B1(n15416), .B2(n13126), .A(n12946), .ZN(n13127) );
  AOI22_X1 U15183 ( .A1(n12947), .A2(n15442), .B1(P3_REG2_REG_26__SCAN_IN), 
        .B2(n15465), .ZN(n12949) );
  NAND2_X1 U15184 ( .A1(n13125), .A2(n13085), .ZN(n12948) );
  OAI211_X1 U15185 ( .C1(n13126), .C2(n12992), .A(n12949), .B(n12948), .ZN(
        n12950) );
  AOI21_X1 U15186 ( .B1(n13127), .B2(n15463), .A(n12950), .ZN(n12951) );
  INV_X1 U15187 ( .A(n12951), .ZN(P3_U3207) );
  INV_X1 U15188 ( .A(n12958), .ZN(n12953) );
  OAI211_X1 U15189 ( .C1(n12953), .C2(n6789), .A(n12952), .B(n15453), .ZN(
        n12955) );
  NAND2_X1 U15190 ( .A1(n12986), .A2(n15447), .ZN(n12954) );
  OAI211_X1 U15191 ( .C1(n12956), .C2(n15450), .A(n12955), .B(n12954), .ZN(
        n13131) );
  INV_X1 U15192 ( .A(n13131), .ZN(n12965) );
  OAI21_X1 U15193 ( .B1(n12959), .B2(n12958), .A(n12957), .ZN(n13132) );
  INV_X1 U15194 ( .A(n12960), .ZN(n13201) );
  AOI22_X1 U15195 ( .A1(n12961), .A2(n15442), .B1(n15465), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12962) );
  OAI21_X1 U15196 ( .B1(n13201), .B2(n13104), .A(n12962), .ZN(n12963) );
  AOI21_X1 U15197 ( .B1(n13132), .B2(n14864), .A(n12963), .ZN(n12964) );
  OAI21_X1 U15198 ( .B1(n12965), .B2(n15465), .A(n12964), .ZN(P3_U3208) );
  XNOR2_X1 U15199 ( .A(n12967), .B(n12966), .ZN(n12973) );
  OAI21_X1 U15200 ( .B1(n12969), .B2(n9063), .A(n12968), .ZN(n13136) );
  OAI22_X1 U15201 ( .A1(n12970), .A2(n15450), .B1(n12997), .B2(n15425), .ZN(
        n12971) );
  AOI21_X1 U15202 ( .B1(n13136), .B2(n15435), .A(n12971), .ZN(n12972) );
  OAI21_X1 U15203 ( .B1(n12973), .B2(n15430), .A(n12972), .ZN(n13135) );
  INV_X1 U15204 ( .A(n13135), .ZN(n12980) );
  INV_X1 U15205 ( .A(n12974), .ZN(n13205) );
  AOI22_X1 U15206 ( .A1(n12975), .A2(n15442), .B1(n15465), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12976) );
  OAI21_X1 U15207 ( .B1(n13205), .B2(n13104), .A(n12976), .ZN(n12977) );
  AOI21_X1 U15208 ( .B1(n13136), .B2(n12978), .A(n12977), .ZN(n12979) );
  OAI21_X1 U15209 ( .B1(n12980), .B2(n15465), .A(n12979), .ZN(P3_U3209) );
  XNOR2_X1 U15210 ( .A(n12981), .B(n12982), .ZN(n13140) );
  XNOR2_X1 U15211 ( .A(n12983), .B(n12982), .ZN(n12984) );
  NAND2_X1 U15212 ( .A1(n12984), .A2(n15453), .ZN(n12988) );
  AOI22_X1 U15213 ( .A1(n12986), .A2(n15398), .B1(n15447), .B2(n12985), .ZN(
        n12987) );
  OAI211_X1 U15214 ( .C1(n15416), .C2(n13140), .A(n12988), .B(n12987), .ZN(
        n13141) );
  AOI22_X1 U15215 ( .A1(n12989), .A2(n15442), .B1(n15465), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U15216 ( .A1(n13139), .A2(n13085), .ZN(n12990) );
  OAI211_X1 U15217 ( .C1(n13140), .C2(n12992), .A(n12991), .B(n12990), .ZN(
        n12993) );
  AOI21_X1 U15218 ( .B1(n13141), .B2(n15463), .A(n12993), .ZN(n12994) );
  INV_X1 U15219 ( .A(n12994), .ZN(P3_U3210) );
  XOR2_X1 U15220 ( .A(n12995), .B(n12999), .Z(n12996) );
  OAI222_X1 U15221 ( .A1(n15450), .A2(n12997), .B1(n15425), .B2(n13018), .C1(
        n15430), .C2(n12996), .ZN(n13145) );
  INV_X1 U15222 ( .A(n13145), .ZN(n13004) );
  XOR2_X1 U15223 ( .A(n12998), .B(n12999), .Z(n13146) );
  AOI22_X1 U15224 ( .A1(n13000), .A2(n15442), .B1(n15465), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n13001) );
  OAI21_X1 U15225 ( .B1(n13213), .B2(n13104), .A(n13001), .ZN(n13002) );
  AOI21_X1 U15226 ( .B1(n13146), .B2(n14864), .A(n13002), .ZN(n13003) );
  OAI21_X1 U15227 ( .B1(n13004), .B2(n15465), .A(n13003), .ZN(P3_U3211) );
  XNOR2_X1 U15228 ( .A(n13005), .B(n13008), .ZN(n13006) );
  OAI222_X1 U15229 ( .A1(n15450), .A2(n13007), .B1(n15425), .B2(n13031), .C1(
        n15430), .C2(n13006), .ZN(n13149) );
  INV_X1 U15230 ( .A(n13149), .ZN(n13015) );
  XNOR2_X1 U15231 ( .A(n13009), .B(n13008), .ZN(n13150) );
  INV_X1 U15232 ( .A(n13010), .ZN(n13217) );
  AOI22_X1 U15233 ( .A1(n15465), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13011), 
        .B2(n15442), .ZN(n13012) );
  OAI21_X1 U15234 ( .B1(n13217), .B2(n13104), .A(n13012), .ZN(n13013) );
  AOI21_X1 U15235 ( .B1(n13150), .B2(n14864), .A(n13013), .ZN(n13014) );
  OAI21_X1 U15236 ( .B1(n13015), .B2(n15465), .A(n13014), .ZN(P3_U3212) );
  XNOR2_X1 U15237 ( .A(n13016), .B(n13020), .ZN(n13017) );
  OAI222_X1 U15238 ( .A1(n15450), .A2(n13018), .B1(n15425), .B2(n13051), .C1(
        n15430), .C2(n13017), .ZN(n13153) );
  INV_X1 U15239 ( .A(n13019), .ZN(n13221) );
  NAND2_X1 U15240 ( .A1(n13021), .A2(n13020), .ZN(n13022) );
  AND2_X1 U15241 ( .A1(n13023), .A2(n13022), .ZN(n13154) );
  NAND2_X1 U15242 ( .A1(n13154), .A2(n14864), .ZN(n13026) );
  AOI22_X1 U15243 ( .A1(n15465), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15442), 
        .B2(n13024), .ZN(n13025) );
  OAI211_X1 U15244 ( .C1(n13221), .C2(n13104), .A(n13026), .B(n13025), .ZN(
        n13027) );
  AOI21_X1 U15245 ( .B1(n13153), .B2(n15463), .A(n13027), .ZN(n13028) );
  INV_X1 U15246 ( .A(n13028), .ZN(P3_U3213) );
  OAI211_X1 U15247 ( .C1(n13030), .C2(n13041), .A(n13029), .B(n15453), .ZN(
        n13034) );
  OAI22_X1 U15248 ( .A1(n13031), .A2(n15450), .B1(n13061), .B2(n15425), .ZN(
        n13032) );
  INV_X1 U15249 ( .A(n13032), .ZN(n13033) );
  AND2_X1 U15250 ( .A1(n13034), .A2(n13033), .ZN(n13160) );
  INV_X1 U15251 ( .A(n13035), .ZN(n13036) );
  OAI22_X1 U15252 ( .A1(n15463), .A2(n13037), .B1(n13036), .B2(n15458), .ZN(
        n13038) );
  AOI21_X1 U15253 ( .B1(n13157), .B2(n13085), .A(n13038), .ZN(n13044) );
  NAND2_X1 U15254 ( .A1(n13039), .A2(n13040), .ZN(n13042) );
  XNOR2_X1 U15255 ( .A(n13042), .B(n13041), .ZN(n13158) );
  NAND2_X1 U15256 ( .A1(n13158), .A2(n14864), .ZN(n13043) );
  OAI211_X1 U15257 ( .C1(n13160), .C2(n15465), .A(n13044), .B(n13043), .ZN(
        P3_U3214) );
  NAND2_X1 U15258 ( .A1(n13045), .A2(n7332), .ZN(n13046) );
  AND2_X1 U15259 ( .A1(n13039), .A2(n13046), .ZN(n13165) );
  INV_X1 U15260 ( .A(n13165), .ZN(n13058) );
  AOI21_X1 U15261 ( .B1(n13049), .B2(n13048), .A(n13047), .ZN(n13050) );
  OAI222_X1 U15262 ( .A1(n15450), .A2(n13051), .B1(n15425), .B2(n13077), .C1(
        n15430), .C2(n13050), .ZN(n13164) );
  NAND2_X1 U15263 ( .A1(n13164), .A2(n15463), .ZN(n13057) );
  INV_X1 U15264 ( .A(n13052), .ZN(n13053) );
  OAI22_X1 U15265 ( .A1(n15463), .A2(n13054), .B1(n13053), .B2(n15458), .ZN(
        n13055) );
  AOI21_X1 U15266 ( .B1(n13163), .B2(n13085), .A(n13055), .ZN(n13056) );
  OAI211_X1 U15267 ( .C1(n15460), .C2(n13058), .A(n13057), .B(n13056), .ZN(
        P3_U3215) );
  XNOR2_X1 U15268 ( .A(n13059), .B(n13066), .ZN(n13060) );
  NAND2_X1 U15269 ( .A1(n13060), .A2(n15453), .ZN(n13065) );
  OAI22_X1 U15270 ( .A1(n13062), .A2(n15425), .B1(n13061), .B2(n15450), .ZN(
        n13063) );
  INV_X1 U15271 ( .A(n13063), .ZN(n13064) );
  NAND2_X1 U15272 ( .A1(n13065), .A2(n13064), .ZN(n13173) );
  INV_X1 U15273 ( .A(n13173), .ZN(n13075) );
  OR2_X1 U15274 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  NAND2_X1 U15275 ( .A1(n13069), .A2(n13068), .ZN(n13169) );
  NOR2_X1 U15276 ( .A1(n13171), .A2(n13104), .ZN(n13073) );
  OAI22_X1 U15277 ( .A1(n15463), .A2(n13071), .B1(n13070), .B2(n15458), .ZN(
        n13072) );
  AOI211_X1 U15278 ( .C1(n13169), .C2(n14864), .A(n13073), .B(n13072), .ZN(
        n13074) );
  OAI21_X1 U15279 ( .B1(n13075), .B2(n15465), .A(n13074), .ZN(P3_U3216) );
  AOI21_X1 U15280 ( .B1(n13076), .B2(n13087), .A(n15430), .ZN(n13081) );
  OAI22_X1 U15281 ( .A1(n13078), .A2(n15425), .B1(n13077), .B2(n15450), .ZN(
        n13079) );
  AOI21_X1 U15282 ( .B1(n13081), .B2(n13080), .A(n13079), .ZN(n13177) );
  OAI22_X1 U15283 ( .A1(n15463), .A2(n13083), .B1(n13082), .B2(n15458), .ZN(
        n13084) );
  AOI21_X1 U15284 ( .B1(n13174), .B2(n13085), .A(n13084), .ZN(n13090) );
  OAI21_X1 U15285 ( .B1(n13088), .B2(n13087), .A(n13086), .ZN(n13175) );
  NAND2_X1 U15286 ( .A1(n13175), .A2(n14864), .ZN(n13089) );
  OAI211_X1 U15287 ( .C1(n13177), .C2(n15465), .A(n13090), .B(n13089), .ZN(
        P3_U3217) );
  NAND2_X1 U15288 ( .A1(n13091), .A2(n13097), .ZN(n13092) );
  NAND2_X1 U15289 ( .A1(n6821), .A2(n13092), .ZN(n13093) );
  NAND2_X1 U15290 ( .A1(n13093), .A2(n15453), .ZN(n13096) );
  AOI22_X1 U15291 ( .A1(n13094), .A2(n15398), .B1(n15447), .B2(n14843), .ZN(
        n13095) );
  NAND2_X1 U15292 ( .A1(n13096), .A2(n13095), .ZN(n13182) );
  INV_X1 U15293 ( .A(n13182), .ZN(n13107) );
  OR2_X1 U15294 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  NAND2_X1 U15295 ( .A1(n13100), .A2(n13099), .ZN(n13179) );
  INV_X1 U15296 ( .A(n13101), .ZN(n13102) );
  AOI22_X1 U15297 ( .A1(n15465), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15442), 
        .B2(n13102), .ZN(n13103) );
  OAI21_X1 U15298 ( .B1(n13178), .B2(n13104), .A(n13103), .ZN(n13105) );
  AOI21_X1 U15299 ( .B1(n13179), .B2(n14864), .A(n13105), .ZN(n13106) );
  OAI21_X1 U15300 ( .B1(n13107), .B2(n15465), .A(n13106), .ZN(P3_U3218) );
  INV_X1 U15301 ( .A(n13168), .ZN(n13110) );
  NAND2_X1 U15302 ( .A1(n13183), .A2(n13110), .ZN(n13108) );
  NAND2_X1 U15303 ( .A1(n13184), .A2(n15532), .ZN(n13112) );
  OAI211_X1 U15304 ( .C1(n15532), .C2(n13109), .A(n13108), .B(n13112), .ZN(
        P3_U3490) );
  NAND2_X1 U15305 ( .A1(n13111), .A2(n13110), .ZN(n13113) );
  OAI211_X1 U15306 ( .C1(n15532), .C2(n9155), .A(n13113), .B(n13112), .ZN(
        P3_U3489) );
  OR2_X1 U15307 ( .A1(n15438), .A2(n13115), .ZN(n13122) );
  NAND2_X1 U15308 ( .A1(n13118), .A2(n15495), .ZN(n13119) );
  INV_X1 U15309 ( .A(n13125), .ZN(n13197) );
  INV_X1 U15310 ( .A(n13126), .ZN(n13128) );
  AOI21_X1 U15311 ( .B1(n15509), .B2(n13128), .A(n13127), .ZN(n13194) );
  MUX2_X1 U15312 ( .A(n13129), .B(n13194), .S(n15532), .Z(n13130) );
  OAI21_X1 U15313 ( .B1(n13197), .B2(n13168), .A(n13130), .ZN(P3_U3485) );
  AOI21_X1 U15314 ( .B1(n15515), .B2(n13132), .A(n13131), .ZN(n13198) );
  MUX2_X1 U15315 ( .A(n13133), .B(n13198), .S(n15532), .Z(n13134) );
  OAI21_X1 U15316 ( .B1(n13201), .B2(n13168), .A(n13134), .ZN(P3_U3484) );
  AOI21_X1 U15317 ( .B1(n15509), .B2(n13136), .A(n13135), .ZN(n13202) );
  MUX2_X1 U15318 ( .A(n13137), .B(n13202), .S(n15532), .Z(n13138) );
  OAI21_X1 U15319 ( .B1(n13205), .B2(n13168), .A(n13138), .ZN(P3_U3483) );
  INV_X1 U15320 ( .A(n13139), .ZN(n13209) );
  INV_X1 U15321 ( .A(n13140), .ZN(n13142) );
  AOI21_X1 U15322 ( .B1(n15509), .B2(n13142), .A(n13141), .ZN(n13206) );
  MUX2_X1 U15323 ( .A(n13143), .B(n13206), .S(n15532), .Z(n13144) );
  OAI21_X1 U15324 ( .B1(n13209), .B2(n13168), .A(n13144), .ZN(P3_U3482) );
  AOI21_X1 U15325 ( .B1(n13146), .B2(n15515), .A(n13145), .ZN(n13210) );
  MUX2_X1 U15326 ( .A(n13147), .B(n13210), .S(n15532), .Z(n13148) );
  OAI21_X1 U15327 ( .B1(n13213), .B2(n13168), .A(n13148), .ZN(P3_U3481) );
  AOI21_X1 U15328 ( .B1(n13150), .B2(n15515), .A(n13149), .ZN(n13214) );
  MUX2_X1 U15329 ( .A(n13151), .B(n13214), .S(n15532), .Z(n13152) );
  OAI21_X1 U15330 ( .B1(n13217), .B2(n13168), .A(n13152), .ZN(P3_U3480) );
  INV_X1 U15331 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13155) );
  AOI21_X1 U15332 ( .B1(n13154), .B2(n15515), .A(n13153), .ZN(n13218) );
  MUX2_X1 U15333 ( .A(n13155), .B(n13218), .S(n15532), .Z(n13156) );
  OAI21_X1 U15334 ( .B1(n13221), .B2(n13168), .A(n13156), .ZN(P3_U3479) );
  INV_X1 U15335 ( .A(n13157), .ZN(n13225) );
  INV_X1 U15336 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U15337 ( .A1(n13158), .A2(n15515), .ZN(n13159) );
  AND2_X1 U15338 ( .A1(n13160), .A2(n13159), .ZN(n13223) );
  MUX2_X1 U15339 ( .A(n13161), .B(n13223), .S(n15532), .Z(n13162) );
  OAI21_X1 U15340 ( .B1(n13225), .B2(n13168), .A(n13162), .ZN(P3_U3478) );
  INV_X1 U15341 ( .A(n13163), .ZN(n13230) );
  AOI21_X1 U15342 ( .B1(n13165), .B2(n15515), .A(n13164), .ZN(n13226) );
  MUX2_X1 U15343 ( .A(n13166), .B(n13226), .S(n15532), .Z(n13167) );
  OAI21_X1 U15344 ( .B1(n13230), .B2(n13168), .A(n13167), .ZN(P3_U3477) );
  NAND2_X1 U15345 ( .A1(n13169), .A2(n15515), .ZN(n13170) );
  OAI21_X1 U15346 ( .B1(n15512), .B2(n13171), .A(n13170), .ZN(n13172) );
  MUX2_X1 U15347 ( .A(n13231), .B(P3_REG1_REG_17__SCAN_IN), .S(n15530), .Z(
        P3_U3476) );
  AOI22_X1 U15348 ( .A1(n13175), .A2(n15515), .B1(n15495), .B2(n13174), .ZN(
        n13176) );
  NAND2_X1 U15349 ( .A1(n13177), .A2(n13176), .ZN(n13232) );
  MUX2_X1 U15350 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13232), .S(n15532), .Z(
        P3_U3475) );
  NOR2_X1 U15351 ( .A1(n13178), .A2(n15512), .ZN(n13181) );
  AND2_X1 U15352 ( .A1(n13179), .A2(n15515), .ZN(n13180) );
  MUX2_X1 U15353 ( .A(n13233), .B(P3_REG1_REG_15__SCAN_IN), .S(n15530), .Z(
        P3_U3474) );
  INV_X1 U15354 ( .A(n13183), .ZN(n13186) );
  NAND2_X1 U15355 ( .A1(n13184), .A2(n15519), .ZN(n13187) );
  NAND2_X1 U15356 ( .A1(n15517), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13185) );
  OAI211_X1 U15357 ( .C1(n13186), .C2(n13229), .A(n13187), .B(n13185), .ZN(
        P3_U3458) );
  NAND2_X1 U15358 ( .A1(n15517), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13188) );
  OAI211_X1 U15359 ( .C1(n13189), .C2(n13229), .A(n13188), .B(n13187), .ZN(
        P3_U3457) );
  INV_X1 U15360 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13192) );
  INV_X1 U15361 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13195) );
  MUX2_X1 U15362 ( .A(n13195), .B(n13194), .S(n15519), .Z(n13196) );
  OAI21_X1 U15363 ( .B1(n13197), .B2(n13229), .A(n13196), .ZN(P3_U3453) );
  INV_X1 U15364 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13199) );
  MUX2_X1 U15365 ( .A(n13199), .B(n13198), .S(n15519), .Z(n13200) );
  OAI21_X1 U15366 ( .B1(n13201), .B2(n13229), .A(n13200), .ZN(P3_U3452) );
  INV_X1 U15367 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13203) );
  MUX2_X1 U15368 ( .A(n13203), .B(n13202), .S(n15519), .Z(n13204) );
  OAI21_X1 U15369 ( .B1(n13205), .B2(n13229), .A(n13204), .ZN(P3_U3451) );
  INV_X1 U15370 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13207) );
  MUX2_X1 U15371 ( .A(n13207), .B(n13206), .S(n15519), .Z(n13208) );
  OAI21_X1 U15372 ( .B1(n13209), .B2(n13229), .A(n13208), .ZN(P3_U3450) );
  INV_X1 U15373 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13211) );
  MUX2_X1 U15374 ( .A(n13211), .B(n13210), .S(n15519), .Z(n13212) );
  OAI21_X1 U15375 ( .B1(n13213), .B2(n13229), .A(n13212), .ZN(P3_U3449) );
  INV_X1 U15376 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13215) );
  MUX2_X1 U15377 ( .A(n13215), .B(n13214), .S(n15519), .Z(n13216) );
  OAI21_X1 U15378 ( .B1(n13217), .B2(n13229), .A(n13216), .ZN(P3_U3448) );
  INV_X1 U15379 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13219) );
  MUX2_X1 U15380 ( .A(n13219), .B(n13218), .S(n15519), .Z(n13220) );
  OAI21_X1 U15381 ( .B1(n13221), .B2(n13229), .A(n13220), .ZN(P3_U3447) );
  MUX2_X1 U15382 ( .A(n13223), .B(n13222), .S(n15517), .Z(n13224) );
  OAI21_X1 U15383 ( .B1(n13225), .B2(n13229), .A(n13224), .ZN(P3_U3446) );
  MUX2_X1 U15384 ( .A(n13227), .B(n13226), .S(n15519), .Z(n13228) );
  OAI21_X1 U15385 ( .B1(n13230), .B2(n13229), .A(n13228), .ZN(P3_U3444) );
  MUX2_X1 U15386 ( .A(n13231), .B(P3_REG0_REG_17__SCAN_IN), .S(n15517), .Z(
        P3_U3441) );
  MUX2_X1 U15387 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13232), .S(n15519), .Z(
        P3_U3438) );
  MUX2_X1 U15388 ( .A(n13233), .B(P3_REG0_REG_15__SCAN_IN), .S(n15517), .Z(
        P3_U3435) );
  MUX2_X1 U15389 ( .A(n13234), .B(P3_D_REG_1__SCAN_IN), .S(n13235), .Z(
        P3_U3377) );
  MUX2_X1 U15390 ( .A(n13236), .B(P3_D_REG_0__SCAN_IN), .S(n13235), .Z(
        P3_U3376) );
  INV_X1 U15391 ( .A(n13237), .ZN(n13242) );
  NOR4_X1 U15392 ( .A1(n13238), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), 
        .A4(n8645), .ZN(n13239) );
  AOI21_X1 U15393 ( .B1(n13240), .B2(SI_31_), .A(n13239), .ZN(n13241) );
  OAI21_X1 U15394 ( .B1(n13242), .B2(n6670), .A(n13241), .ZN(P3_U3264) );
  INV_X1 U15395 ( .A(n13244), .ZN(n13246) );
  OAI222_X1 U15396 ( .A1(n13243), .A2(P3_U3151), .B1(n6670), .B2(n13246), .C1(
        n13245), .C2(n13251), .ZN(P3_U3265) );
  INV_X1 U15397 ( .A(n13247), .ZN(n13250) );
  OAI222_X1 U15398 ( .A1(n13251), .A2(n15597), .B1(n6670), .B2(n13250), .C1(
        P3_U3151), .C2(n13248), .ZN(P3_U3266) );
  XNOR2_X1 U15399 ( .A(n13253), .B(n13252), .ZN(n13258) );
  AOI22_X1 U15400 ( .A1(n13538), .A2(n13336), .B1(n13307), .B2(n13569), .ZN(
        n13606) );
  NOR2_X1 U15401 ( .A1(n13606), .A2(n13339), .ZN(n13256) );
  OAI22_X1 U15402 ( .A1(n13604), .A2(n14911), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13254), .ZN(n13255) );
  AOI211_X1 U15403 ( .C1(n13764), .C2(n14908), .A(n13256), .B(n13255), .ZN(
        n13257) );
  OAI21_X1 U15404 ( .B1(n13258), .B2(n13342), .A(n13257), .ZN(P2_U3186) );
  XNOR2_X1 U15405 ( .A(n13260), .B(n13259), .ZN(n13262) );
  NAND3_X1 U15406 ( .A1(n13262), .A2(n14903), .A3(n13261), .ZN(n13270) );
  INV_X1 U15407 ( .A(n13262), .ZN(n13263) );
  INV_X1 U15408 ( .A(n13561), .ZN(n13529) );
  NAND3_X1 U15409 ( .A1(n13263), .A2(n13313), .A3(n13529), .ZN(n13269) );
  INV_X1 U15410 ( .A(n13559), .ZN(n13525) );
  OAI22_X1 U15411 ( .A1(n13288), .A2(n13326), .B1(n13525), .B2(n13544), .ZN(
        n13791) );
  INV_X1 U15412 ( .A(n13666), .ZN(n13265) );
  OAI22_X1 U15413 ( .A1(n13265), .A2(n14911), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13264), .ZN(n13266) );
  AOI21_X1 U15414 ( .B1(n13791), .B2(n14905), .A(n13266), .ZN(n13268) );
  NAND2_X1 U15415 ( .A1(n7237), .A2(n14908), .ZN(n13267) );
  NAND4_X1 U15416 ( .A1(n13270), .A2(n13269), .A3(n13268), .A4(n13267), .ZN(
        P2_U3188) );
  NAND2_X1 U15417 ( .A1(n13272), .A2(n13271), .ZN(n13274) );
  XOR2_X1 U15418 ( .A(n13274), .B(n13273), .Z(n13278) );
  OAI22_X1 U15419 ( .A1(n13556), .A2(n13326), .B1(n13553), .B2(n13544), .ZN(
        n13717) );
  NAND2_X1 U15420 ( .A1(n13717), .A2(n14905), .ZN(n13275) );
  NAND2_X1 U15421 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13495)
         );
  OAI211_X1 U15422 ( .C1(n14911), .C2(n13722), .A(n13275), .B(n13495), .ZN(
        n13276) );
  AOI21_X1 U15423 ( .B1(n13822), .B2(n14908), .A(n13276), .ZN(n13277) );
  OAI21_X1 U15424 ( .B1(n13278), .B2(n13342), .A(n13277), .ZN(P2_U3191) );
  XNOR2_X1 U15425 ( .A(n13280), .B(n13279), .ZN(n13285) );
  AOI22_X1 U15426 ( .A1(n13559), .A2(n13336), .B1(n13347), .B2(n13307), .ZN(
        n13807) );
  OAI22_X1 U15427 ( .A1(n13807), .A2(n13339), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13281), .ZN(n13283) );
  NOR2_X1 U15428 ( .A1(n13809), .A2(n13330), .ZN(n13282) );
  AOI211_X1 U15429 ( .C1(n13337), .C2(n13696), .A(n13283), .B(n13282), .ZN(
        n13284) );
  OAI21_X1 U15430 ( .B1(n13285), .B2(n13342), .A(n13284), .ZN(P2_U3195) );
  XNOR2_X1 U15431 ( .A(n13287), .B(n13286), .ZN(n13294) );
  OAI22_X1 U15432 ( .A1(n13571), .A2(n13326), .B1(n13288), .B2(n13544), .ZN(
        n13631) );
  INV_X1 U15433 ( .A(n13637), .ZN(n13290) );
  OAI22_X1 U15434 ( .A1(n13290), .A2(n14911), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13289), .ZN(n13291) );
  AOI21_X1 U15435 ( .B1(n13631), .B2(n14905), .A(n13291), .ZN(n13293) );
  NAND2_X1 U15436 ( .A1(n13858), .A2(n14908), .ZN(n13292) );
  OAI211_X1 U15437 ( .C1(n13294), .C2(n13342), .A(n13293), .B(n13292), .ZN(
        P2_U3197) );
  XNOR2_X1 U15438 ( .A(n13296), .B(n13295), .ZN(n13301) );
  OAI22_X1 U15439 ( .A1(n13567), .A2(n13326), .B1(n13561), .B2(n13544), .ZN(
        n13650) );
  OAI22_X1 U15440 ( .A1(n13655), .A2(n14911), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13297), .ZN(n13298) );
  AOI21_X1 U15441 ( .B1(n13650), .B2(n14905), .A(n13298), .ZN(n13300) );
  NAND2_X1 U15442 ( .A1(n13787), .A2(n14908), .ZN(n13299) );
  OAI211_X1 U15443 ( .C1(n13301), .C2(n13342), .A(n13300), .B(n13299), .ZN(
        P2_U3201) );
  INV_X1 U15444 ( .A(n13302), .ZN(n13303) );
  AOI21_X1 U15445 ( .B1(n13305), .B2(n13304), .A(n13303), .ZN(n13312) );
  NOR2_X1 U15446 ( .A1(n14911), .A2(n13306), .ZN(n13310) );
  AOI22_X1 U15447 ( .A1(n13557), .A2(n13336), .B1(n13307), .B2(n13517), .ZN(
        n13814) );
  OAI22_X1 U15448 ( .A1(n13814), .A2(n13339), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13308), .ZN(n13309) );
  AOI211_X1 U15449 ( .C1(n13711), .C2(n14908), .A(n13310), .B(n13309), .ZN(
        n13311) );
  OAI21_X1 U15450 ( .B1(n13312), .B2(n13342), .A(n13311), .ZN(P2_U3205) );
  NAND2_X1 U15451 ( .A1(n13559), .A2(n13313), .ZN(n13317) );
  OR2_X1 U15452 ( .A1(n13314), .A2(n13342), .ZN(n13316) );
  MUX2_X1 U15453 ( .A(n13317), .B(n13316), .S(n13315), .Z(n13321) );
  OAI22_X1 U15454 ( .A1(n13561), .A2(n13326), .B1(n13523), .B2(n13544), .ZN(
        n13801) );
  OAI22_X1 U15455 ( .A1(n13682), .A2(n14911), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13318), .ZN(n13319) );
  AOI21_X1 U15456 ( .B1(n13801), .B2(n14905), .A(n13319), .ZN(n13320) );
  OAI211_X1 U15457 ( .C1(n7236), .C2(n13330), .A(n13321), .B(n13320), .ZN(
        P2_U3207) );
  AOI21_X1 U15458 ( .B1(n13323), .B2(n13322), .A(n13342), .ZN(n13325) );
  NAND2_X1 U15459 ( .A1(n13325), .A2(n13324), .ZN(n13329) );
  OAI22_X1 U15460 ( .A1(n13555), .A2(n13326), .B1(n13549), .B2(n13544), .ZN(
        n13827) );
  AND2_X1 U15461 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15322) );
  NOR2_X1 U15462 ( .A1(n14911), .A2(n13738), .ZN(n13327) );
  AOI211_X1 U15463 ( .C1(n13827), .C2(n14905), .A(n15322), .B(n13327), .ZN(
        n13328) );
  OAI211_X1 U15464 ( .C1(n13744), .C2(n13330), .A(n13329), .B(n13328), .ZN(
        P2_U3210) );
  INV_X1 U15465 ( .A(n13331), .ZN(n13332) );
  AOI21_X1 U15466 ( .B1(n13334), .B2(n13333), .A(n13332), .ZN(n13343) );
  NOR2_X1 U15467 ( .A1(n13567), .A2(n13544), .ZN(n13335) );
  AOI21_X1 U15468 ( .B1(n13537), .B2(n13336), .A(n13335), .ZN(n13771) );
  AOI22_X1 U15469 ( .A1(n13622), .A2(n13337), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13338) );
  OAI21_X1 U15470 ( .B1(n13771), .B2(n13339), .A(n13338), .ZN(n13340) );
  AOI21_X1 U15471 ( .B1(n13854), .B2(n14908), .A(n13340), .ZN(n13341) );
  OAI21_X1 U15472 ( .B1(n13343), .B2(n13342), .A(n13341), .ZN(P2_U3212) );
  MUX2_X1 U15473 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13344), .S(P2_U3947), .Z(
        P2_U3562) );
  MUX2_X1 U15474 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13345), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15475 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13346), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15476 ( .A(n13538), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13356), .Z(
        P2_U3559) );
  MUX2_X1 U15477 ( .A(n13537), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13356), .Z(
        P2_U3558) );
  MUX2_X1 U15478 ( .A(n13569), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13356), .Z(
        P2_U3557) );
  MUX2_X1 U15479 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13532), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15480 ( .A(n13564), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13356), .Z(
        P2_U3555) );
  MUX2_X1 U15481 ( .A(n13529), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13356), .Z(
        P2_U3554) );
  MUX2_X1 U15482 ( .A(n13559), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13356), .Z(
        P2_U3553) );
  MUX2_X1 U15483 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13557), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15484 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13347), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15485 ( .A(n13517), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13356), .Z(
        P2_U3550) );
  MUX2_X1 U15486 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13513), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U15487 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13511), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U15488 ( .A(n13348), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13356), .Z(
        P2_U3547) );
  MUX2_X1 U15489 ( .A(n13349), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13356), .Z(
        P2_U3546) );
  MUX2_X1 U15490 ( .A(n13350), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13356), .Z(
        P2_U3545) );
  MUX2_X1 U15491 ( .A(n13351), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13356), .Z(
        P2_U3544) );
  MUX2_X1 U15492 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13352), .S(P2_U3947), .Z(
        P2_U3543) );
  MUX2_X1 U15493 ( .A(n13353), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13356), .Z(
        P2_U3542) );
  INV_X1 U15494 ( .A(n13354), .ZN(n13355) );
  MUX2_X1 U15495 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13355), .S(P2_U3947), .Z(
        P2_U3541) );
  MUX2_X1 U15496 ( .A(n13357), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13356), .Z(
        P2_U3540) );
  MUX2_X1 U15497 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13358), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U15498 ( .A(n13359), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13356), .Z(
        P2_U3538) );
  MUX2_X1 U15499 ( .A(n13360), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13356), .Z(
        P2_U3537) );
  MUX2_X1 U15500 ( .A(n13361), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13356), .Z(
        P2_U3536) );
  MUX2_X1 U15501 ( .A(n13362), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13356), .Z(
        P2_U3535) );
  MUX2_X1 U15502 ( .A(n8584), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13356), .Z(
        P2_U3534) );
  MUX2_X1 U15503 ( .A(n13363), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13356), .Z(
        P2_U3533) );
  MUX2_X1 U15504 ( .A(n13364), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13356), .Z(
        P2_U3532) );
  MUX2_X1 U15505 ( .A(n8582), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13356), .Z(
        P2_U3531) );
  OAI211_X1 U15506 ( .C1(n13367), .C2(n13366), .A(n15299), .B(n13365), .ZN(
        n13377) );
  AOI22_X1 U15507 ( .A1(n15328), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n13376) );
  MUX2_X1 U15508 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n11176), .S(n13368), .Z(
        n13369) );
  OAI21_X1 U15509 ( .B1(n13370), .B2(n12470), .A(n13369), .ZN(n13371) );
  NAND3_X1 U15510 ( .A1(n15306), .A2(n13372), .A3(n13371), .ZN(n13375) );
  NAND2_X1 U15511 ( .A1(n15310), .A2(n13373), .ZN(n13374) );
  NAND4_X1 U15512 ( .A1(n13377), .A2(n13376), .A3(n13375), .A4(n13374), .ZN(
        P2_U3215) );
  OAI211_X1 U15513 ( .C1(n13380), .C2(n13379), .A(n15299), .B(n13378), .ZN(
        n13390) );
  AND2_X1 U15514 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n13381) );
  AOI21_X1 U15515 ( .B1(n15328), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13381), .ZN(
        n13389) );
  MUX2_X1 U15516 ( .A(n11220), .B(P2_REG2_REG_3__SCAN_IN), .S(n13386), .Z(
        n13383) );
  NAND3_X1 U15517 ( .A1(n13383), .A2(n15240), .A3(n13382), .ZN(n13384) );
  NAND3_X1 U15518 ( .A1(n15306), .A2(n13385), .A3(n13384), .ZN(n13388) );
  NAND2_X1 U15519 ( .A1(n15310), .A2(n13386), .ZN(n13387) );
  NAND4_X1 U15520 ( .A1(n13390), .A2(n13389), .A3(n13388), .A4(n13387), .ZN(
        P2_U3217) );
  OAI211_X1 U15521 ( .C1(n13393), .C2(n13392), .A(n15299), .B(n13391), .ZN(
        n13403) );
  INV_X1 U15522 ( .A(n13394), .ZN(n13395) );
  AOI21_X1 U15523 ( .B1(n15328), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n13395), .ZN(
        n13402) );
  MUX2_X1 U15524 ( .A(n10329), .B(P2_REG2_REG_5__SCAN_IN), .S(n13399), .Z(
        n13396) );
  NAND3_X1 U15525 ( .A1(n15253), .A2(n13397), .A3(n13396), .ZN(n13398) );
  NAND3_X1 U15526 ( .A1(n15306), .A2(n13413), .A3(n13398), .ZN(n13401) );
  NAND2_X1 U15527 ( .A1(n15310), .A2(n13399), .ZN(n13400) );
  NAND4_X1 U15528 ( .A1(n13403), .A2(n13402), .A3(n13401), .A4(n13400), .ZN(
        P2_U3219) );
  NOR2_X1 U15529 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13404), .ZN(n13406) );
  INV_X1 U15530 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14774) );
  NOR2_X1 U15531 ( .A1(n15298), .A2(n14774), .ZN(n13405) );
  AOI211_X1 U15532 ( .C1(n15310), .C2(n13410), .A(n13406), .B(n13405), .ZN(
        n13417) );
  OAI211_X1 U15533 ( .C1(n13409), .C2(n13408), .A(n15299), .B(n13407), .ZN(
        n13416) );
  MUX2_X1 U15534 ( .A(n11210), .B(P2_REG2_REG_6__SCAN_IN), .S(n13410), .Z(
        n13411) );
  NAND3_X1 U15535 ( .A1(n13413), .A2(n13412), .A3(n13411), .ZN(n13414) );
  NAND3_X1 U15536 ( .A1(n15306), .A2(n13427), .A3(n13414), .ZN(n13415) );
  NAND3_X1 U15537 ( .A1(n13417), .A2(n13416), .A3(n13415), .ZN(P2_U3220) );
  INV_X1 U15538 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n13419) );
  OAI21_X1 U15539 ( .B1(n15298), .B2(n13419), .A(n13418), .ZN(n13420) );
  AOI21_X1 U15540 ( .B1(n13424), .B2(n15310), .A(n13420), .ZN(n13431) );
  OAI211_X1 U15541 ( .C1(n13423), .C2(n13422), .A(n15299), .B(n13421), .ZN(
        n13430) );
  MUX2_X1 U15542 ( .A(n11097), .B(P2_REG2_REG_7__SCAN_IN), .S(n13424), .Z(
        n13425) );
  NAND3_X1 U15543 ( .A1(n13427), .A2(n13426), .A3(n13425), .ZN(n13428) );
  NAND3_X1 U15544 ( .A1(n15306), .A2(n13441), .A3(n13428), .ZN(n13429) );
  NAND3_X1 U15545 ( .A1(n13431), .A2(n13430), .A3(n13429), .ZN(P2_U3221) );
  INV_X1 U15546 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n13433) );
  OAI21_X1 U15547 ( .B1(n15298), .B2(n13433), .A(n13432), .ZN(n13434) );
  AOI21_X1 U15548 ( .B1(n13438), .B2(n15310), .A(n13434), .ZN(n13446) );
  OAI211_X1 U15549 ( .C1(n13437), .C2(n13436), .A(n15299), .B(n13435), .ZN(
        n13445) );
  MUX2_X1 U15550 ( .A(n11383), .B(P2_REG2_REG_8__SCAN_IN), .S(n13438), .Z(
        n13439) );
  NAND3_X1 U15551 ( .A1(n13441), .A2(n13440), .A3(n13439), .ZN(n13442) );
  NAND3_X1 U15552 ( .A1(n15306), .A2(n13443), .A3(n13442), .ZN(n13444) );
  NAND3_X1 U15553 ( .A1(n13446), .A2(n13445), .A3(n13444), .ZN(P2_U3222) );
  NOR2_X1 U15554 ( .A1(n15284), .A2(n13448), .ZN(n13449) );
  AOI21_X1 U15555 ( .B1(n15284), .B2(n13448), .A(n13449), .ZN(n15281) );
  NOR2_X1 U15556 ( .A1(n15280), .A2(n15281), .ZN(n15279) );
  NOR2_X1 U15557 ( .A1(n13450), .A2(n13461), .ZN(n13451) );
  XNOR2_X1 U15558 ( .A(n13450), .B(n13461), .ZN(n15290) );
  NOR2_X1 U15559 ( .A1(n8225), .A2(n15290), .ZN(n15289) );
  XNOR2_X1 U15560 ( .A(n13481), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13452) );
  AOI21_X1 U15561 ( .B1(n13453), .B2(n13452), .A(n15319), .ZN(n13454) );
  NAND2_X1 U15562 ( .A1(n13454), .A2(n13483), .ZN(n13471) );
  NAND2_X1 U15563 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14894)
         );
  INV_X1 U15564 ( .A(n14894), .ZN(n13455) );
  AOI21_X1 U15565 ( .B1(n15328), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n13455), 
        .ZN(n13470) );
  NAND2_X1 U15566 ( .A1(n13456), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n13457) );
  NAND2_X1 U15567 ( .A1(n13458), .A2(n13457), .ZN(n13459) );
  NAND2_X1 U15568 ( .A1(n13459), .A2(n15284), .ZN(n15278) );
  NAND2_X1 U15569 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n15275), .ZN(n15274) );
  NAND2_X1 U15570 ( .A1(n15278), .A2(n15274), .ZN(n13460) );
  NAND2_X1 U15571 ( .A1(n15293), .A2(n13460), .ZN(n13462) );
  XNOR2_X1 U15572 ( .A(n13461), .B(n13460), .ZN(n15295) );
  NAND2_X1 U15573 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15295), .ZN(n15294) );
  NAND2_X1 U15574 ( .A1(n13462), .A2(n15294), .ZN(n13467) );
  NAND2_X1 U15575 ( .A1(n13481), .A2(n13463), .ZN(n13464) );
  OAI21_X1 U15576 ( .B1(n13481), .B2(n13463), .A(n13464), .ZN(n13466) );
  NAND2_X1 U15577 ( .A1(n13481), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13465) );
  OAI211_X1 U15578 ( .C1(n13481), .C2(P2_REG2_REG_16__SCAN_IN), .A(n13467), 
        .B(n13465), .ZN(n13474) );
  OAI211_X1 U15579 ( .C1(n13467), .C2(n13466), .A(n13474), .B(n15306), .ZN(
        n13469) );
  NAND2_X1 U15580 ( .A1(n15310), .A2(n13481), .ZN(n13468) );
  NAND4_X1 U15581 ( .A1(n13471), .A2(n13470), .A3(n13469), .A4(n13468), .ZN(
        P2_U3230) );
  INV_X1 U15582 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13473) );
  AOI22_X1 U15583 ( .A1(n15309), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13473), 
        .B2(n13472), .ZN(n15308) );
  OAI21_X1 U15584 ( .B1(n13463), .B2(n13475), .A(n13474), .ZN(n15307) );
  NAND2_X1 U15585 ( .A1(n15308), .A2(n15307), .ZN(n15305) );
  NAND2_X1 U15586 ( .A1(n15309), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13476) );
  AND2_X1 U15587 ( .A1(n15305), .A2(n13476), .ZN(n13478) );
  AND2_X1 U15588 ( .A1(n13478), .A2(n15324), .ZN(n13479) );
  INV_X1 U15589 ( .A(n13479), .ZN(n13477) );
  OAI21_X1 U15590 ( .B1(n13478), .B2(n15324), .A(n13477), .ZN(n15316) );
  NOR2_X1 U15591 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n15316), .ZN(n15315) );
  NOR2_X1 U15592 ( .A1(n15315), .A2(n13479), .ZN(n13480) );
  XOR2_X1 U15593 ( .A(n13480), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13488) );
  NAND2_X1 U15594 ( .A1(n13481), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n13482) );
  NAND2_X1 U15595 ( .A1(n13483), .A2(n13482), .ZN(n15301) );
  INV_X1 U15596 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13484) );
  XNOR2_X1 U15597 ( .A(n15309), .B(n13484), .ZN(n15300) );
  NOR2_X1 U15598 ( .A1(n13485), .A2(n15324), .ZN(n13486) );
  AOI21_X1 U15599 ( .B1(n13485), .B2(n15324), .A(n13486), .ZN(n15317) );
  AND2_X1 U15600 ( .A1(n15317), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n15318) );
  NOR2_X1 U15601 ( .A1(n15318), .A2(n13486), .ZN(n13487) );
  AOI22_X1 U15602 ( .A1(n13488), .A2(n15306), .B1(n13489), .B2(n15299), .ZN(
        n13494) );
  INV_X1 U15603 ( .A(n13488), .ZN(n13491) );
  NOR2_X1 U15604 ( .A1(n13489), .A2(n15319), .ZN(n13490) );
  AOI211_X1 U15605 ( .C1(n15306), .C2(n13491), .A(n15310), .B(n13490), .ZN(
        n13493) );
  MUX2_X1 U15606 ( .A(n13494), .B(n13493), .S(n6686), .Z(n13496) );
  OAI211_X1 U15607 ( .C1(n15298), .C2(n13497), .A(n13496), .B(n13495), .ZN(
        P2_U3233) );
  XNOR2_X1 U15608 ( .A(n13499), .B(n13498), .ZN(n13500) );
  NAND2_X1 U15609 ( .A1(n13753), .A2(n14931), .ZN(n13503) );
  NOR2_X1 U15610 ( .A1(n14919), .A2(n13501), .ZN(n13506) );
  AOI21_X1 U15611 ( .B1(n14935), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13506), 
        .ZN(n13502) );
  OAI211_X1 U15612 ( .C1(n7041), .C2(n13743), .A(n13503), .B(n13502), .ZN(
        P2_U3234) );
  NOR2_X1 U15613 ( .A1(n13504), .A2(n13743), .ZN(n13505) );
  AOI211_X1 U15614 ( .C1(n14935), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13506), 
        .B(n13505), .ZN(n13507) );
  OAI21_X1 U15615 ( .B1(n13713), .B2(n13508), .A(n13507), .ZN(P2_U3235) );
  NAND2_X1 U15616 ( .A1(n13550), .A2(n13511), .ZN(n13512) );
  NAND2_X1 U15617 ( .A1(n13828), .A2(n13553), .ZN(n13514) );
  NAND2_X1 U15618 ( .A1(n13515), .A2(n13514), .ZN(n13716) );
  NAND2_X1 U15619 ( .A1(n13725), .A2(n13517), .ZN(n13516) );
  NAND2_X1 U15620 ( .A1(n13716), .A2(n13516), .ZN(n13519) );
  OR2_X1 U15621 ( .A1(n13725), .A2(n13517), .ZN(n13518) );
  INV_X1 U15622 ( .A(n13520), .ZN(n13691) );
  OAI21_X1 U15623 ( .B1(n13699), .B2(n13523), .A(n13521), .ZN(n13522) );
  NAND2_X1 U15624 ( .A1(n13699), .A2(n13523), .ZN(n13524) );
  NAND2_X1 U15625 ( .A1(n13802), .A2(n13525), .ZN(n13526) );
  NOR2_X1 U15626 ( .A1(n13865), .A2(n13529), .ZN(n13528) );
  NAND2_X1 U15627 ( .A1(n13865), .A2(n13529), .ZN(n13530) );
  OR2_X1 U15628 ( .A1(n13639), .A2(n13532), .ZN(n13533) );
  NAND2_X1 U15629 ( .A1(n13629), .A2(n13533), .ZN(n13615) );
  NAND2_X1 U15630 ( .A1(n13619), .A2(n13569), .ZN(n13534) );
  NAND2_X1 U15631 ( .A1(n13615), .A2(n13534), .ZN(n13536) );
  NAND2_X1 U15632 ( .A1(n13854), .A2(n13571), .ZN(n13535) );
  NAND2_X1 U15633 ( .A1(n13536), .A2(n13535), .ZN(n13601) );
  NAND2_X1 U15634 ( .A1(n13586), .A2(n13585), .ZN(n13584) );
  NAND2_X1 U15635 ( .A1(n13596), .A2(n13538), .ZN(n13539) );
  NAND2_X1 U15636 ( .A1(n13584), .A2(n13539), .ZN(n13540) );
  XNOR2_X1 U15637 ( .A(n13540), .B(n13575), .ZN(n13541) );
  OAI22_X1 U15638 ( .A1(n13545), .A2(n13544), .B1(n13543), .B2(n13542), .ZN(
        n13546) );
  INV_X1 U15639 ( .A(n13546), .ZN(n13547) );
  OR2_X1 U15640 ( .A1(n13550), .A2(n13549), .ZN(n13551) );
  NAND2_X1 U15641 ( .A1(n13552), .A2(n13551), .ZN(n13733) );
  NAND2_X1 U15642 ( .A1(n13744), .A2(n13553), .ZN(n13554) );
  NAND2_X1 U15643 ( .A1(n13731), .A2(n13554), .ZN(n13727) );
  INV_X1 U15644 ( .A(n13689), .ZN(n13692) );
  OR2_X1 U15645 ( .A1(n13699), .A2(n13557), .ZN(n13558) );
  NAND2_X1 U15646 ( .A1(n13865), .A2(n13561), .ZN(n13560) );
  NAND2_X1 U15647 ( .A1(n13667), .A2(n13560), .ZN(n13563) );
  OR2_X1 U15648 ( .A1(n13865), .A2(n13561), .ZN(n13562) );
  NAND2_X1 U15649 ( .A1(n13563), .A2(n13562), .ZN(n13645) );
  NAND2_X1 U15650 ( .A1(n13645), .A2(n13647), .ZN(n13566) );
  NAND2_X1 U15651 ( .A1(n13787), .A2(n13564), .ZN(n13565) );
  NAND2_X1 U15652 ( .A1(n13639), .A2(n13567), .ZN(n13568) );
  NAND2_X1 U15653 ( .A1(n13854), .A2(n13569), .ZN(n13570) );
  NAND2_X1 U15654 ( .A1(n13619), .A2(n13571), .ZN(n13572) );
  INV_X1 U15655 ( .A(n13585), .ZN(n13590) );
  NAND2_X1 U15656 ( .A1(n13591), .A2(n13590), .ZN(n13589) );
  NAND2_X1 U15657 ( .A1(n13589), .A2(n13574), .ZN(n13576) );
  XNOR2_X1 U15658 ( .A(n13576), .B(n13575), .ZN(n13756) );
  OAI211_X1 U15659 ( .C1(n13580), .C2(n13593), .A(n14928), .B(n13577), .ZN(
        n13757) );
  NOR2_X1 U15660 ( .A1(n13757), .A2(n13713), .ZN(n13582) );
  AOI22_X1 U15661 ( .A1(n13578), .A2(n14918), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14935), .ZN(n13579) );
  OAI21_X1 U15662 ( .B1(n13580), .B2(n13743), .A(n13579), .ZN(n13581) );
  AOI211_X1 U15663 ( .C1(n13756), .C2(n14932), .A(n13582), .B(n13581), .ZN(
        n13583) );
  OAI21_X1 U15664 ( .B1(n6804), .B2(n14919), .A(n13583), .ZN(P2_U3236) );
  OAI211_X1 U15665 ( .C1(n13586), .C2(n13585), .A(n13584), .B(n14915), .ZN(
        n13588) );
  OAI21_X1 U15666 ( .B1(n13591), .B2(n13590), .A(n13589), .ZN(n13761) );
  INV_X1 U15667 ( .A(n13761), .ZN(n13599) );
  OAI21_X1 U15668 ( .B1(n13596), .B2(n13602), .A(n14928), .ZN(n13592) );
  NOR2_X1 U15669 ( .A1(n13759), .A2(n13713), .ZN(n13598) );
  AOI22_X1 U15670 ( .A1(n13594), .A2(n14918), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14935), .ZN(n13595) );
  OAI21_X1 U15671 ( .B1(n13596), .B2(n13743), .A(n13595), .ZN(n13597) );
  AOI211_X1 U15672 ( .C1(n13599), .C2(n14932), .A(n13598), .B(n13597), .ZN(
        n13600) );
  OAI21_X1 U15673 ( .B1(n13760), .B2(n14919), .A(n13600), .ZN(P2_U3237) );
  XOR2_X1 U15674 ( .A(n13601), .B(n13611), .Z(n13769) );
  INV_X1 U15675 ( .A(n13621), .ZN(n13603) );
  AOI211_X1 U15676 ( .C1(n13764), .C2(n13603), .A(n13720), .B(n13602), .ZN(
        n13762) );
  INV_X1 U15677 ( .A(n13604), .ZN(n13605) );
  AOI22_X1 U15678 ( .A1(n13605), .A2(n14918), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14935), .ZN(n13608) );
  INV_X1 U15679 ( .A(n13606), .ZN(n13763) );
  NAND2_X1 U15680 ( .A1(n13763), .A2(n13741), .ZN(n13607) );
  OAI211_X1 U15681 ( .C1(n13609), .C2(n13743), .A(n13608), .B(n13607), .ZN(
        n13610) );
  AOI21_X1 U15682 ( .B1(n13762), .B2(n14931), .A(n13610), .ZN(n13614) );
  NAND2_X1 U15683 ( .A1(n13612), .A2(n13611), .ZN(n13765) );
  NAND3_X1 U15684 ( .A1(n13766), .A2(n13765), .A3(n14932), .ZN(n13613) );
  OAI211_X1 U15685 ( .C1(n13769), .C2(n13688), .A(n13614), .B(n13613), .ZN(
        P2_U3238) );
  XNOR2_X1 U15686 ( .A(n13616), .B(n13615), .ZN(n13774) );
  INV_X1 U15687 ( .A(n13774), .ZN(n13628) );
  INV_X1 U15688 ( .A(n13616), .ZN(n13617) );
  XNOR2_X1 U15689 ( .A(n13618), .B(n13617), .ZN(n13770) );
  OAI21_X1 U15690 ( .B1(n13619), .B2(n13641), .A(n14928), .ZN(n13620) );
  OR2_X1 U15691 ( .A1(n13621), .A2(n13620), .ZN(n13772) );
  AOI22_X1 U15692 ( .A1(n13622), .A2(n14918), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14919), .ZN(n13623) );
  OAI21_X1 U15693 ( .B1(n13771), .B2(n14935), .A(n13623), .ZN(n13624) );
  AOI21_X1 U15694 ( .B1(n13854), .B2(n14920), .A(n13624), .ZN(n13625) );
  OAI21_X1 U15695 ( .B1(n13772), .B2(n13713), .A(n13625), .ZN(n13626) );
  AOI21_X1 U15696 ( .B1(n13770), .B2(n14932), .A(n13626), .ZN(n13627) );
  OAI21_X1 U15697 ( .B1(n13628), .B2(n13688), .A(n13627), .ZN(P2_U3239) );
  OAI21_X1 U15698 ( .B1(n13630), .B2(n13633), .A(n13629), .ZN(n13632) );
  AOI21_X1 U15699 ( .B1(n13632), .B2(n14915), .A(n13631), .ZN(n13781) );
  NAND2_X1 U15700 ( .A1(n13634), .A2(n13633), .ZN(n13635) );
  NAND2_X1 U15701 ( .A1(n13636), .A2(n13635), .ZN(n13779) );
  AOI22_X1 U15702 ( .A1(n13637), .A2(n14918), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14919), .ZN(n13638) );
  OAI21_X1 U15703 ( .B1(n13639), .B2(n13743), .A(n13638), .ZN(n13643) );
  OAI21_X1 U15704 ( .B1(n13639), .B2(n13653), .A(n14928), .ZN(n13640) );
  OR2_X1 U15705 ( .A1(n13641), .A2(n13640), .ZN(n13780) );
  NOR2_X1 U15706 ( .A1(n13780), .A2(n13713), .ZN(n13642) );
  AOI211_X1 U15707 ( .C1(n13779), .C2(n14932), .A(n13643), .B(n13642), .ZN(
        n13644) );
  OAI21_X1 U15708 ( .B1(n14935), .B2(n13781), .A(n13644), .ZN(P2_U3240) );
  XNOR2_X1 U15709 ( .A(n13645), .B(n7174), .ZN(n13785) );
  NAND2_X1 U15710 ( .A1(n13647), .A2(n13646), .ZN(n13648) );
  AOI21_X1 U15711 ( .B1(n13649), .B2(n13648), .A(n13806), .ZN(n13651) );
  AOI211_X1 U15712 ( .C1(n13785), .C2(n13652), .A(n13651), .B(n13650), .ZN(
        n13789) );
  INV_X1 U15713 ( .A(n13670), .ZN(n13654) );
  AOI211_X1 U15714 ( .C1(n13787), .C2(n13654), .A(n13720), .B(n13653), .ZN(
        n13786) );
  NAND2_X1 U15715 ( .A1(n13786), .A2(n14931), .ZN(n13658) );
  INV_X1 U15716 ( .A(n13655), .ZN(n13656) );
  AOI22_X1 U15717 ( .A1(n13656), .A2(n14918), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14935), .ZN(n13657) );
  OAI211_X1 U15718 ( .C1(n13659), .C2(n13743), .A(n13658), .B(n13657), .ZN(
        n13660) );
  AOI21_X1 U15719 ( .B1(n13785), .B2(n13661), .A(n13660), .ZN(n13662) );
  OAI21_X1 U15720 ( .B1(n13789), .B2(n14919), .A(n13662), .ZN(P2_U3241) );
  XOR2_X1 U15721 ( .A(n13668), .B(n13663), .Z(n13664) );
  NAND2_X1 U15722 ( .A1(n13664), .A2(n14915), .ZN(n13794) );
  INV_X1 U15723 ( .A(n13794), .ZN(n13665) );
  AOI211_X1 U15724 ( .C1(n14918), .C2(n13666), .A(n13791), .B(n13665), .ZN(
        n13674) );
  XOR2_X1 U15725 ( .A(n13668), .B(n13667), .Z(n13796) );
  OAI21_X1 U15726 ( .B1(n13865), .B2(n13680), .A(n14928), .ZN(n13669) );
  OR2_X1 U15727 ( .A1(n13670), .A2(n13669), .ZN(n13792) );
  AOI22_X1 U15728 ( .A1(n7237), .A2(n14920), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14935), .ZN(n13671) );
  OAI21_X1 U15729 ( .B1(n13792), .B2(n13713), .A(n13671), .ZN(n13672) );
  AOI21_X1 U15730 ( .B1(n13796), .B2(n14932), .A(n13672), .ZN(n13673) );
  OAI21_X1 U15731 ( .B1(n13674), .B2(n14919), .A(n13673), .ZN(P2_U3242) );
  XOR2_X1 U15732 ( .A(n13677), .B(n13675), .Z(n13805) );
  AOI21_X1 U15733 ( .B1(n13677), .B2(n13676), .A(n6753), .ZN(n13799) );
  NAND2_X1 U15734 ( .A1(n13694), .A2(n13802), .ZN(n13678) );
  NAND2_X1 U15735 ( .A1(n13678), .A2(n14928), .ZN(n13679) );
  NOR2_X1 U15736 ( .A1(n13680), .A2(n13679), .ZN(n13800) );
  NAND2_X1 U15737 ( .A1(n13800), .A2(n14931), .ZN(n13685) );
  INV_X1 U15738 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13681) );
  OAI22_X1 U15739 ( .A1(n13682), .A2(n13737), .B1(n13681), .B2(n13741), .ZN(
        n13683) );
  AOI21_X1 U15740 ( .B1(n13801), .B2(n13741), .A(n13683), .ZN(n13684) );
  OAI211_X1 U15741 ( .C1(n7236), .C2(n13743), .A(n13685), .B(n13684), .ZN(
        n13686) );
  AOI21_X1 U15742 ( .B1(n13799), .B2(n14932), .A(n13686), .ZN(n13687) );
  OAI21_X1 U15743 ( .B1(n13805), .B2(n13688), .A(n13687), .ZN(P2_U3243) );
  XNOR2_X1 U15744 ( .A(n13690), .B(n13689), .ZN(n13813) );
  INV_X1 U15745 ( .A(n13703), .ZN(n13705) );
  AOI21_X1 U15746 ( .B1(n13706), .B2(n13705), .A(n13691), .ZN(n13693) );
  XNOR2_X1 U15747 ( .A(n13693), .B(n13692), .ZN(n13811) );
  INV_X1 U15748 ( .A(n13707), .ZN(n13695) );
  OAI211_X1 U15749 ( .C1(n13809), .C2(n13695), .A(n13694), .B(n14928), .ZN(
        n13808) );
  AOI22_X1 U15750 ( .A1(n13696), .A2(n14918), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n14919), .ZN(n13697) );
  OAI21_X1 U15751 ( .B1(n13807), .B2(n14935), .A(n13697), .ZN(n13698) );
  AOI21_X1 U15752 ( .B1(n13699), .B2(n14920), .A(n13698), .ZN(n13700) );
  OAI21_X1 U15753 ( .B1(n13808), .B2(n13713), .A(n13700), .ZN(n13701) );
  AOI21_X1 U15754 ( .B1(n13811), .B2(n13748), .A(n13701), .ZN(n13702) );
  OAI21_X1 U15755 ( .B1(n13813), .B2(n13751), .A(n13702), .ZN(P2_U3244) );
  XNOR2_X1 U15756 ( .A(n13704), .B(n13703), .ZN(n13820) );
  XNOR2_X1 U15757 ( .A(n13706), .B(n13705), .ZN(n13818) );
  OAI211_X1 U15758 ( .C1(n13719), .C2(n13816), .A(n14928), .B(n13707), .ZN(
        n13815) );
  AOI22_X1 U15759 ( .A1(n13708), .A2(n14918), .B1(P2_REG2_REG_20__SCAN_IN), 
        .B2(n14919), .ZN(n13709) );
  OAI21_X1 U15760 ( .B1(n13814), .B2(n14935), .A(n13709), .ZN(n13710) );
  AOI21_X1 U15761 ( .B1(n13711), .B2(n14920), .A(n13710), .ZN(n13712) );
  OAI21_X1 U15762 ( .B1(n13815), .B2(n13713), .A(n13712), .ZN(n13714) );
  AOI21_X1 U15763 ( .B1(n13818), .B2(n13748), .A(n13714), .ZN(n13715) );
  OAI21_X1 U15764 ( .B1(n13820), .B2(n13751), .A(n13715), .ZN(P2_U3245) );
  XNOR2_X1 U15765 ( .A(n13716), .B(n13726), .ZN(n13718) );
  AOI21_X1 U15766 ( .B1(n13718), .B2(n14915), .A(n13717), .ZN(n13823) );
  INV_X1 U15767 ( .A(n13735), .ZN(n13721) );
  AOI211_X1 U15768 ( .C1(n13822), .C2(n13721), .A(n13720), .B(n13719), .ZN(
        n13821) );
  INV_X1 U15769 ( .A(n13722), .ZN(n13723) );
  AOI22_X1 U15770 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(n14919), .B1(n13723), 
        .B2(n14918), .ZN(n13724) );
  OAI21_X1 U15771 ( .B1(n13725), .B2(n13743), .A(n13724), .ZN(n13729) );
  XNOR2_X1 U15772 ( .A(n13727), .B(n13726), .ZN(n13825) );
  NOR2_X1 U15773 ( .A1(n13825), .A2(n13751), .ZN(n13728) );
  AOI211_X1 U15774 ( .C1(n13821), .C2(n14931), .A(n13729), .B(n13728), .ZN(
        n13730) );
  OAI21_X1 U15775 ( .B1(n14919), .B2(n13823), .A(n13730), .ZN(P2_U3246) );
  INV_X1 U15776 ( .A(n13731), .ZN(n13732) );
  AOI21_X1 U15777 ( .B1(n13747), .B2(n13733), .A(n13732), .ZN(n13832) );
  OAI21_X1 U15778 ( .B1(n13744), .B2(n13734), .A(n14928), .ZN(n13736) );
  NOR2_X1 U15779 ( .A1(n13736), .A2(n13735), .ZN(n13826) );
  NOR2_X1 U15780 ( .A1(n13738), .A2(n13737), .ZN(n13740) );
  AND2_X1 U15781 ( .A1(n14919), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13739) );
  AOI211_X1 U15782 ( .C1(n13827), .C2(n13741), .A(n13740), .B(n13739), .ZN(
        n13742) );
  OAI21_X1 U15783 ( .B1(n13744), .B2(n13743), .A(n13742), .ZN(n13745) );
  AOI21_X1 U15784 ( .B1(n13826), .B2(n14931), .A(n13745), .ZN(n13750) );
  XOR2_X1 U15785 ( .A(n13747), .B(n13746), .Z(n13829) );
  NAND2_X1 U15786 ( .A1(n13829), .A2(n13748), .ZN(n13749) );
  OAI211_X1 U15787 ( .C1(n13832), .C2(n13751), .A(n13750), .B(n13749), .ZN(
        P2_U3247) );
  INV_X1 U15788 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13754) );
  NOR2_X1 U15789 ( .A1(n13753), .A2(n13752), .ZN(n13844) );
  MUX2_X1 U15790 ( .A(n13754), .B(n13844), .S(n15391), .Z(n13755) );
  OAI21_X1 U15791 ( .B1(n7041), .B2(n7353), .A(n13755), .ZN(P2_U3530) );
  NAND2_X1 U15792 ( .A1(n13756), .A2(n14941), .ZN(n13758) );
  AOI211_X1 U15793 ( .C1(n15373), .C2(n13764), .A(n13763), .B(n13762), .ZN(
        n13768) );
  NAND3_X1 U15794 ( .A1(n13766), .A2(n14941), .A3(n13765), .ZN(n13767) );
  OAI211_X1 U15795 ( .C1(n13806), .C2(n13769), .A(n13768), .B(n13767), .ZN(
        n13851) );
  MUX2_X1 U15796 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13851), .S(n15391), .Z(
        P2_U3526) );
  NAND2_X1 U15797 ( .A1(n13770), .A2(n14941), .ZN(n13776) );
  NAND2_X1 U15798 ( .A1(n13772), .A2(n13771), .ZN(n13773) );
  AOI21_X1 U15799 ( .B1(n13774), .B2(n14915), .A(n13773), .ZN(n13775) );
  NAND2_X1 U15800 ( .A1(n13776), .A2(n13775), .ZN(n13852) );
  MUX2_X1 U15801 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13852), .S(n15391), .Z(
        n13777) );
  AOI21_X1 U15802 ( .B1(n13837), .B2(n13854), .A(n13777), .ZN(n13778) );
  INV_X1 U15803 ( .A(n13778), .ZN(P2_U3525) );
  NAND2_X1 U15804 ( .A1(n13779), .A2(n14941), .ZN(n13782) );
  NAND3_X1 U15805 ( .A1(n13782), .A2(n13781), .A3(n13780), .ZN(n13856) );
  MUX2_X1 U15806 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13856), .S(n15391), .Z(
        n13783) );
  AOI21_X1 U15807 ( .B1(n13837), .B2(n13858), .A(n13783), .ZN(n13784) );
  INV_X1 U15808 ( .A(n13784), .ZN(P2_U3524) );
  INV_X1 U15809 ( .A(n13785), .ZN(n13790) );
  AOI21_X1 U15810 ( .B1(n15373), .B2(n13787), .A(n13786), .ZN(n13788) );
  OAI211_X1 U15811 ( .C1(n15377), .C2(n13790), .A(n13789), .B(n13788), .ZN(
        n13860) );
  MUX2_X1 U15812 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13860), .S(n15391), .Z(
        P2_U3523) );
  INV_X1 U15813 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13797) );
  INV_X1 U15814 ( .A(n13791), .ZN(n13793) );
  NAND3_X1 U15815 ( .A1(n13794), .A2(n13793), .A3(n13792), .ZN(n13795) );
  AOI21_X1 U15816 ( .B1(n13796), .B2(n14941), .A(n13795), .ZN(n13861) );
  MUX2_X1 U15817 ( .A(n13797), .B(n13861), .S(n15391), .Z(n13798) );
  OAI21_X1 U15818 ( .B1(n13865), .B2(n7353), .A(n13798), .ZN(P2_U3522) );
  NAND2_X1 U15819 ( .A1(n13799), .A2(n14941), .ZN(n13804) );
  AOI211_X1 U15820 ( .C1(n15373), .C2(n13802), .A(n13801), .B(n13800), .ZN(
        n13803) );
  OAI211_X1 U15821 ( .C1(n13806), .C2(n13805), .A(n13804), .B(n13803), .ZN(
        n13866) );
  MUX2_X1 U15822 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13866), .S(n15391), .Z(
        P2_U3521) );
  OAI211_X1 U15823 ( .C1(n13809), .C2(n15381), .A(n13808), .B(n13807), .ZN(
        n13810) );
  AOI21_X1 U15824 ( .B1(n13811), .B2(n14915), .A(n13810), .ZN(n13812) );
  OAI21_X1 U15825 ( .B1(n13813), .B2(n13842), .A(n13812), .ZN(n13867) );
  MUX2_X1 U15826 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13867), .S(n15391), .Z(
        P2_U3520) );
  OAI211_X1 U15827 ( .C1(n13816), .C2(n15381), .A(n13815), .B(n13814), .ZN(
        n13817) );
  AOI21_X1 U15828 ( .B1(n13818), .B2(n14915), .A(n13817), .ZN(n13819) );
  OAI21_X1 U15829 ( .B1(n13820), .B2(n13842), .A(n13819), .ZN(n13868) );
  MUX2_X1 U15830 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13868), .S(n15391), .Z(
        P2_U3519) );
  AOI21_X1 U15831 ( .B1(n15373), .B2(n13822), .A(n13821), .ZN(n13824) );
  OAI211_X1 U15832 ( .C1(n13825), .C2(n13842), .A(n13824), .B(n13823), .ZN(
        n13869) );
  MUX2_X1 U15833 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13869), .S(n15391), .Z(
        P2_U3518) );
  AOI211_X1 U15834 ( .C1(n15373), .C2(n13828), .A(n13827), .B(n13826), .ZN(
        n13831) );
  NAND2_X1 U15835 ( .A1(n13829), .A2(n14915), .ZN(n13830) );
  OAI211_X1 U15836 ( .C1(n13832), .C2(n13842), .A(n13831), .B(n13830), .ZN(
        n13870) );
  MUX2_X1 U15837 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13870), .S(n15391), .Z(
        P2_U3517) );
  OAI211_X1 U15838 ( .C1(n13835), .C2(n13842), .A(n13834), .B(n13833), .ZN(
        n13871) );
  MUX2_X1 U15839 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13871), .S(n15391), .Z(
        n13836) );
  AOI21_X1 U15840 ( .B1(n13837), .B2(n14907), .A(n13836), .ZN(n13838) );
  INV_X1 U15841 ( .A(n13838), .ZN(P2_U3516) );
  AOI21_X1 U15842 ( .B1(n15373), .B2(n14893), .A(n13839), .ZN(n13840) );
  OAI211_X1 U15843 ( .C1(n13843), .C2(n13842), .A(n13841), .B(n13840), .ZN(
        n13875) );
  MUX2_X1 U15844 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13875), .S(n15391), .Z(
        P2_U3515) );
  MUX2_X1 U15845 ( .A(n13845), .B(n13844), .S(n15387), .Z(n13846) );
  OAI21_X1 U15846 ( .B1(n7041), .B2(n13864), .A(n13846), .ZN(P2_U3498) );
  MUX2_X1 U15847 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13851), .S(n15387), .Z(
        P2_U3494) );
  MUX2_X1 U15848 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13852), .S(n15387), .Z(
        n13853) );
  AOI21_X1 U15849 ( .B1(n13873), .B2(n13854), .A(n13853), .ZN(n13855) );
  INV_X1 U15850 ( .A(n13855), .ZN(P2_U3493) );
  MUX2_X1 U15851 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13856), .S(n15387), .Z(
        n13857) );
  AOI21_X1 U15852 ( .B1(n13873), .B2(n13858), .A(n13857), .ZN(n13859) );
  INV_X1 U15853 ( .A(n13859), .ZN(P2_U3492) );
  MUX2_X1 U15854 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13860), .S(n15387), .Z(
        P2_U3491) );
  MUX2_X1 U15855 ( .A(n13862), .B(n13861), .S(n15387), .Z(n13863) );
  OAI21_X1 U15856 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(P2_U3490) );
  MUX2_X1 U15857 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13866), .S(n15387), .Z(
        P2_U3489) );
  MUX2_X1 U15858 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13867), .S(n15387), .Z(
        P2_U3488) );
  MUX2_X1 U15859 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13868), .S(n15387), .Z(
        P2_U3487) );
  MUX2_X1 U15860 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13869), .S(n15387), .Z(
        P2_U3486) );
  MUX2_X1 U15861 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13870), .S(n15387), .Z(
        P2_U3484) );
  MUX2_X1 U15862 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13871), .S(n15387), .Z(
        n13872) );
  AOI21_X1 U15863 ( .B1(n13873), .B2(n14907), .A(n13872), .ZN(n13874) );
  INV_X1 U15864 ( .A(n13874), .ZN(P2_U3481) );
  MUX2_X1 U15865 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13875), .S(n15387), .Z(
        P2_U3478) );
  INV_X1 U15866 ( .A(n13876), .ZN(n14681) );
  INV_X1 U15867 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13878) );
  NAND3_X1 U15868 ( .A1(n13878), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13880) );
  OAI22_X1 U15869 ( .A1(n13877), .A2(n13880), .B1(n13879), .B2(n13894), .ZN(
        n13881) );
  INV_X1 U15870 ( .A(n13881), .ZN(n13882) );
  OAI21_X1 U15871 ( .B1(n14681), .B2(n13883), .A(n13882), .ZN(P2_U3296) );
  INV_X1 U15872 ( .A(n13884), .ZN(n14683) );
  OAI222_X1 U15873 ( .A1(n13892), .A2(n14683), .B1(P2_U3088), .B2(n13885), 
        .C1(n13886), .C2(n13894), .ZN(P2_U3297) );
  INV_X1 U15874 ( .A(n13887), .ZN(n14688) );
  OAI222_X1 U15875 ( .A1(n13889), .A2(P2_U3088), .B1(n13892), .B2(n14688), 
        .C1(n13888), .C2(n13894), .ZN(P2_U3301) );
  INV_X1 U15876 ( .A(n13890), .ZN(n14693) );
  OAI222_X1 U15877 ( .A1(n13894), .A2(n13893), .B1(n13892), .B2(n14693), .C1(
        n13891), .C2(P2_U3088), .ZN(P2_U3302) );
  MUX2_X1 U15878 ( .A(n13895), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15879 ( .A1(n14589), .A2(n14042), .ZN(n13897) );
  NAND2_X1 U15880 ( .A1(n14344), .A2(n6666), .ZN(n13896) );
  NAND2_X1 U15881 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  XNOR2_X1 U15882 ( .A(n13898), .B(n14043), .ZN(n13902) );
  NAND2_X1 U15883 ( .A1(n14589), .A2(n6666), .ZN(n13900) );
  NAND2_X1 U15884 ( .A1(n14344), .A2(n14045), .ZN(n13899) );
  NAND2_X1 U15885 ( .A1(n13900), .A2(n13899), .ZN(n13901) );
  NOR2_X1 U15886 ( .A1(n13902), .A2(n13901), .ZN(n14039) );
  AOI21_X1 U15887 ( .B1(n13902), .B2(n13901), .A(n14039), .ZN(n14004) );
  NOR2_X1 U15888 ( .A1(n14109), .A2(n13940), .ZN(n13903) );
  AOI21_X1 U15889 ( .B1(n14512), .B2(n6666), .A(n13903), .ZN(n13939) );
  NAND2_X1 U15890 ( .A1(n14512), .A2(n14042), .ZN(n13905) );
  INV_X1 U15891 ( .A(n14109), .ZN(n14304) );
  NAND2_X1 U15892 ( .A1(n14304), .A2(n6666), .ZN(n13904) );
  NAND2_X1 U15893 ( .A1(n13905), .A2(n13904), .ZN(n13906) );
  XNOR2_X1 U15894 ( .A(n13906), .B(n14043), .ZN(n13934) );
  NAND2_X1 U15895 ( .A1(n14963), .A2(n14042), .ZN(n13912) );
  OR2_X1 U15896 ( .A1(n14294), .A2(n13941), .ZN(n13911) );
  NAND2_X1 U15897 ( .A1(n13912), .A2(n13911), .ZN(n13913) );
  XNOR2_X1 U15898 ( .A(n13913), .B(n14043), .ZN(n13916) );
  NOR2_X1 U15899 ( .A1(n14294), .A2(n13940), .ZN(n13914) );
  AOI21_X1 U15900 ( .B1(n14963), .B2(n6666), .A(n13914), .ZN(n14151) );
  OAI22_X1 U15901 ( .A1(n14562), .A2(n13942), .B1(n14298), .B2(n13941), .ZN(
        n13917) );
  XOR2_X1 U15902 ( .A(n14043), .B(n13917), .Z(n13919) );
  AOI22_X1 U15903 ( .A1(n14656), .A2(n6666), .B1(n14045), .B2(n14327), .ZN(
        n13918) );
  NAND2_X1 U15904 ( .A1(n13919), .A2(n13918), .ZN(n13920) );
  OAI21_X1 U15905 ( .B1(n13919), .B2(n13918), .A(n13920), .ZN(n14073) );
  INV_X1 U15906 ( .A(n13920), .ZN(n14085) );
  NAND2_X1 U15907 ( .A1(n14650), .A2(n14042), .ZN(n13922) );
  OR2_X1 U15908 ( .A1(n14132), .A2(n13941), .ZN(n13921) );
  NAND2_X1 U15909 ( .A1(n13922), .A2(n13921), .ZN(n13923) );
  XNOR2_X1 U15910 ( .A(n13923), .B(n13985), .ZN(n13925) );
  NOR2_X1 U15911 ( .A1(n14132), .A2(n13940), .ZN(n13924) );
  AOI21_X1 U15912 ( .B1(n14650), .B2(n6666), .A(n13924), .ZN(n13926) );
  NAND2_X1 U15913 ( .A1(n13925), .A2(n13926), .ZN(n13930) );
  INV_X1 U15914 ( .A(n13925), .ZN(n13928) );
  INV_X1 U15915 ( .A(n13926), .ZN(n13927) );
  NAND2_X1 U15916 ( .A1(n13928), .A2(n13927), .ZN(n13929) );
  AND2_X1 U15917 ( .A1(n13930), .A2(n13929), .ZN(n14084) );
  OAI22_X1 U15918 ( .A1(n14529), .A2(n13941), .B1(n14302), .B2(n13940), .ZN(
        n13936) );
  NAND2_X1 U15919 ( .A1(n14646), .A2(n14042), .ZN(n13932) );
  NAND2_X1 U15920 ( .A1(n14330), .A2(n6666), .ZN(n13931) );
  NAND2_X1 U15921 ( .A1(n13932), .A2(n13931), .ZN(n13933) );
  XNOR2_X1 U15922 ( .A(n13933), .B(n14043), .ZN(n13935) );
  XOR2_X1 U15923 ( .A(n13936), .B(n13935), .Z(n14130) );
  NAND2_X1 U15924 ( .A1(n14129), .A2(n14130), .ZN(n14128) );
  XNOR2_X1 U15925 ( .A(n13934), .B(n13939), .ZN(n14032) );
  INV_X1 U15926 ( .A(n13935), .ZN(n13938) );
  INV_X1 U15927 ( .A(n13936), .ZN(n13937) );
  NAND2_X1 U15928 ( .A1(n13938), .A2(n13937), .ZN(n14030) );
  OAI22_X1 U15929 ( .A1(n14634), .A2(n13941), .B1(n14309), .B2(n13940), .ZN(
        n13945) );
  OAI22_X1 U15930 ( .A1(n14634), .A2(n13942), .B1(n14309), .B2(n13941), .ZN(
        n13943) );
  XNOR2_X1 U15931 ( .A(n13943), .B(n14043), .ZN(n13944) );
  XOR2_X1 U15932 ( .A(n13945), .B(n13944), .Z(n14107) );
  NAND2_X1 U15933 ( .A1(n14484), .A2(n14042), .ZN(n13947) );
  NAND2_X1 U15934 ( .A1(n14336), .A2(n6666), .ZN(n13946) );
  NAND2_X1 U15935 ( .A1(n13947), .A2(n13946), .ZN(n13948) );
  XNOR2_X1 U15936 ( .A(n13948), .B(n14043), .ZN(n13952) );
  NAND2_X1 U15937 ( .A1(n14484), .A2(n6666), .ZN(n13950) );
  NAND2_X1 U15938 ( .A1(n14336), .A2(n14045), .ZN(n13949) );
  NAND2_X1 U15939 ( .A1(n13950), .A2(n13949), .ZN(n13951) );
  NOR2_X1 U15940 ( .A1(n13952), .A2(n13951), .ZN(n13953) );
  AOI21_X1 U15941 ( .B1(n13952), .B2(n13951), .A(n13953), .ZN(n14054) );
  INV_X1 U15942 ( .A(n13953), .ZN(n14117) );
  NAND2_X1 U15943 ( .A1(n14461), .A2(n14042), .ZN(n13955) );
  NAND2_X1 U15944 ( .A1(n14311), .A2(n6666), .ZN(n13954) );
  NAND2_X1 U15945 ( .A1(n13955), .A2(n13954), .ZN(n13956) );
  XNOR2_X1 U15946 ( .A(n13956), .B(n13985), .ZN(n13958) );
  AND2_X1 U15947 ( .A1(n14311), .A2(n14045), .ZN(n13957) );
  AOI21_X1 U15948 ( .B1(n14461), .B2(n6666), .A(n13957), .ZN(n13959) );
  NAND2_X1 U15949 ( .A1(n13958), .A2(n13959), .ZN(n13963) );
  INV_X1 U15950 ( .A(n13958), .ZN(n13961) );
  INV_X1 U15951 ( .A(n13959), .ZN(n13960) );
  NAND2_X1 U15952 ( .A1(n13961), .A2(n13960), .ZN(n13962) );
  NAND2_X1 U15953 ( .A1(n13963), .A2(n13962), .ZN(n14116) );
  INV_X1 U15954 ( .A(n13963), .ZN(n14011) );
  NAND2_X1 U15955 ( .A1(n14452), .A2(n14042), .ZN(n13965) );
  NAND2_X1 U15956 ( .A1(n14313), .A2(n6666), .ZN(n13964) );
  NAND2_X1 U15957 ( .A1(n13965), .A2(n13964), .ZN(n13966) );
  XNOR2_X1 U15958 ( .A(n13966), .B(n13985), .ZN(n13968) );
  AND2_X1 U15959 ( .A1(n14313), .A2(n14045), .ZN(n13967) );
  AOI21_X1 U15960 ( .B1(n14452), .B2(n6666), .A(n13967), .ZN(n13969) );
  NAND2_X1 U15961 ( .A1(n13968), .A2(n13969), .ZN(n14096) );
  INV_X1 U15962 ( .A(n13968), .ZN(n13971) );
  INV_X1 U15963 ( .A(n13969), .ZN(n13970) );
  NAND2_X1 U15964 ( .A1(n13971), .A2(n13970), .ZN(n13972) );
  AND2_X1 U15965 ( .A1(n14096), .A2(n13972), .ZN(n14010) );
  NAND2_X1 U15966 ( .A1(n14437), .A2(n14042), .ZN(n13974) );
  NAND2_X1 U15967 ( .A1(n14169), .A2(n6666), .ZN(n13973) );
  NAND2_X1 U15968 ( .A1(n13974), .A2(n13973), .ZN(n13975) );
  XNOR2_X1 U15969 ( .A(n13975), .B(n13985), .ZN(n13977) );
  AND2_X1 U15970 ( .A1(n14169), .A2(n14045), .ZN(n13976) );
  AOI21_X1 U15971 ( .B1(n14437), .B2(n6666), .A(n13976), .ZN(n13978) );
  NAND2_X1 U15972 ( .A1(n13977), .A2(n13978), .ZN(n13982) );
  INV_X1 U15973 ( .A(n13977), .ZN(n13980) );
  INV_X1 U15974 ( .A(n13978), .ZN(n13979) );
  NAND2_X1 U15975 ( .A1(n13980), .A2(n13979), .ZN(n13981) );
  NAND2_X1 U15976 ( .A1(n13982), .A2(n13981), .ZN(n14095) );
  INV_X1 U15977 ( .A(n13982), .ZN(n14065) );
  NAND2_X1 U15978 ( .A1(n14420), .A2(n14042), .ZN(n13984) );
  NAND2_X1 U15979 ( .A1(n14321), .A2(n6666), .ZN(n13983) );
  NAND2_X1 U15980 ( .A1(n13984), .A2(n13983), .ZN(n13986) );
  XNOR2_X1 U15981 ( .A(n13986), .B(n13985), .ZN(n13988) );
  AND2_X1 U15982 ( .A1(n14321), .A2(n14045), .ZN(n13987) );
  AOI21_X1 U15983 ( .B1(n14420), .B2(n6666), .A(n13987), .ZN(n13989) );
  NAND2_X1 U15984 ( .A1(n13988), .A2(n13989), .ZN(n13993) );
  INV_X1 U15985 ( .A(n13988), .ZN(n13991) );
  INV_X1 U15986 ( .A(n13989), .ZN(n13990) );
  NAND2_X1 U15987 ( .A1(n13991), .A2(n13990), .ZN(n13992) );
  AND2_X1 U15988 ( .A1(n13993), .A2(n13992), .ZN(n14064) );
  NAND2_X1 U15989 ( .A1(n14063), .A2(n13993), .ZN(n14140) );
  NAND2_X1 U15990 ( .A1(n14596), .A2(n14042), .ZN(n13995) );
  NAND2_X1 U15991 ( .A1(n14342), .A2(n6666), .ZN(n13994) );
  NAND2_X1 U15992 ( .A1(n13995), .A2(n13994), .ZN(n13996) );
  XNOR2_X1 U15993 ( .A(n13996), .B(n14043), .ZN(n14000) );
  NAND2_X1 U15994 ( .A1(n14596), .A2(n6666), .ZN(n13998) );
  NAND2_X1 U15995 ( .A1(n14342), .A2(n14045), .ZN(n13997) );
  NAND2_X1 U15996 ( .A1(n13998), .A2(n13997), .ZN(n13999) );
  NOR2_X1 U15997 ( .A1(n14000), .A2(n13999), .ZN(n14001) );
  AOI21_X1 U15998 ( .B1(n14000), .B2(n13999), .A(n14001), .ZN(n14141) );
  INV_X1 U15999 ( .A(n14001), .ZN(n14002) );
  NAND2_X1 U16000 ( .A1(n14139), .A2(n14002), .ZN(n14003) );
  NAND2_X1 U16001 ( .A1(n14003), .A2(n14004), .ZN(n14041) );
  OAI21_X1 U16002 ( .B1(n14004), .B2(n14003), .A(n14041), .ZN(n14005) );
  INV_X1 U16003 ( .A(n14005), .ZN(n14009) );
  AOI22_X1 U16004 ( .A1(n14346), .A2(n14281), .B1(n14521), .B2(n14342), .ZN(
        n14381) );
  AOI22_X1 U16005 ( .A1(n14387), .A2(n14124), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14006) );
  OAI21_X1 U16006 ( .B1(n14381), .B2(n14133), .A(n14006), .ZN(n14007) );
  AOI21_X1 U16007 ( .B1(n14589), .B2(n14163), .A(n14007), .ZN(n14008) );
  OAI21_X1 U16008 ( .B1(n14009), .B2(n14165), .A(n14008), .ZN(P1_U3214) );
  INV_X1 U16009 ( .A(n14452), .ZN(n14613) );
  INV_X1 U16010 ( .A(n14097), .ZN(n14013) );
  NOR3_X1 U16011 ( .A1(n14120), .A2(n14011), .A3(n14010), .ZN(n14012) );
  OAI21_X1 U16012 ( .B1(n14013), .B2(n14012), .A(n14142), .ZN(n14018) );
  AND2_X1 U16013 ( .A1(n14311), .A2(n14521), .ZN(n14014) );
  AOI21_X1 U16014 ( .B1(n14169), .B2(n14281), .A(n14014), .ZN(n14611) );
  OAI22_X1 U16015 ( .A1(n14611), .A2(n14133), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14015), .ZN(n14016) );
  AOI21_X1 U16016 ( .B1(n14451), .B2(n14124), .A(n14016), .ZN(n14017) );
  OAI211_X1 U16017 ( .C1(n14613), .C2(n14150), .A(n14018), .B(n14017), .ZN(
        P1_U3216) );
  AOI21_X1 U16018 ( .B1(n14020), .B2(n14019), .A(n14165), .ZN(n14022) );
  NAND2_X1 U16019 ( .A1(n14022), .A2(n14021), .ZN(n14029) );
  OR2_X1 U16020 ( .A1(n14023), .A2(n14156), .ZN(n14025) );
  NAND2_X1 U16021 ( .A1(n14181), .A2(n14521), .ZN(n14024) );
  NAND2_X1 U16022 ( .A1(n14025), .A2(n14024), .ZN(n15092) );
  AOI22_X1 U16023 ( .A1(n14163), .A2(n14026), .B1(n14159), .B2(n15092), .ZN(
        n14028) );
  MUX2_X1 U16024 ( .A(n14161), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n14027) );
  NAND3_X1 U16025 ( .A1(n14029), .A2(n14028), .A3(n14027), .ZN(P1_U3218) );
  INV_X1 U16026 ( .A(n14512), .ZN(n14638) );
  AND2_X1 U16027 ( .A1(n14128), .A2(n14030), .ZN(n14033) );
  OAI211_X1 U16028 ( .C1(n14033), .C2(n14032), .A(n14142), .B(n14031), .ZN(
        n14038) );
  INV_X1 U16029 ( .A(n14509), .ZN(n14036) );
  AND2_X1 U16030 ( .A1(n14330), .A2(n14521), .ZN(n14034) );
  AOI21_X1 U16031 ( .B1(n14334), .B2(n14281), .A(n14034), .ZN(n14637) );
  NAND2_X1 U16032 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14273)
         );
  OAI21_X1 U16033 ( .B1(n14637), .B2(n14133), .A(n14273), .ZN(n14035) );
  AOI21_X1 U16034 ( .B1(n14036), .B2(n14124), .A(n14035), .ZN(n14037) );
  OAI211_X1 U16035 ( .C1(n14638), .C2(n14150), .A(n14038), .B(n14037), .ZN(
        P1_U3219) );
  INV_X1 U16036 ( .A(n14039), .ZN(n14040) );
  NAND2_X1 U16037 ( .A1(n14041), .A2(n14040), .ZN(n14049) );
  AOI22_X1 U16038 ( .A1(n14583), .A2(n14042), .B1(n6666), .B2(n14346), .ZN(
        n14044) );
  XNOR2_X1 U16039 ( .A(n14044), .B(n14043), .ZN(n14047) );
  AOI22_X1 U16040 ( .A1(n14583), .A2(n6666), .B1(n14045), .B2(n14346), .ZN(
        n14046) );
  XNOR2_X1 U16041 ( .A(n14047), .B(n14046), .ZN(n14048) );
  XNOR2_X1 U16042 ( .A(n14049), .B(n14048), .ZN(n14053) );
  AOI22_X1 U16043 ( .A1(n14168), .A2(n14281), .B1(n14521), .B2(n14344), .ZN(
        n14366) );
  AOI22_X1 U16044 ( .A1(n14371), .A2(n14124), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14050) );
  OAI21_X1 U16045 ( .B1(n14366), .B2(n14133), .A(n14050), .ZN(n14051) );
  AOI21_X1 U16046 ( .B1(n14583), .B2(n14163), .A(n14051), .ZN(n14052) );
  OAI21_X1 U16047 ( .B1(n14053), .B2(n14165), .A(n14052), .ZN(P1_U3220) );
  INV_X1 U16048 ( .A(n14484), .ZN(n14627) );
  OAI21_X1 U16049 ( .B1(n14055), .B2(n14054), .A(n14118), .ZN(n14056) );
  NAND2_X1 U16050 ( .A1(n14056), .A2(n14142), .ZN(n14061) );
  AND2_X1 U16051 ( .A1(n14334), .A2(n14521), .ZN(n14057) );
  AOI21_X1 U16052 ( .B1(n14311), .B2(n14281), .A(n14057), .ZN(n14475) );
  OAI22_X1 U16053 ( .A1(n14475), .A2(n14133), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14058), .ZN(n14059) );
  AOI21_X1 U16054 ( .B1(n14483), .B2(n14124), .A(n14059), .ZN(n14060) );
  OAI211_X1 U16055 ( .C1(n14627), .C2(n14150), .A(n14061), .B(n14060), .ZN(
        P1_U3223) );
  INV_X1 U16056 ( .A(n14062), .ZN(n14106) );
  NAND2_X1 U16057 ( .A1(n14420), .A2(n15192), .ZN(n14604) );
  INV_X1 U16058 ( .A(n14063), .ZN(n14067) );
  NOR3_X1 U16059 ( .A1(n14099), .A2(n14065), .A3(n14064), .ZN(n14066) );
  OAI21_X1 U16060 ( .B1(n14067), .B2(n14066), .A(n14142), .ZN(n14072) );
  INV_X1 U16061 ( .A(n14342), .ZN(n14343) );
  OAI22_X1 U16062 ( .A1(n14343), .A2(n14156), .B1(n14315), .B2(n14357), .ZN(
        n14415) );
  INV_X1 U16063 ( .A(n14419), .ZN(n14069) );
  OAI22_X1 U16064 ( .A1(n14069), .A2(n14161), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14068), .ZN(n14070) );
  AOI21_X1 U16065 ( .B1(n14415), .B2(n14159), .A(n14070), .ZN(n14071) );
  OAI211_X1 U16066 ( .C1(n14106), .C2(n14604), .A(n14072), .B(n14071), .ZN(
        P1_U3225) );
  AOI21_X1 U16067 ( .B1(n14074), .B2(n14073), .A(n14086), .ZN(n14082) );
  OR2_X1 U16068 ( .A1(n14132), .A2(n14156), .ZN(n14076) );
  OR2_X1 U16069 ( .A1(n14294), .A2(n14357), .ZN(n14075) );
  AND2_X1 U16070 ( .A1(n14076), .A2(n14075), .ZN(n14554) );
  INV_X1 U16071 ( .A(n14077), .ZN(n14560) );
  NAND2_X1 U16072 ( .A1(n14124), .A2(n14560), .ZN(n14079) );
  OAI211_X1 U16073 ( .C1(n14554), .C2(n14133), .A(n14079), .B(n14078), .ZN(
        n14080) );
  AOI21_X1 U16074 ( .B1(n14656), .B2(n14163), .A(n14080), .ZN(n14081) );
  OAI21_X1 U16075 ( .B1(n14082), .B2(n14165), .A(n14081), .ZN(P1_U3226) );
  INV_X1 U16076 ( .A(n14650), .ZN(n14545) );
  INV_X1 U16077 ( .A(n14083), .ZN(n14088) );
  NOR3_X1 U16078 ( .A1(n14086), .A2(n14085), .A3(n14084), .ZN(n14087) );
  OAI21_X1 U16079 ( .B1(n14088), .B2(n14087), .A(n14142), .ZN(n14094) );
  OR2_X1 U16080 ( .A1(n14298), .A2(n14357), .ZN(n14090) );
  NAND2_X1 U16081 ( .A1(n14330), .A2(n14281), .ZN(n14089) );
  NAND2_X1 U16082 ( .A1(n14090), .A2(n14089), .ZN(n14538) );
  NOR2_X1 U16083 ( .A1(n14091), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14225) );
  NOR2_X1 U16084 ( .A1(n14161), .A2(n14542), .ZN(n14092) );
  AOI211_X1 U16085 ( .C1(n14159), .C2(n14538), .A(n14225), .B(n14092), .ZN(
        n14093) );
  OAI211_X1 U16086 ( .C1(n14545), .C2(n14150), .A(n14094), .B(n14093), .ZN(
        P1_U3228) );
  NAND2_X1 U16087 ( .A1(n14437), .A2(n15192), .ZN(n14609) );
  AND3_X1 U16088 ( .A1(n14097), .A2(n14096), .A3(n14095), .ZN(n14098) );
  OAI21_X1 U16089 ( .B1(n14099), .B2(n14098), .A(n14142), .ZN(n14105) );
  INV_X1 U16090 ( .A(n14100), .ZN(n14436) );
  AND2_X1 U16091 ( .A1(n14313), .A2(n14521), .ZN(n14101) );
  AOI21_X1 U16092 ( .B1(n14321), .B2(n14281), .A(n14101), .ZN(n14430) );
  OAI22_X1 U16093 ( .A1(n14430), .A2(n14133), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14102), .ZN(n14103) );
  AOI21_X1 U16094 ( .B1(n14436), .B2(n14124), .A(n14103), .ZN(n14104) );
  OAI211_X1 U16095 ( .C1(n14106), .C2(n14609), .A(n14105), .B(n14104), .ZN(
        P1_U3229) );
  XNOR2_X1 U16096 ( .A(n14108), .B(n14107), .ZN(n14115) );
  NOR2_X1 U16097 ( .A1(n14161), .A2(n14493), .ZN(n14113) );
  NOR2_X1 U16098 ( .A1(n14109), .A2(n14357), .ZN(n14110) );
  AOI21_X1 U16099 ( .B1(n14336), .B2(n14281), .A(n14110), .ZN(n14491) );
  OAI22_X1 U16100 ( .A1(n14491), .A2(n14133), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14111), .ZN(n14112) );
  AOI211_X1 U16101 ( .C1(n14499), .C2(n14163), .A(n14113), .B(n14112), .ZN(
        n14114) );
  OAI21_X1 U16102 ( .B1(n14115), .B2(n14165), .A(n14114), .ZN(P1_U3233) );
  AND3_X1 U16103 ( .A1(n14118), .A2(n14117), .A3(n14116), .ZN(n14119) );
  OAI21_X1 U16104 ( .B1(n14120), .B2(n14119), .A(n14142), .ZN(n14127) );
  INV_X1 U16105 ( .A(n14462), .ZN(n14125) );
  AND2_X1 U16106 ( .A1(n14336), .A2(n14521), .ZN(n14121) );
  AOI21_X1 U16107 ( .B1(n14313), .B2(n14281), .A(n14121), .ZN(n14618) );
  OAI22_X1 U16108 ( .A1(n14618), .A2(n14133), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14122), .ZN(n14123) );
  AOI21_X1 U16109 ( .B1(n14125), .B2(n14124), .A(n14123), .ZN(n14126) );
  OAI211_X1 U16110 ( .C1(n14150), .C2(n6906), .A(n14127), .B(n14126), .ZN(
        P1_U3235) );
  OAI21_X1 U16111 ( .B1(n14130), .B2(n14129), .A(n14128), .ZN(n14131) );
  NAND2_X1 U16112 ( .A1(n14131), .A2(n14142), .ZN(n14138) );
  INV_X1 U16113 ( .A(n14132), .ZN(n14522) );
  NAND2_X1 U16114 ( .A1(n14304), .A2(n14281), .ZN(n14523) );
  NAND2_X1 U16115 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14242)
         );
  OAI21_X1 U16116 ( .B1(n14523), .B2(n14133), .A(n14242), .ZN(n14135) );
  NOR2_X1 U16117 ( .A1(n14161), .A2(n14530), .ZN(n14134) );
  AOI211_X1 U16118 ( .C1(n14136), .C2(n14522), .A(n14135), .B(n14134), .ZN(
        n14137) );
  OAI211_X1 U16119 ( .C1(n14529), .C2(n14150), .A(n14138), .B(n14137), .ZN(
        P1_U3238) );
  INV_X1 U16120 ( .A(n14596), .ZN(n14407) );
  OAI21_X1 U16121 ( .B1(n14141), .B2(n14140), .A(n14139), .ZN(n14143) );
  NAND2_X1 U16122 ( .A1(n14143), .A2(n14142), .ZN(n14149) );
  NAND2_X1 U16123 ( .A1(n14344), .A2(n14281), .ZN(n14145) );
  NAND2_X1 U16124 ( .A1(n14321), .A2(n14521), .ZN(n14144) );
  NAND2_X1 U16125 ( .A1(n14145), .A2(n14144), .ZN(n14595) );
  OAI22_X1 U16126 ( .A1(n14403), .A2(n14161), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14146), .ZN(n14147) );
  AOI21_X1 U16127 ( .B1(n14595), .B2(n14159), .A(n14147), .ZN(n14148) );
  OAI211_X1 U16128 ( .C1(n14407), .C2(n14150), .A(n14149), .B(n14148), .ZN(
        P1_U3240) );
  AOI21_X1 U16129 ( .B1(n7386), .B2(n14152), .A(n14151), .ZN(n14153) );
  AOI21_X1 U16130 ( .B1(n14154), .B2(n7386), .A(n14153), .ZN(n14166) );
  NAND2_X1 U16131 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15066)
         );
  OR2_X1 U16132 ( .A1(n14155), .A2(n14357), .ZN(n14158) );
  OR2_X1 U16133 ( .A1(n14298), .A2(n14156), .ZN(n14157) );
  NAND2_X1 U16134 ( .A1(n14158), .A2(n14157), .ZN(n14953) );
  NAND2_X1 U16135 ( .A1(n14159), .A2(n14953), .ZN(n14160) );
  OAI211_X1 U16136 ( .C1(n14161), .C2(n14955), .A(n15066), .B(n14160), .ZN(
        n14162) );
  AOI21_X1 U16137 ( .B1(n14963), .B2(n14163), .A(n14162), .ZN(n14164) );
  OAI21_X1 U16138 ( .B1(n14166), .B2(n14165), .A(n14164), .ZN(P1_U3241) );
  MUX2_X1 U16139 ( .A(n14283), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14180), .Z(
        P1_U3591) );
  MUX2_X1 U16140 ( .A(n14167), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14180), .Z(
        P1_U3590) );
  MUX2_X1 U16141 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14168), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16142 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14346), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16143 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14344), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16144 ( .A(n14342), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14180), .Z(
        P1_U3586) );
  MUX2_X1 U16145 ( .A(n14321), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14180), .Z(
        P1_U3585) );
  MUX2_X1 U16146 ( .A(n14169), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14180), .Z(
        P1_U3584) );
  MUX2_X1 U16147 ( .A(n14313), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14180), .Z(
        P1_U3583) );
  MUX2_X1 U16148 ( .A(n14311), .B(P1_DATAO_REG_22__SCAN_IN), .S(n14180), .Z(
        P1_U3582) );
  MUX2_X1 U16149 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14336), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16150 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14334), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16151 ( .A(n14304), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14180), .Z(
        P1_U3579) );
  MUX2_X1 U16152 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14330), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16153 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14522), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16154 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14327), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16155 ( .A(n14170), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14180), .Z(
        P1_U3573) );
  MUX2_X1 U16156 ( .A(n14171), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14180), .Z(
        P1_U3572) );
  MUX2_X1 U16157 ( .A(n14172), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14180), .Z(
        P1_U3571) );
  MUX2_X1 U16158 ( .A(n14173), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14180), .Z(
        P1_U3570) );
  MUX2_X1 U16159 ( .A(n14174), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14180), .Z(
        P1_U3569) );
  MUX2_X1 U16160 ( .A(n14175), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14180), .Z(
        P1_U3568) );
  MUX2_X1 U16161 ( .A(n14176), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14180), .Z(
        P1_U3567) );
  MUX2_X1 U16162 ( .A(n14177), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14180), .Z(
        P1_U3566) );
  MUX2_X1 U16163 ( .A(n14178), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14180), .Z(
        P1_U3565) );
  MUX2_X1 U16164 ( .A(n14179), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14180), .Z(
        P1_U3563) );
  MUX2_X1 U16165 ( .A(n14181), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14180), .Z(
        P1_U3562) );
  MUX2_X1 U16166 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14182), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16167 ( .C1(n14185), .C2(n14184), .A(n15059), .B(n14183), .ZN(
        n14192) );
  NAND2_X1 U16168 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14194) );
  OAI211_X1 U16169 ( .C1(n10286), .C2(n14187), .A(n15046), .B(n14186), .ZN(
        n14191) );
  NAND2_X1 U16170 ( .A1(n15039), .A2(n14188), .ZN(n14190) );
  AOI22_X1 U16171 ( .A1(n15027), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14189) );
  NAND4_X1 U16172 ( .A1(n14192), .A2(n14191), .A3(n14190), .A4(n14189), .ZN(
        P1_U3244) );
  MUX2_X1 U16173 ( .A(n14194), .B(n14193), .S(n15020), .Z(n14199) );
  NAND2_X1 U16174 ( .A1(n14279), .A2(n14195), .ZN(n14196) );
  NAND2_X1 U16175 ( .A1(n14197), .A2(n14196), .ZN(n15021) );
  NAND2_X1 U16176 ( .A1(n15021), .A2(n14198), .ZN(n15024) );
  OAI211_X1 U16177 ( .C1(n14199), .C2(n10107), .A(P1_U4016), .B(n15024), .ZN(
        n15049) );
  AOI22_X1 U16178 ( .A1(n15027), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14211) );
  OAI21_X1 U16179 ( .B1(n14202), .B2(n14201), .A(n14200), .ZN(n14206) );
  XNOR2_X1 U16180 ( .A(n14204), .B(n14203), .ZN(n14205) );
  OAI22_X1 U16181 ( .A1(n15036), .A2(n14206), .B1(n15055), .B2(n14205), .ZN(
        n14207) );
  INV_X1 U16182 ( .A(n14207), .ZN(n14210) );
  OR2_X1 U16183 ( .A1(n15064), .A2(n14208), .ZN(n14209) );
  NAND4_X1 U16184 ( .A1(n15049), .A2(n14211), .A3(n14210), .A4(n14209), .ZN(
        P1_U3245) );
  OAI211_X1 U16185 ( .C1(n14213), .C2(n14212), .A(n15059), .B(n15033), .ZN(
        n14223) );
  MUX2_X1 U16186 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14214), .S(n14218), .Z(
        n14217) );
  INV_X1 U16187 ( .A(n14215), .ZN(n14216) );
  OAI211_X1 U16188 ( .C1(n14217), .C2(n14216), .A(n15046), .B(n15043), .ZN(
        n14222) );
  NAND2_X1 U16189 ( .A1(n15039), .A2(n14218), .ZN(n14221) );
  AND2_X1 U16190 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14219) );
  AOI21_X1 U16191 ( .B1(n15027), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14219), .ZN(
        n14220) );
  NAND4_X1 U16192 ( .A1(n14223), .A2(n14222), .A3(n14221), .A4(n14220), .ZN(
        P1_U3246) );
  NOR2_X1 U16193 ( .A1(n15064), .A2(n14246), .ZN(n14224) );
  AOI211_X1 U16194 ( .C1(n15027), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n14225), 
        .B(n14224), .ZN(n14241) );
  NAND2_X1 U16195 ( .A1(n14246), .A2(n14227), .ZN(n14226) );
  OAI21_X1 U16196 ( .B1(n14246), .B2(n14227), .A(n14226), .ZN(n14228) );
  INV_X1 U16197 ( .A(n14228), .ZN(n14232) );
  OAI21_X1 U16198 ( .B1(n14230), .B2(n12030), .A(n14229), .ZN(n14231) );
  NAND2_X1 U16199 ( .A1(n14232), .A2(n14231), .ZN(n14245) );
  OAI211_X1 U16200 ( .C1(n14232), .C2(n14231), .A(n15046), .B(n14245), .ZN(
        n14240) );
  XNOR2_X1 U16201 ( .A(n14246), .B(n14235), .ZN(n14236) );
  NOR2_X1 U16202 ( .A1(n14237), .A2(n14236), .ZN(n14248) );
  AOI211_X1 U16203 ( .C1(n14237), .C2(n14236), .A(n14248), .B(n15036), .ZN(
        n14238) );
  INV_X1 U16204 ( .A(n14238), .ZN(n14239) );
  NAND3_X1 U16205 ( .A1(n14241), .A2(n14240), .A3(n14239), .ZN(P1_U3260) );
  INV_X1 U16206 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14243) );
  OAI21_X1 U16207 ( .B1(n15068), .B2(n14243), .A(n14242), .ZN(n14244) );
  AOI21_X1 U16208 ( .B1(n14263), .B2(n15039), .A(n14244), .ZN(n14256) );
  OAI21_X1 U16209 ( .B1(n14227), .B2(n14246), .A(n14245), .ZN(n14262) );
  XNOR2_X1 U16210 ( .A(n14257), .B(n14262), .ZN(n14247) );
  NAND2_X1 U16211 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14247), .ZN(n14265) );
  OAI211_X1 U16212 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14247), .A(n15046), 
        .B(n14265), .ZN(n14255) );
  INV_X1 U16213 ( .A(n14250), .ZN(n14253) );
  INV_X1 U16214 ( .A(n14260), .ZN(n14252) );
  OAI211_X1 U16215 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14253), .A(n15059), 
        .B(n14252), .ZN(n14254) );
  NAND3_X1 U16216 ( .A1(n14256), .A2(n14255), .A3(n14254), .ZN(P1_U3261) );
  NOR2_X1 U16217 ( .A1(n14258), .A2(n14257), .ZN(n14259) );
  XNOR2_X1 U16218 ( .A(n14261), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14270) );
  INV_X1 U16219 ( .A(n14270), .ZN(n14268) );
  NAND2_X1 U16220 ( .A1(n14263), .A2(n14262), .ZN(n14264) );
  NAND2_X1 U16221 ( .A1(n14265), .A2(n14264), .ZN(n14266) );
  XOR2_X1 U16222 ( .A(n14266), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14269) );
  OAI21_X1 U16223 ( .B1(n14269), .B2(n15055), .A(n15064), .ZN(n14267) );
  AOI21_X1 U16224 ( .B1(n14268), .B2(n15059), .A(n14267), .ZN(n14272) );
  AOI22_X1 U16225 ( .A1(n14270), .A2(n15059), .B1(n15046), .B2(n14269), .ZN(
        n14271) );
  OAI211_X1 U16226 ( .C1(n7690), .C2(n15068), .A(n14274), .B(n14273), .ZN(
        P1_U3262) );
  INV_X1 U16227 ( .A(n14573), .ZN(n14276) );
  INV_X1 U16228 ( .A(n14589), .ZN(n14389) );
  INV_X1 U16229 ( .A(n14420), .ZN(n14418) );
  NAND2_X1 U16230 ( .A1(n14562), .A2(n14557), .ZN(n14558) );
  OR2_X2 U16231 ( .A1(n14495), .A2(n14484), .ZN(n14481) );
  NAND2_X1 U16232 ( .A1(n14389), .A2(n14401), .ZN(n14384) );
  XNOR2_X1 U16233 ( .A(n14277), .B(n14284), .ZN(n14278) );
  NAND2_X1 U16234 ( .A1(n14278), .A2(n15143), .ZN(n14568) );
  NAND2_X1 U16235 ( .A1(n14279), .A2(P1_B_REG_SCAN_IN), .ZN(n14280) );
  NAND2_X1 U16236 ( .A1(n14281), .A2(n14280), .ZN(n14351) );
  INV_X1 U16237 ( .A(n14351), .ZN(n14282) );
  NAND2_X1 U16238 ( .A1(n14283), .A2(n14282), .ZN(n14571) );
  NOR2_X1 U16239 ( .A1(n15096), .A2(n14571), .ZN(n14287) );
  INV_X1 U16240 ( .A(n14284), .ZN(n14569) );
  NOR2_X1 U16241 ( .A1(n14569), .A2(n15098), .ZN(n14285) );
  AOI211_X1 U16242 ( .C1(n15108), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14287), 
        .B(n14285), .ZN(n14286) );
  OAI21_X1 U16243 ( .B1(n14568), .B2(n14496), .A(n14286), .ZN(P1_U3263) );
  XNOR2_X1 U16244 ( .A(n14573), .B(n14349), .ZN(n14570) );
  NAND2_X1 U16245 ( .A1(n14570), .A2(n14550), .ZN(n14289) );
  AOI21_X1 U16246 ( .B1(n15096), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14287), 
        .ZN(n14288) );
  OAI211_X1 U16247 ( .C1(n14573), .C2(n15098), .A(n14289), .B(n14288), .ZN(
        P1_U3264) );
  NAND2_X1 U16248 ( .A1(n14292), .A2(n14291), .ZN(n14293) );
  INV_X1 U16249 ( .A(n14961), .ZN(n14325) );
  INV_X1 U16250 ( .A(n14294), .ZN(n14295) );
  OR2_X1 U16251 ( .A1(n14963), .A2(n14295), .ZN(n14296) );
  AND2_X1 U16252 ( .A1(n14562), .A2(n14298), .ZN(n14297) );
  OR2_X1 U16253 ( .A1(n14562), .A2(n14298), .ZN(n14299) );
  NAND2_X1 U16254 ( .A1(n14650), .A2(n14522), .ZN(n14301) );
  NAND2_X1 U16255 ( .A1(n14529), .A2(n14302), .ZN(n14303) );
  OR2_X1 U16256 ( .A1(n14512), .A2(n14304), .ZN(n14305) );
  INV_X1 U16257 ( .A(n14500), .ZN(n14307) );
  OR2_X1 U16258 ( .A1(n14634), .A2(n14309), .ZN(n14310) );
  INV_X1 U16259 ( .A(n14338), .ZN(n14468) );
  OR2_X1 U16260 ( .A1(n14461), .A2(n14311), .ZN(n14312) );
  NAND2_X1 U16261 ( .A1(n14452), .A2(n14313), .ZN(n14314) );
  NAND2_X1 U16262 ( .A1(n14420), .A2(n14321), .ZN(n14316) );
  NAND2_X1 U16263 ( .A1(n14596), .A2(n14342), .ZN(n14318) );
  INV_X1 U16264 ( .A(n14379), .ZN(n14391) );
  INV_X1 U16265 ( .A(n14321), .ZN(n14341) );
  INV_X1 U16266 ( .A(n14563), .ZN(n14552) );
  OR2_X1 U16267 ( .A1(n14562), .A2(n14327), .ZN(n14328) );
  NAND2_X1 U16268 ( .A1(n14529), .A2(n14330), .ZN(n14331) );
  NAND2_X1 U16269 ( .A1(n14634), .A2(n14334), .ZN(n14335) );
  NAND2_X1 U16270 ( .A1(n14429), .A2(n14428), .ZN(n14427) );
  INV_X1 U16271 ( .A(n14583), .ZN(n14345) );
  NOR2_X1 U16272 ( .A1(n14345), .A2(n14346), .ZN(n14347) );
  INV_X1 U16273 ( .A(n14346), .ZN(n14358) );
  NOR2_X1 U16274 ( .A1(n14578), .A2(n14350), .ZN(n14363) );
  NOR2_X1 U16275 ( .A1(n14352), .A2(n14351), .ZN(n14575) );
  INV_X1 U16276 ( .A(n14575), .ZN(n14354) );
  OAI22_X1 U16277 ( .A1(n14355), .A2(n15094), .B1(n14354), .B2(n14353), .ZN(
        n14356) );
  AOI21_X1 U16278 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n15108), .A(n14356), 
        .ZN(n14360) );
  NOR2_X1 U16279 ( .A1(n14358), .A2(n14357), .ZN(n14574) );
  NAND2_X1 U16280 ( .A1(n14574), .A2(n14532), .ZN(n14359) );
  OAI211_X1 U16281 ( .C1(n14361), .C2(n15098), .A(n14360), .B(n14359), .ZN(
        n14362) );
  AOI211_X1 U16282 ( .C1(n14579), .C2(n14516), .A(n14363), .B(n14362), .ZN(
        n14364) );
  OAI21_X1 U16283 ( .B1(n14580), .B2(n14564), .A(n14364), .ZN(P1_U3356) );
  XNOR2_X1 U16284 ( .A(n14365), .B(n14375), .ZN(n14368) );
  INV_X1 U16285 ( .A(n14366), .ZN(n14367) );
  AND2_X1 U16286 ( .A1(n14384), .A2(n14583), .ZN(n14369) );
  AOI22_X1 U16287 ( .A1(n14371), .A2(n14956), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15096), .ZN(n14373) );
  NAND2_X1 U16288 ( .A1(n14583), .A2(n14958), .ZN(n14372) );
  OAI211_X1 U16289 ( .C1(n14586), .C2(n14496), .A(n14373), .B(n14372), .ZN(
        n14374) );
  INV_X1 U16290 ( .A(n14374), .ZN(n14378) );
  NAND2_X1 U16291 ( .A1(n14376), .A2(n14375), .ZN(n14581) );
  NAND3_X1 U16292 ( .A1(n14582), .A2(n14967), .A3(n14581), .ZN(n14377) );
  OAI211_X1 U16293 ( .C1(n14587), .C2(n15096), .A(n14378), .B(n14377), .ZN(
        P1_U3265) );
  XNOR2_X1 U16294 ( .A(n14380), .B(n14379), .ZN(n14383) );
  INV_X1 U16295 ( .A(n14381), .ZN(n14382) );
  AOI21_X1 U16296 ( .B1(n14383), .B2(n15189), .A(n14382), .ZN(n14591) );
  INV_X1 U16297 ( .A(n14401), .ZN(n14386) );
  INV_X1 U16298 ( .A(n14384), .ZN(n14385) );
  AOI211_X1 U16299 ( .C1(n14589), .C2(n14386), .A(n15205), .B(n14385), .ZN(
        n14588) );
  AOI22_X1 U16300 ( .A1(n14387), .A2(n14956), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15096), .ZN(n14388) );
  OAI21_X1 U16301 ( .B1(n14389), .B2(n15098), .A(n14388), .ZN(n14393) );
  AOI21_X1 U16302 ( .B1(n14391), .B2(n14390), .A(n6748), .ZN(n14592) );
  NOR2_X1 U16303 ( .A1(n14592), .A2(n14564), .ZN(n14392) );
  AOI211_X1 U16304 ( .C1(n14588), .C2(n15104), .A(n14393), .B(n14392), .ZN(
        n14394) );
  OAI21_X1 U16305 ( .B1(n14591), .B2(n15096), .A(n14394), .ZN(P1_U3266) );
  XNOR2_X1 U16306 ( .A(n14395), .B(n14397), .ZN(n14593) );
  OAI21_X1 U16307 ( .B1(n14398), .B2(n14397), .A(n14396), .ZN(n14599) );
  NOR2_X1 U16308 ( .A1(n14599), .A2(n14564), .ZN(n14409) );
  NAND2_X1 U16309 ( .A1(n14596), .A2(n14417), .ZN(n14399) );
  NAND2_X1 U16310 ( .A1(n14399), .A2(n15143), .ZN(n14400) );
  NOR2_X1 U16311 ( .A1(n14401), .A2(n14400), .ZN(n14594) );
  NAND2_X1 U16312 ( .A1(n14594), .A2(n15104), .ZN(n14406) );
  INV_X1 U16313 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14402) );
  OAI22_X1 U16314 ( .A1(n14403), .A2(n15094), .B1(n14402), .B2(n14532), .ZN(
        n14404) );
  AOI21_X1 U16315 ( .B1(n14595), .B2(n14532), .A(n14404), .ZN(n14405) );
  OAI211_X1 U16316 ( .C1(n14407), .C2(n15098), .A(n14406), .B(n14405), .ZN(
        n14408) );
  AOI211_X1 U16317 ( .C1(n14593), .C2(n14516), .A(n14409), .B(n14408), .ZN(
        n14410) );
  INV_X1 U16318 ( .A(n14410), .ZN(P1_U3267) );
  AOI21_X1 U16319 ( .B1(n14413), .B2(n14412), .A(n14411), .ZN(n14414) );
  NOR2_X1 U16320 ( .A1(n14414), .A2(n15089), .ZN(n14416) );
  NOR2_X1 U16321 ( .A1(n14416), .A2(n14415), .ZN(n14605) );
  OAI211_X1 U16322 ( .C1(n14418), .C2(n14433), .A(n15143), .B(n14417), .ZN(
        n14602) );
  AOI22_X1 U16323 ( .A1(n14419), .A2(n14956), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15096), .ZN(n14422) );
  NAND2_X1 U16324 ( .A1(n14420), .A2(n14958), .ZN(n14421) );
  OAI211_X1 U16325 ( .C1(n14602), .C2(n14496), .A(n14422), .B(n14421), .ZN(
        n14423) );
  INV_X1 U16326 ( .A(n14423), .ZN(n14426) );
  NAND2_X1 U16327 ( .A1(n6782), .A2(n14424), .ZN(n14601) );
  NAND3_X1 U16328 ( .A1(n14601), .A2(n14967), .A3(n14600), .ZN(n14425) );
  OAI211_X1 U16329 ( .C1(n14605), .C2(n15096), .A(n14426), .B(n14425), .ZN(
        P1_U3268) );
  OAI211_X1 U16330 ( .C1(n14429), .C2(n14428), .A(n14427), .B(n15189), .ZN(
        n14431) );
  OAI21_X1 U16331 ( .B1(n6712), .B2(n14432), .A(n7603), .ZN(n14606) );
  INV_X1 U16332 ( .A(n14433), .ZN(n14434) );
  OAI211_X1 U16333 ( .C1(n14435), .C2(n6904), .A(n14434), .B(n15143), .ZN(
        n14607) );
  AOI22_X1 U16334 ( .A1(n14436), .A2(n14956), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15096), .ZN(n14439) );
  NAND2_X1 U16335 ( .A1(n14437), .A2(n14958), .ZN(n14438) );
  OAI211_X1 U16336 ( .C1(n14607), .C2(n14496), .A(n14439), .B(n14438), .ZN(
        n14440) );
  AOI21_X1 U16337 ( .B1(n14606), .B2(n14967), .A(n14440), .ZN(n14441) );
  OAI21_X1 U16338 ( .B1(n14610), .B2(n15108), .A(n14441), .ZN(P1_U3269) );
  AOI21_X1 U16339 ( .B1(n14443), .B2(n14442), .A(n6766), .ZN(n14617) );
  INV_X1 U16340 ( .A(n14516), .ZN(n14472) );
  INV_X1 U16341 ( .A(n14444), .ZN(n14445) );
  AOI21_X1 U16342 ( .B1(n7475), .B2(n14446), .A(n14445), .ZN(n14615) );
  INV_X1 U16343 ( .A(n14611), .ZN(n14450) );
  OAI211_X1 U16344 ( .C1(n14613), .C2(n14460), .A(n15143), .B(n14447), .ZN(
        n14612) );
  NOR2_X1 U16345 ( .A1(n14612), .A2(n14448), .ZN(n14449) );
  AOI211_X1 U16346 ( .C1(n14956), .C2(n14451), .A(n14450), .B(n14449), .ZN(
        n14454) );
  AOI22_X1 U16347 ( .A1(n14452), .A2(n14958), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15096), .ZN(n14453) );
  OAI21_X1 U16348 ( .B1(n14454), .B2(n15096), .A(n14453), .ZN(n14455) );
  AOI21_X1 U16349 ( .B1(n14615), .B2(n14967), .A(n14455), .ZN(n14456) );
  OAI21_X1 U16350 ( .B1(n14617), .B2(n14472), .A(n14456), .ZN(P1_U3270) );
  XNOR2_X1 U16351 ( .A(n14457), .B(n14468), .ZN(n14623) );
  NAND2_X1 U16352 ( .A1(n14461), .A2(n14481), .ZN(n14458) );
  NAND2_X1 U16353 ( .A1(n14458), .A2(n15143), .ZN(n14459) );
  NOR2_X1 U16354 ( .A1(n14460), .A2(n14459), .ZN(n14620) );
  NAND2_X1 U16355 ( .A1(n14461), .A2(n14958), .ZN(n14466) );
  OAI22_X1 U16356 ( .A1(n14618), .A2(n15096), .B1(n14462), .B2(n15094), .ZN(
        n14463) );
  INV_X1 U16357 ( .A(n14463), .ZN(n14465) );
  NAND2_X1 U16358 ( .A1(n15096), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n14464) );
  NAND3_X1 U16359 ( .A1(n14466), .A2(n14465), .A3(n14464), .ZN(n14467) );
  AOI21_X1 U16360 ( .B1(n14620), .B2(n15104), .A(n14467), .ZN(n14471) );
  XNOR2_X1 U16361 ( .A(n14469), .B(n14468), .ZN(n14621) );
  NAND2_X1 U16362 ( .A1(n14621), .A2(n14967), .ZN(n14470) );
  OAI211_X1 U16363 ( .C1(n14623), .C2(n14472), .A(n14471), .B(n14470), .ZN(
        P1_U3271) );
  XNOR2_X1 U16364 ( .A(n14473), .B(n7605), .ZN(n14474) );
  NAND2_X1 U16365 ( .A1(n14474), .A2(n15189), .ZN(n14476) );
  NAND2_X1 U16366 ( .A1(n14476), .A2(n14475), .ZN(n14629) );
  INV_X1 U16367 ( .A(n14629), .ZN(n14489) );
  NAND2_X1 U16368 ( .A1(n14478), .A2(n14477), .ZN(n14479) );
  NAND2_X1 U16369 ( .A1(n14480), .A2(n14479), .ZN(n14624) );
  AOI21_X1 U16370 ( .B1(n14495), .B2(n14484), .A(n15205), .ZN(n14482) );
  NAND2_X1 U16371 ( .A1(n14482), .A2(n14481), .ZN(n14625) );
  AOI22_X1 U16372 ( .A1(n15096), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14483), 
        .B2(n14956), .ZN(n14486) );
  NAND2_X1 U16373 ( .A1(n14484), .A2(n14958), .ZN(n14485) );
  OAI211_X1 U16374 ( .C1(n14625), .C2(n14496), .A(n14486), .B(n14485), .ZN(
        n14487) );
  AOI21_X1 U16375 ( .B1(n14624), .B2(n14967), .A(n14487), .ZN(n14488) );
  OAI21_X1 U16376 ( .B1(n14489), .B2(n15108), .A(n14488), .ZN(P1_U3272) );
  OAI211_X1 U16377 ( .C1(n7801), .C2(n14500), .A(n14490), .B(n15189), .ZN(
        n14492) );
  NAND2_X1 U16378 ( .A1(n14492), .A2(n14491), .ZN(n14636) );
  INV_X1 U16379 ( .A(n14636), .ZN(n14504) );
  INV_X1 U16380 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14494) );
  OAI22_X1 U16381 ( .A1(n14532), .A2(n14494), .B1(n14493), .B2(n15094), .ZN(
        n14498) );
  OAI211_X1 U16382 ( .C1(n14508), .C2(n14634), .A(n15143), .B(n14495), .ZN(
        n14632) );
  NOR2_X1 U16383 ( .A1(n14632), .A2(n14496), .ZN(n14497) );
  AOI211_X1 U16384 ( .C1(n14958), .C2(n14499), .A(n14498), .B(n14497), .ZN(
        n14503) );
  NAND2_X1 U16385 ( .A1(n7063), .A2(n14500), .ZN(n14630) );
  NAND3_X1 U16386 ( .A1(n14631), .A2(n14630), .A3(n14967), .ZN(n14502) );
  OAI211_X1 U16387 ( .C1(n14504), .C2(n15108), .A(n14503), .B(n14502), .ZN(
        P1_U3273) );
  XNOR2_X1 U16388 ( .A(n14505), .B(n14507), .ZN(n14643) );
  OAI21_X1 U16389 ( .B1(n6751), .B2(n14507), .A(n14506), .ZN(n14641) );
  AOI211_X1 U16390 ( .C1(n14512), .C2(n14527), .A(n15205), .B(n14508), .ZN(
        n14639) );
  OAI21_X1 U16391 ( .B1(n14509), .B2(n15094), .A(n14637), .ZN(n14510) );
  AOI21_X1 U16392 ( .B1(n14639), .B2(n14511), .A(n14510), .ZN(n14514) );
  AOI22_X1 U16393 ( .A1(n14512), .A2(n14958), .B1(P1_REG2_REG_19__SCAN_IN), 
        .B2(n15096), .ZN(n14513) );
  OAI21_X1 U16394 ( .B1(n14514), .B2(n15108), .A(n14513), .ZN(n14515) );
  AOI21_X1 U16395 ( .B1(n14516), .B2(n14641), .A(n14515), .ZN(n14517) );
  OAI21_X1 U16396 ( .B1(n14643), .B2(n14564), .A(n14517), .ZN(P1_U3274) );
  XNOR2_X1 U16397 ( .A(n14518), .B(n14520), .ZN(n14644) );
  XNOR2_X1 U16398 ( .A(n14519), .B(n14520), .ZN(n14525) );
  NAND2_X1 U16399 ( .A1(n14522), .A2(n14521), .ZN(n14524) );
  OAI211_X1 U16400 ( .C1(n14525), .C2(n15089), .A(n14524), .B(n14523), .ZN(
        n14526) );
  AOI21_X1 U16401 ( .B1(n15093), .B2(n14644), .A(n14526), .ZN(n14648) );
  INV_X1 U16402 ( .A(n14527), .ZN(n14528) );
  AOI211_X1 U16403 ( .C1(n14646), .C2(n14541), .A(n15205), .B(n14528), .ZN(
        n14645) );
  NOR2_X1 U16404 ( .A1(n14529), .A2(n15098), .ZN(n14534) );
  OAI22_X1 U16405 ( .A1(n14532), .A2(n14531), .B1(n14530), .B2(n15094), .ZN(
        n14533) );
  AOI211_X1 U16406 ( .C1(n14645), .C2(n15104), .A(n14534), .B(n14533), .ZN(
        n14536) );
  NAND2_X1 U16407 ( .A1(n14644), .A2(n15105), .ZN(n14535) );
  OAI211_X1 U16408 ( .C1(n14648), .C2(n15096), .A(n14536), .B(n14535), .ZN(
        P1_U3275) );
  AOI21_X1 U16409 ( .B1(n14537), .B2(n14546), .A(n15089), .ZN(n14540) );
  AOI21_X1 U16410 ( .B1(n14540), .B2(n14539), .A(n14538), .ZN(n14653) );
  AOI21_X1 U16411 ( .B1(n14650), .B2(n14558), .A(n7286), .ZN(n14651) );
  INV_X1 U16412 ( .A(n14542), .ZN(n14543) );
  AOI22_X1 U16413 ( .A1(n15108), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14543), 
        .B2(n14956), .ZN(n14544) );
  OAI21_X1 U16414 ( .B1(n14545), .B2(n15098), .A(n14544), .ZN(n14549) );
  XNOR2_X1 U16415 ( .A(n14547), .B(n14546), .ZN(n14654) );
  NOR2_X1 U16416 ( .A1(n14654), .A2(n14564), .ZN(n14548) );
  AOI211_X1 U16417 ( .C1(n14651), .C2(n14550), .A(n14549), .B(n14548), .ZN(
        n14551) );
  OAI21_X1 U16418 ( .B1(n15096), .B2(n14653), .A(n14551), .ZN(P1_U3276) );
  XNOR2_X1 U16419 ( .A(n14553), .B(n14552), .ZN(n14556) );
  INV_X1 U16420 ( .A(n14554), .ZN(n14555) );
  AOI21_X1 U16421 ( .B1(n14556), .B2(n15189), .A(n14555), .ZN(n14658) );
  INV_X1 U16422 ( .A(n14557), .ZN(n14964) );
  INV_X1 U16423 ( .A(n14558), .ZN(n14559) );
  AOI211_X1 U16424 ( .C1(n14656), .C2(n14964), .A(n15205), .B(n14559), .ZN(
        n14655) );
  AOI22_X1 U16425 ( .A1(n15096), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n14560), 
        .B2(n14956), .ZN(n14561) );
  OAI21_X1 U16426 ( .B1(n14562), .B2(n15098), .A(n14561), .ZN(n14566) );
  NOR2_X1 U16427 ( .A1(n14659), .A2(n14564), .ZN(n14565) );
  AOI211_X1 U16428 ( .C1(n14655), .C2(n15104), .A(n14566), .B(n14565), .ZN(
        n14567) );
  OAI21_X1 U16429 ( .B1(n15108), .B2(n14658), .A(n14567), .ZN(P1_U3277) );
  NAND2_X1 U16430 ( .A1(n14570), .A2(n15143), .ZN(n14572) );
  OAI211_X1 U16431 ( .C1(n14573), .C2(n15213), .A(n14572), .B(n14571), .ZN(
        n14661) );
  MUX2_X1 U16432 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14661), .S(n15233), .Z(
        P1_U3558) );
  AOI211_X1 U16433 ( .C1(n14576), .C2(n15192), .A(n14575), .B(n14574), .ZN(
        n14577) );
  MUX2_X1 U16434 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14662), .S(n15233), .Z(
        P1_U3557) );
  NAND3_X1 U16435 ( .A1(n14582), .A2(n15218), .A3(n14581), .ZN(n14585) );
  NAND2_X1 U16436 ( .A1(n14583), .A2(n15192), .ZN(n14584) );
  MUX2_X1 U16437 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14663), .S(n15233), .Z(
        P1_U3556) );
  AOI21_X1 U16438 ( .B1(n14589), .B2(n15192), .A(n14588), .ZN(n14590) );
  OAI211_X1 U16439 ( .C1(n15176), .C2(n14592), .A(n14591), .B(n14590), .ZN(
        n14664) );
  MUX2_X1 U16440 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14664), .S(n15233), .Z(
        P1_U3555) );
  NAND2_X1 U16441 ( .A1(n14593), .A2(n15189), .ZN(n14598) );
  AOI211_X1 U16442 ( .C1(n14596), .C2(n15192), .A(n14595), .B(n14594), .ZN(
        n14597) );
  OAI211_X1 U16443 ( .C1(n15176), .C2(n14599), .A(n14598), .B(n14597), .ZN(
        n14665) );
  MUX2_X1 U16444 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14665), .S(n15233), .Z(
        P1_U3554) );
  NAND3_X1 U16445 ( .A1(n14601), .A2(n15218), .A3(n14600), .ZN(n14603) );
  NAND4_X1 U16446 ( .A1(n14605), .A2(n14604), .A3(n14603), .A4(n14602), .ZN(
        n14666) );
  MUX2_X1 U16447 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14666), .S(n15233), .Z(
        P1_U3553) );
  NAND2_X1 U16448 ( .A1(n14606), .A2(n15218), .ZN(n14608) );
  NAND4_X1 U16449 ( .A1(n14610), .A2(n14609), .A3(n14608), .A4(n14607), .ZN(
        n14667) );
  MUX2_X1 U16450 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14667), .S(n15233), .Z(
        P1_U3552) );
  OAI211_X1 U16451 ( .C1(n14613), .C2(n15213), .A(n14612), .B(n14611), .ZN(
        n14614) );
  AOI21_X1 U16452 ( .B1(n14615), .B2(n15218), .A(n14614), .ZN(n14616) );
  OAI21_X1 U16453 ( .B1(n14617), .B2(n15089), .A(n14616), .ZN(n14668) );
  MUX2_X1 U16454 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14668), .S(n15233), .Z(
        P1_U3551) );
  OAI21_X1 U16455 ( .B1(n6906), .B2(n15213), .A(n14618), .ZN(n14619) );
  AOI211_X1 U16456 ( .C1(n14621), .C2(n15218), .A(n14620), .B(n14619), .ZN(
        n14622) );
  OAI21_X1 U16457 ( .B1(n14623), .B2(n15089), .A(n14622), .ZN(n14669) );
  MUX2_X1 U16458 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14669), .S(n15233), .Z(
        P1_U3550) );
  NAND2_X1 U16459 ( .A1(n14624), .A2(n15218), .ZN(n14626) );
  OAI211_X1 U16460 ( .C1(n14627), .C2(n15213), .A(n14626), .B(n14625), .ZN(
        n14628) );
  MUX2_X1 U16461 ( .A(n14670), .B(P1_REG1_REG_21__SCAN_IN), .S(n15231), .Z(
        P1_U3549) );
  NAND3_X1 U16462 ( .A1(n14631), .A2(n14630), .A3(n15218), .ZN(n14633) );
  OAI211_X1 U16463 ( .C1(n14634), .C2(n15213), .A(n14633), .B(n14632), .ZN(
        n14635) );
  MUX2_X1 U16464 ( .A(n14671), .B(P1_REG1_REG_20__SCAN_IN), .S(n15231), .Z(
        P1_U3548) );
  OAI21_X1 U16465 ( .B1(n14638), .B2(n15213), .A(n14637), .ZN(n14640) );
  AOI211_X1 U16466 ( .C1(n14641), .C2(n15189), .A(n14640), .B(n14639), .ZN(
        n14642) );
  OAI21_X1 U16467 ( .B1(n15176), .B2(n14643), .A(n14642), .ZN(n14672) );
  MUX2_X1 U16468 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14672), .S(n15233), .Z(
        P1_U3547) );
  INV_X1 U16469 ( .A(n14644), .ZN(n14649) );
  AOI21_X1 U16470 ( .B1(n14646), .B2(n15192), .A(n14645), .ZN(n14647) );
  OAI211_X1 U16471 ( .C1(n14649), .C2(n15197), .A(n14648), .B(n14647), .ZN(
        n14673) );
  MUX2_X1 U16472 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14673), .S(n15233), .Z(
        P1_U3546) );
  AOI22_X1 U16473 ( .A1(n14651), .A2(n15143), .B1(n14650), .B2(n15192), .ZN(
        n14652) );
  OAI211_X1 U16474 ( .C1(n15176), .C2(n14654), .A(n14653), .B(n14652), .ZN(
        n14674) );
  MUX2_X1 U16475 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14674), .S(n15233), .Z(
        P1_U3545) );
  AOI21_X1 U16476 ( .B1(n14656), .B2(n15192), .A(n14655), .ZN(n14657) );
  OAI211_X1 U16477 ( .C1(n15176), .C2(n14659), .A(n14658), .B(n14657), .ZN(
        n14675) );
  MUX2_X1 U16478 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14675), .S(n15233), .Z(
        P1_U3544) );
  MUX2_X1 U16479 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14660), .S(n15221), .Z(
        P1_U3527) );
  MUX2_X1 U16480 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14661), .S(n15221), .Z(
        P1_U3526) );
  MUX2_X1 U16481 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14662), .S(n15221), .Z(
        P1_U3525) );
  MUX2_X1 U16482 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14663), .S(n15221), .Z(
        P1_U3524) );
  MUX2_X1 U16483 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14664), .S(n15221), .Z(
        P1_U3523) );
  MUX2_X1 U16484 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14665), .S(n15221), .Z(
        P1_U3522) );
  MUX2_X1 U16485 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14666), .S(n15221), .Z(
        P1_U3521) );
  MUX2_X1 U16486 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14667), .S(n15221), .Z(
        P1_U3520) );
  MUX2_X1 U16487 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14668), .S(n15221), .Z(
        P1_U3519) );
  MUX2_X1 U16488 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14669), .S(n15221), .Z(
        P1_U3518) );
  MUX2_X1 U16489 ( .A(n14670), .B(P1_REG0_REG_21__SCAN_IN), .S(n15219), .Z(
        P1_U3517) );
  MUX2_X1 U16490 ( .A(n14671), .B(P1_REG0_REG_20__SCAN_IN), .S(n15219), .Z(
        P1_U3516) );
  MUX2_X1 U16491 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14672), .S(n15221), .Z(
        P1_U3515) );
  MUX2_X1 U16492 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14673), .S(n15221), .Z(
        P1_U3513) );
  MUX2_X1 U16493 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14674), .S(n15221), .Z(
        P1_U3510) );
  MUX2_X1 U16494 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14675), .S(n15221), .Z(
        P1_U3507) );
  NOR4_X1 U16495 ( .A1(n14677), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14676), .A4(
        P1_U3086), .ZN(n14678) );
  AOI21_X1 U16496 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14679), .A(n14678), 
        .ZN(n14680) );
  OAI21_X1 U16497 ( .B1(n14681), .B2(n14694), .A(n14680), .ZN(P1_U3324) );
  OAI222_X1 U16498 ( .A1(n15020), .A2(P1_U3086), .B1(n14694), .B2(n14686), 
        .C1(n14685), .C2(n14691), .ZN(P1_U3328) );
  OAI222_X1 U16499 ( .A1(P1_U3086), .A2(n14689), .B1(n14694), .B2(n14688), 
        .C1(n14687), .C2(n14691), .ZN(P1_U3329) );
  INV_X1 U16500 ( .A(n14690), .ZN(n14695) );
  OAI222_X1 U16501 ( .A1(n14695), .A2(P1_U3086), .B1(n14694), .B2(n14693), 
        .C1(n14692), .C2(n14691), .ZN(P1_U3330) );
  MUX2_X1 U16502 ( .A(n14697), .B(n14696), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16503 ( .A(n14698), .ZN(n14699) );
  MUX2_X1 U16504 ( .A(n14699), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16505 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15069) );
  NOR2_X1 U16506 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15069), .ZN(n14732) );
  INV_X1 U16507 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14731) );
  XNOR2_X1 U16508 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14791) );
  INV_X1 U16509 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14729) );
  INV_X1 U16510 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14726) );
  XNOR2_X1 U16511 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n14784) );
  INV_X1 U16512 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15852) );
  XNOR2_X1 U16513 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), 
        .ZN(n14751) );
  INV_X1 U16514 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15822) );
  XNOR2_X1 U16515 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n14753) );
  INV_X1 U16516 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14713) );
  XNOR2_X1 U16517 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14772) );
  NAND2_X1 U16518 ( .A1(n14757), .A2(n14758), .ZN(n14701) );
  NAND2_X1 U16519 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14702), .ZN(n14704) );
  INV_X1 U16520 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14703) );
  NAND2_X1 U16521 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14705), .ZN(n14707) );
  INV_X1 U16522 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15052) );
  NAND2_X1 U16523 ( .A1(n14755), .A2(n15052), .ZN(n14706) );
  NAND2_X1 U16524 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14708), .ZN(n14711) );
  INV_X1 U16525 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14709) );
  NAND2_X1 U16526 ( .A1(n14768), .A2(n14709), .ZN(n14710) );
  NAND2_X1 U16527 ( .A1(n14772), .A2(n14773), .ZN(n14712) );
  NAND2_X1 U16528 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14714), .ZN(n14717) );
  XOR2_X1 U16529 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14714), .Z(n14777) );
  INV_X1 U16530 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14715) );
  NAND2_X1 U16531 ( .A1(n14777), .A2(n14715), .ZN(n14716) );
  NAND2_X1 U16532 ( .A1(n14717), .A2(n14716), .ZN(n14754) );
  NAND2_X1 U16533 ( .A1(n14753), .A2(n14754), .ZN(n14718) );
  NAND2_X1 U16534 ( .A1(n14751), .A2(n14752), .ZN(n14719) );
  OAI21_X1 U16535 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15852), .A(n14719), .ZN(
        n14720) );
  INV_X1 U16536 ( .A(n14720), .ZN(n14721) );
  XNOR2_X1 U16537 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(P3_ADDR_REG_11__SCAN_IN), 
        .ZN(n14746) );
  NAND2_X1 U16538 ( .A1(n14747), .A2(n14746), .ZN(n14723) );
  NAND2_X1 U16539 ( .A1(n14784), .A2(n14785), .ZN(n14725) );
  NAND2_X1 U16540 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14727), .ZN(n14728) );
  NAND2_X1 U16541 ( .A1(n14791), .A2(n14790), .ZN(n14730) );
  OAI22_X1 U16542 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14743), .B1(n14732), 
        .B2(n14744), .ZN(n14733) );
  NOR2_X1 U16543 ( .A1(n14733), .A2(n12016), .ZN(n14735) );
  XOR2_X1 U16544 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n14733), .Z(n14793) );
  NOR2_X1 U16545 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14793), .ZN(n14734) );
  NOR2_X1 U16546 ( .A1(n14735), .A2(n14734), .ZN(n14736) );
  INV_X1 U16547 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14737) );
  NAND2_X1 U16548 ( .A1(n14736), .A2(n14737), .ZN(n14740) );
  XNOR2_X1 U16549 ( .A(n14737), .B(n14736), .ZN(n14796) );
  OR2_X1 U16550 ( .A1(n14738), .A2(n14796), .ZN(n14739) );
  NAND2_X1 U16551 ( .A1(n14740), .A2(n14739), .ZN(n15533) );
  NOR2_X1 U16552 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15536), .ZN(n14741) );
  AOI21_X1 U16553 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15536), .A(n14741), 
        .ZN(n15534) );
  XOR2_X1 U16554 ( .A(n15533), .B(n15534), .Z(n15919) );
  NOR2_X1 U16555 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14743), .ZN(n14742) );
  AOI21_X1 U16556 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n14743), .A(n14742), 
        .ZN(n14745) );
  XNOR2_X1 U16557 ( .A(n14745), .B(n14744), .ZN(n15012) );
  XOR2_X1 U16558 ( .A(n14747), .B(n14746), .Z(n14996) );
  NOR2_X1 U16559 ( .A1(n14749), .A2(n14748), .ZN(n14750) );
  XNOR2_X1 U16560 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14750), .ZN(n14782) );
  XOR2_X1 U16561 ( .A(n14752), .B(n14751), .Z(n14811) );
  XOR2_X1 U16562 ( .A(n14754), .B(n14753), .Z(n14807) );
  AND2_X1 U16563 ( .A1(n14766), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n14767) );
  XNOR2_X1 U16564 ( .A(n14756), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15934) );
  XOR2_X1 U16565 ( .A(n14758), .B(n14757), .Z(n14801) );
  INV_X1 U16566 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14762) );
  NOR2_X1 U16567 ( .A1(n14761), .A2(n14762), .ZN(n14763) );
  AOI21_X1 U16568 ( .B1(n15861), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n14759), .ZN(
        n15928) );
  INV_X1 U16569 ( .A(n15928), .ZN(n14760) );
  NAND2_X1 U16570 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n14760), .ZN(n15938) );
  XNOR2_X1 U16571 ( .A(n14762), .B(n14761), .ZN(n15937) );
  NOR2_X1 U16572 ( .A1(n15938), .A2(n15937), .ZN(n15936) );
  NOR2_X1 U16573 ( .A1(n14801), .A2(n14800), .ZN(n14764) );
  NAND2_X1 U16574 ( .A1(n14801), .A2(n14800), .ZN(n14799) );
  NAND2_X1 U16575 ( .A1(n15934), .A2(n15933), .ZN(n14765) );
  NOR2_X1 U16576 ( .A1(n15934), .A2(n15933), .ZN(n15932) );
  NOR2_X1 U16577 ( .A1(n15924), .A2(n15923), .ZN(n15922) );
  XNOR2_X1 U16578 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14768), .ZN(n14770) );
  NAND2_X1 U16579 ( .A1(n14769), .A2(n14770), .ZN(n14771) );
  INV_X1 U16580 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15926) );
  NOR2_X1 U16581 ( .A1(n14775), .A2(n14774), .ZN(n14776) );
  XOR2_X1 U16582 ( .A(n14773), .B(n14772), .Z(n14805) );
  NAND2_X1 U16583 ( .A1(n14778), .A2(n13419), .ZN(n14779) );
  XNOR2_X1 U16584 ( .A(n14777), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15931) );
  NAND2_X1 U16585 ( .A1(n14807), .A2(n14808), .ZN(n14806) );
  INV_X1 U16586 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14818) );
  NAND2_X1 U16587 ( .A1(n14996), .A2(n14995), .ZN(n14783) );
  XOR2_X1 U16588 ( .A(n14785), .B(n14784), .Z(n14999) );
  XOR2_X1 U16589 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .Z(n14786) );
  XOR2_X1 U16590 ( .A(n14787), .B(n14786), .Z(n14788) );
  INV_X1 U16591 ( .A(n15003), .ZN(n15004) );
  INV_X1 U16592 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15006) );
  NAND2_X1 U16593 ( .A1(n14789), .A2(n14788), .ZN(n15005) );
  NAND2_X1 U16594 ( .A1(n15006), .A2(n15005), .ZN(n15002) );
  XNOR2_X1 U16595 ( .A(n14791), .B(n14790), .ZN(n15008) );
  NOR2_X1 U16596 ( .A1(n15009), .A2(n15008), .ZN(n14792) );
  NAND2_X1 U16597 ( .A1(n15009), .A2(n15008), .ZN(n15007) );
  XOR2_X1 U16598 ( .A(n14794), .B(n14793), .Z(n15016) );
  NAND2_X1 U16599 ( .A1(n15017), .A2(n15016), .ZN(n14795) );
  XNOR2_X1 U16600 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14796), .ZN(n14828) );
  NOR2_X1 U16601 ( .A1(n14829), .A2(n14828), .ZN(n14797) );
  NAND2_X1 U16602 ( .A1(n14829), .A2(n14828), .ZN(n14827) );
  AOI21_X1 U16603 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14798) );
  OAI21_X1 U16604 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14798), 
        .ZN(U28) );
  OAI21_X1 U16605 ( .B1(n14801), .B2(n14800), .A(n14799), .ZN(n14802) );
  XNOR2_X1 U16606 ( .A(n14802), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16607 ( .B1(n14805), .B2(n14804), .A(n14803), .ZN(SUB_1596_U57) );
  OAI21_X1 U16608 ( .B1(n14808), .B2(n14807), .A(n14806), .ZN(n14809) );
  XNOR2_X1 U16609 ( .A(n14809), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  OAI21_X1 U16610 ( .B1(n14812), .B2(n14811), .A(n14810), .ZN(n14813) );
  XNOR2_X1 U16611 ( .A(n14813), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  OAI222_X1 U16612 ( .A1(n14818), .A2(n14817), .B1(n14818), .B2(n14816), .C1(
        n14815), .C2(n14814), .ZN(SUB_1596_U70) );
  NAND2_X1 U16613 ( .A1(n14819), .A2(n15192), .ZN(n14820) );
  OAI211_X1 U16614 ( .C1(n14822), .C2(n15197), .A(n14821), .B(n14820), .ZN(
        n14823) );
  NOR2_X1 U16615 ( .A1(n14824), .A2(n14823), .ZN(n14826) );
  INV_X1 U16616 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14825) );
  AOI22_X1 U16617 ( .A1(n15221), .A2(n14826), .B1(n14825), .B2(n15219), .ZN(
        P1_U3495) );
  AOI22_X1 U16618 ( .A1(n15233), .A2(n14826), .B1(n9752), .B2(n15231), .ZN(
        P1_U3540) );
  OAI21_X1 U16619 ( .B1(n14829), .B2(n14828), .A(n14827), .ZN(n14830) );
  XNOR2_X1 U16620 ( .A(n14830), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  XNOR2_X1 U16621 ( .A(n14832), .B(n14831), .ZN(n14834) );
  AOI222_X1 U16622 ( .A1(n15453), .A2(n14834), .B1(n14833), .B2(n15398), .C1(
        n14856), .C2(n15447), .ZN(n14867) );
  AOI22_X1 U16623 ( .A1(n15465), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15442), 
        .B2(n14835), .ZN(n14840) );
  XNOR2_X1 U16624 ( .A(n14837), .B(n14836), .ZN(n14870) );
  NOR2_X1 U16625 ( .A1(n14838), .A2(n15512), .ZN(n14869) );
  AOI22_X1 U16626 ( .A1(n14870), .A2(n14864), .B1(n14869), .B2(n15419), .ZN(
        n14839) );
  OAI211_X1 U16627 ( .C1(n15465), .C2(n14867), .A(n14840), .B(n14839), .ZN(
        P3_U3219) );
  XNOR2_X1 U16628 ( .A(n6827), .B(n14841), .ZN(n14842) );
  NAND2_X1 U16629 ( .A1(n14842), .A2(n15453), .ZN(n14846) );
  AOI22_X1 U16630 ( .A1(n14844), .A2(n15447), .B1(n15398), .B2(n14843), .ZN(
        n14845) );
  NAND2_X1 U16631 ( .A1(n14846), .A2(n14845), .ZN(n14874) );
  OAI22_X1 U16632 ( .A1(n8876), .A2(n15463), .B1(n15458), .B2(n14847), .ZN(
        n14853) );
  XNOR2_X1 U16633 ( .A(n14849), .B(n14848), .ZN(n14871) );
  AND2_X1 U16634 ( .A1(n14850), .A2(n15495), .ZN(n14872) );
  AOI22_X1 U16635 ( .A1(n14871), .A2(n14864), .B1(n14872), .B2(n15419), .ZN(
        n14851) );
  INV_X1 U16636 ( .A(n14851), .ZN(n14852) );
  AOI211_X1 U16637 ( .C1(n15463), .C2(n14874), .A(n14853), .B(n14852), .ZN(
        n14854) );
  INV_X1 U16638 ( .A(n14854), .ZN(P3_U3220) );
  XOR2_X1 U16639 ( .A(n14861), .B(n14855), .Z(n14858) );
  AOI222_X1 U16640 ( .A1(n15453), .A2(n14858), .B1(n14857), .B2(n15447), .C1(
        n14856), .C2(n15398), .ZN(n14875) );
  AOI22_X1 U16641 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n15465), .B1(n15442), 
        .B2(n14859), .ZN(n14866) );
  OAI21_X1 U16642 ( .B1(n14862), .B2(n14861), .A(n14860), .ZN(n14878) );
  NOR2_X1 U16643 ( .A1(n14863), .A2(n15512), .ZN(n14877) );
  AOI22_X1 U16644 ( .A1(n14878), .A2(n14864), .B1(n14877), .B2(n15419), .ZN(
        n14865) );
  OAI211_X1 U16645 ( .C1(n15465), .C2(n14875), .A(n14866), .B(n14865), .ZN(
        P3_U3221) );
  INV_X1 U16646 ( .A(n14867), .ZN(n14868) );
  AOI211_X1 U16647 ( .C1(n15515), .C2(n14870), .A(n14869), .B(n14868), .ZN(
        n14882) );
  AOI22_X1 U16648 ( .A1(n15532), .A2(n14882), .B1(n8896), .B2(n15530), .ZN(
        P3_U3473) );
  AND2_X1 U16649 ( .A1(n14871), .A2(n15515), .ZN(n14873) );
  NOR3_X1 U16650 ( .A1(n14874), .A2(n14873), .A3(n14872), .ZN(n14884) );
  AOI22_X1 U16651 ( .A1(n15532), .A2(n14884), .B1(n8877), .B2(n15530), .ZN(
        P3_U3472) );
  INV_X1 U16652 ( .A(n14875), .ZN(n14876) );
  AOI211_X1 U16653 ( .C1(n15515), .C2(n14878), .A(n14877), .B(n14876), .ZN(
        n14885) );
  AOI22_X1 U16654 ( .A1(n15532), .A2(n14885), .B1(n11946), .B2(n15530), .ZN(
        P3_U3471) );
  AOI211_X1 U16655 ( .C1(n15515), .C2(n14881), .A(n14880), .B(n14879), .ZN(
        n14887) );
  AOI22_X1 U16656 ( .A1(n15532), .A2(n14887), .B1(n8828), .B2(n15530), .ZN(
        P3_U3470) );
  AOI22_X1 U16657 ( .A1(n15519), .A2(n14882), .B1(n8895), .B2(n15517), .ZN(
        P3_U3432) );
  INV_X1 U16658 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14883) );
  AOI22_X1 U16659 ( .A1(n15519), .A2(n14884), .B1(n14883), .B2(n15517), .ZN(
        P3_U3429) );
  AOI22_X1 U16660 ( .A1(n15519), .A2(n14885), .B1(n8858), .B2(n15517), .ZN(
        P3_U3426) );
  INV_X1 U16661 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14886) );
  AOI22_X1 U16662 ( .A1(n15519), .A2(n14887), .B1(n14886), .B2(n15517), .ZN(
        P3_U3423) );
  NAND2_X1 U16663 ( .A1(n14889), .A2(n14888), .ZN(n14890) );
  NAND2_X1 U16664 ( .A1(n14900), .A2(n14890), .ZN(n14891) );
  AOI222_X1 U16665 ( .A1(n14908), .A2(n14893), .B1(n14892), .B2(n14905), .C1(
        n14891), .C2(n14903), .ZN(n14895) );
  OAI211_X1 U16666 ( .C1(n14911), .C2(n14896), .A(n14895), .B(n14894), .ZN(
        P2_U3198) );
  INV_X1 U16667 ( .A(n14897), .ZN(n14899) );
  NAND3_X1 U16668 ( .A1(n14900), .A2(n14899), .A3(n14898), .ZN(n14901) );
  NAND2_X1 U16669 ( .A1(n14902), .A2(n14901), .ZN(n14904) );
  AOI222_X1 U16670 ( .A1(n14908), .A2(n14907), .B1(n14906), .B2(n14905), .C1(
        n14904), .C2(n14903), .ZN(n14909) );
  NAND2_X1 U16671 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n15313)
         );
  OAI211_X1 U16672 ( .C1(n14911), .C2(n14910), .A(n14909), .B(n15313), .ZN(
        P2_U3200) );
  XNOR2_X1 U16673 ( .A(n14913), .B(n14912), .ZN(n14916) );
  AOI21_X1 U16674 ( .B1(n14916), .B2(n14915), .A(n14914), .ZN(n14938) );
  AOI222_X1 U16675 ( .A1(n14921), .A2(n14920), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n14919), .C1(n14918), .C2(n14917), .ZN(n14934) );
  INV_X1 U16676 ( .A(n14922), .ZN(n14923) );
  AOI21_X1 U16677 ( .B1(n14925), .B2(n14924), .A(n14923), .ZN(n14942) );
  INV_X1 U16678 ( .A(n14926), .ZN(n14929) );
  OAI211_X1 U16679 ( .C1(n14937), .C2(n14929), .A(n14928), .B(n14927), .ZN(
        n14936) );
  INV_X1 U16680 ( .A(n14936), .ZN(n14930) );
  AOI22_X1 U16681 ( .A1(n14942), .A2(n14932), .B1(n14931), .B2(n14930), .ZN(
        n14933) );
  OAI211_X1 U16682 ( .C1(n14935), .C2(n14938), .A(n14934), .B(n14933), .ZN(
        P2_U3251) );
  OAI21_X1 U16683 ( .B1(n14937), .B2(n15381), .A(n14936), .ZN(n14940) );
  INV_X1 U16684 ( .A(n14938), .ZN(n14939) );
  AOI211_X1 U16685 ( .C1(n14942), .C2(n14941), .A(n14940), .B(n14939), .ZN(
        n14949) );
  AOI22_X1 U16686 ( .A1(n15391), .A2(n14949), .B1(n13448), .B2(n15389), .ZN(
        P2_U3513) );
  INV_X1 U16687 ( .A(n14943), .ZN(n14948) );
  OAI21_X1 U16688 ( .B1(n14945), .B2(n15381), .A(n14944), .ZN(n14947) );
  AOI22_X1 U16689 ( .A1(n15391), .A2(n14951), .B1(n10828), .B2(n15389), .ZN(
        P2_U3511) );
  AOI22_X1 U16690 ( .A1(n15387), .A2(n14949), .B1(n8205), .B2(n15386), .ZN(
        P2_U3472) );
  INV_X1 U16691 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14950) );
  AOI22_X1 U16692 ( .A1(n15387), .A2(n14951), .B1(n14950), .B2(n15386), .ZN(
        P2_U3466) );
  XNOR2_X1 U16693 ( .A(n14952), .B(n14961), .ZN(n14954) );
  AOI21_X1 U16694 ( .B1(n14954), .B2(n15189), .A(n14953), .ZN(n14972) );
  INV_X1 U16695 ( .A(n14955), .ZN(n14957) );
  AOI222_X1 U16696 ( .A1(n14963), .A2(n14958), .B1(n14957), .B2(n14956), .C1(
        P1_REG2_REG_15__SCAN_IN), .C2(n15108), .ZN(n14969) );
  INV_X1 U16697 ( .A(n14959), .ZN(n14962) );
  OAI21_X1 U16698 ( .B1(n14962), .B2(n14961), .A(n14960), .ZN(n14975) );
  INV_X1 U16699 ( .A(n14963), .ZN(n14971) );
  OAI211_X1 U16700 ( .C1(n14971), .C2(n14965), .A(n14964), .B(n15143), .ZN(
        n14970) );
  INV_X1 U16701 ( .A(n14970), .ZN(n14966) );
  AOI22_X1 U16702 ( .A1(n14975), .A2(n14967), .B1(n15104), .B2(n14966), .ZN(
        n14968) );
  OAI211_X1 U16703 ( .C1(n15108), .C2(n14972), .A(n14969), .B(n14968), .ZN(
        P1_U3278) );
  OAI21_X1 U16704 ( .B1(n14971), .B2(n15213), .A(n14970), .ZN(n14974) );
  INV_X1 U16705 ( .A(n14972), .ZN(n14973) );
  AOI211_X1 U16706 ( .C1(n15218), .C2(n14975), .A(n14974), .B(n14973), .ZN(
        n14989) );
  AOI22_X1 U16707 ( .A1(n15233), .A2(n14989), .B1(n9799), .B2(n15231), .ZN(
        P1_U3543) );
  INV_X1 U16708 ( .A(n14976), .ZN(n14978) );
  OAI21_X1 U16709 ( .B1(n14978), .B2(n15213), .A(n14977), .ZN(n14979) );
  AOI21_X1 U16710 ( .B1(n14980), .B2(n15218), .A(n14979), .ZN(n14981) );
  AND2_X1 U16711 ( .A1(n14982), .A2(n14981), .ZN(n14991) );
  AOI22_X1 U16712 ( .A1(n15233), .A2(n14991), .B1(n11248), .B2(n15231), .ZN(
        P1_U3541) );
  OAI21_X1 U16713 ( .B1(n14984), .B2(n15213), .A(n14983), .ZN(n14985) );
  AOI21_X1 U16714 ( .B1(n14986), .B2(n15218), .A(n14985), .ZN(n14987) );
  AND2_X1 U16715 ( .A1(n14988), .A2(n14987), .ZN(n14993) );
  AOI22_X1 U16716 ( .A1(n15233), .A2(n14993), .B1(n10594), .B2(n15231), .ZN(
        P1_U3539) );
  AOI22_X1 U16717 ( .A1(n15221), .A2(n14989), .B1(n9794), .B2(n15219), .ZN(
        P1_U3504) );
  INV_X1 U16718 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14990) );
  AOI22_X1 U16719 ( .A1(n15221), .A2(n14991), .B1(n14990), .B2(n15219), .ZN(
        P1_U3498) );
  INV_X1 U16720 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U16721 ( .A1(n15221), .A2(n14993), .B1(n14992), .B2(n15219), .ZN(
        P1_U3492) );
  AOI21_X1 U16722 ( .B1(n14996), .B2(n14995), .A(n14994), .ZN(n14997) );
  XOR2_X1 U16723 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14997), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16724 ( .B1(n15000), .B2(n14999), .A(n14998), .ZN(n15001) );
  XNOR2_X1 U16725 ( .A(n15001), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  OAI222_X1 U16726 ( .A1(n15006), .A2(n15005), .B1(n15006), .B2(n15004), .C1(
        n15003), .C2(n15002), .ZN(SUB_1596_U67) );
  OAI21_X1 U16727 ( .B1(n15009), .B2(n15008), .A(n15007), .ZN(n15010) );
  XNOR2_X1 U16728 ( .A(n15010), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U16729 ( .B1(n15013), .B2(n15012), .A(n15011), .ZN(n15014) );
  XNOR2_X1 U16730 ( .A(n15014), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  AOI21_X1 U16731 ( .B1(n15017), .B2(n15016), .A(n15015), .ZN(n15018) );
  XOR2_X1 U16732 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n15018), .Z(SUB_1596_U64)
         );
  AND2_X1 U16733 ( .A1(n15020), .A2(n15019), .ZN(n15023) );
  NOR2_X1 U16734 ( .A1(n15021), .A2(n15023), .ZN(n15022) );
  MUX2_X1 U16735 ( .A(n15023), .B(n15022), .S(P1_IR_REG_0__SCAN_IN), .Z(n15026) );
  INV_X1 U16736 ( .A(n15024), .ZN(n15025) );
  OR2_X1 U16737 ( .A1(n15026), .A2(n15025), .ZN(n15029) );
  AOI22_X1 U16738 ( .A1(n15027), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15028) );
  OAI21_X1 U16739 ( .B1(n15030), .B2(n15029), .A(n15028), .ZN(P1_U3243) );
  AND3_X1 U16740 ( .A1(n15033), .A2(n15032), .A3(n15031), .ZN(n15034) );
  NOR3_X1 U16741 ( .A1(n15036), .A2(n15035), .A3(n15034), .ZN(n15037) );
  AOI21_X1 U16742 ( .B1(n15039), .B2(n15038), .A(n15037), .ZN(n15048) );
  INV_X1 U16743 ( .A(n15040), .ZN(n15045) );
  NAND3_X1 U16744 ( .A1(n15043), .A2(n15042), .A3(n15041), .ZN(n15044) );
  NAND3_X1 U16745 ( .A1(n15046), .A2(n15045), .A3(n15044), .ZN(n15047) );
  AND3_X1 U16746 ( .A1(n15049), .A2(n15048), .A3(n15047), .ZN(n15051) );
  NAND2_X1 U16747 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15050) );
  OAI211_X1 U16748 ( .C1(n15052), .C2(n15068), .A(n15051), .B(n15050), .ZN(
        P1_U3247) );
  AOI21_X1 U16749 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n15054), .A(n15053), 
        .ZN(n15056) );
  OR2_X1 U16750 ( .A1(n15056), .A2(n15055), .ZN(n15062) );
  OAI21_X1 U16751 ( .B1(n15058), .B2(n9799), .A(n15057), .ZN(n15060) );
  NAND2_X1 U16752 ( .A1(n15060), .A2(n15059), .ZN(n15061) );
  OAI211_X1 U16753 ( .C1(n15064), .C2(n15063), .A(n15062), .B(n15061), .ZN(
        n15065) );
  INV_X1 U16754 ( .A(n15065), .ZN(n15067) );
  OAI211_X1 U16755 ( .C1(n15069), .C2(n15068), .A(n15067), .B(n15066), .ZN(
        P1_U3258) );
  XNOR2_X1 U16756 ( .A(n15070), .B(n15071), .ZN(n15075) );
  XNOR2_X1 U16757 ( .A(n15072), .B(n15071), .ZN(n15196) );
  OAI21_X1 U16758 ( .B1(n15196), .B2(n15187), .A(n15073), .ZN(n15074) );
  AOI21_X1 U16759 ( .B1(n15189), .B2(n15075), .A(n15074), .ZN(n15195) );
  INV_X1 U16760 ( .A(n15193), .ZN(n15079) );
  NOR2_X1 U16761 ( .A1(n15094), .A2(n15076), .ZN(n15077) );
  AOI21_X1 U16762 ( .B1(n15108), .B2(P1_REG2_REG_7__SCAN_IN), .A(n15077), .ZN(
        n15078) );
  OAI21_X1 U16763 ( .B1(n15098), .B2(n15079), .A(n15078), .ZN(n15080) );
  INV_X1 U16764 ( .A(n15080), .ZN(n15085) );
  INV_X1 U16765 ( .A(n15196), .ZN(n15083) );
  AOI211_X1 U16766 ( .C1(n15193), .C2(n15082), .A(n15205), .B(n15081), .ZN(
        n15191) );
  AOI22_X1 U16767 ( .A1(n15083), .A2(n15105), .B1(n15104), .B2(n15191), .ZN(
        n15084) );
  OAI211_X1 U16768 ( .C1(n15108), .C2(n15195), .A(n15085), .B(n15084), .ZN(
        P1_U3286) );
  XNOR2_X1 U16769 ( .A(n15086), .B(n15088), .ZN(n15163) );
  XNOR2_X1 U16770 ( .A(n15088), .B(n15087), .ZN(n15090) );
  NOR2_X1 U16771 ( .A1(n15090), .A2(n15089), .ZN(n15091) );
  AOI211_X1 U16772 ( .C1(n15093), .C2(n15163), .A(n15092), .B(n15091), .ZN(
        n15160) );
  NOR2_X1 U16773 ( .A1(n15094), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n15095) );
  AOI21_X1 U16774 ( .B1(n15096), .B2(P1_REG2_REG_3__SCAN_IN), .A(n15095), .ZN(
        n15097) );
  OAI21_X1 U16775 ( .B1(n15098), .B2(n15159), .A(n15097), .ZN(n15099) );
  INV_X1 U16776 ( .A(n15099), .ZN(n15107) );
  INV_X1 U16777 ( .A(n15101), .ZN(n15102) );
  OAI211_X1 U16778 ( .C1(n15159), .C2(n6902), .A(n15102), .B(n15143), .ZN(
        n15158) );
  INV_X1 U16779 ( .A(n15158), .ZN(n15103) );
  AOI22_X1 U16780 ( .A1(n15163), .A2(n15105), .B1(n15104), .B2(n15103), .ZN(
        n15106) );
  OAI211_X1 U16781 ( .C1(n15108), .C2(n15160), .A(n15107), .B(n15106), .ZN(
        P1_U3290) );
  INV_X1 U16782 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15109) );
  NOR2_X1 U16783 ( .A1(n15139), .A2(n15109), .ZN(P1_U3294) );
  INV_X1 U16784 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15110) );
  NOR2_X1 U16785 ( .A1(n15139), .A2(n15110), .ZN(P1_U3295) );
  INV_X1 U16786 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15111) );
  NOR2_X1 U16787 ( .A1(n15139), .A2(n15111), .ZN(P1_U3296) );
  INV_X1 U16788 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15112) );
  NOR2_X1 U16789 ( .A1(n15139), .A2(n15112), .ZN(P1_U3297) );
  INV_X1 U16790 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15113) );
  NOR2_X1 U16791 ( .A1(n15139), .A2(n15113), .ZN(P1_U3298) );
  INV_X1 U16792 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15114) );
  NOR2_X1 U16793 ( .A1(n15139), .A2(n15114), .ZN(P1_U3299) );
  INV_X1 U16794 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15115) );
  NOR2_X1 U16795 ( .A1(n15139), .A2(n15115), .ZN(P1_U3300) );
  INV_X1 U16796 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15116) );
  NOR2_X1 U16797 ( .A1(n15139), .A2(n15116), .ZN(P1_U3301) );
  INV_X1 U16798 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15117) );
  NOR2_X1 U16799 ( .A1(n15139), .A2(n15117), .ZN(P1_U3302) );
  INV_X1 U16800 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15118) );
  NOR2_X1 U16801 ( .A1(n15139), .A2(n15118), .ZN(P1_U3303) );
  INV_X1 U16802 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15119) );
  NOR2_X1 U16803 ( .A1(n15139), .A2(n15119), .ZN(P1_U3304) );
  INV_X1 U16804 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15120) );
  NOR2_X1 U16805 ( .A1(n15139), .A2(n15120), .ZN(P1_U3305) );
  INV_X1 U16806 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15121) );
  NOR2_X1 U16807 ( .A1(n15139), .A2(n15121), .ZN(P1_U3306) );
  INV_X1 U16808 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15122) );
  NOR2_X1 U16809 ( .A1(n15139), .A2(n15122), .ZN(P1_U3307) );
  INV_X1 U16810 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15123) );
  NOR2_X1 U16811 ( .A1(n15139), .A2(n15123), .ZN(P1_U3308) );
  INV_X1 U16812 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15124) );
  NOR2_X1 U16813 ( .A1(n15139), .A2(n15124), .ZN(P1_U3309) );
  INV_X1 U16814 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15125) );
  NOR2_X1 U16815 ( .A1(n15139), .A2(n15125), .ZN(P1_U3310) );
  INV_X1 U16816 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15126) );
  NOR2_X1 U16817 ( .A1(n15139), .A2(n15126), .ZN(P1_U3311) );
  INV_X1 U16818 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U16819 ( .A1(n15139), .A2(n15127), .ZN(P1_U3312) );
  INV_X1 U16820 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15128) );
  NOR2_X1 U16821 ( .A1(n15139), .A2(n15128), .ZN(P1_U3313) );
  INV_X1 U16822 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15129) );
  NOR2_X1 U16823 ( .A1(n15139), .A2(n15129), .ZN(P1_U3314) );
  INV_X1 U16824 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15130) );
  NOR2_X1 U16825 ( .A1(n15139), .A2(n15130), .ZN(P1_U3315) );
  INV_X1 U16826 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15131) );
  NOR2_X1 U16827 ( .A1(n15139), .A2(n15131), .ZN(P1_U3316) );
  INV_X1 U16828 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15132) );
  NOR2_X1 U16829 ( .A1(n15139), .A2(n15132), .ZN(P1_U3317) );
  INV_X1 U16830 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15133) );
  NOR2_X1 U16831 ( .A1(n15139), .A2(n15133), .ZN(P1_U3318) );
  INV_X1 U16832 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15134) );
  NOR2_X1 U16833 ( .A1(n15139), .A2(n15134), .ZN(P1_U3319) );
  NOR2_X1 U16834 ( .A1(n15139), .A2(n15135), .ZN(P1_U3320) );
  NOR2_X1 U16835 ( .A1(n15139), .A2(n15136), .ZN(P1_U3321) );
  NOR2_X1 U16836 ( .A1(n15139), .A2(n15137), .ZN(P1_U3322) );
  NOR2_X1 U16837 ( .A1(n15139), .A2(n15138), .ZN(P1_U3323) );
  INV_X1 U16838 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15140) );
  AOI22_X1 U16839 ( .A1(n15221), .A2(n15141), .B1(n15140), .B2(n15219), .ZN(
        P1_U3459) );
  AOI22_X1 U16840 ( .A1(n15144), .A2(n15143), .B1(n15142), .B2(n15192), .ZN(
        n15145) );
  OAI211_X1 U16841 ( .C1(n15197), .C2(n15147), .A(n15146), .B(n15145), .ZN(
        n15148) );
  INV_X1 U16842 ( .A(n15148), .ZN(n15222) );
  INV_X1 U16843 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15149) );
  AOI22_X1 U16844 ( .A1(n15221), .A2(n15222), .B1(n15149), .B2(n15219), .ZN(
        P1_U3462) );
  NOR2_X1 U16845 ( .A1(n15153), .A2(n15187), .ZN(n15155) );
  AOI21_X1 U16846 ( .B1(n7010), .B2(n15192), .A(n15150), .ZN(n15152) );
  OAI211_X1 U16847 ( .C1(n15153), .C2(n15197), .A(n15152), .B(n15151), .ZN(
        n15154) );
  AOI211_X1 U16848 ( .C1(n15156), .C2(n15189), .A(n15155), .B(n15154), .ZN(
        n15223) );
  INV_X1 U16849 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15157) );
  AOI22_X1 U16850 ( .A1(n15221), .A2(n15223), .B1(n15157), .B2(n15219), .ZN(
        P1_U3465) );
  INV_X1 U16851 ( .A(n15197), .ZN(n15210) );
  OAI21_X1 U16852 ( .B1(n15159), .B2(n15213), .A(n15158), .ZN(n15162) );
  INV_X1 U16853 ( .A(n15160), .ZN(n15161) );
  AOI211_X1 U16854 ( .C1(n15210), .C2(n15163), .A(n15162), .B(n15161), .ZN(
        n15224) );
  INV_X1 U16855 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U16856 ( .A1(n15221), .A2(n15224), .B1(n15164), .B2(n15219), .ZN(
        P1_U3468) );
  OAI211_X1 U16857 ( .C1(n15167), .C2(n15213), .A(n15166), .B(n15165), .ZN(
        n15170) );
  NOR2_X1 U16858 ( .A1(n15168), .A2(n15176), .ZN(n15169) );
  AOI211_X1 U16859 ( .C1(n15189), .C2(n15171), .A(n15170), .B(n15169), .ZN(
        n15225) );
  AOI22_X1 U16860 ( .A1(n15221), .A2(n15225), .B1(n9620), .B2(n15219), .ZN(
        P1_U3471) );
  NOR2_X1 U16861 ( .A1(n15173), .A2(n15172), .ZN(n15175) );
  OAI211_X1 U16862 ( .C1(n15177), .C2(n15176), .A(n15175), .B(n15174), .ZN(
        n15179) );
  NOR2_X1 U16863 ( .A1(n15179), .A2(n15178), .ZN(n15226) );
  INV_X1 U16864 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15180) );
  AOI22_X1 U16865 ( .A1(n15221), .A2(n15226), .B1(n15180), .B2(n15219), .ZN(
        P1_U3474) );
  OAI211_X1 U16866 ( .C1(n7284), .C2(n15213), .A(n15182), .B(n15181), .ZN(
        n15183) );
  AOI21_X1 U16867 ( .B1(n15184), .B2(n15210), .A(n15183), .ZN(n15185) );
  OAI21_X1 U16868 ( .B1(n15187), .B2(n15186), .A(n15185), .ZN(n15188) );
  AOI21_X1 U16869 ( .B1(n15190), .B2(n15189), .A(n15188), .ZN(n15227) );
  AOI22_X1 U16870 ( .A1(n15221), .A2(n15227), .B1(n9646), .B2(n15219), .ZN(
        P1_U3477) );
  AOI21_X1 U16871 ( .B1(n15193), .B2(n15192), .A(n15191), .ZN(n15194) );
  OAI211_X1 U16872 ( .C1(n15197), .C2(n15196), .A(n15195), .B(n15194), .ZN(
        n15198) );
  INV_X1 U16873 ( .A(n15198), .ZN(n15228) );
  INV_X1 U16874 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15199) );
  AOI22_X1 U16875 ( .A1(n15221), .A2(n15228), .B1(n15199), .B2(n15219), .ZN(
        P1_U3480) );
  OAI21_X1 U16876 ( .B1(n15201), .B2(n15213), .A(n15200), .ZN(n15203) );
  AOI211_X1 U16877 ( .C1(n15204), .C2(n15218), .A(n15203), .B(n15202), .ZN(
        n15229) );
  AOI22_X1 U16878 ( .A1(n15221), .A2(n15229), .B1(n9681), .B2(n15219), .ZN(
        P1_U3483) );
  OAI22_X1 U16879 ( .A1(n15206), .A2(n15205), .B1(n7087), .B2(n15213), .ZN(
        n15208) );
  AOI211_X1 U16880 ( .C1(n15210), .C2(n15209), .A(n15208), .B(n15207), .ZN(
        n15230) );
  INV_X1 U16881 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15211) );
  AOI22_X1 U16882 ( .A1(n15221), .A2(n15230), .B1(n15211), .B2(n15219), .ZN(
        P1_U3486) );
  OAI21_X1 U16883 ( .B1(n15214), .B2(n15213), .A(n15212), .ZN(n15216) );
  AOI211_X1 U16884 ( .C1(n15218), .C2(n15217), .A(n15216), .B(n15215), .ZN(
        n15232) );
  INV_X1 U16885 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15220) );
  AOI22_X1 U16886 ( .A1(n15221), .A2(n15232), .B1(n15220), .B2(n15219), .ZN(
        P1_U3489) );
  AOI22_X1 U16887 ( .A1(n15233), .A2(n15222), .B1(n9572), .B2(n15231), .ZN(
        P1_U3529) );
  AOI22_X1 U16888 ( .A1(n15233), .A2(n15223), .B1(n10280), .B2(n15231), .ZN(
        P1_U3530) );
  AOI22_X1 U16889 ( .A1(n15233), .A2(n15224), .B1(n9597), .B2(n15231), .ZN(
        P1_U3531) );
  AOI22_X1 U16890 ( .A1(n15233), .A2(n15225), .B1(n10281), .B2(n15231), .ZN(
        P1_U3532) );
  AOI22_X1 U16891 ( .A1(n15233), .A2(n15226), .B1(n10282), .B2(n15231), .ZN(
        P1_U3533) );
  AOI22_X1 U16892 ( .A1(n15233), .A2(n15227), .B1(n10278), .B2(n15231), .ZN(
        P1_U3534) );
  AOI22_X1 U16893 ( .A1(n15233), .A2(n15228), .B1(n10359), .B2(n15231), .ZN(
        P1_U3535) );
  AOI22_X1 U16894 ( .A1(n15233), .A2(n15229), .B1(n10415), .B2(n15231), .ZN(
        P1_U3536) );
  AOI22_X1 U16895 ( .A1(n15233), .A2(n15230), .B1(n10435), .B2(n15231), .ZN(
        P1_U3537) );
  AOI22_X1 U16896 ( .A1(n15233), .A2(n15232), .B1(n10480), .B2(n15231), .ZN(
        P1_U3538) );
  OAI211_X1 U16897 ( .C1(n15236), .C2(n15235), .A(n15299), .B(n15234), .ZN(
        n15237) );
  INV_X1 U16898 ( .A(n15237), .ZN(n15238) );
  AOI21_X1 U16899 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .A(n15238), 
        .ZN(n15245) );
  AOI22_X1 U16900 ( .A1(n15310), .A2(n15239), .B1(n15328), .B2(
        P2_ADDR_REG_2__SCAN_IN), .ZN(n15244) );
  OAI211_X1 U16901 ( .C1(n15242), .C2(n15241), .A(n15306), .B(n15240), .ZN(
        n15243) );
  NAND3_X1 U16902 ( .A1(n15245), .A2(n15244), .A3(n15243), .ZN(P2_U3216) );
  OAI211_X1 U16903 ( .C1(n15248), .C2(n15247), .A(n15299), .B(n15246), .ZN(
        n15252) );
  INV_X1 U16904 ( .A(n15249), .ZN(n15250) );
  AOI22_X1 U16905 ( .A1(n15310), .A2(n15250), .B1(n15328), .B2(
        P2_ADDR_REG_4__SCAN_IN), .ZN(n15251) );
  AND2_X1 U16906 ( .A1(n15252), .A2(n15251), .ZN(n15258) );
  NAND2_X1 U16907 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n15257) );
  OAI211_X1 U16908 ( .C1(n15255), .C2(n15254), .A(n15306), .B(n15253), .ZN(
        n15256) );
  NAND3_X1 U16909 ( .A1(n15258), .A2(n15257), .A3(n15256), .ZN(P2_U3218) );
  AOI22_X1 U16910 ( .A1(n15310), .A2(n15259), .B1(n15328), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n15273) );
  INV_X1 U16911 ( .A(n15260), .ZN(n15261) );
  AOI21_X1 U16912 ( .B1(n15263), .B2(n15262), .A(n15261), .ZN(n15264) );
  OR2_X1 U16913 ( .A1(n15264), .A2(n15330), .ZN(n15271) );
  INV_X1 U16914 ( .A(n15265), .ZN(n15266) );
  AOI21_X1 U16915 ( .B1(n15268), .B2(n15267), .A(n15266), .ZN(n15269) );
  OR2_X1 U16916 ( .A1(n15269), .A2(n15319), .ZN(n15270) );
  NAND4_X1 U16917 ( .A1(n15273), .A2(n15272), .A3(n15271), .A4(n15270), .ZN(
        P2_U3223) );
  INV_X1 U16918 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15287) );
  INV_X1 U16919 ( .A(n15274), .ZN(n15277) );
  AOI21_X1 U16920 ( .B1(n15278), .B2(n15275), .A(P2_REG2_REG_14__SCAN_IN), 
        .ZN(n15276) );
  AOI211_X1 U16921 ( .C1(n15278), .C2(n15277), .A(n15276), .B(n15330), .ZN(
        n15283) );
  AOI211_X1 U16922 ( .C1(n15281), .C2(n15280), .A(n15319), .B(n15279), .ZN(
        n15282) );
  AOI211_X1 U16923 ( .C1(n15310), .C2(n15284), .A(n15283), .B(n15282), .ZN(
        n15286) );
  NAND2_X1 U16924 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15285)
         );
  OAI211_X1 U16925 ( .C1(n15287), .C2(n15298), .A(n15286), .B(n15285), .ZN(
        P2_U3228) );
  NOR2_X1 U16926 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15288), .ZN(n15292) );
  AOI211_X1 U16927 ( .C1(n15290), .C2(n8225), .A(n15289), .B(n15319), .ZN(
        n15291) );
  AOI211_X1 U16928 ( .C1(n15310), .C2(n15293), .A(n15292), .B(n15291), .ZN(
        n15297) );
  OAI211_X1 U16929 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15295), .A(n15306), 
        .B(n15294), .ZN(n15296) );
  OAI211_X1 U16930 ( .C1(n15298), .C2(n7293), .A(n15297), .B(n15296), .ZN(
        P2_U3229) );
  OAI21_X1 U16931 ( .B1(n15301), .B2(n15300), .A(n15299), .ZN(n15303) );
  NOR2_X1 U16932 ( .A1(n15303), .A2(n15302), .ZN(n15304) );
  AOI21_X1 U16933 ( .B1(n15328), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n15304), 
        .ZN(n15314) );
  OAI211_X1 U16934 ( .C1(n15308), .C2(n15307), .A(n15306), .B(n15305), .ZN(
        n15312) );
  NAND2_X1 U16935 ( .A1(n15310), .A2(n15309), .ZN(n15311) );
  NAND4_X1 U16936 ( .A1(n15314), .A2(n15313), .A3(n15312), .A4(n15311), .ZN(
        P2_U3231) );
  AOI21_X1 U16937 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n15316), .A(n15315), 
        .ZN(n15331) );
  INV_X1 U16938 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15321) );
  INV_X1 U16939 ( .A(n15317), .ZN(n15320) );
  AOI211_X1 U16940 ( .C1(n15321), .C2(n15320), .A(n15319), .B(n15318), .ZN(
        n15327) );
  INV_X1 U16941 ( .A(n15322), .ZN(n15323) );
  OAI21_X1 U16942 ( .B1(n15325), .B2(n15324), .A(n15323), .ZN(n15326) );
  AOI211_X1 U16943 ( .C1(n15328), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n15327), 
        .B(n15326), .ZN(n15329) );
  OAI21_X1 U16944 ( .B1(n15331), .B2(n15330), .A(n15329), .ZN(P2_U3232) );
  NOR2_X1 U16945 ( .A1(n15332), .A2(n15365), .ZN(n15360) );
  INV_X1 U16946 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U16947 ( .A1(n15364), .A2(n15333), .ZN(P2_U3266) );
  INV_X1 U16948 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15334) );
  NOR2_X1 U16949 ( .A1(n15364), .A2(n15334), .ZN(P2_U3267) );
  INV_X1 U16950 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U16951 ( .A1(n15364), .A2(n15335), .ZN(P2_U3268) );
  INV_X1 U16952 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15336) );
  NOR2_X1 U16953 ( .A1(n15360), .A2(n15336), .ZN(P2_U3269) );
  INV_X1 U16954 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15337) );
  NOR2_X1 U16955 ( .A1(n15360), .A2(n15337), .ZN(P2_U3270) );
  INV_X1 U16956 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15338) );
  NOR2_X1 U16957 ( .A1(n15360), .A2(n15338), .ZN(P2_U3271) );
  INV_X1 U16958 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15339) );
  NOR2_X1 U16959 ( .A1(n15360), .A2(n15339), .ZN(P2_U3272) );
  INV_X1 U16960 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15340) );
  NOR2_X1 U16961 ( .A1(n15360), .A2(n15340), .ZN(P2_U3273) );
  INV_X1 U16962 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15341) );
  NOR2_X1 U16963 ( .A1(n15360), .A2(n15341), .ZN(P2_U3274) );
  INV_X1 U16964 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15342) );
  NOR2_X1 U16965 ( .A1(n15360), .A2(n15342), .ZN(P2_U3275) );
  INV_X1 U16966 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15343) );
  NOR2_X1 U16967 ( .A1(n15360), .A2(n15343), .ZN(P2_U3276) );
  INV_X1 U16968 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15344) );
  NOR2_X1 U16969 ( .A1(n15360), .A2(n15344), .ZN(P2_U3277) );
  INV_X1 U16970 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15345) );
  NOR2_X1 U16971 ( .A1(n15364), .A2(n15345), .ZN(P2_U3278) );
  INV_X1 U16972 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15346) );
  NOR2_X1 U16973 ( .A1(n15364), .A2(n15346), .ZN(P2_U3279) );
  INV_X1 U16974 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15347) );
  NOR2_X1 U16975 ( .A1(n15364), .A2(n15347), .ZN(P2_U3280) );
  INV_X1 U16976 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15348) );
  NOR2_X1 U16977 ( .A1(n15364), .A2(n15348), .ZN(P2_U3281) );
  INV_X1 U16978 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U16979 ( .A1(n15364), .A2(n15349), .ZN(P2_U3282) );
  INV_X1 U16980 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15350) );
  NOR2_X1 U16981 ( .A1(n15364), .A2(n15350), .ZN(P2_U3283) );
  INV_X1 U16982 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15351) );
  NOR2_X1 U16983 ( .A1(n15364), .A2(n15351), .ZN(P2_U3284) );
  INV_X1 U16984 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15352) );
  NOR2_X1 U16985 ( .A1(n15364), .A2(n15352), .ZN(P2_U3285) );
  INV_X1 U16986 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15353) );
  NOR2_X1 U16987 ( .A1(n15364), .A2(n15353), .ZN(P2_U3286) );
  INV_X1 U16988 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15354) );
  NOR2_X1 U16989 ( .A1(n15364), .A2(n15354), .ZN(P2_U3287) );
  INV_X1 U16990 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15355) );
  NOR2_X1 U16991 ( .A1(n15364), .A2(n15355), .ZN(P2_U3288) );
  INV_X1 U16992 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15356) );
  NOR2_X1 U16993 ( .A1(n15364), .A2(n15356), .ZN(P2_U3289) );
  INV_X1 U16994 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15357) );
  NOR2_X1 U16995 ( .A1(n15360), .A2(n15357), .ZN(P2_U3290) );
  INV_X1 U16996 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15358) );
  NOR2_X1 U16997 ( .A1(n15364), .A2(n15358), .ZN(P2_U3291) );
  INV_X1 U16998 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15359) );
  NOR2_X1 U16999 ( .A1(n15360), .A2(n15359), .ZN(P2_U3292) );
  INV_X1 U17000 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15361) );
  NOR2_X1 U17001 ( .A1(n15364), .A2(n15361), .ZN(P2_U3293) );
  INV_X1 U17002 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15362) );
  NOR2_X1 U17003 ( .A1(n15364), .A2(n15362), .ZN(P2_U3294) );
  INV_X1 U17004 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15363) );
  NOR2_X1 U17005 ( .A1(n15364), .A2(n15363), .ZN(P2_U3295) );
  INV_X1 U17006 ( .A(n15365), .ZN(n15370) );
  AOI22_X1 U17007 ( .A1(n15370), .A2(n15367), .B1(n15366), .B2(n15365), .ZN(
        P2_U3416) );
  OAI21_X1 U17008 ( .B1(n15370), .B2(n15369), .A(n15368), .ZN(P2_U3417) );
  AOI21_X1 U17009 ( .B1(n15373), .B2(n15372), .A(n15371), .ZN(n15374) );
  OAI211_X1 U17010 ( .C1(n15377), .C2(n15376), .A(n15375), .B(n15374), .ZN(
        n15378) );
  INV_X1 U17011 ( .A(n15378), .ZN(n15388) );
  AOI22_X1 U17012 ( .A1(n15387), .A2(n15388), .B1(n8081), .B2(n15386), .ZN(
        P2_U3454) );
  INV_X1 U17013 ( .A(n15379), .ZN(n15385) );
  OAI21_X1 U17014 ( .B1(n15382), .B2(n15381), .A(n15380), .ZN(n15384) );
  AOI22_X1 U17015 ( .A1(n15387), .A2(n15390), .B1(n7887), .B2(n15386), .ZN(
        P2_U3460) );
  AOI22_X1 U17016 ( .A1(n15391), .A2(n15388), .B1(n10314), .B2(n15389), .ZN(
        P2_U3507) );
  AOI22_X1 U17017 ( .A1(n15391), .A2(n15390), .B1(n10303), .B2(n15389), .ZN(
        P2_U3509) );
  NOR2_X1 U17018 ( .A1(P3_U3897), .A2(n15392), .ZN(P3_U3150) );
  XNOR2_X1 U17019 ( .A(n15393), .B(n15396), .ZN(n15503) );
  AOI21_X1 U17020 ( .B1(n15396), .B2(n15395), .A(n15394), .ZN(n15402) );
  AOI22_X1 U17021 ( .A1(n15399), .A2(n15447), .B1(n15398), .B2(n15397), .ZN(
        n15401) );
  NAND2_X1 U17022 ( .A1(n15503), .A2(n15435), .ZN(n15400) );
  OAI211_X1 U17023 ( .C1(n15402), .C2(n15430), .A(n15401), .B(n15400), .ZN(
        n15501) );
  AOI21_X1 U17024 ( .B1(n15439), .B2(n15503), .A(n15501), .ZN(n15406) );
  NOR2_X1 U17025 ( .A1(n15403), .A2(n15512), .ZN(n15502) );
  AOI22_X1 U17026 ( .A1(n15419), .A2(n15502), .B1(n15442), .B2(n15404), .ZN(
        n15405) );
  OAI221_X1 U17027 ( .B1(n15465), .B2(n15406), .C1(n15463), .C2(n11009), .A(
        n15405), .ZN(P3_U3225) );
  XNOR2_X1 U17028 ( .A(n15407), .B(n15412), .ZN(n15417) );
  INV_X1 U17029 ( .A(n15417), .ZN(n15477) );
  OAI22_X1 U17030 ( .A1(n15408), .A2(n15450), .B1(n15451), .B2(n15425), .ZN(
        n15409) );
  INV_X1 U17031 ( .A(n15409), .ZN(n15415) );
  AND2_X1 U17032 ( .A1(n15432), .A2(n15410), .ZN(n15413) );
  OAI211_X1 U17033 ( .C1(n15413), .C2(n15412), .A(n15411), .B(n15453), .ZN(
        n15414) );
  OAI211_X1 U17034 ( .C1(n15417), .C2(n15416), .A(n15415), .B(n15414), .ZN(
        n15475) );
  AOI21_X1 U17035 ( .B1(n15439), .B2(n15477), .A(n15475), .ZN(n15421) );
  NOR2_X1 U17036 ( .A1(n15418), .A2(n15512), .ZN(n15476) );
  AOI22_X1 U17037 ( .A1(n15476), .A2(n15419), .B1(n15442), .B2(n15581), .ZN(
        n15420) );
  OAI221_X1 U17038 ( .B1(n15465), .B2(n15421), .C1(n15463), .C2(n10760), .A(
        n15420), .ZN(P3_U3230) );
  OAI21_X1 U17039 ( .B1(n15423), .B2(n15429), .A(n15422), .ZN(n15473) );
  OAI22_X1 U17040 ( .A1(n15426), .A2(n15425), .B1(n15424), .B2(n15450), .ZN(
        n15434) );
  NAND3_X1 U17041 ( .A1(n15427), .A2(n15429), .A3(n15428), .ZN(n15431) );
  AOI21_X1 U17042 ( .B1(n15432), .B2(n15431), .A(n15430), .ZN(n15433) );
  AOI211_X1 U17043 ( .C1(n15435), .C2(n15473), .A(n15434), .B(n15433), .ZN(
        n15436) );
  INV_X1 U17044 ( .A(n15436), .ZN(n15471) );
  NOR2_X1 U17045 ( .A1(n15437), .A2(n15512), .ZN(n15472) );
  AOI22_X1 U17046 ( .A1(n15473), .A2(n15439), .B1(n15472), .B2(n15438), .ZN(
        n15440) );
  INV_X1 U17047 ( .A(n15440), .ZN(n15441) );
  AOI211_X1 U17048 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15442), .A(n15471), .B(
        n15441), .ZN(n15443) );
  AOI22_X1 U17049 ( .A1(n15465), .A2(n10667), .B1(n15443), .B2(n15463), .ZN(
        P3_U3231) );
  NAND2_X1 U17050 ( .A1(n15444), .A2(n15495), .ZN(n15468) );
  OR2_X1 U17051 ( .A1(n11570), .A2(n15445), .ZN(n15446) );
  NAND2_X1 U17052 ( .A1(n15427), .A2(n15446), .ZN(n15454) );
  NAND2_X1 U17053 ( .A1(n15448), .A2(n15447), .ZN(n15449) );
  OAI21_X1 U17054 ( .B1(n15451), .B2(n15450), .A(n15449), .ZN(n15452) );
  AOI21_X1 U17055 ( .B1(n15454), .B2(n15453), .A(n15452), .ZN(n15470) );
  OAI21_X1 U17056 ( .B1(n15455), .B2(n15468), .A(n15470), .ZN(n15456) );
  INV_X1 U17057 ( .A(n15456), .ZN(n15464) );
  XNOR2_X1 U17058 ( .A(n11570), .B(n15457), .ZN(n15467) );
  OAI22_X1 U17059 ( .A1(n15467), .A2(n15460), .B1(n15459), .B2(n15458), .ZN(
        n15461) );
  INV_X1 U17060 ( .A(n15461), .ZN(n15462) );
  OAI221_X1 U17061 ( .B1(n15465), .B2(n15464), .C1(n15463), .C2(n8662), .A(
        n15462), .ZN(P3_U3232) );
  OR2_X1 U17062 ( .A1(n15467), .A2(n15466), .ZN(n15469) );
  AND3_X1 U17063 ( .A1(n15470), .A2(n15469), .A3(n15468), .ZN(n15520) );
  AOI22_X1 U17064 ( .A1(n15519), .A2(n15520), .B1(n7000), .B2(n15517), .ZN(
        P3_U3393) );
  AOI211_X1 U17065 ( .C1(n15509), .C2(n15473), .A(n15472), .B(n15471), .ZN(
        n15521) );
  INV_X1 U17066 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15474) );
  AOI22_X1 U17067 ( .A1(n15519), .A2(n15521), .B1(n15474), .B2(n15517), .ZN(
        P3_U3396) );
  AOI211_X1 U17068 ( .C1(n15477), .C2(n15509), .A(n15476), .B(n15475), .ZN(
        n15522) );
  INV_X1 U17069 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U17070 ( .A1(n15519), .A2(n15522), .B1(n15478), .B2(n15517), .ZN(
        P3_U3399) );
  INV_X1 U17071 ( .A(n15479), .ZN(n15481) );
  AOI211_X1 U17072 ( .C1(n15509), .C2(n15482), .A(n15481), .B(n15480), .ZN(
        n15523) );
  INV_X1 U17073 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U17074 ( .A1(n15519), .A2(n15523), .B1(n15483), .B2(n15517), .ZN(
        P3_U3402) );
  AOI21_X1 U17075 ( .B1(n15485), .B2(n15509), .A(n15484), .ZN(n15486) );
  AND2_X1 U17076 ( .A1(n15487), .A2(n15486), .ZN(n15524) );
  INV_X1 U17077 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15488) );
  AOI22_X1 U17078 ( .A1(n15519), .A2(n15524), .B1(n15488), .B2(n15517), .ZN(
        P3_U3405) );
  INV_X1 U17079 ( .A(n15489), .ZN(n15492) );
  AND2_X1 U17080 ( .A1(n15490), .A2(n15509), .ZN(n15491) );
  NOR3_X1 U17081 ( .A1(n15493), .A2(n15492), .A3(n15491), .ZN(n15525) );
  INV_X1 U17082 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15494) );
  AOI22_X1 U17083 ( .A1(n15519), .A2(n15525), .B1(n15494), .B2(n15517), .ZN(
        P3_U3408) );
  AOI22_X1 U17084 ( .A1(n15497), .A2(n15509), .B1(n15496), .B2(n15495), .ZN(
        n15498) );
  AND2_X1 U17085 ( .A1(n15499), .A2(n15498), .ZN(n15527) );
  INV_X1 U17086 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U17087 ( .A1(n15519), .A2(n15527), .B1(n15500), .B2(n15517), .ZN(
        P3_U3411) );
  AOI211_X1 U17088 ( .C1(n15503), .C2(n15509), .A(n15502), .B(n15501), .ZN(
        n15528) );
  INV_X1 U17089 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U17090 ( .A1(n15519), .A2(n15528), .B1(n15504), .B2(n15517), .ZN(
        P3_U3414) );
  INV_X1 U17091 ( .A(n15505), .ZN(n15506) );
  AOI211_X1 U17092 ( .C1(n15509), .C2(n15508), .A(n15507), .B(n15506), .ZN(
        n15529) );
  INV_X1 U17093 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15510) );
  AOI22_X1 U17094 ( .A1(n15519), .A2(n15529), .B1(n15510), .B2(n15517), .ZN(
        P3_U3417) );
  OAI21_X1 U17095 ( .B1(n15513), .B2(n15512), .A(n15511), .ZN(n15514) );
  AOI21_X1 U17096 ( .B1(n15516), .B2(n15515), .A(n15514), .ZN(n15531) );
  INV_X1 U17097 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U17098 ( .A1(n15519), .A2(n15531), .B1(n15518), .B2(n15517), .ZN(
        P3_U3420) );
  AOI22_X1 U17099 ( .A1(n15532), .A2(n15520), .B1(n8663), .B2(n15530), .ZN(
        P3_U3460) );
  AOI22_X1 U17100 ( .A1(n15532), .A2(n15521), .B1(n10666), .B2(n15530), .ZN(
        P3_U3461) );
  AOI22_X1 U17101 ( .A1(n15532), .A2(n15522), .B1(n10759), .B2(n15530), .ZN(
        P3_U3462) );
  AOI22_X1 U17102 ( .A1(n15532), .A2(n15523), .B1(n10764), .B2(n15530), .ZN(
        P3_U3463) );
  AOI22_X1 U17103 ( .A1(n15532), .A2(n15524), .B1(n10770), .B2(n15530), .ZN(
        P3_U3464) );
  AOI22_X1 U17104 ( .A1(n15532), .A2(n15525), .B1(n10946), .B2(n15530), .ZN(
        P3_U3465) );
  AOI22_X1 U17105 ( .A1(n15532), .A2(n15527), .B1(n15526), .B2(n15530), .ZN(
        P3_U3466) );
  AOI22_X1 U17106 ( .A1(n15532), .A2(n15528), .B1(n11022), .B2(n15530), .ZN(
        P3_U3467) );
  AOI22_X1 U17107 ( .A1(n15532), .A2(n15529), .B1(n11155), .B2(n15530), .ZN(
        P3_U3468) );
  AOI22_X1 U17108 ( .A1(n15532), .A2(n15531), .B1(n11440), .B2(n15530), .ZN(
        P3_U3469) );
  NAND2_X1 U17109 ( .A1(n15534), .A2(n15533), .ZN(n15535) );
  OAI21_X1 U17110 ( .B1(n15536), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n15535), 
        .ZN(n15921) );
  OAI22_X1 U17111 ( .A1(P3_DATAO_REG_2__SCAN_IN), .A2(keyinput_g94), .B1(
        P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .ZN(n15537) );
  AOI221_X1 U17112 ( .B1(P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_g94), .C1(
        keyinput_g79), .C2(P3_DATAO_REG_17__SCAN_IN), .A(n15537), .ZN(n15544)
         );
  OAI22_X1 U17113 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_g124), .B1(
        P3_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .ZN(n15538) );
  AOI221_X1 U17114 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_g124), .C1(
        keyinput_g80), .C2(P3_DATAO_REG_16__SCAN_IN), .A(n15538), .ZN(n15543)
         );
  OAI22_X1 U17115 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        keyinput_g120), .B2(P1_IR_REG_13__SCAN_IN), .ZN(n15539) );
  AOI221_X1 U17116 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_g120), .A(n15539), .ZN(n15542) );
  OAI22_X1 U17117 ( .A1(SI_15_), .A2(keyinput_g17), .B1(keyinput_g25), .B2(
        SI_7_), .ZN(n15540) );
  AOI221_X1 U17118 ( .B1(SI_15_), .B2(keyinput_g17), .C1(SI_7_), .C2(
        keyinput_g25), .A(n15540), .ZN(n15541) );
  NAND4_X1 U17119 ( .A1(n15544), .A2(n15543), .A3(n15542), .A4(n15541), .ZN(
        n15677) );
  AOI22_X1 U17120 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        P3_WR_REG_SCAN_IN), .B2(keyinput_g0), .ZN(n15545) );
  OAI221_X1 U17121 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        P3_WR_REG_SCAN_IN), .C2(keyinput_g0), .A(n15545), .ZN(n15552) );
  AOI22_X1 U17122 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_g112), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n15546) );
  OAI221_X1 U17123 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_g112), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n15546), .ZN(n15551)
         );
  AOI22_X1 U17124 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n15547) );
  OAI221_X1 U17125 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n15547), .ZN(n15550)
         );
  AOI22_X1 U17126 ( .A1(SI_20_), .A2(keyinput_g12), .B1(P3_STATE_REG_SCAN_IN), 
        .B2(keyinput_g34), .ZN(n15548) );
  OAI221_X1 U17127 ( .B1(SI_20_), .B2(keyinput_g12), .C1(P3_STATE_REG_SCAN_IN), 
        .C2(keyinput_g34), .A(n15548), .ZN(n15549) );
  NOR4_X1 U17128 ( .A1(n15552), .A2(n15551), .A3(n15550), .A4(n15549), .ZN(
        n15570) );
  AOI22_X1 U17129 ( .A1(P3_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .ZN(n15553) );
  OAI221_X1 U17130 ( .B1(P3_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_g45), .A(n15553), .ZN(n15560)
         );
  AOI22_X1 U17131 ( .A1(P3_DATAO_REG_24__SCAN_IN), .A2(keyinput_g72), .B1(
        P3_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n15554) );
  OAI221_X1 U17132 ( .B1(P3_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n15554), .ZN(n15559) );
  AOI22_X1 U17133 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        P3_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .ZN(n15555) );
  OAI221_X1 U17134 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        P3_DATAO_REG_26__SCAN_IN), .C2(keyinput_g70), .A(n15555), .ZN(n15558)
         );
  AOI22_X1 U17135 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(keyinput_g100), .B1(
        P3_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .ZN(n15556) );
  OAI221_X1 U17136 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(keyinput_g100), .C1(
        P3_REG3_REG_5__SCAN_IN), .C2(keyinput_g49), .A(n15556), .ZN(n15557) );
  NOR4_X1 U17137 ( .A1(n15560), .A2(n15559), .A3(n15558), .A4(n15557), .ZN(
        n15569) );
  OAI22_X1 U17138 ( .A1(SI_5_), .A2(keyinput_g27), .B1(P3_ADDR_REG_7__SCAN_IN), 
        .B2(keyinput_g104), .ZN(n15561) );
  AOI221_X1 U17139 ( .B1(SI_5_), .B2(keyinput_g27), .C1(keyinput_g104), .C2(
        P3_ADDR_REG_7__SCAN_IN), .A(n15561), .ZN(n15567) );
  OAI22_X1 U17140 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        P3_DATAO_REG_22__SCAN_IN), .B2(keyinput_g74), .ZN(n15562) );
  AOI221_X1 U17141 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        keyinput_g74), .C2(P3_DATAO_REG_22__SCAN_IN), .A(n15562), .ZN(n15566)
         );
  OAI22_X1 U17142 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_g127), .B1(
        P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_g99), .ZN(n15563) );
  AOI221_X1 U17143 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_g127), .C1(
        keyinput_g99), .C2(P3_ADDR_REG_2__SCAN_IN), .A(n15563), .ZN(n15565) );
  XNOR2_X1 U17144 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g113), .ZN(n15564)
         );
  AND4_X1 U17145 ( .A1(n15567), .A2(n15566), .A3(n15565), .A4(n15564), .ZN(
        n15568) );
  NAND3_X1 U17146 ( .A1(n15570), .A2(n15569), .A3(n15568), .ZN(n15676) );
  AOI22_X1 U17147 ( .A1(P3_DATAO_REG_31__SCAN_IN), .A2(keyinput_g65), .B1(
        P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n15571) );
  OAI221_X1 U17148 ( .B1(P3_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n15571), .ZN(n15579)
         );
  AOI22_X1 U17149 ( .A1(n15880), .A2(keyinput_g96), .B1(n15895), .B2(
        keyinput_g13), .ZN(n15572) );
  OAI221_X1 U17150 ( .B1(n15880), .B2(keyinput_g96), .C1(n15895), .C2(
        keyinput_g13), .A(n15572), .ZN(n15578) );
  AOI22_X1 U17151 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g110), .B1(SI_21_), 
        .B2(keyinput_g11), .ZN(n15573) );
  OAI221_X1 U17152 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g110), .C1(SI_21_), .C2(keyinput_g11), .A(n15573), .ZN(n15577) );
  XNOR2_X1 U17153 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g119), .ZN(n15575)
         );
  XNOR2_X1 U17154 ( .A(SI_18_), .B(keyinput_g14), .ZN(n15574) );
  NAND2_X1 U17155 ( .A1(n15575), .A2(n15574), .ZN(n15576) );
  NOR4_X1 U17156 ( .A1(n15579), .A2(n15578), .A3(n15577), .A4(n15576), .ZN(
        n15623) );
  AOI22_X1 U17157 ( .A1(n15581), .A2(keyinput_g40), .B1(keyinput_g101), .B2(
        n15887), .ZN(n15580) );
  OAI221_X1 U17158 ( .B1(n15581), .B2(keyinput_g40), .C1(n15887), .C2(
        keyinput_g101), .A(n15580), .ZN(n15593) );
  AOI22_X1 U17159 ( .A1(n15584), .A2(keyinput_g77), .B1(n15583), .B2(
        keyinput_g83), .ZN(n15582) );
  OAI221_X1 U17160 ( .B1(n15584), .B2(keyinput_g77), .C1(n15583), .C2(
        keyinput_g83), .A(n15582), .ZN(n15592) );
  AOI22_X1 U17161 ( .A1(n15587), .A2(keyinput_g35), .B1(keyinput_g28), .B2(
        n15586), .ZN(n15585) );
  OAI221_X1 U17162 ( .B1(n15587), .B2(keyinput_g35), .C1(n15586), .C2(
        keyinput_g28), .A(n15585), .ZN(n15591) );
  XNOR2_X1 U17163 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g111), .ZN(n15589)
         );
  XNOR2_X1 U17164 ( .A(SI_17_), .B(keyinput_g15), .ZN(n15588) );
  NAND2_X1 U17165 ( .A1(n15589), .A2(n15588), .ZN(n15590) );
  NOR4_X1 U17166 ( .A1(n15593), .A2(n15592), .A3(n15591), .A4(n15590), .ZN(
        n15622) );
  AOI22_X1 U17167 ( .A1(n15812), .A2(keyinput_g62), .B1(keyinput_g16), .B2(
        n15595), .ZN(n15594) );
  OAI221_X1 U17168 ( .B1(n15812), .B2(keyinput_g62), .C1(n15595), .C2(
        keyinput_g16), .A(n15594), .ZN(n15606) );
  AOI22_X1 U17169 ( .A1(n15598), .A2(keyinput_g52), .B1(keyinput_g3), .B2(
        n15597), .ZN(n15596) );
  OAI221_X1 U17170 ( .B1(n15598), .B2(keyinput_g52), .C1(n15597), .C2(
        keyinput_g3), .A(n15596), .ZN(n15605) );
  INV_X1 U17171 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15853) );
  AOI22_X1 U17172 ( .A1(n15600), .A2(keyinput_g37), .B1(n15853), .B2(
        keyinput_g47), .ZN(n15599) );
  OAI221_X1 U17173 ( .B1(n15600), .B2(keyinput_g37), .C1(n15853), .C2(
        keyinput_g47), .A(n15599), .ZN(n15604) );
  XOR2_X1 U17174 ( .A(n8790), .B(keyinput_g53), .Z(n15602) );
  XNOR2_X1 U17175 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_g121), .ZN(n15601)
         );
  NAND2_X1 U17176 ( .A1(n15602), .A2(n15601), .ZN(n15603) );
  NOR4_X1 U17177 ( .A1(n15606), .A2(n15605), .A3(n15604), .A4(n15603), .ZN(
        n15621) );
  AOI22_X1 U17178 ( .A1(n15809), .A2(keyinput_g73), .B1(n15608), .B2(
        keyinput_g66), .ZN(n15607) );
  OAI221_X1 U17179 ( .B1(n15809), .B2(keyinput_g73), .C1(n15608), .C2(
        keyinput_g66), .A(n15607), .ZN(n15619) );
  AOI22_X1 U17180 ( .A1(n15832), .A2(keyinput_g92), .B1(n15610), .B2(
        keyinput_g89), .ZN(n15609) );
  OAI221_X1 U17181 ( .B1(n15832), .B2(keyinput_g92), .C1(n15610), .C2(
        keyinput_g89), .A(n15609), .ZN(n15618) );
  AOI22_X1 U17182 ( .A1(n15613), .A2(keyinput_g8), .B1(keyinput_g31), .B2(
        n15612), .ZN(n15611) );
  OAI221_X1 U17183 ( .B1(n15613), .B2(keyinput_g8), .C1(n15612), .C2(
        keyinput_g31), .A(n15611), .ZN(n15617) );
  XNOR2_X1 U17184 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g107), .ZN(n15615)
         );
  XNOR2_X1 U17185 ( .A(SI_13_), .B(keyinput_g19), .ZN(n15614) );
  NAND2_X1 U17186 ( .A1(n15615), .A2(n15614), .ZN(n15616) );
  NOR4_X1 U17187 ( .A1(n15619), .A2(n15618), .A3(n15617), .A4(n15616), .ZN(
        n15620) );
  NAND4_X1 U17188 ( .A1(n15623), .A2(n15622), .A3(n15621), .A4(n15620), .ZN(
        n15675) );
  AOI22_X1 U17189 ( .A1(n15625), .A2(keyinput_g50), .B1(keyinput_g105), .B2(
        n15822), .ZN(n15624) );
  OAI221_X1 U17190 ( .B1(n15625), .B2(keyinput_g50), .C1(n15822), .C2(
        keyinput_g105), .A(n15624), .ZN(n15634) );
  INV_X1 U17191 ( .A(SI_31_), .ZN(n15627) );
  AOI22_X1 U17192 ( .A1(n15814), .A2(keyinput_g20), .B1(keyinput_g1), .B2(
        n15627), .ZN(n15626) );
  OAI221_X1 U17193 ( .B1(n15814), .B2(keyinput_g20), .C1(n15627), .C2(
        keyinput_g1), .A(n15626), .ZN(n15633) );
  INV_X1 U17194 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15790) );
  AOI22_X1 U17195 ( .A1(n15864), .A2(keyinput_g98), .B1(n15790), .B2(
        keyinput_g55), .ZN(n15628) );
  OAI221_X1 U17196 ( .B1(n15864), .B2(keyinput_g98), .C1(n15790), .C2(
        keyinput_g55), .A(n15628), .ZN(n15632) );
  XNOR2_X1 U17197 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g118), .ZN(n15630)
         );
  XNOR2_X1 U17198 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_g116), .ZN(n15629)
         );
  NAND2_X1 U17199 ( .A1(n15630), .A2(n15629), .ZN(n15631) );
  NOR4_X1 U17200 ( .A1(n15634), .A2(n15633), .A3(n15632), .A4(n15631), .ZN(
        n15673) );
  INV_X1 U17201 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15637) );
  AOI22_X1 U17202 ( .A1(n15637), .A2(keyinput_g57), .B1(keyinput_g84), .B2(
        n15636), .ZN(n15635) );
  OAI221_X1 U17203 ( .B1(n15637), .B2(keyinput_g57), .C1(n15636), .C2(
        keyinput_g84), .A(n15635), .ZN(n15645) );
  INV_X1 U17204 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n15826) );
  AOI22_X1 U17205 ( .A1(n9689), .A2(keyinput_g114), .B1(n15826), .B2(
        keyinput_g122), .ZN(n15638) );
  OAI221_X1 U17206 ( .B1(n9689), .B2(keyinput_g114), .C1(n15826), .C2(
        keyinput_g122), .A(n15638), .ZN(n15644) );
  AOI22_X1 U17207 ( .A1(n15866), .A2(keyinput_g95), .B1(n15861), .B2(
        keyinput_g97), .ZN(n15639) );
  OAI221_X1 U17208 ( .B1(n15866), .B2(keyinput_g95), .C1(n15861), .C2(
        keyinput_g97), .A(n15639), .ZN(n15643) );
  AOI22_X1 U17209 ( .A1(n15641), .A2(keyinput_g71), .B1(n15823), .B2(
        keyinput_g22), .ZN(n15640) );
  OAI221_X1 U17210 ( .B1(n15641), .B2(keyinput_g71), .C1(n15823), .C2(
        keyinput_g22), .A(n15640), .ZN(n15642) );
  NOR4_X1 U17211 ( .A1(n15645), .A2(n15644), .A3(n15643), .A4(n15642), .ZN(
        n15672) );
  INV_X1 U17212 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n15859) );
  AOI22_X1 U17213 ( .A1(n15850), .A2(keyinput_g93), .B1(keyinput_g67), .B2(
        n15859), .ZN(n15646) );
  OAI221_X1 U17214 ( .B1(n15850), .B2(keyinput_g93), .C1(n15859), .C2(
        keyinput_g67), .A(n15646), .ZN(n15649) );
  XNOR2_X1 U17215 ( .A(n15647), .B(keyinput_g90), .ZN(n15648) );
  NOR2_X1 U17216 ( .A1(n15649), .A2(n15648), .ZN(n15658) );
  AOI22_X1 U17217 ( .A1(n15459), .A2(keyinput_g44), .B1(n15789), .B2(
        keyinput_g23), .ZN(n15650) );
  OAI221_X1 U17218 ( .B1(n15459), .B2(keyinput_g44), .C1(n15789), .C2(
        keyinput_g23), .A(n15650), .ZN(n15651) );
  INV_X1 U17219 ( .A(n15651), .ZN(n15657) );
  AOI22_X1 U17220 ( .A1(n15653), .A2(keyinput_g36), .B1(keyinput_g106), .B2(
        n15852), .ZN(n15652) );
  OAI221_X1 U17221 ( .B1(n15653), .B2(keyinput_g36), .C1(n15852), .C2(
        keyinput_g106), .A(n15652), .ZN(n15654) );
  INV_X1 U17222 ( .A(n15654), .ZN(n15656) );
  XNOR2_X1 U17223 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_g126), .ZN(n15655)
         );
  AND4_X1 U17224 ( .A1(n15658), .A2(n15657), .A3(n15656), .A4(n15655), .ZN(
        n15671) );
  INV_X1 U17225 ( .A(SI_22_), .ZN(n15660) );
  AOI22_X1 U17226 ( .A1(n15660), .A2(keyinput_g10), .B1(n15849), .B2(
        keyinput_g39), .ZN(n15659) );
  OAI221_X1 U17227 ( .B1(n15660), .B2(keyinput_g10), .C1(n15849), .C2(
        keyinput_g39), .A(n15659), .ZN(n15669) );
  AOI22_X1 U17228 ( .A1(n10135), .A2(keyinput_g32), .B1(n15662), .B2(
        keyinput_g9), .ZN(n15661) );
  OAI221_X1 U17229 ( .B1(n10135), .B2(keyinput_g32), .C1(n15662), .C2(
        keyinput_g9), .A(n15661), .ZN(n15668) );
  AOI22_X1 U17230 ( .A1(n15810), .A2(keyinput_g87), .B1(n15664), .B2(
        keyinput_g76), .ZN(n15663) );
  OAI221_X1 U17231 ( .B1(n15810), .B2(keyinput_g87), .C1(n15664), .C2(
        keyinput_g76), .A(n15663), .ZN(n15667) );
  AOI22_X1 U17232 ( .A1(n7067), .A2(keyinput_g29), .B1(keyinput_g6), .B2(
        n15877), .ZN(n15665) );
  OAI221_X1 U17233 ( .B1(n7067), .B2(keyinput_g29), .C1(n15877), .C2(
        keyinput_g6), .A(n15665), .ZN(n15666) );
  NOR4_X1 U17234 ( .A1(n15669), .A2(n15668), .A3(n15667), .A4(n15666), .ZN(
        n15670) );
  NAND4_X1 U17235 ( .A1(n15673), .A2(n15672), .A3(n15671), .A4(n15670), .ZN(
        n15674) );
  NOR4_X1 U17236 ( .A1(n15677), .A2(n15676), .A3(n15675), .A4(n15674), .ZN(
        n15914) );
  OAI22_X1 U17237 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_g123), .ZN(n15678) );
  AOI221_X1 U17238 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        keyinput_g123), .C2(P1_IR_REG_16__SCAN_IN), .A(n15678), .ZN(n15685) );
  OAI22_X1 U17239 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g109), .B1(
        P3_DATAO_REG_5__SCAN_IN), .B2(keyinput_g91), .ZN(n15679) );
  AOI221_X1 U17240 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g109), .C1(
        keyinput_g91), .C2(P3_DATAO_REG_5__SCAN_IN), .A(n15679), .ZN(n15684)
         );
  OAI22_X1 U17241 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(keyinput_g103), .B1(
        P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .ZN(n15680) );
  AOI221_X1 U17242 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(keyinput_g103), .C1(
        keyinput_g85), .C2(P3_DATAO_REG_11__SCAN_IN), .A(n15680), .ZN(n15683)
         );
  OAI22_X1 U17243 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        P3_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .ZN(n15681) );
  AOI221_X1 U17244 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        keyinput_g82), .C2(P3_DATAO_REG_14__SCAN_IN), .A(n15681), .ZN(n15682)
         );
  NAND4_X1 U17245 ( .A1(n15685), .A2(n15684), .A3(n15683), .A4(n15682), .ZN(
        n15713) );
  OAI22_X1 U17246 ( .A1(SI_27_), .A2(keyinput_g5), .B1(keyinput_g108), .B2(
        P1_IR_REG_1__SCAN_IN), .ZN(n15686) );
  AOI221_X1 U17247 ( .B1(SI_27_), .B2(keyinput_g5), .C1(P1_IR_REG_1__SCAN_IN), 
        .C2(keyinput_g108), .A(n15686), .ZN(n15693) );
  OAI22_X1 U17248 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_g102), .ZN(n15687) );
  AOI221_X1 U17249 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        keyinput_g102), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n15687), .ZN(n15692)
         );
  OAI22_X1 U17250 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(SI_2_), .B2(keyinput_g30), .ZN(n15688) );
  AOI221_X1 U17251 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        keyinput_g30), .C2(SI_2_), .A(n15688), .ZN(n15691) );
  OAI22_X1 U17252 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        keyinput_g24), .B2(SI_8_), .ZN(n15689) );
  AOI221_X1 U17253 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        SI_8_), .C2(keyinput_g24), .A(n15689), .ZN(n15690) );
  NAND4_X1 U17254 ( .A1(n15693), .A2(n15692), .A3(n15691), .A4(n15690), .ZN(
        n15712) );
  OAI22_X1 U17255 ( .A1(P3_B_REG_SCAN_IN), .A2(keyinput_g64), .B1(keyinput_g43), .B2(P3_REG3_REG_8__SCAN_IN), .ZN(n15694) );
  AOI221_X1 U17256 ( .B1(P3_B_REG_SCAN_IN), .B2(keyinput_g64), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput_g43), .A(n15694), .ZN(n15701) );
  OAI22_X1 U17257 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_g117), .B1(
        P3_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .ZN(n15695) );
  AOI221_X1 U17258 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_g117), .C1(
        keyinput_g69), .C2(P3_DATAO_REG_27__SCAN_IN), .A(n15695), .ZN(n15700)
         );
  OAI22_X1 U17259 ( .A1(SI_28_), .A2(keyinput_g4), .B1(SI_11_), .B2(
        keyinput_g21), .ZN(n15696) );
  AOI221_X1 U17260 ( .B1(SI_28_), .B2(keyinput_g4), .C1(keyinput_g21), .C2(
        SI_11_), .A(n15696), .ZN(n15699) );
  OAI22_X1 U17261 ( .A1(SI_14_), .A2(keyinput_g18), .B1(
        P3_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .ZN(n15697) );
  AOI221_X1 U17262 ( .B1(SI_14_), .B2(keyinput_g18), .C1(keyinput_g78), .C2(
        P3_DATAO_REG_18__SCAN_IN), .A(n15697), .ZN(n15698) );
  NAND4_X1 U17263 ( .A1(n15701), .A2(n15700), .A3(n15699), .A4(n15698), .ZN(
        n15711) );
  OAI22_X1 U17264 ( .A1(SI_25_), .A2(keyinput_g7), .B1(P3_RD_REG_SCAN_IN), 
        .B2(keyinput_g33), .ZN(n15702) );
  AOI221_X1 U17265 ( .B1(SI_25_), .B2(keyinput_g7), .C1(keyinput_g33), .C2(
        P3_RD_REG_SCAN_IN), .A(n15702), .ZN(n15709) );
  OAI22_X1 U17266 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        keyinput_g125), .B2(P1_IR_REG_18__SCAN_IN), .ZN(n15703) );
  AOI221_X1 U17267 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_g125), .A(n15703), .ZN(n15708) );
  OAI22_X1 U17268 ( .A1(SI_6_), .A2(keyinput_g26), .B1(keyinput_g2), .B2(
        SI_30_), .ZN(n15704) );
  AOI221_X1 U17269 ( .B1(SI_6_), .B2(keyinput_g26), .C1(SI_30_), .C2(
        keyinput_g2), .A(n15704), .ZN(n15707) );
  OAI22_X1 U17270 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_g115), .B1(
        P3_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .ZN(n15705) );
  AOI221_X1 U17271 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_g115), .C1(
        keyinput_g68), .C2(P3_DATAO_REG_28__SCAN_IN), .A(n15705), .ZN(n15706)
         );
  NAND4_X1 U17272 ( .A1(n15709), .A2(n15708), .A3(n15707), .A4(n15706), .ZN(
        n15710) );
  NOR4_X1 U17273 ( .A1(n15713), .A2(n15712), .A3(n15711), .A4(n15710), .ZN(
        n15913) );
  XOR2_X1 U17274 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_f76), .Z(n15720)
         );
  AOI22_X1 U17275 ( .A1(keyinput_f72), .A2(P3_DATAO_REG_24__SCAN_IN), .B1(
        keyinput_f83), .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n15714) );
  OAI221_X1 U17276 ( .B1(keyinput_f72), .B2(P3_DATAO_REG_24__SCAN_IN), .C1(
        keyinput_f83), .C2(P3_DATAO_REG_13__SCAN_IN), .A(n15714), .ZN(n15719)
         );
  AOI22_X1 U17277 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(SI_13_), .B2(keyinput_f19), .ZN(n15715) );
  OAI221_X1 U17278 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        SI_13_), .C2(keyinput_f19), .A(n15715), .ZN(n15718) );
  AOI22_X1 U17279 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_f124), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_f126), .ZN(n15716) );
  OAI221_X1 U17280 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_f124), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_f126), .A(n15716), .ZN(n15717) );
  NOR4_X1 U17281 ( .A1(n15720), .A2(n15719), .A3(n15718), .A4(n15717), .ZN(
        n15748) );
  AOI22_X1 U17282 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n15721) );
  OAI221_X1 U17283 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n15721), .ZN(n15728)
         );
  AOI22_X1 U17284 ( .A1(keyinput_f0), .A2(P3_WR_REG_SCAN_IN), .B1(SI_18_), 
        .B2(keyinput_f14), .ZN(n15722) );
  OAI221_X1 U17285 ( .B1(keyinput_f0), .B2(P3_WR_REG_SCAN_IN), .C1(SI_18_), 
        .C2(keyinput_f14), .A(n15722), .ZN(n15727) );
  AOI22_X1 U17286 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_f127), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .ZN(n15723) );
  OAI221_X1 U17287 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_f127), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n15723), .ZN(n15726) );
  AOI22_X1 U17288 ( .A1(keyinput_f88), .A2(P3_DATAO_REG_8__SCAN_IN), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n15724) );
  OAI221_X1 U17289 ( .B1(keyinput_f88), .B2(P3_DATAO_REG_8__SCAN_IN), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n15724), .ZN(n15725)
         );
  NOR4_X1 U17290 ( .A1(n15728), .A2(n15727), .A3(n15726), .A4(n15725), .ZN(
        n15747) );
  AOI22_X1 U17291 ( .A1(SI_11_), .A2(keyinput_f21), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n15729) );
  OAI221_X1 U17292 ( .B1(SI_11_), .B2(keyinput_f21), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n15729), .ZN(n15736)
         );
  AOI22_X1 U17293 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_f117), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n15730) );
  OAI221_X1 U17294 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_f117), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n15730), .ZN(n15735)
         );
  AOI22_X1 U17295 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_f114), .B1(SI_17_), 
        .B2(keyinput_f15), .ZN(n15731) );
  OAI221_X1 U17296 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_f114), .C1(SI_17_), .C2(keyinput_f15), .A(n15731), .ZN(n15734) );
  AOI22_X1 U17297 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_f107), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput_f116), .ZN(n15732) );
  OAI221_X1 U17298 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_f107), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_f116), .A(n15732), .ZN(n15733) );
  NOR4_X1 U17299 ( .A1(n15736), .A2(n15735), .A3(n15734), .A4(n15733), .ZN(
        n15746) );
  AOI22_X1 U17300 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f115), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_f119), .ZN(n15737) );
  OAI221_X1 U17301 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f115), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_f119), .A(n15737), .ZN(n15744) );
  AOI22_X1 U17302 ( .A1(keyinput_f80), .A2(P3_DATAO_REG_16__SCAN_IN), .B1(
        SI_31_), .B2(keyinput_f1), .ZN(n15738) );
  OAI221_X1 U17303 ( .B1(keyinput_f80), .B2(P3_DATAO_REG_16__SCAN_IN), .C1(
        SI_31_), .C2(keyinput_f1), .A(n15738), .ZN(n15743) );
  AOI22_X1 U17304 ( .A1(keyinput_f91), .A2(P3_DATAO_REG_5__SCAN_IN), .B1(
        P3_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .ZN(n15739) );
  OAI221_X1 U17305 ( .B1(keyinput_f91), .B2(P3_DATAO_REG_5__SCAN_IN), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n15739), .ZN(n15742)
         );
  AOI22_X1 U17306 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(keyinput_f100), .B1(SI_1_), .B2(keyinput_f31), .ZN(n15740) );
  OAI221_X1 U17307 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(keyinput_f100), .C1(
        SI_1_), .C2(keyinput_f31), .A(n15740), .ZN(n15741) );
  NOR4_X1 U17308 ( .A1(n15744), .A2(n15743), .A3(n15742), .A4(n15741), .ZN(
        n15745) );
  NAND4_X1 U17309 ( .A1(n15748), .A2(n15747), .A3(n15746), .A4(n15745), .ZN(
        n15907) );
  AOI22_X1 U17310 ( .A1(keyinput_f90), .A2(P3_DATAO_REG_6__SCAN_IN), .B1(
        keyinput_f77), .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n15749) );
  OAI221_X1 U17311 ( .B1(keyinput_f90), .B2(P3_DATAO_REG_6__SCAN_IN), .C1(
        keyinput_f77), .C2(P3_DATAO_REG_19__SCAN_IN), .A(n15749), .ZN(n15756)
         );
  AOI22_X1 U17312 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_4_), .B2(
        keyinput_f28), .ZN(n15750) );
  OAI221_X1 U17313 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_4_), .C2(
        keyinput_f28), .A(n15750), .ZN(n15755) );
  AOI22_X1 U17314 ( .A1(SI_21_), .A2(keyinput_f11), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n15751) );
  OAI221_X1 U17315 ( .B1(SI_21_), .B2(keyinput_f11), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n15751), .ZN(n15754)
         );
  AOI22_X1 U17316 ( .A1(keyinput_f71), .A2(P3_DATAO_REG_25__SCAN_IN), .B1(
        P3_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n15752) );
  OAI221_X1 U17317 ( .B1(keyinput_f71), .B2(P3_DATAO_REG_25__SCAN_IN), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_f56), .A(n15752), .ZN(n15753)
         );
  NOR4_X1 U17318 ( .A1(n15756), .A2(n15755), .A3(n15754), .A4(n15753), .ZN(
        n15784) );
  AOI22_X1 U17319 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P3_REG3_REG_8__SCAN_IN), 
        .B2(keyinput_f43), .ZN(n15757) );
  OAI221_X1 U17320 ( .B1(SI_23_), .B2(keyinput_f9), .C1(P3_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n15757), .ZN(n15764) );
  AOI22_X1 U17321 ( .A1(keyinput_f65), .A2(P3_DATAO_REG_31__SCAN_IN), .B1(
        P3_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n15758) );
  OAI221_X1 U17322 ( .B1(keyinput_f65), .B2(P3_DATAO_REG_31__SCAN_IN), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n15758), .ZN(n15763) );
  AOI22_X1 U17323 ( .A1(keyinput_f84), .A2(P3_DATAO_REG_12__SCAN_IN), .B1(
        keyinput_f89), .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n15759) );
  OAI221_X1 U17324 ( .B1(keyinput_f84), .B2(P3_DATAO_REG_12__SCAN_IN), .C1(
        keyinput_f89), .C2(P3_DATAO_REG_7__SCAN_IN), .A(n15759), .ZN(n15762)
         );
  AOI22_X1 U17325 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(keyinput_f103), .B1(SI_7_), .B2(keyinput_f25), .ZN(n15760) );
  OAI221_X1 U17326 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(keyinput_f103), .C1(
        SI_7_), .C2(keyinput_f25), .A(n15760), .ZN(n15761) );
  NOR4_X1 U17327 ( .A1(n15764), .A2(n15763), .A3(n15762), .A4(n15761), .ZN(
        n15783) );
  AOI22_X1 U17328 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(keyinput_f102), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .ZN(n15765) );
  OAI221_X1 U17329 ( .B1(P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_f102), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n15765), .ZN(n15772) );
  AOI22_X1 U17330 ( .A1(keyinput_f94), .A2(P3_DATAO_REG_2__SCAN_IN), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_f112), .ZN(n15766) );
  OAI221_X1 U17331 ( .B1(keyinput_f94), .B2(P3_DATAO_REG_2__SCAN_IN), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_f112), .A(n15766), .ZN(n15771) );
  AOI22_X1 U17332 ( .A1(keyinput_f85), .A2(P3_DATAO_REG_11__SCAN_IN), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_f110), .ZN(n15767) );
  OAI221_X1 U17333 ( .B1(keyinput_f85), .B2(P3_DATAO_REG_11__SCAN_IN), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput_f110), .A(n15767), .ZN(n15770) );
  AOI22_X1 U17334 ( .A1(keyinput_f69), .A2(P3_DATAO_REG_27__SCAN_IN), .B1(
        P3_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .ZN(n15768) );
  OAI221_X1 U17335 ( .B1(keyinput_f69), .B2(P3_DATAO_REG_27__SCAN_IN), .C1(
        P3_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n15768), .ZN(n15769) );
  NOR4_X1 U17336 ( .A1(n15772), .A2(n15771), .A3(n15770), .A4(n15769), .ZN(
        n15782) );
  AOI22_X1 U17337 ( .A1(SI_22_), .A2(keyinput_f10), .B1(SI_29_), .B2(
        keyinput_f3), .ZN(n15773) );
  OAI221_X1 U17338 ( .B1(SI_22_), .B2(keyinput_f10), .C1(SI_29_), .C2(
        keyinput_f3), .A(n15773), .ZN(n15780) );
  AOI22_X1 U17339 ( .A1(keyinput_f66), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput_f113), .ZN(n15774) );
  OAI221_X1 U17340 ( .B1(keyinput_f66), .B2(P3_DATAO_REG_30__SCAN_IN), .C1(
        P1_IR_REG_6__SCAN_IN), .C2(keyinput_f113), .A(n15774), .ZN(n15779) );
  AOI22_X1 U17341 ( .A1(SI_27_), .A2(keyinput_f5), .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n15775) );
  OAI221_X1 U17342 ( .B1(SI_27_), .B2(keyinput_f5), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n15775), .ZN(n15778)
         );
  AOI22_X1 U17343 ( .A1(keyinput_f70), .A2(P3_DATAO_REG_26__SCAN_IN), .B1(
        P1_IR_REG_1__SCAN_IN), .B2(keyinput_f108), .ZN(n15776) );
  OAI221_X1 U17344 ( .B1(keyinput_f70), .B2(P3_DATAO_REG_26__SCAN_IN), .C1(
        P1_IR_REG_1__SCAN_IN), .C2(keyinput_f108), .A(n15776), .ZN(n15777) );
  NOR4_X1 U17345 ( .A1(n15780), .A2(n15779), .A3(n15778), .A4(n15777), .ZN(
        n15781) );
  NAND4_X1 U17346 ( .A1(n15784), .A2(n15783), .A3(n15782), .A4(n15781), .ZN(
        n15906) );
  AOI22_X1 U17347 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_f125), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n15785) );
  OAI221_X1 U17348 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_f125), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n15785), .ZN(n15794)
         );
  AOI22_X1 U17349 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f118), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_f120), .ZN(n15786) );
  OAI221_X1 U17350 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f118), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_f120), .A(n15786), .ZN(n15793) );
  AOI22_X1 U17351 ( .A1(SI_24_), .A2(keyinput_f8), .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n15787) );
  OAI221_X1 U17352 ( .B1(SI_24_), .B2(keyinput_f8), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n15787), .ZN(n15792)
         );
  AOI22_X1 U17353 ( .A1(n15790), .A2(keyinput_f55), .B1(keyinput_f23), .B2(
        n15789), .ZN(n15788) );
  OAI221_X1 U17354 ( .B1(n15790), .B2(keyinput_f55), .C1(n15789), .C2(
        keyinput_f23), .A(n15788), .ZN(n15791) );
  NOR4_X1 U17355 ( .A1(n15794), .A2(n15793), .A3(n15792), .A4(n15791), .ZN(
        n15841) );
  AOI22_X1 U17356 ( .A1(n15797), .A2(keyinput_f58), .B1(keyinput_f75), .B2(
        n15796), .ZN(n15795) );
  OAI221_X1 U17357 ( .B1(n15797), .B2(keyinput_f58), .C1(n15796), .C2(
        keyinput_f75), .A(n15795), .ZN(n15807) );
  AOI22_X1 U17358 ( .A1(n15800), .A2(keyinput_f24), .B1(n15799), .B2(
        keyinput_f4), .ZN(n15798) );
  OAI221_X1 U17359 ( .B1(n15800), .B2(keyinput_f24), .C1(n15799), .C2(
        keyinput_f4), .A(n15798), .ZN(n15806) );
  XOR2_X1 U17360 ( .A(n9529), .B(keyinput_f109), .Z(n15804) );
  XNOR2_X1 U17361 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_f123), .ZN(n15803)
         );
  XNOR2_X1 U17362 ( .A(SI_2_), .B(keyinput_f30), .ZN(n15802) );
  XNOR2_X1 U17363 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_f54), .ZN(n15801)
         );
  NAND4_X1 U17364 ( .A1(n15804), .A2(n15803), .A3(n15802), .A4(n15801), .ZN(
        n15805) );
  NOR3_X1 U17365 ( .A1(n15807), .A2(n15806), .A3(n15805), .ZN(n15840) );
  AOI22_X1 U17366 ( .A1(n15810), .A2(keyinput_f87), .B1(keyinput_f73), .B2(
        n15809), .ZN(n15808) );
  OAI221_X1 U17367 ( .B1(n15810), .B2(keyinput_f87), .C1(n15809), .C2(
        keyinput_f73), .A(n15808), .ZN(n15820) );
  AOI22_X1 U17368 ( .A1(n15812), .A2(keyinput_f62), .B1(keyinput_f32), .B2(
        n10135), .ZN(n15811) );
  OAI221_X1 U17369 ( .B1(n15812), .B2(keyinput_f62), .C1(n10135), .C2(
        keyinput_f32), .A(n15811), .ZN(n15819) );
  AOI22_X1 U17370 ( .A1(n8790), .A2(keyinput_f53), .B1(keyinput_f20), .B2(
        n15814), .ZN(n15813) );
  OAI221_X1 U17371 ( .B1(n8790), .B2(keyinput_f53), .C1(n15814), .C2(
        keyinput_f20), .A(n15813), .ZN(n15818) );
  XNOR2_X1 U17372 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f111), .ZN(n15816)
         );
  XNOR2_X1 U17373 ( .A(SI_16_), .B(keyinput_f16), .ZN(n15815) );
  NAND2_X1 U17374 ( .A1(n15816), .A2(n15815), .ZN(n15817) );
  NOR4_X1 U17375 ( .A1(n15820), .A2(n15819), .A3(n15818), .A4(n15817), .ZN(
        n15839) );
  AOI22_X1 U17376 ( .A1(n15823), .A2(keyinput_f22), .B1(keyinput_f105), .B2(
        n15822), .ZN(n15821) );
  OAI221_X1 U17377 ( .B1(n15823), .B2(keyinput_f22), .C1(n15822), .C2(
        keyinput_f105), .A(n15821), .ZN(n15830) );
  AOI22_X1 U17378 ( .A1(n15826), .A2(keyinput_f122), .B1(n15825), .B2(
        keyinput_f64), .ZN(n15824) );
  OAI221_X1 U17379 ( .B1(n15826), .B2(keyinput_f122), .C1(n15825), .C2(
        keyinput_f64), .A(n15824), .ZN(n15829) );
  XNOR2_X1 U17380 ( .A(n15827), .B(keyinput_f121), .ZN(n15828) );
  OR3_X1 U17381 ( .A1(n15830), .A2(n15829), .A3(n15828), .ZN(n15837) );
  AOI22_X1 U17382 ( .A1(n15833), .A2(keyinput_f86), .B1(keyinput_f92), .B2(
        n15832), .ZN(n15831) );
  OAI221_X1 U17383 ( .B1(n15833), .B2(keyinput_f86), .C1(n15832), .C2(
        keyinput_f92), .A(n15831), .ZN(n15836) );
  XNOR2_X1 U17384 ( .A(n15834), .B(keyinput_f82), .ZN(n15835) );
  NOR3_X1 U17385 ( .A1(n15837), .A2(n15836), .A3(n15835), .ZN(n15838) );
  NAND4_X1 U17386 ( .A1(n15841), .A2(n15840), .A3(n15839), .A4(n15838), .ZN(
        n15905) );
  AOI22_X1 U17387 ( .A1(n15844), .A2(keyinput_f12), .B1(n15843), .B2(
        keyinput_f26), .ZN(n15842) );
  OAI221_X1 U17388 ( .B1(n15844), .B2(keyinput_f12), .C1(n15843), .C2(
        keyinput_f26), .A(n15842), .ZN(n15857) );
  AOI22_X1 U17389 ( .A1(n15847), .A2(keyinput_f51), .B1(keyinput_f7), .B2(
        n15846), .ZN(n15845) );
  OAI221_X1 U17390 ( .B1(n15847), .B2(keyinput_f51), .C1(n15846), .C2(
        keyinput_f7), .A(n15845), .ZN(n15856) );
  AOI22_X1 U17391 ( .A1(n15850), .A2(keyinput_f93), .B1(n15849), .B2(
        keyinput_f39), .ZN(n15848) );
  OAI221_X1 U17392 ( .B1(n15850), .B2(keyinput_f93), .C1(n15849), .C2(
        keyinput_f39), .A(n15848), .ZN(n15855) );
  AOI22_X1 U17393 ( .A1(n15853), .A2(keyinput_f47), .B1(keyinput_f106), .B2(
        n15852), .ZN(n15851) );
  OAI221_X1 U17394 ( .B1(n15853), .B2(keyinput_f47), .C1(n15852), .C2(
        keyinput_f106), .A(n15851), .ZN(n15854) );
  NOR4_X1 U17395 ( .A1(n15857), .A2(n15856), .A3(n15855), .A4(n15854), .ZN(
        n15903) );
  AOI22_X1 U17396 ( .A1(P3_U3151), .A2(keyinput_f34), .B1(keyinput_f67), .B2(
        n15859), .ZN(n15858) );
  OAI221_X1 U17397 ( .B1(P3_U3151), .B2(keyinput_f34), .C1(n15859), .C2(
        keyinput_f67), .A(n15858), .ZN(n15871) );
  AOI22_X1 U17398 ( .A1(n8720), .A2(keyinput_f49), .B1(keyinput_f97), .B2(
        n15861), .ZN(n15860) );
  OAI221_X1 U17399 ( .B1(n8720), .B2(keyinput_f49), .C1(n15861), .C2(
        keyinput_f97), .A(n15860), .ZN(n15870) );
  INV_X1 U17400 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15863) );
  AOI22_X1 U17401 ( .A1(n15864), .A2(keyinput_f98), .B1(n15863), .B2(
        keyinput_f38), .ZN(n15862) );
  OAI221_X1 U17402 ( .B1(n15864), .B2(keyinput_f98), .C1(n15863), .C2(
        keyinput_f38), .A(n15862), .ZN(n15869) );
  AOI22_X1 U17403 ( .A1(n15867), .A2(keyinput_f27), .B1(keyinput_f95), .B2(
        n15866), .ZN(n15865) );
  OAI221_X1 U17404 ( .B1(n15867), .B2(keyinput_f27), .C1(n15866), .C2(
        keyinput_f95), .A(n15865), .ZN(n15868) );
  NOR4_X1 U17405 ( .A1(n15871), .A2(n15870), .A3(n15869), .A4(n15868), .ZN(
        n15902) );
  AOI22_X1 U17406 ( .A1(n15873), .A2(keyinput_f18), .B1(n9017), .B2(
        keyinput_f45), .ZN(n15872) );
  OAI221_X1 U17407 ( .B1(n15873), .B2(keyinput_f18), .C1(n9017), .C2(
        keyinput_f45), .A(n15872), .ZN(n15884) );
  AOI22_X1 U17408 ( .A1(n15875), .A2(keyinput_f17), .B1(keyinput_f104), .B2(
        n10962), .ZN(n15874) );
  OAI221_X1 U17409 ( .B1(n15875), .B2(keyinput_f17), .C1(n10962), .C2(
        keyinput_f104), .A(n15874), .ZN(n15883) );
  AOI22_X1 U17410 ( .A1(n7067), .A2(keyinput_f29), .B1(keyinput_f6), .B2(
        n15877), .ZN(n15876) );
  OAI221_X1 U17411 ( .B1(n7067), .B2(keyinput_f29), .C1(n15877), .C2(
        keyinput_f6), .A(n15876), .ZN(n15882) );
  AOI22_X1 U17412 ( .A1(n15880), .A2(keyinput_f96), .B1(keyinput_f68), .B2(
        n15879), .ZN(n15878) );
  OAI221_X1 U17413 ( .B1(n15880), .B2(keyinput_f96), .C1(n15879), .C2(
        keyinput_f68), .A(n15878), .ZN(n15881) );
  NOR4_X1 U17414 ( .A1(n15884), .A2(n15883), .A3(n15882), .A4(n15881), .ZN(
        n15901) );
  AOI22_X1 U17415 ( .A1(n15887), .A2(keyinput_f101), .B1(keyinput_f33), .B2(
        n15886), .ZN(n15885) );
  OAI221_X1 U17416 ( .B1(n15887), .B2(keyinput_f101), .C1(n15886), .C2(
        keyinput_f33), .A(n15885), .ZN(n15899) );
  AOI22_X1 U17417 ( .A1(n15890), .A2(keyinput_f74), .B1(keyinput_f79), .B2(
        n15889), .ZN(n15888) );
  OAI221_X1 U17418 ( .B1(n15890), .B2(keyinput_f74), .C1(n15889), .C2(
        keyinput_f79), .A(n15888), .ZN(n15898) );
  AOI22_X1 U17419 ( .A1(n15892), .A2(keyinput_f78), .B1(n8670), .B2(
        keyinput_f59), .ZN(n15891) );
  OAI221_X1 U17420 ( .B1(n15892), .B2(keyinput_f78), .C1(n8670), .C2(
        keyinput_f59), .A(n15891), .ZN(n15897) );
  AOI22_X1 U17421 ( .A1(n15895), .A2(keyinput_f13), .B1(keyinput_f99), .B2(
        n15894), .ZN(n15893) );
  OAI221_X1 U17422 ( .B1(n15895), .B2(keyinput_f13), .C1(n15894), .C2(
        keyinput_f99), .A(n15893), .ZN(n15896) );
  NOR4_X1 U17423 ( .A1(n15899), .A2(n15898), .A3(n15897), .A4(n15896), .ZN(
        n15900) );
  NAND4_X1 U17424 ( .A1(n15903), .A2(n15902), .A3(n15901), .A4(n15900), .ZN(
        n15904) );
  OR4_X1 U17425 ( .A1(n15907), .A2(n15906), .A3(n15905), .A4(n15904), .ZN(
        n15909) );
  AOI21_X1 U17426 ( .B1(keyinput_f81), .B2(n15909), .A(keyinput_g81), .ZN(
        n15911) );
  INV_X1 U17427 ( .A(keyinput_f81), .ZN(n15908) );
  AOI21_X1 U17428 ( .B1(n15909), .B2(n15908), .A(P3_DATAO_REG_15__SCAN_IN), 
        .ZN(n15910) );
  AOI22_X1 U17429 ( .A1(P3_DATAO_REG_15__SCAN_IN), .A2(n15911), .B1(
        keyinput_g81), .B2(n15910), .ZN(n15912) );
  AOI21_X1 U17430 ( .B1(n15914), .B2(n15913), .A(n15912), .ZN(n15917) );
  XNOR2_X1 U17431 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15915) );
  XNOR2_X1 U17432 ( .A(n7690), .B(n15915), .ZN(n15916) );
  XNOR2_X1 U17433 ( .A(n15917), .B(n15916), .ZN(n15920) );
  AOI21_X1 U17434 ( .B1(n15924), .B2(n15923), .A(n15922), .ZN(SUB_1596_U59) );
  OAI21_X1 U17435 ( .B1(n15927), .B2(n15926), .A(n15925), .ZN(SUB_1596_U58) );
  XNOR2_X1 U17436 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15928), .ZN(SUB_1596_U53)
         );
  OAI21_X1 U17437 ( .B1(n15931), .B2(n15930), .A(n15929), .ZN(SUB_1596_U56) );
  AOI21_X1 U17438 ( .B1(n15934), .B2(n15933), .A(n15932), .ZN(n15935) );
  XOR2_X1 U17439 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15935), .Z(SUB_1596_U60) );
  AOI21_X1 U17440 ( .B1(n15938), .B2(n15937), .A(n15936), .ZN(SUB_1596_U5) );
  INV_X1 U7504 ( .A(n13243), .ZN(n7296) );
  CLKBUF_X1 U7505 ( .A(n9154), .Z(n7003) );
  INV_X1 U7614 ( .A(n7914), .ZN(n8150) );
  INV_X1 U9668 ( .A(n12445), .ZN(n9550) );
  NAND2_X1 U9944 ( .A1(n9550), .A2(n7588), .ZN(n9886) );
endmodule

