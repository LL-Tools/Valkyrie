

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979;

  NAND2_X1 U4780 ( .A1(n6045), .A2(n6044), .ZN(n6253) );
  INV_X2 U4781 ( .A(n5653), .ZN(n7320) );
  INV_X1 U4782 ( .A(n5450), .ZN(n7522) );
  CLKBUF_X1 U4783 ( .A(n5566), .Z(n4277) );
  CLKBUF_X2 U4784 ( .A(n5566), .Z(n4278) );
  NAND3_X1 U4785 ( .A1(n5109), .A2(n5107), .A3(n5108), .ZN(n8702) );
  NAND2_X2 U4786 ( .A1(n5212), .A2(n8934), .ZN(n9652) );
  BUF_X2 U4787 ( .A(n8679), .Z(n4280) );
  INV_X1 U4788 ( .A(n5281), .ZN(n5881) );
  NAND2_X1 U4789 ( .A1(n5112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U4790 ( .A1(n4309), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4846) );
  NOR2_X2 U4791 ( .A1(n5051), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5078) );
  CLKBUF_X1 U4792 ( .A(n8669), .Z(n4275) );
  NOR2_X1 U4793 ( .A1(n5527), .A2(n5526), .ZN(n8669) );
  OR2_X1 U4794 ( .A1(n7619), .A2(n7618), .ZN(n7631) );
  INV_X1 U4795 ( .A(n7690), .ZN(n7671) );
  OR2_X1 U4796 ( .A1(n5279), .A2(n5653), .ZN(n5282) );
  INV_X1 U4797 ( .A(n7319), .ZN(n7289) );
  NAND2_X1 U4798 ( .A1(n5881), .A2(n5231), .ZN(n7318) );
  NAND2_X1 U4799 ( .A1(n5466), .A2(n7532), .ZN(n5718) );
  INV_X2 U4800 ( .A(n4287), .ZN(n7473) );
  INV_X1 U4801 ( .A(n7286), .ZN(n7322) );
  INV_X1 U4802 ( .A(n8687), .ZN(n7086) );
  INV_X1 U4803 ( .A(n5554), .ZN(n6486) );
  NOR2_X1 U4805 ( .A1(n7354), .A2(n8495), .ZN(n7355) );
  INV_X1 U4806 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8522) );
  AND3_X1 U4807 ( .A1(n5517), .A2(n5516), .A3(n5515), .ZN(n9683) );
  NAND2_X1 U4808 ( .A1(n5073), .A2(n5072), .ZN(n5084) );
  AND2_X1 U4809 ( .A1(n7449), .A2(n7669), .ZN(n8102) );
  NAND2_X1 U4810 ( .A1(n4842), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4844) );
  INV_X1 U4811 ( .A(n7738), .ZN(n6642) );
  INV_X1 U4812 ( .A(n9654), .ZN(n8701) );
  AOI21_X1 U4813 ( .B1(n9232), .B2(n5254), .A(n5259), .ZN(n9242) );
  INV_X1 U4814 ( .A(n9188), .ZN(n9638) );
  OAI21_X1 U4815 ( .B1(n4923), .B2(n4922), .A(n4921), .ZN(n9006) );
  OR2_X1 U4818 ( .A1(n8945), .A2(n8944), .ZN(n4276) );
  INV_X4 U4819 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4911) );
  NOR2_X4 U4820 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4771) );
  OAI22_X2 U4824 ( .A1(n5169), .A2(n5168), .B1(n6053), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n5163) );
  INV_X2 U4825 ( .A(n6526), .ZN(n9850) );
  NAND2_X1 U4826 ( .A1(n7556), .A2(n7554), .ZN(n5470) );
  NAND2_X2 U4827 ( .A1(n4860), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4857) );
  NAND2_X2 U4828 ( .A1(n8523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5114) );
  OAI21_X2 U4829 ( .B1(n9412), .B2(P1_IR_REG_29__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5098) );
  XNOR2_X2 U4830 ( .A(n4983), .B(SI_2_), .ZN(n4981) );
  NAND2_X1 U4831 ( .A1(n5120), .A2(n5451), .ZN(n5566) );
  OAI21_X2 U4832 ( .B1(n6253), .B2(n6252), .A(n6251), .ZN(n6259) );
  XNOR2_X2 U4833 ( .A(n4844), .B(n4843), .ZN(n7333) );
  XNOR2_X2 U4834 ( .A(n5380), .B(n5382), .ZN(n5383) );
  INV_X2 U4835 ( .A(n6985), .ZN(n5450) );
  BUF_X4 U4836 ( .A(n5580), .Z(n4279) );
  NAND2_X1 U4837 ( .A1(n4582), .A2(n4587), .ZN(n7915) );
  NAND2_X1 U4838 ( .A1(n7438), .A2(n7437), .ZN(n8432) );
  MUX2_X1 U4839 ( .A(n7602), .B(n7601), .S(n7690), .Z(n7603) );
  INV_X1 U4840 ( .A(n8696), .ZN(n9518) );
  NAND2_X1 U4841 ( .A1(n6814), .A2(n6813), .ZN(n8495) );
  NAND2_X1 U4842 ( .A1(n6709), .A2(n6708), .ZN(n9523) );
  NAND2_X1 U4843 ( .A1(n6451), .A2(n6450), .ZN(n6491) );
  XNOR2_X1 U4844 ( .A(n5084), .B(n4828), .ZN(n6384) );
  NAND2_X1 U4845 ( .A1(n7583), .A2(n7584), .ZN(n7706) );
  AND2_X2 U4846 ( .A1(n4726), .A2(n9652), .ZN(n7286) );
  NOR2_X2 U4847 ( .A1(n8702), .A2(n8701), .ZN(n8886) );
  NAND4_X1 U4848 ( .A1(n5478), .A2(n5477), .A3(n5476), .A4(n5475), .ZN(n7940)
         );
  INV_X4 U4849 ( .A(n5255), .ZN(n8683) );
  CLKBUF_X2 U4850 ( .A(n5425), .Z(n7167) );
  CLKBUF_X1 U4851 ( .A(n5513), .Z(n8687) );
  BUF_X1 U4853 ( .A(n5285), .Z(n5846) );
  CLKBUF_X1 U4854 ( .A(n8995), .Z(n4283) );
  AOI21_X1 U4855 ( .B1(n4619), .B2(n4618), .A(n7679), .ZN(n7686) );
  OAI21_X1 U4856 ( .B1(n7915), .B2(n7787), .A(n7786), .ZN(n7788) );
  AOI21_X1 U4857 ( .B1(n8090), .B2(n9776), .A(n8089), .ZN(n8428) );
  AOI21_X1 U4858 ( .B1(n4779), .B2(n4783), .A(n4366), .ZN(n4777) );
  NOR2_X1 U4859 ( .A1(n8070), .A2(n8415), .ZN(n8063) );
  OR2_X1 U4860 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  NAND2_X1 U4861 ( .A1(n7234), .A2(n7233), .ZN(n8662) );
  AND2_X1 U4862 ( .A1(n4460), .A2(n4458), .ZN(n9214) );
  AOI21_X1 U4863 ( .B1(n4762), .B2(n4760), .A(n4335), .ZN(n4759) );
  OAI21_X1 U4864 ( .B1(n8369), .B2(n8368), .A(n7627), .ZN(n8350) );
  AOI21_X1 U4865 ( .B1(n9378), .B2(n8959), .A(n7095), .ZN(n9238) );
  NAND2_X1 U4866 ( .A1(n6695), .A2(n6692), .ZN(n6742) );
  OR2_X1 U4867 ( .A1(n8170), .A2(n8030), .ZN(n4823) );
  NAND2_X1 U4868 ( .A1(n7387), .A2(n7386), .ZN(n8457) );
  INV_X1 U4869 ( .A(n9264), .ZN(n9378) );
  INV_X1 U4870 ( .A(n6562), .ZN(n4281) );
  NAND2_X1 U4871 ( .A1(n6714), .A2(n8789), .ZN(n8786) );
  NAND2_X1 U4872 ( .A1(n4416), .A2(n4415), .ZN(n7354) );
  NAND2_X1 U4873 ( .A1(n7082), .A2(n7081), .ZN(n9313) );
  NAND2_X1 U4874 ( .A1(n5845), .A2(n5844), .ZN(n6068) );
  AOI21_X1 U4875 ( .B1(n4553), .B2(n4551), .A(n4550), .ZN(n4549) );
  NAND2_X1 U4876 ( .A1(n6559), .A2(n6558), .ZN(n6836) );
  AOI21_X1 U4877 ( .B1(n6287), .B2(n4322), .A(n4475), .ZN(n6426) );
  NAND2_X1 U4878 ( .A1(n6586), .A2(n6585), .ZN(n6670) );
  AND2_X1 U4879 ( .A1(n8782), .A2(n8773), .ZN(n8881) );
  NAND2_X1 U4880 ( .A1(n4496), .A2(n4494), .ZN(n5614) );
  INV_X1 U4881 ( .A(n6356), .ZN(n4415) );
  AND2_X1 U4882 ( .A1(n7596), .A2(n7592), .ZN(n7708) );
  NAND2_X1 U4883 ( .A1(n6334), .A2(n6333), .ZN(n6471) );
  NAND2_X1 U4884 ( .A1(n4487), .A2(n8708), .ZN(n8755) );
  AND2_X1 U4885 ( .A1(n7588), .A2(n7589), .ZN(n7709) );
  AND2_X2 U4886 ( .A1(n6103), .A2(n9792), .ZN(n8399) );
  AND2_X2 U4887 ( .A1(n5894), .A2(n9306), .ZN(n9660) );
  INV_X1 U4888 ( .A(n5998), .ZN(n9856) );
  AND2_X2 U4889 ( .A1(n9805), .A2(n9804), .ZN(n9826) );
  NAND2_X1 U4890 ( .A1(n4630), .A2(n5818), .ZN(n5998) );
  INV_X2 U4891 ( .A(n5725), .ZN(n5560) );
  INV_X1 U4892 ( .A(n5801), .ZN(n6198) );
  NAND2_X1 U4893 ( .A1(n5573), .A2(n4399), .ZN(n5798) );
  NAND2_X4 U4894 ( .A1(n5986), .A2(n5543), .ZN(n5554) );
  AND4_X1 U4895 ( .A1(n5536), .A2(n5535), .A3(n5534), .A4(n5533), .ZN(n6120)
         );
  OAI211_X1 U4896 ( .C1(n6007), .C2(n6015), .A(n6009), .B(n4694), .ZN(n7904)
         );
  AND3_X1 U4897 ( .A1(n5724), .A2(n5723), .A3(n5722), .ZN(n5801) );
  NAND4_X2 U4898 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n8970)
         );
  CLKBUF_X2 U4899 ( .A(n5718), .Z(n4287) );
  AND4_X1 U4900 ( .A1(n5464), .A2(n5463), .A3(n5462), .A4(n5461), .ZN(n5786)
         );
  AND2_X2 U4901 ( .A1(n4946), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  CLKBUF_X1 U4902 ( .A(n5718), .Z(n4288) );
  NAND4_X1 U4903 ( .A1(n6026), .A2(n6025), .A3(n6024), .A4(n6023), .ZN(n7935)
         );
  NAND2_X1 U4904 ( .A1(n8995), .A2(n8991), .ZN(n5285) );
  NAND2_X1 U4905 ( .A1(n7796), .A2(n5103), .ZN(n5300) );
  AND2_X1 U4906 ( .A1(n7796), .A2(n7363), .ZN(n5299) );
  NAND2_X1 U4907 ( .A1(n5102), .A2(n5103), .ZN(n5425) );
  INV_X1 U4908 ( .A(n8679), .ZN(n4284) );
  XNOR2_X1 U4909 ( .A(n5059), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U4910 ( .A1(n5066), .A2(n5112), .ZN(n8009) );
  XNOR2_X1 U4911 ( .A(n4443), .B(n4863), .ZN(n8995) );
  XNOR2_X1 U4912 ( .A(n5098), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5102) );
  XNOR2_X1 U4913 ( .A(n5099), .B(n5097), .ZN(n7363) );
  NAND2_X1 U4914 ( .A1(n9412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5099) );
  XNOR2_X1 U4915 ( .A(n5043), .B(SI_7_), .ZN(n5040) );
  OR2_X1 U4916 ( .A1(n9007), .A2(n4951), .ZN(n9008) );
  MUX2_X1 U4917 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5065), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5066) );
  NAND2_X1 U4918 ( .A1(n4444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4443) );
  AND2_X1 U4919 ( .A1(n5272), .A2(n5271), .ZN(n5438) );
  OR2_X1 U4920 ( .A1(n5115), .A2(n8522), .ZN(n5117) );
  AOI21_X1 U4921 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n8973), .A(n8982), .ZN(
        n9007) );
  NAND2_X2 U4922 ( .A1(n4968), .A2(P2_U3152), .ZN(n7800) );
  INV_X8 U4923 ( .A(n4968), .ZN(n7532) );
  NAND2_X2 U4924 ( .A1(n4968), .A2(P1_U3084), .ZN(n7361) );
  AND4_X1 U4925 ( .A1(n4869), .A2(n4815), .A3(n4868), .A4(n4867), .ZN(n4824)
         );
  NAND2_X1 U4926 ( .A1(n4845), .A2(n4747), .ZN(n4746) );
  INV_X4 U4927 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4928 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5637) );
  INV_X1 U4929 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5634) );
  INV_X1 U4930 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4887) );
  INV_X1 U4931 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4891) );
  INV_X1 U4932 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5271) );
  INV_X1 U4933 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4845) );
  INV_X1 U4934 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5436) );
  INV_X1 U4935 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4747) );
  INV_X1 U4936 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8199) );
  INV_X4 U4937 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4938 ( .A(n7319), .ZN(n4282) );
  AOI21_X2 U4939 ( .B1(n8314), .B2(n8323), .A(n8029), .ZN(n8165) );
  OAI21_X2 U4940 ( .B1(n8331), .B2(n8028), .A(n4360), .ZN(n8314) );
  NAND4_X4 U4941 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n5380)
         );
  OR2_X2 U4942 ( .A1(n9368), .A2(n9242), .ZN(n8830) );
  OAI21_X2 U4943 ( .B1(n8326), .B2(n8452), .A(n8031), .ZN(n8146) );
  AND2_X2 U4944 ( .A1(n7231), .A2(n7232), .ZN(n7228) );
  NAND2_X2 U4945 ( .A1(n7225), .A2(n7224), .ZN(n7231) );
  NOR2_X2 U4947 ( .A1(n9118), .A2(n9117), .ZN(n9116) );
  NOR2_X2 U4948 ( .A1(n9137), .A2(n8743), .ZN(n9118) );
  AOI21_X2 U4949 ( .B1(n8023), .B2(n8022), .A(n8021), .ZN(n8389) );
  NAND2_X2 U4950 ( .A1(n6967), .A2(n6966), .ZN(n8023) );
  NAND2_X1 U4951 ( .A1(n5102), .A2(n7363), .ZN(n8679) );
  NAND2_X2 U4952 ( .A1(n8643), .A2(n8642), .ZN(n8648) );
  BUF_X8 U4953 ( .A(n7290), .Z(n4285) );
  NAND2_X2 U4954 ( .A1(n7259), .A2(n7258), .ZN(n8644) );
  INV_X1 U4955 ( .A(n8952), .ZN(n5212) );
  XNOR2_X2 U4956 ( .A(n4846), .B(n4845), .ZN(n6764) );
  INV_X1 U4957 ( .A(n5299), .ZN(n4286) );
  OAI22_X2 U4958 ( .A1(n6320), .A2(n4330), .B1(n4695), .B2(n4295), .ZN(n6400)
         );
  OAI211_X2 U4959 ( .C1(n5466), .C2(n5559), .A(n5558), .B(n5557), .ZN(n6526)
         );
  AOI211_X1 U4960 ( .C1(n6526), .C2(n6525), .A(n6524), .B(n9902), .ZN(n9848)
         );
  XNOR2_X2 U4961 ( .A(n5063), .B(n4813), .ZN(n5310) );
  OAI21_X1 U4962 ( .B1(n7674), .B2(n7673), .A(n4623), .ZN(n4622) );
  AND2_X1 U4963 ( .A1(n7694), .A2(n7672), .ZN(n4623) );
  NOR2_X1 U4964 ( .A1(n9167), .A2(n4485), .ZN(n4484) );
  INV_X1 U4965 ( .A(n8845), .ZN(n4485) );
  AND2_X1 U4966 ( .A1(n4765), .A2(n4342), .ZN(n4762) );
  AOI21_X1 U4967 ( .B1(n4742), .B2(n4740), .A(n4332), .ZN(n4739) );
  INV_X1 U4968 ( .A(n4743), .ZN(n4740) );
  NOR2_X1 U4969 ( .A1(n8881), .A2(n4731), .ZN(n4730) );
  INV_X1 U4970 ( .A(n6420), .ZN(n4731) );
  INV_X1 U4971 ( .A(n4746), .ZN(n4745) );
  INV_X1 U4972 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4865) );
  NOR2_X1 U4973 ( .A1(n4327), .A2(n4290), .ZN(n4618) );
  NAND2_X1 U4974 ( .A1(n5090), .A2(n5089), .ZN(n5139) );
  NAND2_X1 U4975 ( .A1(n5075), .A2(n8256), .ZN(n5085) );
  NAND2_X1 U4976 ( .A1(n6367), .A2(n6368), .ZN(n4558) );
  AND2_X1 U4977 ( .A1(n4567), .A2(n4565), .ZN(n7766) );
  AND2_X1 U4978 ( .A1(n4566), .A2(n4343), .ZN(n4565) );
  AND2_X1 U4979 ( .A1(n5365), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4653) );
  OR2_X1 U4980 ( .A1(n8426), .A2(n8036), .ZN(n7696) );
  NOR2_X1 U4981 ( .A1(n8332), .A2(n4326), .ZN(n4678) );
  OR2_X1 U4982 ( .A1(n8474), .A2(n8385), .ZN(n7627) );
  NOR2_X1 U4983 ( .A1(n6491), .A2(n6471), .ZN(n4419) );
  NAND2_X1 U4984 ( .A1(n4392), .A2(n7567), .ZN(n4391) );
  INV_X1 U4985 ( .A(n5988), .ZN(n4392) );
  NAND2_X1 U4986 ( .A1(n5458), .A2(n5459), .ZN(n7556) );
  NAND2_X1 U4987 ( .A1(n5545), .A2(n6266), .ZN(n7554) );
  NAND2_X1 U4988 ( .A1(n4380), .A2(n4361), .ZN(n8868) );
  NAND2_X1 U4989 ( .A1(n8867), .A2(n4381), .ZN(n4380) );
  AND2_X1 U4990 ( .A1(n9319), .A2(n9102), .ZN(n8938) );
  NAND2_X1 U4991 ( .A1(n9105), .A2(n8684), .ZN(n8939) );
  INV_X1 U4992 ( .A(n4463), .ZN(n4459) );
  OR2_X1 U4993 ( .A1(n9313), .A2(n9290), .ZN(n8811) );
  AOI21_X1 U4994 ( .B1(n6647), .B2(n6601), .A(n6600), .ZN(n6712) );
  AND2_X1 U4995 ( .A1(n8891), .A2(n6205), .ZN(n4735) );
  XNOR2_X1 U4996 ( .A(n7529), .B(n7528), .ZN(n7526) );
  NAND2_X1 U4997 ( .A1(n4530), .A2(n4363), .ZN(n6939) );
  NAND2_X1 U4998 ( .A1(n6763), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U4999 ( .A1(n4537), .A2(n4535), .ZN(n4534) );
  AOI21_X1 U5000 ( .B1(n4527), .B2(n6623), .A(n4365), .ZN(n4526) );
  NOR2_X1 U5001 ( .A1(n6258), .A2(n4528), .ZN(n4527) );
  NOR2_X1 U5002 ( .A1(n5262), .A2(n4505), .ZN(n4504) );
  INV_X1 U5003 ( .A(n5180), .ZN(n4505) );
  NAND2_X1 U5004 ( .A1(n4561), .A2(n4560), .ZN(n4559) );
  INV_X1 U5005 ( .A(n6129), .ZN(n4560) );
  AND2_X1 U5006 ( .A1(n4559), .A2(n4558), .ZN(n4555) );
  NAND2_X1 U5007 ( .A1(n4554), .A2(n4558), .ZN(n4553) );
  INV_X1 U5008 ( .A(n4556), .ZN(n4554) );
  AOI21_X1 U5009 ( .B1(n6131), .B2(n4559), .A(n4557), .ZN(n4556) );
  INV_X1 U5010 ( .A(n6369), .ZN(n4557) );
  INV_X1 U5011 ( .A(n5330), .ZN(n4651) );
  INV_X1 U5012 ( .A(n4633), .ZN(n7999) );
  NAND2_X1 U5013 ( .A1(n8063), .A2(n8410), .ZN(n8045) );
  INV_X1 U5014 ( .A(n8102), .ZN(n4688) );
  INV_X1 U5015 ( .A(n4398), .ZN(n4397) );
  OAI21_X1 U5016 ( .B1(n4291), .B2(n7665), .A(n4687), .ZN(n4398) );
  NAND2_X1 U5017 ( .A1(n7695), .A2(n4689), .ZN(n4687) );
  NAND2_X1 U5018 ( .A1(n7696), .A2(n7449), .ZN(n4689) );
  NAND2_X1 U5019 ( .A1(n8129), .A2(n7435), .ZN(n8119) );
  AND2_X1 U5020 ( .A1(n8120), .A2(n8118), .ZN(n7435) );
  NAND2_X1 U5021 ( .A1(n8171), .A2(n7416), .ZN(n8155) );
  AND2_X1 U5022 ( .A1(n8156), .A2(n8157), .ZN(n7416) );
  INV_X1 U5023 ( .A(n8028), .ZN(n8332) );
  NAND2_X1 U5024 ( .A1(n7355), .A2(n4325), .ZN(n8363) );
  INV_X1 U5025 ( .A(n8474), .ZN(n4420) );
  NAND2_X1 U5026 ( .A1(n4419), .A2(n9896), .ZN(n4418) );
  NOR2_X1 U5027 ( .A1(n4873), .A2(n4328), .ZN(n4814) );
  INV_X1 U5028 ( .A(n4581), .ZN(n4580) );
  OAI21_X1 U5029 ( .B1(n5442), .B2(n8522), .A(n5445), .ZN(n4581) );
  AND4_X1 U5030 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n6277)
         );
  AND2_X1 U5031 ( .A1(n8850), .A2(n9155), .ZN(n4483) );
  XNOR2_X1 U5032 ( .A(n9342), .B(n9142), .ZN(n9155) );
  AND4_X1 U5033 ( .A1(n7150), .A2(n7149), .A3(n7148), .A4(n7147), .ZN(n9161)
         );
  INV_X1 U5034 ( .A(n4767), .ZN(n4760) );
  AOI21_X1 U5035 ( .B1(n4767), .B2(n9225), .A(n4766), .ZN(n4765) );
  NOR2_X1 U5036 ( .A1(n9363), .A2(n9207), .ZN(n4766) );
  NOR2_X1 U5037 ( .A1(n4744), .A2(n6867), .ZN(n4743) );
  INV_X1 U5038 ( .A(n6765), .ZN(n4744) );
  AOI21_X1 U5039 ( .B1(n4300), .B2(n4730), .A(n4331), .ZN(n4729) );
  NAND2_X1 U5040 ( .A1(n6421), .A2(n4730), .ZN(n4728) );
  NAND2_X1 U5041 ( .A1(n6426), .A2(n8773), .ZN(n6647) );
  NAND2_X1 U5042 ( .A1(n5285), .A2(n7532), .ZN(n6051) );
  INV_X1 U5043 ( .A(n9105), .ZN(n9319) );
  NAND2_X1 U5044 ( .A1(n7206), .A2(n9617), .ZN(n7212) );
  OR2_X1 U5045 ( .A1(n8869), .A2(n8946), .ZN(n9693) );
  XNOR2_X1 U5046 ( .A(n7535), .B(n7534), .ZN(n8676) );
  OR2_X1 U5047 ( .A1(n4864), .A2(n4933), .ZN(n4442) );
  NOR2_X1 U5048 ( .A1(n4926), .A2(n4435), .ZN(n9005) );
  NAND2_X1 U5049 ( .A1(n9558), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4435) );
  NAND2_X1 U5050 ( .A1(n7652), .A2(n7671), .ZN(n4610) );
  NAND2_X1 U5051 ( .A1(n7655), .A2(n8156), .ZN(n4608) );
  INV_X1 U5052 ( .A(n7659), .ZN(n4604) );
  INV_X1 U5053 ( .A(n7693), .ZN(n4672) );
  OR2_X1 U5054 ( .A1(n8344), .A2(n8353), .ZN(n7649) );
  AND2_X1 U5055 ( .A1(n8866), .A2(n7204), .ZN(n4381) );
  NOR2_X1 U5056 ( .A1(n9373), .A2(n9378), .ZN(n4451) );
  AND2_X1 U5057 ( .A1(n4499), .A2(n4820), .ZN(n4498) );
  NAND2_X1 U5058 ( .A1(n4502), .A2(n4500), .ZN(n4499) );
  INV_X1 U5059 ( .A(n4504), .ZN(n4500) );
  INV_X1 U5060 ( .A(n4502), .ZN(n4501) );
  NAND2_X1 U5061 ( .A1(n5048), .A2(n5047), .ZN(n5072) );
  NAND2_X1 U5062 ( .A1(n4586), .A2(n7842), .ZN(n4585) );
  AND2_X1 U5063 ( .A1(n8405), .A2(n7540), .ZN(n7682) );
  AND2_X1 U5064 ( .A1(n8410), .A2(n8058), .ZN(n7678) );
  INV_X1 U5065 ( .A(n7928), .ZN(n8036) );
  NOR2_X1 U5066 ( .A1(n8447), .A2(n8440), .ZN(n4412) );
  AND2_X1 U5067 ( .A1(n7649), .A2(n7384), .ZN(n8028) );
  NAND2_X1 U5068 ( .A1(n6983), .A2(n6982), .ZN(n7018) );
  NOR2_X1 U5069 ( .A1(n4683), .A2(n7614), .ZN(n4682) );
  INV_X1 U5070 ( .A(n4685), .ZN(n4683) );
  NAND2_X1 U5071 ( .A1(n8495), .A2(n6932), .ZN(n4685) );
  AND2_X1 U5072 ( .A1(n6837), .A2(n7711), .ZN(n4809) );
  OR2_X1 U5073 ( .A1(n6836), .A2(n6862), .ZN(n7612) );
  OR2_X1 U5074 ( .A1(n7882), .A2(n6803), .ZN(n7606) );
  INV_X1 U5075 ( .A(n4789), .ZN(n8331) );
  OAI21_X1 U5076 ( .B1(n8348), .B2(n4791), .A(n4790), .ZN(n4789) );
  NAND2_X1 U5077 ( .A1(n8467), .A2(n8027), .ZN(n4790) );
  NOR2_X1 U5078 ( .A1(n8467), .A2(n8027), .ZN(n4791) );
  AND2_X1 U5079 ( .A1(n4987), .A2(n4774), .ZN(n4773) );
  INV_X1 U5080 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4774) );
  INV_X1 U5081 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4775) );
  INV_X1 U5082 ( .A(n6741), .ZN(n4721) );
  INV_X1 U5083 ( .A(n6692), .ZN(n4717) );
  INV_X1 U5084 ( .A(n7224), .ZN(n4722) );
  XNOR2_X1 U5085 ( .A(n5291), .B(n5653), .ZN(n5294) );
  NAND2_X1 U5086 ( .A1(n7250), .A2(n7249), .ZN(n7256) );
  NOR2_X1 U5087 ( .A1(n7281), .A2(n8634), .ZN(n4712) );
  NAND2_X1 U5088 ( .A1(n7204), .A2(n4489), .ZN(n8914) );
  NOR3_X1 U5089 ( .A1(n9117), .A2(n4492), .A3(n9139), .ZN(n4489) );
  INV_X1 U5090 ( .A(n7363), .ZN(n5103) );
  INV_X1 U5091 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4833) );
  OR2_X1 U5092 ( .A1(n9325), .A2(n9115), .ZN(n8870) );
  OR2_X1 U5093 ( .A1(n9357), .A2(n9216), .ZN(n8844) );
  INV_X1 U5094 ( .A(n4464), .ZN(n4462) );
  INV_X1 U5095 ( .A(n4479), .ZN(n4478) );
  XNOR2_X1 U5096 ( .A(n8970), .B(n9683), .ZN(n8889) );
  NAND2_X1 U5097 ( .A1(n6121), .A2(n5923), .ZN(n5886) );
  AND2_X1 U5098 ( .A1(n8702), .A2(n9654), .ZN(n5381) );
  INV_X1 U5099 ( .A(n9176), .ZN(n9173) );
  AND2_X1 U5100 ( .A1(n9192), .A2(n9197), .ZN(n9186) );
  NAND2_X1 U5101 ( .A1(n9287), .A2(n8809), .ZN(n9272) );
  NAND2_X1 U5102 ( .A1(n5212), .A2(n9638), .ZN(n8869) );
  AOI21_X1 U5103 ( .B1(n4539), .B2(n6900), .A(n4538), .ZN(n4537) );
  INV_X1 U5104 ( .A(n6909), .ZN(n4538) );
  NOR2_X1 U5105 ( .A1(n6910), .A2(n4540), .ZN(n4539) );
  INV_X1 U5106 ( .A(n6899), .ZN(n4540) );
  AND2_X1 U5107 ( .A1(n6272), .A2(n6257), .ZN(n6258) );
  NAND2_X1 U5108 ( .A1(n4510), .A2(n4509), .ZN(n6042) );
  AOI21_X1 U5109 ( .B1(n4299), .B2(n4511), .A(n4364), .ZN(n4509) );
  AOI21_X1 U5110 ( .B1(n5686), .B2(n4515), .A(n4514), .ZN(n4513) );
  INV_X1 U5111 ( .A(n5622), .ZN(n4515) );
  INV_X1 U5112 ( .A(n5688), .ZN(n4514) );
  NAND2_X1 U5113 ( .A1(n5622), .A2(n5621), .ZN(n5631) );
  AOI21_X1 U5114 ( .B1(n4506), .B2(n4504), .A(n4503), .ZN(n4502) );
  INV_X1 U5115 ( .A(n5261), .ZN(n4503) );
  NAND2_X1 U5116 ( .A1(n5179), .A2(SI_11_), .ZN(n5180) );
  NAND2_X1 U5117 ( .A1(n5261), .A2(n5185), .ZN(n5262) );
  INV_X1 U5118 ( .A(n5177), .ZN(n4506) );
  NAND2_X1 U5119 ( .A1(n5140), .A2(n5139), .ZN(n5181) );
  INV_X1 U5120 ( .A(n5040), .ZN(n5041) );
  NAND2_X1 U5121 ( .A1(n5216), .A2(n4611), .ZN(n4973) );
  AND2_X1 U5122 ( .A1(n6926), .A2(n6860), .ZN(n4600) );
  AND2_X1 U5123 ( .A1(n6929), .A2(n4321), .ZN(n4598) );
  NAND2_X1 U5124 ( .A1(n7869), .A2(n4302), .ZN(n7820) );
  INV_X1 U5125 ( .A(n7768), .ZN(n4588) );
  OR2_X1 U5126 ( .A1(n7388), .A2(n7864), .ZN(n7402) );
  NOR2_X1 U5127 ( .A1(n4818), .A2(n4572), .ZN(n4571) );
  INV_X1 U5128 ( .A(n7890), .ZN(n4572) );
  NAND2_X1 U5129 ( .A1(n4574), .A2(n4570), .ZN(n4569) );
  NAND2_X1 U5130 ( .A1(n7760), .A2(n4575), .ZN(n4570) );
  AOI22_X1 U5131 ( .A1(n7877), .A2(n7878), .B1(n6796), .B2(n6795), .ZN(n6800)
         );
  OAI21_X1 U5132 ( .B1(n6861), .B2(n4597), .A(n4595), .ZN(n7031) );
  INV_X1 U5133 ( .A(n4598), .ZN(n4597) );
  AOI21_X1 U5134 ( .B1(n4598), .B2(n4596), .A(n6995), .ZN(n4595) );
  INV_X1 U5135 ( .A(n4600), .ZN(n4596) );
  OR2_X1 U5136 ( .A1(n7420), .A2(n7824), .ZN(n7428) );
  INV_X1 U5137 ( .A(n6373), .ZN(n4550) );
  INV_X1 U5138 ( .A(n4555), .ZN(n4551) );
  INV_X1 U5139 ( .A(n4553), .ZN(n4552) );
  NAND2_X1 U5140 ( .A1(n4592), .A2(n4591), .ZN(n4589) );
  OR2_X1 U5141 ( .A1(n4279), .A2(n7907), .ZN(n5826) );
  NOR2_X1 U5142 ( .A1(n9439), .A2(n4644), .ZN(n9438) );
  NAND2_X1 U5143 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n4644) );
  NOR2_X1 U5144 ( .A1(n9438), .A2(n4643), .ZN(n9452) );
  NOR2_X1 U5145 ( .A1(n5314), .A2(n6265), .ZN(n4643) );
  OR2_X1 U5146 ( .A1(n9452), .A2(n9451), .ZN(n4642) );
  AOI21_X1 U5147 ( .B1(n5365), .B2(P2_REG1_REG_3__SCAN_IN), .A(n5354), .ZN(
        n5318) );
  AOI21_X1 U5148 ( .B1(n4651), .B2(n4653), .A(n4315), .ZN(n4649) );
  AND2_X1 U5149 ( .A1(n5078), .A2(n4544), .ZN(n5272) );
  NOR2_X1 U5150 ( .A1(n5189), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n4544) );
  INV_X1 U5151 ( .A(n9498), .ZN(n8016) );
  AOI21_X1 U5152 ( .B1(n8119), .B2(n4397), .A(n4395), .ZN(n4394) );
  NAND2_X1 U5153 ( .A1(n4396), .A2(n8076), .ZN(n4395) );
  NAND2_X1 U5154 ( .A1(n4397), .A2(n4291), .ZN(n4396) );
  XNOR2_X1 U5155 ( .A(n8420), .B(n8057), .ZN(n8076) );
  NAND2_X1 U5156 ( .A1(n8086), .A2(n8036), .ZN(n4788) );
  AND2_X1 U5157 ( .A1(n8103), .A2(n8102), .ZN(n8106) );
  NAND2_X1 U5158 ( .A1(n7696), .A2(n7695), .ZN(n8088) );
  AOI21_X1 U5159 ( .B1(n4803), .B2(n8130), .A(n4805), .ZN(n4801) );
  INV_X1 U5160 ( .A(n4803), .ZN(n4802) );
  OR2_X1 U5161 ( .A1(n8139), .A2(n8034), .ZN(n4816) );
  NOR2_X1 U5162 ( .A1(n8120), .A2(n4804), .ZN(n4803) );
  INV_X1 U5163 ( .A(n4816), .ZN(n4804) );
  NAND2_X1 U5164 ( .A1(n8155), .A2(n4817), .ZN(n8129) );
  NAND2_X1 U5165 ( .A1(n8350), .A2(n7645), .ZN(n4674) );
  OR2_X1 U5166 ( .A1(n8350), .A2(n8351), .ZN(n4680) );
  NAND2_X1 U5167 ( .A1(n8365), .A2(n4792), .ZN(n8348) );
  OR2_X1 U5168 ( .A1(n8474), .A2(n8026), .ZN(n4792) );
  OR2_X1 U5169 ( .A1(n7348), .A2(n7714), .ZN(n4686) );
  AND2_X1 U5170 ( .A1(n4686), .A2(n4685), .ZN(n6826) );
  NAND2_X1 U5171 ( .A1(n6815), .A2(n7612), .ZN(n7348) );
  NOR2_X1 U5172 ( .A1(n4418), .A2(n6836), .ZN(n4416) );
  NAND2_X1 U5173 ( .A1(n6447), .A2(n4665), .ZN(n4664) );
  NOR2_X1 U5174 ( .A1(n9773), .A2(n4666), .ZN(n4665) );
  INV_X1 U5175 ( .A(n7592), .ZN(n4666) );
  NAND2_X1 U5176 ( .A1(n6476), .A2(n7711), .ZN(n6556) );
  INV_X1 U5177 ( .A(n6336), .ZN(n4798) );
  NOR2_X1 U5178 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  NAND2_X1 U5179 ( .A1(n4391), .A2(n4390), .ZN(n4393) );
  AND2_X1 U5180 ( .A1(n4822), .A2(n7574), .ZN(n4390) );
  INV_X1 U5181 ( .A(n8371), .ZN(n9776) );
  AND2_X1 U5182 ( .A1(n7543), .A2(n5542), .ZN(n8371) );
  NAND2_X1 U5183 ( .A1(n7452), .A2(n7451), .ZN(n8426) );
  AND2_X1 U5184 ( .A1(n5468), .A2(n5469), .ZN(n9500) );
  AND2_X1 U5185 ( .A1(n4824), .A2(n4811), .ZN(n4810) );
  NOR2_X1 U5186 ( .A1(n4872), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U5187 ( .A1(n5062), .A2(n4813), .ZN(n4812) );
  INV_X1 U5188 ( .A(n4872), .ZN(n4405) );
  NAND2_X1 U5189 ( .A1(n5448), .A2(n5447), .ZN(n7549) );
  NAND2_X1 U5190 ( .A1(n4576), .A2(n4580), .ZN(n5448) );
  OR2_X1 U5191 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  NOR2_X1 U5192 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4770) );
  NAND2_X1 U5193 ( .A1(n6544), .A2(n6543), .ZN(n6546) );
  NAND2_X1 U5194 ( .A1(n7472), .A2(n6383), .ZN(n4493) );
  INV_X1 U5195 ( .A(n6073), .ZN(n6071) );
  AND2_X1 U5196 ( .A1(n5230), .A2(n5229), .ZN(n5235) );
  NAND2_X1 U5197 ( .A1(n4703), .A2(n8566), .ZN(n4709) );
  NAND2_X1 U5198 ( .A1(n4708), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U5199 ( .A1(n7286), .A2(n4725), .ZN(n5423) );
  INV_X1 U5200 ( .A(n6121), .ZN(n4725) );
  AND4_X1 U5201 ( .A1(n7140), .A2(n7139), .A3(n7138), .A4(n7137), .ZN(n8957)
         );
  AND4_X1 U5202 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n6403)
         );
  NOR2_X1 U5203 ( .A1(n9020), .A2(n4314), .ZN(n9570) );
  NOR2_X1 U5204 ( .A1(n9570), .A2(n9569), .ZN(n9568) );
  INV_X1 U5205 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4693) );
  AND2_X1 U5206 ( .A1(n9122), .A2(n4450), .ZN(n4449) );
  NOR2_X1 U5207 ( .A1(n9325), .A2(n9337), .ZN(n4450) );
  INV_X1 U5208 ( .A(n9148), .ZN(n4447) );
  NAND2_X1 U5209 ( .A1(n8689), .A2(n8688), .ZN(n9108) );
  NAND2_X1 U5210 ( .A1(n8865), .A2(n8864), .ZN(n9117) );
  AND2_X1 U5211 ( .A1(n9173), .A2(n9186), .ZN(n9171) );
  NAND2_X1 U5212 ( .A1(n9153), .A2(n9171), .ZN(n9148) );
  AOI21_X1 U5213 ( .B1(n4313), .B2(n4759), .A(n4757), .ZN(n4756) );
  NAND2_X1 U5214 ( .A1(n8850), .A2(n8848), .ZN(n9167) );
  AND4_X1 U5215 ( .A1(n7130), .A2(n7129), .A3(n7128), .A4(n7127), .ZN(n9201)
         );
  AOI21_X1 U5216 ( .B1(n9214), .B2(n9213), .A(n7201), .ZN(n9204) );
  NOR2_X1 U5217 ( .A1(n9357), .A2(n9217), .ZN(n9197) );
  NOR2_X1 U5218 ( .A1(n4769), .A2(n7109), .ZN(n4767) );
  AND2_X1 U5219 ( .A1(n8836), .A2(n8692), .ZN(n9213) );
  NAND2_X1 U5220 ( .A1(n4465), .A2(n4466), .ZN(n4464) );
  NAND2_X1 U5221 ( .A1(n4305), .A2(n4466), .ZN(n4463) );
  AND2_X1 U5222 ( .A1(n8830), .A2(n8691), .ZN(n9225) );
  NAND2_X1 U5223 ( .A1(n4294), .A2(n7094), .ZN(n4749) );
  OR2_X1 U5224 ( .A1(n9254), .A2(n9253), .ZN(n4467) );
  AND2_X1 U5225 ( .A1(n9384), .A2(n8960), .ZN(n7094) );
  NOR2_X1 U5226 ( .A1(n9273), .A2(n4753), .ZN(n4752) );
  AND4_X1 U5227 ( .A1(n6886), .A2(n6885), .A3(n6884), .A4(n6883), .ZN(n9290)
         );
  NAND2_X1 U5228 ( .A1(n6876), .A2(n6875), .ZN(n7197) );
  NAND2_X1 U5229 ( .A1(n4737), .A2(n4736), .ZN(n9315) );
  AOI21_X1 U5230 ( .B1(n4739), .B2(n4741), .A(n4334), .ZN(n4736) );
  AOI21_X1 U5231 ( .B1(n4743), .B2(n6766), .A(n4336), .ZN(n4742) );
  AND2_X1 U5232 ( .A1(n6587), .A2(n4729), .ZN(n4727) );
  NOR2_X1 U5233 ( .A1(n4481), .A2(n4480), .ZN(n4479) );
  NAND2_X1 U5234 ( .A1(n6287), .A2(n8718), .ZN(n8922) );
  OAI21_X1 U5235 ( .B1(n6206), .B2(n4734), .A(n4732), .ZN(n6279) );
  INV_X1 U5236 ( .A(n4733), .ZN(n4732) );
  INV_X1 U5237 ( .A(n5846), .ZN(n7085) );
  NAND2_X1 U5238 ( .A1(n6206), .A2(n4735), .ZN(n6276) );
  AND4_X1 U5239 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n6274)
         );
  NOR2_X1 U5240 ( .A1(n5922), .A2(n5923), .ZN(n6115) );
  AND2_X1 U5241 ( .A1(n5387), .A2(n8949), .ZN(n9614) );
  INV_X1 U5242 ( .A(n9295), .ZN(n9625) );
  NAND2_X1 U5243 ( .A1(n7142), .A2(n7141), .ZN(n9342) );
  INV_X1 U5244 ( .A(n9249), .ZN(n9373) );
  INV_X1 U5245 ( .A(n8672), .ZN(n9511) );
  INV_X1 U5246 ( .A(n6211), .ZN(n9704) );
  OR2_X1 U5247 ( .A1(n5020), .A2(n7333), .ZN(n9664) );
  XNOR2_X1 U5248 ( .A(n7526), .B(SI_30_), .ZN(n8685) );
  XNOR2_X1 U5249 ( .A(n7187), .B(n7186), .ZN(n7489) );
  NAND2_X1 U5250 ( .A1(n7500), .A2(n7498), .ZN(n7187) );
  XNOR2_X1 U5251 ( .A(n6950), .B(n7178), .ZN(n7472) );
  NAND2_X1 U5252 ( .A1(n7503), .A2(n7184), .ZN(n6950) );
  OAI21_X1 U5253 ( .B1(n6901), .B2(n6900), .A(n6899), .ZN(n6911) );
  NAND2_X1 U5254 ( .A1(n4520), .A2(n4521), .ZN(n6761) );
  AOI21_X1 U5255 ( .B1(n4523), .B2(n4529), .A(n4522), .ZN(n4521) );
  INV_X1 U5256 ( .A(n6631), .ZN(n4522) );
  AND2_X2 U5257 ( .A1(n4860), .A2(n4861), .ZN(n8917) );
  XNOR2_X1 U5258 ( .A(n6626), .B(n6623), .ZN(n7398) );
  NAND2_X1 U5259 ( .A1(n6273), .A2(n6272), .ZN(n6626) );
  NOR2_X1 U5260 ( .A1(n5466), .A2(n5574), .ZN(n4400) );
  NAND2_X1 U5261 ( .A1(n4324), .A2(n4426), .ZN(n4425) );
  NAND2_X1 U5262 ( .A1(n7010), .A2(n7009), .ZN(n8477) );
  NOR2_X1 U5263 ( .A1(n5729), .A2(n5728), .ZN(n5816) );
  OR2_X1 U5264 ( .A1(n6015), .A2(n5556), .ZN(n5557) );
  NAND2_X1 U5265 ( .A1(n7730), .A2(n4376), .ZN(n4403) );
  AND2_X1 U5266 ( .A1(n7732), .A2(n4617), .ZN(n4404) );
  INV_X1 U5267 ( .A(n5314), .ZN(n9443) );
  AND2_X1 U5268 ( .A1(n4642), .A2(n4641), .ZN(n5362) );
  NAND2_X1 U5269 ( .A1(n9455), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4641) );
  OAI22_X1 U5270 ( .A1(n8005), .A2(n9449), .B1(n9753), .B2(n8004), .ZN(n4658)
         );
  NAND2_X1 U5271 ( .A1(n8002), .A2(n4661), .ZN(n4660) );
  INV_X1 U5272 ( .A(n4662), .ZN(n4661) );
  OAI21_X1 U5273 ( .B1(n8003), .B2(n9753), .A(n9751), .ZN(n4662) );
  NAND2_X1 U5274 ( .A1(n5720), .A2(n5404), .ZN(n4694) );
  OAI22_X1 U5275 ( .A1(n5817), .A2(n6015), .B1(n5466), .B2(n5819), .ZN(n4631)
         );
  CLKBUF_X1 U5276 ( .A(n7549), .Z(n8375) );
  NAND2_X1 U5277 ( .A1(n7310), .A2(n7311), .ZN(n7312) );
  INV_X1 U5278 ( .A(n9192), .ZN(n9352) );
  AND4_X1 U5279 ( .A1(n6410), .A2(n6409), .A3(n6408), .A4(n6407), .ZN(n6679)
         );
  NAND2_X1 U5280 ( .A1(n4303), .A2(n9188), .ZN(n4519) );
  OAI21_X1 U5281 ( .B1(n4318), .B2(n8946), .A(n4517), .ZN(n4516) );
  NAND2_X1 U5282 ( .A1(n8947), .A2(n8948), .ZN(n4517) );
  INV_X1 U5283 ( .A(n9201), .ZN(n9166) );
  OAI21_X1 U5284 ( .B1(n9005), .B2(n9000), .A(n4927), .ZN(n9003) );
  CLKBUF_X1 U5285 ( .A(n4852), .Z(n4938) );
  XNOR2_X1 U5286 ( .A(n9042), .B(n9048), .ZN(n4945) );
  AOI21_X1 U5287 ( .B1(n9096), .B2(n9587), .A(n9579), .ZN(n4438) );
  NAND2_X1 U5288 ( .A1(n8677), .A2(n4819), .ZN(n9105) );
  NAND2_X1 U5289 ( .A1(n8676), .A2(n6383), .ZN(n8677) );
  INV_X1 U5290 ( .A(n9342), .ZN(n9153) );
  NAND2_X1 U5291 ( .A1(n9327), .A2(n9326), .ZN(n9328) );
  INV_X1 U5292 ( .A(n9324), .ZN(n9327) );
  INV_X1 U5293 ( .A(n4470), .ZN(n4469) );
  NAND2_X1 U5294 ( .A1(n4864), .A2(n4865), .ZN(n4444) );
  AND2_X1 U5295 ( .A1(n7612), .A2(n7690), .ZN(n4629) );
  NOR2_X1 U5296 ( .A1(n4627), .A2(n7690), .ZN(n4626) );
  INV_X1 U5297 ( .A(n7609), .ZN(n4627) );
  NAND2_X1 U5298 ( .A1(n8130), .A2(n7658), .ZN(n4606) );
  OAI21_X1 U5299 ( .B1(n4605), .B2(n4604), .A(n7671), .ZN(n4603) );
  INV_X1 U5300 ( .A(n7836), .ZN(n4568) );
  NAND2_X1 U5301 ( .A1(n7675), .A2(n7690), .ZN(n4620) );
  NOR2_X1 U5302 ( .A1(n4563), .A2(n4568), .ZN(n4562) );
  INV_X1 U5303 ( .A(n4571), .ZN(n4563) );
  OR2_X1 U5304 ( .A1(n4569), .A2(n4568), .ZN(n4566) );
  INV_X1 U5305 ( .A(n4670), .ZN(n4669) );
  OAI21_X1 U5306 ( .B1(n7676), .B2(n4671), .A(n7516), .ZN(n4670) );
  NAND2_X1 U5307 ( .A1(n7497), .A2(n4672), .ZN(n4671) );
  NAND2_X1 U5308 ( .A1(n4669), .A2(n4673), .ZN(n4668) );
  NAND2_X1 U5309 ( .A1(n7694), .A2(n7497), .ZN(n4673) );
  OR2_X1 U5310 ( .A1(n8016), .A2(n7539), .ZN(n7683) );
  INV_X1 U5311 ( .A(n4678), .ZN(n4676) );
  INV_X1 U5312 ( .A(n7276), .ZN(n4711) );
  OR2_X1 U5313 ( .A1(n9530), .A2(n6687), .ZN(n8781) );
  NOR3_X1 U5314 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .A3(
        P1_IR_REG_14__SCAN_IN), .ZN(n4840) );
  INV_X1 U5315 ( .A(n4539), .ZN(n4535) );
  NOR2_X1 U5316 ( .A1(n4536), .A2(n4532), .ZN(n4531) );
  INV_X1 U5317 ( .A(n6762), .ZN(n4532) );
  INV_X1 U5318 ( .A(n4537), .ZN(n4536) );
  INV_X1 U5319 ( .A(n6272), .ZN(n4528) );
  INV_X1 U5320 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4692) );
  AND2_X1 U5321 ( .A1(n7687), .A2(n7685), .ZN(n7680) );
  NAND2_X1 U5322 ( .A1(n4636), .A2(n4635), .ZN(n4634) );
  NAND2_X1 U5323 ( .A1(n7985), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4635) );
  INV_X1 U5324 ( .A(n7979), .ZN(n4636) );
  NAND2_X1 U5325 ( .A1(n4634), .A2(n7995), .ZN(n4633) );
  OR2_X1 U5326 ( .A1(n8435), .A2(n8035), .ZN(n7665) );
  NOR2_X1 U5327 ( .A1(n8435), .A2(n8132), .ZN(n4805) );
  NOR2_X1 U5328 ( .A1(n4422), .A2(n8477), .ZN(n4421) );
  INV_X1 U5329 ( .A(n4423), .ZN(n4422) );
  OR2_X1 U5330 ( .A1(n8482), .A2(n8387), .ZN(n7630) );
  NOR2_X1 U5331 ( .A1(n8482), .A2(n8488), .ZN(n4423) );
  OR2_X1 U5332 ( .A1(n6342), .A2(n6341), .ZN(n6458) );
  OAI211_X1 U5333 ( .C1(n6336), .C2(n4794), .A(n4793), .B(n6472), .ZN(n9761)
         );
  NAND3_X1 U5334 ( .A1(n6093), .A2(n4797), .A3(n6092), .ZN(n4794) );
  NAND2_X1 U5335 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5734) );
  NAND2_X1 U5336 ( .A1(n7940), .A2(n9850), .ZN(n7698) );
  NAND2_X1 U5337 ( .A1(n8166), .A2(n4408), .ZN(n8100) );
  NOR2_X1 U5338 ( .A1(n4410), .A2(n8432), .ZN(n4408) );
  AOI21_X1 U5339 ( .B1(n8350), .B2(n4677), .A(n4406), .ZN(n8172) );
  AND2_X1 U5340 ( .A1(n4679), .A2(n7645), .ZN(n4677) );
  NAND2_X1 U5341 ( .A1(n4675), .A2(n7653), .ZN(n4406) );
  NAND2_X1 U5342 ( .A1(n4679), .A2(n4676), .ZN(n4675) );
  OR2_X1 U5343 ( .A1(n5993), .A2(n5998), .ZN(n6105) );
  AND3_X1 U5344 ( .A1(n9850), .A2(n6266), .A3(n9843), .ZN(n6524) );
  NAND2_X1 U5345 ( .A1(n4579), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U5346 ( .A1(n5953), .A2(n5442), .ZN(n4579) );
  INV_X1 U5347 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5188) );
  INV_X1 U5348 ( .A(n8565), .ZN(n4710) );
  INV_X1 U5349 ( .A(n8621), .ZN(n4708) );
  INV_X1 U5350 ( .A(n8566), .ZN(n4706) );
  INV_X1 U5351 ( .A(n8860), .ZN(n8743) );
  NAND2_X1 U5352 ( .A1(n4493), .A2(n7173), .ZN(n8864) );
  NAND2_X1 U5353 ( .A1(n9332), .A2(n9136), .ZN(n8865) );
  NAND2_X1 U5354 ( .A1(n4491), .A2(n4490), .ZN(n8860) );
  NOR2_X1 U5355 ( .A1(n9352), .A2(n9166), .ZN(n4757) );
  INV_X1 U5356 ( .A(n4742), .ZN(n4741) );
  NAND2_X1 U5357 ( .A1(n9511), .A2(n4456), .ZN(n4455) );
  NOR2_X1 U5358 ( .A1(n6721), .A2(n8208), .ZN(n6775) );
  NOR2_X1 U5359 ( .A1(n8696), .A2(n9523), .ZN(n4456) );
  INV_X1 U5360 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6289) );
  NOR2_X1 U5361 ( .A1(n6290), .A2(n6289), .ZN(n6405) );
  INV_X1 U5362 ( .A(n6275), .ZN(n4734) );
  NAND2_X1 U5363 ( .A1(n5663), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U5364 ( .A1(n8969), .A2(n5901), .ZN(n8754) );
  NAND2_X1 U5365 ( .A1(n9279), .A2(n4451), .ZN(n9243) );
  NAND2_X1 U5366 ( .A1(n9279), .A2(n9264), .ZN(n9257) );
  NAND2_X1 U5367 ( .A1(n7182), .A2(n7181), .ZN(n7500) );
  NAND2_X1 U5368 ( .A1(n7182), .A2(n7180), .ZN(n7503) );
  NAND2_X1 U5369 ( .A1(n6939), .A2(n6938), .ZN(n7182) );
  INV_X1 U5370 ( .A(n6639), .ZN(n4524) );
  NAND2_X1 U5371 ( .A1(n5686), .A2(n4512), .ZN(n4511) );
  INV_X1 U5372 ( .A(n5631), .ZN(n4512) );
  NAND2_X1 U5373 ( .A1(n5619), .A2(n5618), .ZN(n5622) );
  XNOR2_X1 U5374 ( .A(n5615), .B(SI_14_), .ZN(n5612) );
  AOI21_X1 U5375 ( .B1(n4498), .B2(n4501), .A(n4495), .ZN(n4494) );
  INV_X1 U5376 ( .A(n5276), .ZN(n4495) );
  AND2_X1 U5377 ( .A1(n5139), .A2(n5092), .ZN(n4826) );
  AND2_X1 U5378 ( .A1(n5085), .A2(n5077), .ZN(n4828) );
  NAND2_X1 U5379 ( .A1(n5072), .A2(n5050), .ZN(n5070) );
  NAND2_X1 U5380 ( .A1(n5032), .A2(n5031), .ZN(n5042) );
  OAI21_X1 U5381 ( .B1(n4968), .B2(n4508), .A(n4507), .ZN(n5008) );
  AOI21_X1 U5382 ( .B1(n7891), .B2(n7890), .A(n4573), .ZN(n7830) );
  AND2_X1 U5383 ( .A1(n7781), .A2(n7780), .ZN(n7808) );
  NAND2_X1 U5384 ( .A1(n7532), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4426) );
  XNOR2_X1 U5385 ( .A(n5554), .B(n6266), .ZN(n5546) );
  INV_X1 U5386 ( .A(n7931), .ZN(n6932) );
  NAND2_X1 U5387 ( .A1(n7401), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7411) );
  INV_X1 U5388 ( .A(n7402), .ZN(n7401) );
  NAND2_X1 U5389 ( .A1(n7871), .A2(n7870), .ZN(n7869) );
  INV_X1 U5390 ( .A(n5728), .ZN(n4593) );
  NAND2_X1 U5391 ( .A1(n5814), .A2(n6005), .ZN(n4594) );
  NAND2_X1 U5392 ( .A1(n4586), .A2(n7842), .ZN(n4587) );
  AND2_X1 U5393 ( .A1(n5590), .A2(n9804), .ZN(n5587) );
  INV_X1 U5394 ( .A(n4278), .ZN(n7490) );
  OR2_X1 U5395 ( .A1(n4279), .A2(n5995), .ZN(n5738) );
  OAI21_X1 U5396 ( .B1(n9443), .B2(P2_REG2_REG_1__SCAN_IN), .A(n5326), .ZN(
        n9439) );
  AOI21_X1 U5397 ( .B1(n9455), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9446), .ZN(
        n5353) );
  OR2_X1 U5398 ( .A1(n5360), .A2(n4653), .ZN(n4652) );
  AOI21_X1 U5399 ( .B1(n5378), .B2(P2_REG1_REG_5__SCAN_IN), .A(n5369), .ZN(
        n5340) );
  OR2_X1 U5400 ( .A1(n5340), .A2(n5339), .ZN(n5396) );
  OR2_X1 U5401 ( .A1(n5973), .A2(n4358), .ZN(n4640) );
  NAND2_X1 U5402 ( .A1(n4640), .A2(n4639), .ZN(n4638) );
  INV_X1 U5403 ( .A(n5974), .ZN(n4639) );
  AOI21_X1 U5404 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6449), .A(n6309), .ZN(
        n6311) );
  AOI21_X1 U5405 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n6849), .A(n6843), .ZN(
        n6846) );
  NOR2_X1 U5406 ( .A1(n6848), .A2(n4368), .ZN(n6852) );
  NAND2_X1 U5407 ( .A1(n6852), .A2(n6851), .ZN(n6953) );
  NAND2_X1 U5408 ( .A1(n6953), .A2(n4655), .ZN(n7952) );
  NAND2_X1 U5409 ( .A1(n6854), .A2(n6833), .ZN(n4655) );
  NOR2_X1 U5410 ( .A1(n7944), .A2(n7945), .ZN(n7948) );
  NAND2_X1 U5411 ( .A1(n7948), .A2(n7947), .ZN(n7963) );
  OAI21_X1 U5412 ( .B1(n4634), .B2(n7995), .A(n4633), .ZN(n7980) );
  NOR2_X1 U5413 ( .A1(n8045), .A2(n8016), .ZN(n8015) );
  AOI21_X1 U5414 ( .B1(n4782), .B2(n4780), .A(n8053), .ZN(n4779) );
  INV_X1 U5415 ( .A(n4784), .ZN(n4780) );
  NAND2_X1 U5416 ( .A1(n8074), .A2(n4787), .ZN(n4786) );
  NOR2_X1 U5417 ( .A1(n8076), .A2(n4785), .ZN(n4784) );
  INV_X1 U5418 ( .A(n8088), .ZN(n4785) );
  NOR2_X1 U5419 ( .A1(n8100), .A2(n8426), .ZN(n8091) );
  NAND2_X1 U5420 ( .A1(n7427), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7441) );
  NAND2_X1 U5421 ( .A1(n8166), .A2(n4412), .ZN(n8134) );
  OR2_X1 U5422 ( .A1(n8447), .A2(n8032), .ZN(n8128) );
  NAND2_X1 U5423 ( .A1(n8166), .A2(n8153), .ZN(n8147) );
  INV_X1 U5424 ( .A(n8033), .ZN(n8156) );
  AND2_X1 U5425 ( .A1(n8457), .A2(n8174), .ZN(n8029) );
  OR2_X1 U5426 ( .A1(n8317), .A2(n8457), .ZN(n8315) );
  NAND2_X1 U5427 ( .A1(n7375), .A2(n7374), .ZN(n7388) );
  OR2_X1 U5428 ( .A1(n7018), .A2(n7042), .ZN(n7378) );
  NOR2_X1 U5429 ( .A1(n8363), .A2(n8467), .ZN(n8354) );
  NAND2_X1 U5430 ( .A1(n7627), .A2(n7638), .ZN(n8368) );
  NAND2_X1 U5431 ( .A1(n7355), .A2(n4421), .ZN(n8395) );
  AND2_X1 U5432 ( .A1(n8024), .A2(n7697), .ZN(n8388) );
  AOI21_X1 U5433 ( .B1(n7715), .B2(n4682), .A(n4333), .ZN(n4684) );
  NAND2_X1 U5434 ( .A1(n7355), .A2(n4423), .ZN(n8393) );
  NAND2_X1 U5435 ( .A1(n6819), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6981) );
  NAND2_X1 U5436 ( .A1(n6456), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6566) );
  INV_X1 U5437 ( .A(n6458), .ZN(n6456) );
  INV_X1 U5438 ( .A(n6837), .ZN(n4807) );
  OAI21_X1 U5439 ( .B1(n4389), .B2(n4337), .A(n7610), .ZN(n6562) );
  INV_X1 U5440 ( .A(n4664), .ZN(n4389) );
  INV_X1 U5441 ( .A(n7599), .ZN(n4663) );
  NAND2_X1 U5442 ( .A1(n4281), .A2(n4388), .ZN(n6815) );
  NOR2_X1 U5443 ( .A1(n6356), .A2(n4417), .ZN(n9763) );
  INV_X1 U5444 ( .A(n4419), .ZN(n4417) );
  NOR2_X1 U5445 ( .A1(n6356), .A2(n6471), .ZN(n9765) );
  NAND2_X1 U5446 ( .A1(n6447), .A2(n7592), .ZN(n9774) );
  AND2_X1 U5447 ( .A1(n7599), .A2(n7595), .ZN(n9777) );
  NAND2_X1 U5448 ( .A1(n6137), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6342) );
  INV_X1 U5449 ( .A(n6138), .ZN(n6137) );
  OR2_X1 U5450 ( .A1(n6029), .A2(n6028), .ZN(n6138) );
  NOR2_X1 U5451 ( .A1(n6105), .A2(n7904), .ZN(n6189) );
  NAND2_X1 U5452 ( .A1(n4391), .A2(n7574), .ZN(n6097) );
  NAND2_X1 U5453 ( .A1(n5980), .A2(n5979), .ZN(n6090) );
  OR2_X1 U5454 ( .A1(n5985), .A2(n5984), .ZN(n6103) );
  NAND2_X1 U5455 ( .A1(n7557), .A2(n7698), .ZN(n6527) );
  OR2_X1 U5456 ( .A1(n5786), .A2(n9843), .ZN(n5467) );
  AND2_X1 U5457 ( .A1(n5502), .A2(n5496), .ZN(n9803) );
  INV_X1 U5458 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5116) );
  AND2_X1 U5459 ( .A1(n5437), .A2(n5439), .ZN(n4601) );
  NAND2_X1 U5460 ( .A1(n5078), .A2(n5093), .ZN(n4545) );
  NOR2_X1 U5461 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4543) );
  NOR2_X1 U5462 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4542) );
  NOR2_X1 U5463 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4541) );
  NOR2_X1 U5464 ( .A1(n5775), .A2(n5774), .ZN(n5856) );
  OAI21_X1 U5465 ( .B1(n6695), .B2(n4720), .A(n4715), .ZN(n8538) );
  AND2_X1 U5466 ( .A1(n4716), .A2(n4346), .ZN(n4715) );
  NAND2_X1 U5467 ( .A1(n4719), .A2(n4717), .ZN(n4716) );
  INV_X1 U5468 ( .A(n7295), .ZN(n8556) );
  NAND2_X1 U5469 ( .A1(n5856), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6077) );
  INV_X1 U5470 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6076) );
  OR2_X1 U5471 ( .A1(n6077), .A2(n6076), .ZN(n6290) );
  INV_X1 U5472 ( .A(n8594), .ZN(n4714) );
  INV_X1 U5473 ( .A(n5512), .ZN(n4701) );
  AND2_X1 U5474 ( .A1(n4696), .A2(n6397), .ZN(n4695) );
  NAND2_X1 U5475 ( .A1(n6400), .A2(n6401), .ZN(n6544) );
  OR3_X1 U5476 ( .A1(n6605), .A2(n6603), .A3(n6604), .ZN(n6721) );
  NOR2_X1 U5477 ( .A1(n7103), .A2(n8635), .ZN(n7113) );
  CLKBUF_X1 U5478 ( .A(n6673), .Z(n6545) );
  AND2_X1 U5479 ( .A1(n5525), .A2(n9665), .ZN(n5879) );
  AND2_X1 U5480 ( .A1(n7301), .A2(n7300), .ZN(n7302) );
  INV_X1 U5481 ( .A(n7319), .ZN(n4726) );
  AND2_X1 U5482 ( .A1(n8918), .A2(n8934), .ZN(n8941) );
  NOR2_X1 U5483 ( .A1(n8914), .A2(n8913), .ZN(n8915) );
  INV_X1 U5484 ( .A(n8938), .ZN(n8877) );
  OR2_X1 U5485 ( .A1(n4280), .A2(n8999), .ZN(n5415) );
  AOI21_X1 U5486 ( .B1(n4953), .B2(P1_REG1_REG_2__SCAN_IN), .A(n4952), .ZN(
        n9430) );
  NAND2_X1 U5487 ( .A1(n5159), .A2(n5152), .ZN(n5151) );
  NAND2_X1 U5488 ( .A1(n5242), .A2(n5241), .ZN(n5240) );
  NAND2_X1 U5489 ( .A1(n5240), .A2(n4386), .ZN(n9031) );
  OR2_X1 U5490 ( .A1(n6385), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4386) );
  AOI21_X1 U5491 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6385), .A(n5245), .ZN(
        n9034) );
  NAND2_X1 U5492 ( .A1(n9584), .A2(n9585), .ZN(n9583) );
  OR2_X1 U5493 ( .A1(n4902), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n4899) );
  NAND2_X1 U5494 ( .A1(n9581), .A2(n9582), .ZN(n9580) );
  NAND2_X1 U5495 ( .A1(n9583), .A2(n4387), .ZN(n5701) );
  OR2_X1 U5496 ( .A1(n9578), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4387) );
  NOR2_X1 U5497 ( .A1(n5705), .A2(n4430), .ZN(n5937) );
  AND2_X1 U5498 ( .A1(n6590), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4430) );
  INV_X1 U5499 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4830) );
  AOI21_X1 U5500 ( .B1(n9077), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9073), .ZN(
        n9074) );
  INV_X1 U5501 ( .A(n4449), .ZN(n4448) );
  NOR2_X1 U5502 ( .A1(n9131), .A2(n9332), .ZN(n9121) );
  NAND2_X1 U5503 ( .A1(n8859), .A2(n8860), .ZN(n9139) );
  OR2_X1 U5504 ( .A1(n9148), .A2(n9337), .ZN(n9131) );
  AOI22_X1 U5505 ( .A1(n9146), .A2(n7151), .B1(n9142), .B2(n9342), .ZN(n9129)
         );
  NAND2_X1 U5506 ( .A1(n5957), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7145) );
  INV_X1 U5507 ( .A(n7135), .ZN(n5957) );
  INV_X1 U5508 ( .A(n7114), .ZN(n7126) );
  NAND2_X1 U5509 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n7126), .ZN(n7135) );
  NAND2_X1 U5510 ( .A1(n9279), .A2(n4329), .ZN(n9217) );
  AOI21_X1 U5511 ( .B1(n4459), .B2(n9225), .A(n7200), .ZN(n4458) );
  OR2_X1 U5512 ( .A1(n7055), .A2(n5252), .ZN(n7103) );
  NAND2_X1 U5513 ( .A1(n7091), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7065) );
  NOR2_X1 U5514 ( .A1(n4292), .A2(n9390), .ZN(n9294) );
  AND2_X1 U5515 ( .A1(n9294), .A2(n9278), .ZN(n9279) );
  OR2_X1 U5516 ( .A1(n9390), .A2(n9304), .ZN(n4754) );
  AND2_X1 U5517 ( .A1(n8816), .A2(n8751), .ZN(n9273) );
  NOR2_X1 U5518 ( .A1(n7070), .A2(n7069), .ZN(n7089) );
  AND2_X1 U5519 ( .A1(n7078), .A2(n7077), .ZN(n7243) );
  INV_X1 U5520 ( .A(n4472), .ZN(n4471) );
  OAI21_X1 U5521 ( .B1(n6875), .B2(n4473), .A(n8811), .ZN(n4472) );
  OR2_X1 U5522 ( .A1(n7198), .A2(n4474), .ZN(n4473) );
  INV_X1 U5523 ( .A(n8907), .ZN(n9286) );
  AOI21_X1 U5524 ( .B1(n9315), .B2(n8906), .A(n7083), .ZN(n9285) );
  NAND2_X1 U5525 ( .A1(n6775), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6881) );
  OR2_X1 U5526 ( .A1(n6881), .A2(n6880), .ZN(n7070) );
  NOR2_X1 U5527 ( .A1(n6732), .A2(n4454), .ZN(n6891) );
  INV_X1 U5528 ( .A(n4456), .ZN(n4454) );
  NOR2_X1 U5529 ( .A1(n6732), .A2(n9523), .ZN(n6784) );
  OR2_X1 U5530 ( .A1(n6653), .A2(n9530), .ZN(n6732) );
  NAND2_X1 U5531 ( .A1(n6427), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6605) );
  NOR2_X1 U5532 ( .A1(n9607), .A2(n6582), .ZN(n6654) );
  NAND2_X1 U5533 ( .A1(n4477), .A2(n4476), .ZN(n4475) );
  NAND2_X1 U5534 ( .A1(n8777), .A2(n4478), .ZN(n4477) );
  NAND2_X1 U5535 ( .A1(n6208), .A2(n4297), .ZN(n9606) );
  NAND2_X1 U5536 ( .A1(n6208), .A2(n4296), .ZN(n9624) );
  OAI21_X1 U5537 ( .B1(n6215), .B2(n8713), .A(n8710), .ZN(n6286) );
  AND2_X1 U5538 ( .A1(n6208), .A2(n9704), .ZN(n9626) );
  AND2_X1 U5539 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5663) );
  NAND2_X1 U5540 ( .A1(n8711), .A2(n8754), .ZN(n8890) );
  INV_X1 U5541 ( .A(n5885), .ZN(n8888) );
  OR2_X1 U5542 ( .A1(n6051), .A2(n5556), .ZN(n5420) );
  INV_X1 U5543 ( .A(n5382), .ZN(n9634) );
  NAND2_X1 U5544 ( .A1(n5382), .A2(n8701), .ZN(n5922) );
  NAND2_X1 U5545 ( .A1(n7112), .A2(n7111), .ZN(n9357) );
  INV_X1 U5546 ( .A(n9689), .ZN(n9723) );
  XNOR2_X1 U5547 ( .A(n7182), .B(n7180), .ZN(n7462) );
  NAND2_X1 U5548 ( .A1(n4533), .A2(n4537), .ZN(n6917) );
  NAND2_X1 U5549 ( .A1(n6901), .A2(n4539), .ZN(n4533) );
  NAND2_X1 U5550 ( .A1(n4525), .A2(n4526), .ZN(n6640) );
  OR2_X1 U5551 ( .A1(n6259), .A2(n4529), .ZN(n4525) );
  CLKBUF_X1 U5552 ( .A(n4942), .Z(n5641) );
  NAND2_X1 U5553 ( .A1(n4497), .A2(n4502), .ZN(n5275) );
  OAI21_X1 U5554 ( .B1(n5181), .B2(n4506), .A(n5180), .ZN(n5263) );
  OR3_X1 U5555 ( .A1(n4904), .A2(P1_IR_REG_8__SCAN_IN), .A3(
        P1_IR_REG_9__SCAN_IN), .ZN(n4902) );
  XNOR2_X1 U5556 ( .A(n5008), .B(n8293), .ZN(n5010) );
  INV_X1 U5557 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4916) );
  NAND2_X1 U5558 ( .A1(n4385), .A2(n4994), .ZN(n4999) );
  NAND2_X1 U5559 ( .A1(n4975), .A2(n4974), .ZN(n4982) );
  XNOR2_X1 U5560 ( .A(n4973), .B(n4970), .ZN(n4972) );
  NAND2_X1 U5561 ( .A1(n4599), .A2(n4598), .ZN(n6996) );
  AND2_X1 U5562 ( .A1(n4599), .A2(n4321), .ZN(n6928) );
  NAND2_X1 U5563 ( .A1(n6861), .A2(n4600), .ZN(n4599) );
  NAND2_X1 U5564 ( .A1(n7419), .A2(n7418), .ZN(n8440) );
  NAND2_X1 U5565 ( .A1(n4547), .A2(n4546), .ZN(n6793) );
  NAND2_X1 U5566 ( .A1(n7475), .A2(n7474), .ZN(n8415) );
  OAI21_X1 U5567 ( .B1(n6132), .B2(n6131), .A(n4559), .ZN(n6370) );
  NOR2_X1 U5568 ( .A1(n5604), .A2(n5605), .ZN(n5603) );
  NAND2_X1 U5569 ( .A1(n7891), .A2(n4571), .ZN(n4564) );
  NAND2_X1 U5570 ( .A1(n7400), .A2(n7399), .ZN(n8452) );
  OR2_X1 U5571 ( .A1(n7029), .A2(n7035), .ZN(n7037) );
  OAI21_X1 U5572 ( .B1(n6132), .B2(n4552), .A(n4549), .ZN(n6485) );
  NAND2_X1 U5573 ( .A1(n4548), .A2(n4553), .ZN(n6374) );
  NAND2_X1 U5574 ( .A1(n6132), .A2(n4555), .ZN(n4548) );
  AND2_X1 U5575 ( .A1(n6861), .A2(n6860), .ZN(n6927) );
  AND2_X1 U5576 ( .A1(n5593), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7885) );
  NAND4_X1 U5577 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(n7936)
         );
  NAND2_X1 U5578 ( .A1(n5450), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5455) );
  XNOR2_X1 U5579 ( .A(n9443), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9436) );
  INV_X1 U5580 ( .A(n4642), .ZN(n9450) );
  XNOR2_X1 U5581 ( .A(n4980), .B(P2_IR_REG_3__SCAN_IN), .ZN(n5365) );
  AND2_X1 U5582 ( .A1(n4652), .A2(n4651), .ZN(n5344) );
  NAND2_X1 U5583 ( .A1(n4648), .A2(n4650), .ZN(n4647) );
  INV_X1 U5584 ( .A(n4649), .ZN(n4648) );
  NAND2_X1 U5585 ( .A1(n5360), .A2(n4651), .ZN(n4646) );
  INV_X1 U5586 ( .A(n4638), .ZN(n6176) );
  INV_X1 U5587 ( .A(n4640), .ZN(n5975) );
  NOR2_X1 U5588 ( .A1(n6179), .A2(n6178), .ZN(n6304) );
  AND2_X1 U5589 ( .A1(n4638), .A2(n4637), .ZN(n6179) );
  NAND2_X1 U5590 ( .A1(n6332), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4637) );
  AND2_X1 U5591 ( .A1(n6512), .A2(n6511), .ZN(n6848) );
  XNOR2_X1 U5592 ( .A(n7952), .B(n4654), .ZN(n6954) );
  INV_X1 U5593 ( .A(n7953), .ZN(n4654) );
  NAND2_X1 U5594 ( .A1(n7538), .A2(n7537), .ZN(n8405) );
  XNOR2_X1 U5595 ( .A(n8015), .B(n4407), .ZN(n8407) );
  INV_X1 U5596 ( .A(n8405), .ZN(n4407) );
  AND2_X1 U5597 ( .A1(n7513), .A2(n7512), .ZN(n9498) );
  AOI21_X1 U5598 ( .B1(n7489), .B2(n6133), .A(n7488), .ZN(n8410) );
  AOI21_X1 U5599 ( .B1(n8062), .B2(n9776), .A(n8061), .ZN(n8418) );
  NAND2_X1 U5600 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  OAI21_X1 U5601 ( .B1(n8119), .B2(n4291), .A(n4397), .ZN(n8077) );
  INV_X1 U5602 ( .A(n8076), .ZN(n4382) );
  INV_X1 U5603 ( .A(n4788), .ZN(n4781) );
  NOR2_X1 U5604 ( .A1(n8106), .A2(n7663), .ZN(n8087) );
  NAND2_X1 U5605 ( .A1(n8442), .A2(n4816), .ZN(n8113) );
  AND2_X1 U5606 ( .A1(n8442), .A2(n4803), .ZN(n8112) );
  NAND2_X1 U5607 ( .A1(n8142), .A2(n8141), .ZN(n8442) );
  AND2_X1 U5608 ( .A1(n4680), .A2(n7645), .ZN(n8333) );
  NAND2_X1 U5609 ( .A1(n7372), .A2(n7371), .ZN(n8344) );
  NAND2_X1 U5610 ( .A1(n7041), .A2(n7040), .ZN(n8474) );
  NAND2_X1 U5611 ( .A1(n4686), .A2(n4293), .ZN(n6978) );
  NAND2_X1 U5612 ( .A1(n4415), .A2(n4414), .ZN(n6574) );
  INV_X1 U5613 ( .A(n4418), .ZN(n4414) );
  NAND2_X1 U5614 ( .A1(n6556), .A2(n4316), .ZN(n6838) );
  NAND2_X1 U5615 ( .A1(n4664), .A2(n7599), .ZN(n6561) );
  AND2_X1 U5616 ( .A1(n4796), .A2(n4795), .ZN(n6473) );
  AND2_X1 U5617 ( .A1(n4393), .A2(n4298), .ZN(n6185) );
  INV_X1 U5618 ( .A(n5798), .ZN(n9796) );
  OR2_X1 U5619 ( .A1(n5598), .A2(n5588), .ZN(n9792) );
  INV_X1 U5620 ( .A(n9795), .ZN(n8380) );
  INV_X1 U5621 ( .A(n8014), .ZN(n9767) );
  NAND2_X1 U5622 ( .A1(n5064), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U5623 ( .A1(n4578), .A2(n4577), .ZN(n5444) );
  AOI21_X1 U5624 ( .B1(n4580), .B2(n8522), .A(n8522), .ZN(n4577) );
  AND2_X1 U5625 ( .A1(n5438), .A2(n5437), .ZN(n5628) );
  AND2_X1 U5626 ( .A1(n4771), .A2(n4770), .ZN(n4772) );
  INV_X1 U5627 ( .A(n4771), .ZN(n5004) );
  XNOR2_X1 U5628 ( .A(n4988), .B(n4987), .ZN(n5559) );
  NAND2_X1 U5629 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4976) );
  OAI22_X1 U5630 ( .A1(n6068), .A2(n4724), .B1(n6066), .B2(n4723), .ZN(n6073)
         );
  INV_X1 U5631 ( .A(n6067), .ZN(n4723) );
  NOR2_X1 U5632 ( .A1(n6067), .A2(n6069), .ZN(n4724) );
  NAND2_X1 U5633 ( .A1(n8538), .A2(n8537), .ZN(n8541) );
  NOR2_X1 U5634 ( .A1(n8530), .A2(n7315), .ZN(n7316) );
  NAND2_X1 U5635 ( .A1(n6320), .A2(n4295), .ZN(n6399) );
  NAND2_X1 U5636 ( .A1(n6320), .A2(n6319), .ZN(n4698) );
  NAND2_X1 U5637 ( .A1(n8662), .A2(n8658), .ZN(n8593) );
  INV_X1 U5638 ( .A(n5658), .ZN(n5659) );
  OR2_X1 U5639 ( .A1(n5222), .A2(n8949), .ZN(n8664) );
  AND2_X1 U5640 ( .A1(n5301), .A2(n8949), .ZN(n8666) );
  NAND2_X1 U5641 ( .A1(n7261), .A2(n4709), .ZN(n8620) );
  NAND2_X1 U5642 ( .A1(n4713), .A2(n7280), .ZN(n8631) );
  OR2_X1 U5643 ( .A1(n4713), .A2(n7280), .ZN(n8632) );
  AND2_X1 U5644 ( .A1(n5432), .A2(n9689), .ZN(n8671) );
  AND4_X1 U5645 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(n9115)
         );
  NAND2_X1 U5646 ( .A1(n5255), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5427) );
  OR2_X1 U5647 ( .A1(n5300), .A2(n5223), .ZN(n5224) );
  OR2_X1 U5648 ( .A1(n4280), .A2(n5100), .ZN(n5109) );
  NAND2_X1 U5649 ( .A1(n9003), .A2(n4319), .ZN(n9426) );
  NAND2_X1 U5650 ( .A1(n9426), .A2(n9425), .ZN(n9424) );
  NOR2_X1 U5651 ( .A1(n5128), .A2(n5127), .ZN(n5126) );
  NOR2_X1 U5652 ( .A1(n9568), .A2(n4929), .ZN(n5134) );
  NAND2_X1 U5653 ( .A1(n5134), .A2(n5133), .ZN(n5132) );
  NOR2_X1 U5654 ( .A1(n5247), .A2(n5246), .ZN(n5245) );
  NAND2_X1 U5655 ( .A1(n5151), .A2(n4429), .ZN(n5247) );
  OR2_X1 U5656 ( .A1(n6281), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4429) );
  NOR2_X1 U5657 ( .A1(n5707), .A2(n5706), .ZN(n5705) );
  NAND2_X1 U5658 ( .A1(n9580), .A2(n4431), .ZN(n5707) );
  OR2_X1 U5659 ( .A1(n9578), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4431) );
  NOR2_X1 U5660 ( .A1(n4945), .A2(n8200), .ZN(n9043) );
  NOR2_X1 U5661 ( .A1(n9050), .A2(n9049), .ZN(n9053) );
  NAND2_X1 U5662 ( .A1(n4434), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4433) );
  NAND2_X1 U5663 ( .A1(n9044), .A2(n4434), .ZN(n4432) );
  INV_X1 U5664 ( .A(n9046), .ZN(n4434) );
  NOR2_X1 U5665 ( .A1(n9593), .A2(n4693), .ZN(n4441) );
  INV_X1 U5666 ( .A(n9098), .ZN(n4440) );
  NAND2_X1 U5667 ( .A1(n4447), .A2(n4312), .ZN(n9099) );
  INV_X1 U5668 ( .A(n9108), .ZN(n9322) );
  XNOR2_X1 U5669 ( .A(n7190), .B(n8912), .ZN(n9330) );
  AND2_X1 U5670 ( .A1(n4482), .A2(n8850), .ZN(n9156) );
  AND3_X1 U5671 ( .A1(n9148), .A2(n9147), .A3(n9625), .ZN(n9341) );
  NAND2_X1 U5672 ( .A1(n7133), .A2(n7132), .ZN(n9176) );
  NAND2_X1 U5673 ( .A1(n9180), .A2(n8845), .ZN(n9163) );
  AND2_X1 U5674 ( .A1(n7124), .A2(n7123), .ZN(n9192) );
  NAND2_X1 U5675 ( .A1(n4755), .A2(n4759), .ZN(n9179) );
  OR2_X1 U5676 ( .A1(n9226), .A2(n4761), .ZN(n4755) );
  NAND2_X1 U5677 ( .A1(n4763), .A2(n4765), .ZN(n9196) );
  NAND2_X1 U5678 ( .A1(n9226), .A2(n4767), .ZN(n4763) );
  NAND2_X1 U5679 ( .A1(n4764), .A2(n4768), .ZN(n9212) );
  INV_X1 U5680 ( .A(n4769), .ZN(n4768) );
  OR2_X1 U5681 ( .A1(n9226), .A2(n9225), .ZN(n4764) );
  NAND2_X1 U5682 ( .A1(n4457), .A2(n4463), .ZN(n9228) );
  OR2_X1 U5683 ( .A1(n9254), .A2(n4464), .ZN(n4457) );
  AND2_X1 U5684 ( .A1(n7053), .A2(n7052), .ZN(n9249) );
  AND2_X1 U5685 ( .A1(n4467), .A2(n8818), .ZN(n9240) );
  INV_X1 U5686 ( .A(n7094), .ZN(n4750) );
  NAND2_X1 U5687 ( .A1(n7088), .A2(n7087), .ZN(n9384) );
  INV_X1 U5688 ( .A(n7243), .ZN(n9390) );
  NAND2_X1 U5689 ( .A1(n7197), .A2(n8805), .ZN(n9302) );
  NAND2_X1 U5690 ( .A1(n4738), .A2(n4742), .ZN(n7079) );
  NAND2_X1 U5691 ( .A1(n6767), .A2(n4743), .ZN(n4738) );
  NAND2_X1 U5692 ( .A1(n6871), .A2(n6870), .ZN(n8672) );
  NAND2_X1 U5693 ( .A1(n4728), .A2(n4729), .ZN(n6644) );
  NAND2_X1 U5694 ( .A1(n8922), .A2(n4479), .ZN(n9595) );
  NAND2_X1 U5695 ( .A1(n6276), .A2(n6275), .ZN(n9623) );
  INV_X1 U5696 ( .A(n9263), .ZN(n9620) );
  OR2_X1 U5697 ( .A1(n9693), .A2(n5880), .ZN(n9306) );
  AND2_X1 U5698 ( .A1(n9323), .A2(n9693), .ZN(n9659) );
  AND2_X1 U5699 ( .A1(n5022), .A2(n5021), .ZN(n9393) );
  NOR2_X1 U5700 ( .A1(n5523), .A2(P1_U3084), .ZN(n9665) );
  INV_X1 U5701 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5097) );
  AND2_X1 U5702 ( .A1(n4865), .A2(n4863), .ZN(n4488) );
  INV_X1 U5703 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5055) );
  NOR2_X1 U5704 ( .A1(n9490), .A2(n9971), .ZN(n9957) );
  NOR2_X1 U5705 ( .A1(n5816), .A2(n5815), .ZN(n6006) );
  AOI21_X1 U5706 ( .B1(n9755), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8006), .ZN(
        n4656) );
  NAND2_X1 U5707 ( .A1(n4660), .A2(n7370), .ZN(n4659) );
  AOI21_X1 U5708 ( .B1(n4518), .B2(n8946), .A(n4516), .ZN(n8955) );
  NOR2_X1 U5709 ( .A1(n4441), .A2(n4440), .ZN(n4439) );
  NAND2_X1 U5710 ( .A1(n4437), .A2(n9638), .ZN(n4436) );
  NAND2_X1 U5711 ( .A1(n4338), .A2(n4377), .ZN(n9399) );
  INV_X1 U5712 ( .A(n9328), .ZN(n4377) );
  OAI21_X1 U5713 ( .B1(n4338), .B2(n9727), .A(n4468), .ZN(P1_U3520) );
  AOI21_X1 U5714 ( .B1(n9328), .B2(n9729), .A(n4375), .ZN(n4468) );
  AND2_X1 U5715 ( .A1(n7102), .A2(n7101), .ZN(n9222) );
  INV_X1 U5716 ( .A(n9222), .ZN(n9363) );
  OR2_X1 U5717 ( .A1(n7677), .A2(n7678), .ZN(n4290) );
  OR2_X1 U5718 ( .A1(n7461), .A2(n4688), .ZN(n4291) );
  OR3_X1 U5719 ( .A1(n6732), .A2(n9313), .A3(n4455), .ZN(n4292) );
  AND2_X1 U5720 ( .A1(n7715), .A2(n4685), .ZN(n4293) );
  NAND2_X1 U5721 ( .A1(n7277), .A2(n7276), .ZN(n4713) );
  OR2_X1 U5722 ( .A1(n8415), .A2(n8037), .ZN(n7694) );
  OR2_X1 U5723 ( .A1(n9378), .A2(n8959), .ZN(n4294) );
  AND2_X1 U5724 ( .A1(n6322), .A2(n6319), .ZN(n4295) );
  AND2_X1 U5725 ( .A1(n9711), .A2(n9704), .ZN(n4296) );
  AND2_X1 U5726 ( .A1(n4296), .A2(n4446), .ZN(n4297) );
  OR2_X1 U5727 ( .A1(n4307), .A2(n7568), .ZN(n4298) );
  INV_X1 U5728 ( .A(n8766), .ZN(n4480) );
  AND2_X1 U5729 ( .A1(n4513), .A2(n5944), .ZN(n4299) );
  OR2_X1 U5730 ( .A1(n8894), .A2(n4317), .ZN(n4300) );
  INV_X1 U5731 ( .A(n9253), .ZN(n4465) );
  NOR2_X1 U5732 ( .A1(n4712), .A2(n4711), .ZN(n4301) );
  BUF_X1 U5733 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9558) );
  NAND2_X1 U5734 ( .A1(n7368), .A2(n7367), .ZN(n8467) );
  INV_X1 U5735 ( .A(n4783), .ZN(n4782) );
  OAI21_X1 U5736 ( .B1(n8076), .B2(n4788), .A(n4786), .ZN(n4783) );
  NAND2_X1 U5737 ( .A1(n6818), .A2(n6817), .ZN(n8488) );
  AND2_X1 U5738 ( .A1(n7767), .A2(n4588), .ZN(n4302) );
  NOR2_X1 U5739 ( .A1(n8941), .A2(n8937), .ZN(n4303) );
  AND2_X1 U5740 ( .A1(n4451), .A2(n9235), .ZN(n4304) );
  NAND2_X1 U5741 ( .A1(n8817), .A2(n8818), .ZN(n4305) );
  AND2_X1 U5742 ( .A1(n4297), .A2(n4445), .ZN(n4306) );
  AND4_X1 U5743 ( .A1(n7162), .A2(n7161), .A3(n7160), .A4(n7159), .ZN(n7327)
         );
  INV_X1 U5744 ( .A(n7327), .ZN(n4490) );
  NAND2_X1 U5745 ( .A1(n4493), .A2(n7174), .ZN(n9332) );
  AND2_X1 U5746 ( .A1(n6227), .A2(n6094), .ZN(n4307) );
  INV_X2 U5747 ( .A(n5300), .ZN(n5255) );
  INV_X1 U5748 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4813) );
  AND2_X1 U5749 ( .A1(n4674), .A2(n4678), .ZN(n4308) );
  OR2_X1 U5750 ( .A1(n4849), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4309) );
  OR2_X1 U5751 ( .A1(n9192), .A2(n9201), .ZN(n4310) );
  NAND2_X1 U5752 ( .A1(n6004), .A2(n6003), .ZN(n4311) );
  NOR2_X1 U5753 ( .A1(n5544), .A2(n9844), .ZN(n5725) );
  AND2_X1 U5754 ( .A1(n9322), .A2(n4449), .ZN(n4312) );
  XNOR2_X1 U5755 ( .A(n5178), .B(SI_11_), .ZN(n5177) );
  AND2_X1 U5756 ( .A1(n4775), .A2(n9758), .ZN(n4977) );
  AND2_X1 U5757 ( .A1(n4761), .A2(n4310), .ZN(n4313) );
  INV_X1 U5758 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5093) );
  INV_X1 U5759 ( .A(n5459), .ZN(n6266) );
  NAND2_X1 U5760 ( .A1(n4427), .A2(n4424), .ZN(n5459) );
  INV_X1 U5761 ( .A(n8776), .ZN(n4481) );
  AND2_X1 U5762 ( .A1(n9017), .A2(n8220), .ZN(n4314) );
  AND2_X1 U5763 ( .A1(n5721), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4315) );
  AND2_X1 U5764 ( .A1(n7712), .A2(n6555), .ZN(n4316) );
  NAND2_X1 U5765 ( .A1(n7797), .A2(n5118), .ZN(n6985) );
  NOR2_X1 U5766 ( .A1(n9601), .A2(n8966), .ZN(n4317) );
  OR2_X1 U5767 ( .A1(n8947), .A2(n9188), .ZN(n4318) );
  OR2_X1 U5768 ( .A1(n9006), .A2(n8999), .ZN(n4319) );
  NAND2_X1 U5769 ( .A1(n7099), .A2(n7098), .ZN(n9368) );
  NAND2_X1 U5770 ( .A1(n7426), .A2(n7425), .ZN(n8435) );
  INV_X1 U5771 ( .A(n8435), .ZN(n4411) );
  OR3_X1 U5772 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4320) );
  NAND2_X1 U5773 ( .A1(n6925), .A2(n6924), .ZN(n4321) );
  INV_X1 U5774 ( .A(n8850), .ZN(n8842) );
  OR2_X1 U5775 ( .A1(n9176), .A2(n8957), .ZN(n8850) );
  NAND2_X1 U5776 ( .A1(n7410), .A2(n7409), .ZN(n8447) );
  AND2_X1 U5777 ( .A1(n8777), .A2(n8718), .ZN(n4322) );
  NAND4_X1 U5778 ( .A1(n4771), .A2(n4543), .A3(n4542), .A4(n4541), .ZN(n5051)
         );
  NOR2_X1 U5779 ( .A1(n4288), .A2(n5572), .ZN(n4323) );
  OR2_X1 U5780 ( .A1(n5456), .A2(n7532), .ZN(n4324) );
  AND2_X1 U5781 ( .A1(n4421), .A2(n4420), .ZN(n4325) );
  AND2_X1 U5782 ( .A1(n8351), .A2(n7645), .ZN(n4326) );
  NAND2_X1 U5783 ( .A1(n6770), .A2(n6769), .ZN(n8696) );
  INV_X1 U5784 ( .A(n8130), .ZN(n8141) );
  AND2_X1 U5785 ( .A1(n7659), .A2(n8118), .ZN(n8130) );
  INV_X1 U5786 ( .A(n8883), .ZN(n4476) );
  NAND2_X1 U5787 ( .A1(n6972), .A2(n6971), .ZN(n8482) );
  INV_X1 U5788 ( .A(n4605), .ZN(n8120) );
  NAND2_X1 U5789 ( .A1(n7660), .A2(n7665), .ZN(n4605) );
  AND2_X1 U5790 ( .A1(n7676), .A2(n7690), .ZN(n4327) );
  NAND2_X1 U5791 ( .A1(n8166), .A2(n4409), .ZN(n4413) );
  INV_X1 U5792 ( .A(n4818), .ZN(n4574) );
  AND2_X1 U5793 ( .A1(n7063), .A2(n7062), .ZN(n9264) );
  OR2_X1 U5794 ( .A1(n4872), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4328) );
  OR2_X1 U5795 ( .A1(n8432), .A2(n7855), .ZN(n7449) );
  NAND2_X1 U5796 ( .A1(n7189), .A2(n7188), .ZN(n9325) );
  AND2_X1 U5797 ( .A1(n4304), .A2(n9222), .ZN(n4329) );
  OR2_X1 U5798 ( .A1(n8457), .A2(n8335), .ZN(n7653) );
  AND2_X1 U5799 ( .A1(n4695), .A2(n6322), .ZN(n4330) );
  NOR2_X1 U5800 ( .A1(n6582), .A2(n9597), .ZN(n4331) );
  INV_X1 U5801 ( .A(n4575), .ZN(n4573) );
  NAND2_X1 U5802 ( .A1(n7747), .A2(n7748), .ZN(n4575) );
  INV_X1 U5803 ( .A(n4410), .ZN(n4409) );
  NAND2_X1 U5804 ( .A1(n4412), .A2(n4411), .ZN(n4410) );
  NOR2_X1 U5805 ( .A1(n8672), .A2(n9303), .ZN(n4332) );
  NOR2_X1 U5806 ( .A1(n8488), .A2(n7001), .ZN(n4333) );
  NOR2_X1 U5807 ( .A1(n9511), .A2(n8544), .ZN(n4334) );
  NOR2_X1 U5808 ( .A1(n9200), .A2(n9216), .ZN(n4335) );
  NOR2_X1 U5809 ( .A1(n9518), .A2(n8695), .ZN(n4336) );
  INV_X1 U5810 ( .A(n4720), .ZN(n4719) );
  OR2_X1 U5811 ( .A1(n7216), .A2(n4721), .ZN(n4720) );
  OR2_X1 U5812 ( .A1(n6560), .A2(n4663), .ZN(n4337) );
  AND2_X1 U5813 ( .A1(n7212), .A2(n4469), .ZN(n4338) );
  NOR2_X1 U5814 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4339) );
  AND2_X1 U5815 ( .A1(n4759), .A2(n4310), .ZN(n4340) );
  AND2_X1 U5816 ( .A1(n5652), .A2(n5651), .ZN(n4341) );
  OR2_X1 U5817 ( .A1(n9357), .A2(n9183), .ZN(n4342) );
  OR2_X1 U5818 ( .A1(n7763), .A2(n7762), .ZN(n4343) );
  AND2_X1 U5819 ( .A1(n9249), .A2(n8958), .ZN(n8880) );
  INV_X1 U5820 ( .A(n8880), .ZN(n4466) );
  AND2_X1 U5821 ( .A1(n8708), .A2(n8711), .ZN(n4344) );
  AND2_X1 U5822 ( .A1(n4752), .A2(n4294), .ZN(n4345) );
  INV_X1 U5823 ( .A(n9332), .ZN(n9122) );
  INV_X1 U5824 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4933) );
  AND2_X1 U5825 ( .A1(n4722), .A2(n7215), .ZN(n4346) );
  AND2_X1 U5826 ( .A1(n4651), .A2(n4650), .ZN(n4347) );
  AND2_X1 U5827 ( .A1(n9286), .A2(n8812), .ZN(n4348) );
  AND2_X1 U5828 ( .A1(n7525), .A2(n4668), .ZN(n4349) );
  AND2_X1 U5829 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4350) );
  AND2_X1 U5830 ( .A1(n8857), .A2(n9130), .ZN(n4351) );
  AND2_X1 U5831 ( .A1(n4601), .A2(n5440), .ZN(n4352) );
  AND2_X1 U5832 ( .A1(n4298), .A2(n7582), .ZN(n4353) );
  AND2_X1 U5833 ( .A1(n4339), .A2(n4745), .ZN(n4354) );
  AND2_X1 U5834 ( .A1(n4773), .A2(n4775), .ZN(n4355) );
  XNOR2_X1 U5835 ( .A(n5444), .B(n5443), .ZN(n5468) );
  OAI22_X1 U5836 ( .A1(n7745), .A2(n7744), .B1(n7742), .B2(n7743), .ZN(n7891)
         );
  NAND2_X1 U5837 ( .A1(n7153), .A2(n7152), .ZN(n9337) );
  INV_X1 U5838 ( .A(n9337), .ZN(n4491) );
  INV_X1 U5839 ( .A(n8805), .ZN(n4474) );
  INV_X1 U5840 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4508) );
  NAND2_X1 U5841 ( .A1(n5441), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5953) );
  OAI21_X1 U5842 ( .B1(n6767), .B2(n6766), .A(n6765), .ZN(n6868) );
  NAND2_X1 U5843 ( .A1(n6742), .A2(n6741), .ZN(n7217) );
  AND2_X1 U5844 ( .A1(n4751), .A2(n4750), .ZN(n4356) );
  NAND2_X1 U5845 ( .A1(n4564), .A2(n4569), .ZN(n4357) );
  AND2_X1 U5846 ( .A1(n6134), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4358) );
  AND2_X1 U5847 ( .A1(n8634), .A2(n7281), .ZN(n4359) );
  NAND2_X1 U5848 ( .A1(n7464), .A2(n7463), .ZN(n8420) );
  INV_X1 U5849 ( .A(n8420), .ZN(n8074) );
  NAND2_X1 U5850 ( .A1(n8366), .A2(n8368), .ZN(n8365) );
  OR2_X1 U5851 ( .A1(n8465), .A2(n8353), .ZN(n4360) );
  OR2_X1 U5852 ( .A1(n8930), .A2(n8874), .ZN(n4361) );
  NAND2_X1 U5853 ( .A1(n5438), .A2(n4601), .ZN(n5695) );
  NOR2_X1 U5854 ( .A1(n9043), .A2(n9044), .ZN(n4362) );
  NAND2_X1 U5855 ( .A1(n9279), .A2(n4304), .ZN(n4452) );
  NAND2_X1 U5856 ( .A1(n6623), .A2(n6272), .ZN(n4529) );
  AND2_X1 U5857 ( .A1(n4534), .A2(n6916), .ZN(n4363) );
  AND2_X1 U5858 ( .A1(n4526), .A2(n4524), .ZN(n4523) );
  INV_X1 U5859 ( .A(n7843), .ZN(n4586) );
  NAND2_X1 U5860 ( .A1(n7084), .A2(n4752), .ZN(n4751) );
  AND2_X1 U5861 ( .A1(n5946), .A2(SI_17_), .ZN(n4364) );
  AND2_X1 U5862 ( .A1(n6625), .A2(SI_21_), .ZN(n4365) );
  AND2_X1 U5863 ( .A1(n8066), .A2(n8037), .ZN(n4366) );
  OR2_X1 U5864 ( .A1(n7842), .A2(n4586), .ZN(n4367) );
  NAND2_X1 U5865 ( .A1(n5589), .A2(n9792), .ZN(n7903) );
  OR2_X2 U5866 ( .A1(n7549), .A2(n7548), .ZN(n7690) );
  INV_X1 U5867 ( .A(n4279), .ZN(n5731) );
  AND2_X1 U5868 ( .A1(n6849), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4368) );
  NAND2_X1 U5869 ( .A1(n4702), .A2(n5512), .ZN(n5649) );
  OAI21_X1 U5870 ( .B1(n6421), .B2(n4300), .A(n6420), .ZN(n6583) );
  AND2_X1 U5871 ( .A1(n7346), .A2(n7615), .ZN(n6839) );
  NAND2_X1 U5872 ( .A1(n7355), .A2(n6973), .ZN(n4369) );
  INV_X1 U5873 ( .A(n4453), .ZN(n9309) );
  NOR2_X1 U5874 ( .A1(n6732), .A2(n4455), .ZN(n4453) );
  AND2_X1 U5875 ( .A1(n8922), .A2(n8766), .ZN(n4370) );
  INV_X1 U5876 ( .A(n6337), .ZN(n4799) );
  NAND2_X1 U5877 ( .A1(n7612), .A2(n7609), .ZN(n7712) );
  INV_X1 U5878 ( .A(n7712), .ZN(n4388) );
  AND2_X1 U5879 ( .A1(n6206), .A2(n6205), .ZN(n4371) );
  AND2_X1 U5880 ( .A1(n6556), .A2(n6555), .ZN(n4372) );
  INV_X1 U5881 ( .A(n9601), .ZN(n4445) );
  INV_X1 U5882 ( .A(n7939), .ZN(n4401) );
  INV_X1 U5883 ( .A(n6417), .ZN(n4446) );
  NAND4_X1 U5884 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .ZN(n7937)
         );
  INV_X1 U5885 ( .A(n7937), .ZN(n4632) );
  OR2_X1 U5886 ( .A1(n7549), .A2(n6642), .ZN(n5542) );
  AND2_X1 U5887 ( .A1(n4646), .A2(n4649), .ZN(n4373) );
  AND2_X1 U5888 ( .A1(n7546), .A2(n9844), .ZN(n4374) );
  AND2_X1 U5889 ( .A1(n9727), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4375) );
  AND2_X1 U5890 ( .A1(n7547), .A2(n5468), .ZN(n4376) );
  INV_X1 U5891 ( .A(n5545), .ZN(n5458) );
  NOR2_X1 U5892 ( .A1(n9235), .A2(n9242), .ZN(n4769) );
  NAND2_X2 U5893 ( .A1(n6673), .A2(n6672), .ZN(n6695) );
  NOR2_X2 U5894 ( .A1(n9202), .A2(n7202), .ZN(n9182) );
  NAND2_X1 U5895 ( .A1(n9225), .A2(n4462), .ZN(n4461) );
  NAND2_X1 U5896 ( .A1(n4486), .A2(n4483), .ZN(n9154) );
  AOI22_X1 U5897 ( .A1(n9129), .A2(n9139), .B1(n7327), .B2(n4491), .ZN(n9114)
         );
  NOR2_X1 U5898 ( .A1(n9138), .A2(n9139), .ZN(n9137) );
  NAND2_X1 U5899 ( .A1(n4658), .A2(n8375), .ZN(n4657) );
  NAND3_X2 U5900 ( .A1(n4836), .A2(n4915), .A3(n4835), .ZN(n4852) );
  NAND2_X2 U5901 ( .A1(n8661), .A2(n8660), .ZN(n8658) );
  NAND2_X2 U5902 ( .A1(n6071), .A2(n6070), .ZN(n6320) );
  NAND2_X1 U5903 ( .A1(n8648), .A2(n8644), .ZN(n8564) );
  NAND2_X1 U5904 ( .A1(n4378), .A2(n8814), .ZN(n8821) );
  NAND2_X1 U5905 ( .A1(n8813), .A2(n4348), .ZN(n4378) );
  NAND2_X1 U5906 ( .A1(n4379), .A2(n4985), .ZN(n4612) );
  INV_X1 U5907 ( .A(n4981), .ZN(n4379) );
  MUX2_X2 U5908 ( .A(n8853), .B(n8852), .S(n8869), .Z(n8854) );
  NAND2_X1 U5909 ( .A1(n8858), .A2(n4351), .ZN(n8863) );
  MUX2_X2 U5910 ( .A(n8839), .B(n8838), .S(n8869), .Z(n8847) );
  MUX2_X2 U5911 ( .A(n8825), .B(n8824), .S(n8869), .Z(n8833) );
  OAI211_X1 U5912 ( .C1(n8943), .C2(n9188), .A(n4276), .B(n4519), .ZN(n4518)
         );
  OAI22_X4 U5913 ( .A1(n8097), .A2(n8102), .B1(n8122), .B2(n8432), .ZN(n8085)
         );
  OR2_X1 U5914 ( .A1(n7935), .A2(n6222), .ZN(n6226) );
  INV_X1 U5915 ( .A(n4814), .ZN(n5112) );
  NAND2_X1 U5916 ( .A1(n4778), .A2(n4782), .ZN(n8054) );
  NAND2_X1 U5917 ( .A1(n4806), .A2(n4808), .ZN(n7347) );
  NAND2_X1 U5918 ( .A1(n5293), .A2(n5292), .ZN(n5412) );
  AOI22_X2 U5919 ( .A1(n8146), .A2(n8033), .B1(n8153), .B2(n8032), .ZN(n8142)
         );
  OAI21_X2 U5920 ( .B1(n8142), .B2(n4802), .A(n4801), .ZN(n4800) );
  NAND2_X4 U5921 ( .A1(n5231), .A2(n5281), .ZN(n7319) );
  NAND2_X1 U5922 ( .A1(n7347), .A2(n7714), .ZN(n7346) );
  XNOR2_X1 U5923 ( .A(n4383), .B(n4382), .ZN(n8424) );
  AOI21_X1 U5924 ( .B1(n8085), .B2(n8088), .A(n4781), .ZN(n4383) );
  NAND2_X1 U5925 ( .A1(n4718), .A2(n7215), .ZN(n7225) );
  NAND2_X1 U5926 ( .A1(n7613), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U5927 ( .A1(n4621), .A2(n4620), .ZN(n4619) );
  NAND2_X1 U5928 ( .A1(n7662), .A2(n4829), .ZN(n7666) );
  NAND2_X1 U5929 ( .A1(n7691), .A2(n7690), .ZN(n4616) );
  OAI21_X1 U5930 ( .B1(n4607), .B2(n4606), .A(n4603), .ZN(n4602) );
  OAI21_X1 U5931 ( .B1(n7668), .B2(n7690), .A(n7667), .ZN(n4384) );
  AOI21_X1 U5932 ( .B1(n7651), .B2(n7690), .A(n7656), .ZN(n4609) );
  NAND2_X1 U5933 ( .A1(n7608), .A2(n4626), .ZN(n4625) );
  AOI22_X1 U5934 ( .A1(n4384), .A2(n7695), .B1(n7670), .B2(n7690), .ZN(n7674)
         );
  NAND3_X1 U5935 ( .A1(n4612), .A2(n4613), .A3(n4990), .ZN(n4385) );
  MUX2_X1 U5936 ( .A(n7641), .B(n7640), .S(n7671), .Z(n7646) );
  AOI21_X1 U5937 ( .B1(n4610), .B2(n4609), .A(n4608), .ZN(n4607) );
  NAND2_X1 U5938 ( .A1(n4622), .A2(n7693), .ZN(n4621) );
  NAND2_X1 U5939 ( .A1(n4624), .A2(n7617), .ZN(n7619) );
  NAND2_X1 U5940 ( .A1(n4402), .A2(n7733), .ZN(n7740) );
  NAND2_X1 U5941 ( .A1(n4616), .A2(n4615), .ZN(n7730) );
  NAND2_X1 U5942 ( .A1(n4602), .A2(n7660), .ZN(n7662) );
  INV_X1 U5943 ( .A(n4762), .ZN(n4761) );
  OAI21_X1 U5944 ( .B1(n9330), .B2(n9659), .A(n7211), .ZN(n4470) );
  NAND2_X1 U5945 ( .A1(n4758), .A2(n4756), .ZN(n9168) );
  OAI21_X2 U5946 ( .B1(n5614), .B2(n5613), .A(n5617), .ZN(n5632) );
  OAI21_X1 U5947 ( .B1(n9095), .B2(n9094), .A(n4438), .ZN(n4437) );
  OAI211_X1 U5948 ( .C1(n9097), .C2(n9638), .A(n4439), .B(n4436), .ZN(P1_U3260) );
  XNOR2_X2 U5949 ( .A(n4925), .B(n4924), .ZN(n8977) );
  NAND2_X1 U5950 ( .A1(n7338), .A2(n7337), .ZN(n7336) );
  NAND2_X1 U5951 ( .A1(n6742), .A2(n4719), .ZN(n4718) );
  NAND2_X1 U5952 ( .A1(n4393), .A2(n4353), .ZN(n6349) );
  NAND2_X1 U5953 ( .A1(n8119), .A2(n7665), .ZN(n8103) );
  INV_X1 U5954 ( .A(n4394), .ZN(n8075) );
  NAND2_X1 U5955 ( .A1(n7573), .A2(n7566), .ZN(n7700) );
  NAND2_X1 U5956 ( .A1(n4401), .A2(n5798), .ZN(n7566) );
  NOR2_X1 U5957 ( .A1(n4323), .A2(n4400), .ZN(n4399) );
  NAND3_X1 U5958 ( .A1(n7731), .A2(n4404), .A3(n4403), .ZN(n4402) );
  NAND2_X1 U5959 ( .A1(n4824), .A2(n5078), .ZN(n4873) );
  NAND3_X1 U5960 ( .A1(n4824), .A2(n4405), .A3(n5078), .ZN(n5064) );
  INV_X1 U5961 ( .A(n4413), .ZN(n8114) );
  NAND2_X1 U5962 ( .A1(n5466), .A2(n4425), .ZN(n4424) );
  INV_X1 U5963 ( .A(n5466), .ZN(n5720) );
  NAND3_X1 U5964 ( .A1(n8009), .A2(n5310), .A3(n9443), .ZN(n4427) );
  NAND2_X1 U5965 ( .A1(n5466), .A2(n4968), .ZN(n6015) );
  NAND2_X1 U5966 ( .A1(n6524), .A2(n9796), .ZN(n5803) );
  INV_X1 U5967 ( .A(n5803), .ZN(n4428) );
  NAND2_X1 U5968 ( .A1(n4428), .A2(n5801), .ZN(n5993) );
  NAND2_X1 U5969 ( .A1(n6266), .A2(n9843), .ZN(n6525) );
  OAI21_X1 U5970 ( .B1(n4945), .B2(n4433), .A(n4432), .ZN(n9060) );
  XNOR2_X2 U5971 ( .A(n4442), .B(n4865), .ZN(n8991) );
  NAND2_X1 U5972 ( .A1(n4306), .A2(n6208), .ZN(n9607) );
  NOR2_X1 U5973 ( .A1(n9148), .A2(n4448), .ZN(n9107) );
  INV_X1 U5974 ( .A(n4452), .ZN(n9231) );
  AND3_X2 U5975 ( .A1(n5288), .A2(n5286), .A3(n5287), .ZN(n5382) );
  OR2_X1 U5976 ( .A1(n9254), .A2(n4461), .ZN(n4460) );
  INV_X1 U5977 ( .A(n4467), .ZN(n9252) );
  NAND2_X1 U5978 ( .A1(n7212), .A2(n7211), .ZN(n9329) );
  OAI21_X2 U5979 ( .B1(n6876), .B2(n4473), .A(n4471), .ZN(n9287) );
  NAND2_X1 U5980 ( .A1(n9180), .A2(n4484), .ZN(n4486) );
  CLKBUF_X1 U5981 ( .A(n4486), .Z(n4482) );
  INV_X1 U5982 ( .A(n4482), .ZN(n9162) );
  NAND2_X1 U5983 ( .A1(n4487), .A2(n4344), .ZN(n8757) );
  NAND2_X1 U5984 ( .A1(n6118), .A2(n6119), .ZN(n4487) );
  NAND2_X1 U5985 ( .A1(n4864), .A2(n4488), .ZN(n9412) );
  NAND2_X1 U5986 ( .A1(n7290), .A2(n8702), .ZN(n5234) );
  NAND4_X1 U5987 ( .A1(n8911), .A2(n9155), .A3(n8910), .A4(n9181), .ZN(n4492)
         );
  NAND2_X1 U5988 ( .A1(n5181), .A2(n4498), .ZN(n4496) );
  NAND2_X1 U5989 ( .A1(n5181), .A2(n4504), .ZN(n4497) );
  NAND2_X1 U5990 ( .A1(n4968), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U5991 ( .A1(n5632), .A2(n4299), .ZN(n4510) );
  OAI21_X1 U5992 ( .B1(n5632), .B2(n4511), .A(n4513), .ZN(n5947) );
  OAI21_X1 U5993 ( .B1(n5632), .B2(n5631), .A(n5622), .ZN(n5687) );
  NAND2_X1 U5994 ( .A1(n6259), .A2(n4523), .ZN(n4520) );
  NAND2_X1 U5995 ( .A1(n6259), .A2(n6258), .ZN(n6273) );
  NAND2_X1 U5996 ( .A1(n6763), .A2(n6762), .ZN(n6901) );
  NAND2_X1 U5997 ( .A1(n4545), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U5998 ( .A1(n6132), .A2(n4549), .ZN(n4547) );
  AOI21_X1 U5999 ( .B1(n4549), .B2(n4552), .A(n6484), .ZN(n4546) );
  INV_X1 U6000 ( .A(n6130), .ZN(n4561) );
  NAND2_X1 U6001 ( .A1(n7891), .A2(n4562), .ZN(n4567) );
  OR2_X1 U6002 ( .A1(n5953), .A2(n8522), .ZN(n4576) );
  NAND2_X1 U6003 ( .A1(n5953), .A2(n4580), .ZN(n4578) );
  NAND2_X1 U6004 ( .A1(n7775), .A2(n4583), .ZN(n4582) );
  NAND2_X1 U6005 ( .A1(n4584), .A2(n4585), .ZN(n4583) );
  NAND2_X1 U6006 ( .A1(n7774), .A2(n4367), .ZN(n4584) );
  NAND2_X1 U6007 ( .A1(n7775), .A2(n7774), .ZN(n7845) );
  NAND2_X1 U6008 ( .A1(n7869), .A2(n7767), .ZN(n7769) );
  OAI21_X1 U6009 ( .B1(n4592), .B2(n5729), .A(n4591), .ZN(n7899) );
  NAND3_X1 U6010 ( .A1(n4590), .A2(n4589), .A3(n7900), .ZN(n7898) );
  NAND2_X1 U6011 ( .A1(n5729), .A2(n4591), .ZN(n4590) );
  NAND2_X1 U6012 ( .A1(n4594), .A2(n4311), .ZN(n4591) );
  NAND2_X1 U6013 ( .A1(n4593), .A2(n4311), .ZN(n4592) );
  NAND2_X1 U6014 ( .A1(n5438), .A2(n4352), .ZN(n5441) );
  INV_X2 U6015 ( .A(n4986), .ZN(n4968) );
  NAND2_X2 U6016 ( .A1(n4691), .A2(n4690), .ZN(n4986) );
  NAND3_X1 U6017 ( .A1(n4691), .A2(n4350), .A3(n4690), .ZN(n4611) );
  NAND3_X1 U6018 ( .A1(n4985), .A2(n4975), .A3(n4974), .ZN(n4613) );
  NAND2_X1 U6019 ( .A1(n4614), .A2(n4985), .ZN(n4991) );
  NAND2_X1 U6020 ( .A1(n4982), .A2(n4981), .ZN(n4614) );
  NAND2_X1 U6021 ( .A1(n7692), .A2(n7671), .ZN(n4615) );
  NAND3_X1 U6022 ( .A1(n4616), .A2(n4615), .A3(n4374), .ZN(n4617) );
  NAND3_X1 U6023 ( .A1(n4628), .A2(n4625), .A3(n7614), .ZN(n4624) );
  NAND2_X1 U6024 ( .A1(n4632), .A2(n5998), .ZN(n7568) );
  INV_X1 U6025 ( .A(n4631), .ZN(n4630) );
  MUX2_X1 U6026 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n5473), .S(n5559), .Z(n9451)
         );
  NAND2_X1 U6027 ( .A1(n4645), .A2(n4647), .ZN(n5374) );
  NAND2_X1 U6028 ( .A1(n5360), .A2(n4347), .ZN(n4645) );
  INV_X1 U6029 ( .A(n4652), .ZN(n5331) );
  INV_X1 U6030 ( .A(n5375), .ZN(n4650) );
  NAND3_X1 U6031 ( .A1(n4659), .A2(n4657), .A3(n4656), .ZN(P2_U3264) );
  NAND2_X1 U6032 ( .A1(n8172), .A2(n8173), .ZN(n8171) );
  NAND2_X1 U6033 ( .A1(n4667), .A2(n4349), .ZN(n7541) );
  NAND2_X1 U6034 ( .A1(n8056), .A2(n4669), .ZN(n4667) );
  AOI21_X1 U6035 ( .B1(n8056), .B2(n7693), .A(n7676), .ZN(n8039) );
  NOR2_X1 U6036 ( .A1(n8323), .A2(n8322), .ZN(n4679) );
  INV_X1 U6037 ( .A(n4680), .ZN(n8349) );
  NAND2_X1 U6038 ( .A1(n7348), .A2(n4293), .ZN(n4681) );
  NAND2_X1 U6039 ( .A1(n4681), .A2(n4684), .ZN(n6979) );
  INV_X1 U6040 ( .A(n4686), .ZN(n7350) );
  NAND3_X1 U6041 ( .A1(n4966), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4690) );
  NAND3_X1 U6042 ( .A1(n4967), .A2(n4693), .A3(n4692), .ZN(n4691) );
  XNOR2_X1 U6043 ( .A(n5028), .B(n5027), .ZN(n6007) );
  AOI21_X2 U6044 ( .B1(n5014), .B2(n5013), .A(n4825), .ZN(n5028) );
  NAND2_X1 U6045 ( .A1(n4697), .A2(n6323), .ZN(n4696) );
  INV_X1 U6046 ( .A(n6319), .ZN(n4697) );
  NAND2_X1 U6047 ( .A1(n4698), .A2(n6323), .ZN(n6398) );
  NAND3_X1 U6048 ( .A1(n5508), .A2(n5648), .A3(n5507), .ZN(n4699) );
  NAND2_X1 U6049 ( .A1(n5508), .A2(n5507), .ZN(n4702) );
  NAND2_X1 U6050 ( .A1(n4700), .A2(n4699), .ZN(n5657) );
  AOI21_X1 U6051 ( .B1(n4701), .B2(n5648), .A(n4341), .ZN(n4700) );
  NAND4_X1 U6052 ( .A1(n8648), .A2(n8644), .A3(n4710), .A4(n4708), .ZN(n4707)
         );
  NAND3_X1 U6053 ( .A1(n8648), .A2(n8644), .A3(n4710), .ZN(n4703) );
  NAND2_X1 U6054 ( .A1(n7261), .A2(n4704), .ZN(n8624) );
  NAND2_X1 U6055 ( .A1(n4707), .A2(n4705), .ZN(n4704) );
  AOI21_X2 U6056 ( .B1(n7277), .B2(n4301), .A(n4359), .ZN(n8550) );
  OAI21_X2 U6057 ( .B1(n4849), .B2(n4746), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4848) );
  NAND2_X1 U6058 ( .A1(n4728), .A2(n4727), .ZN(n6646) );
  OAI21_X1 U6059 ( .B1(n4735), .B2(n4734), .A(n9622), .ZN(n4733) );
  NAND2_X1 U6060 ( .A1(n6767), .A2(n4739), .ZN(n4737) );
  NAND2_X1 U6061 ( .A1(n4841), .A2(n4821), .ZN(n4849) );
  AND3_X2 U6062 ( .A1(n4841), .A2(n4821), .A3(n4354), .ZN(n4864) );
  NAND2_X1 U6063 ( .A1(n7084), .A2(n4345), .ZN(n4748) );
  NAND2_X1 U6064 ( .A1(n4748), .A2(n4749), .ZN(n7095) );
  NAND2_X1 U6065 ( .A1(n7084), .A2(n4754), .ZN(n9267) );
  INV_X1 U6066 ( .A(n4751), .ZN(n9387) );
  INV_X1 U6067 ( .A(n4754), .ZN(n4753) );
  NAND2_X1 U6068 ( .A1(n9226), .A2(n4340), .ZN(n4758) );
  AND2_X1 U6069 ( .A1(n4772), .A2(n4355), .ZN(n5033) );
  NAND3_X1 U6070 ( .A1(n4773), .A2(n9758), .A3(n4775), .ZN(n5005) );
  NAND2_X1 U6071 ( .A1(n4776), .A2(n4777), .ZN(n8038) );
  NAND2_X1 U6072 ( .A1(n8085), .A2(n4779), .ZN(n4776) );
  NAND2_X1 U6073 ( .A1(n8085), .A2(n4784), .ZN(n4778) );
  INV_X1 U6074 ( .A(n8057), .ZN(n4787) );
  NAND2_X1 U6075 ( .A1(n6093), .A2(n6092), .ZN(n6337) );
  NAND2_X1 U6076 ( .A1(n6340), .A2(n4797), .ZN(n4793) );
  NAND2_X1 U6077 ( .A1(n4799), .A2(n4798), .ZN(n4795) );
  INV_X1 U6078 ( .A(n6340), .ZN(n4796) );
  INV_X1 U6079 ( .A(n7708), .ZN(n4797) );
  INV_X2 U6080 ( .A(n4800), .ZN(n8097) );
  NAND2_X1 U6081 ( .A1(n6476), .A2(n4809), .ZN(n4808) );
  OR2_X1 U6082 ( .A1(n4316), .A2(n4807), .ZN(n4806) );
  AND2_X1 U6083 ( .A1(n5078), .A2(n4810), .ZN(n5115) );
  INV_X1 U6084 ( .A(n5078), .ZN(n5079) );
  NAND2_X4 U6085 ( .A1(n9646), .A2(n5280), .ZN(n9323) );
  AOI21_X2 U6086 ( .B1(n5212), .B2(n5281), .A(n9638), .ZN(n5280) );
  NAND2_X1 U6087 ( .A1(n5450), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5461) );
  INV_X1 U6088 ( .A(n5923), .ZN(n9677) );
  NAND2_X1 U6089 ( .A1(n5468), .A2(n7549), .ZN(n5544) );
  INV_X1 U6090 ( .A(n5468), .ZN(n7729) );
  INV_X1 U6091 ( .A(n5295), .ZN(n5293) );
  XNOR2_X1 U6092 ( .A(n8056), .B(n8055), .ZN(n8062) );
  INV_X1 U6093 ( .A(n5294), .ZN(n5292) );
  NOR2_X1 U6094 ( .A1(n9204), .A2(n9203), .ZN(n9202) );
  AOI21_X2 U6095 ( .B1(n8528), .B2(n7317), .A(n7316), .ZN(n7326) );
  AOI22_X1 U6096 ( .A1(n8582), .A2(n8583), .B1(n7308), .B2(n7307), .ZN(n7338)
         );
  INV_X1 U6097 ( .A(n5102), .ZN(n7796) );
  AND2_X1 U6098 ( .A1(n5385), .A2(n5384), .ZN(n9289) );
  AND4_X1 U6099 ( .A1(n5439), .A2(n5271), .A3(n5187), .A4(n5637), .ZN(n4815)
         );
  AND2_X1 U6100 ( .A1(n8130), .A2(n8128), .ZN(n4817) );
  NOR2_X1 U6101 ( .A1(n7759), .A2(n7758), .ZN(n4818) );
  OR2_X1 U6102 ( .A1(n8687), .A2(n5125), .ZN(n4819) );
  AND2_X1 U6103 ( .A1(n5276), .A2(n5269), .ZN(n4820) );
  AND4_X1 U6104 ( .A1(n4840), .A2(n4839), .A3(n4838), .A4(n4837), .ZN(n4821)
         );
  NOR2_X1 U6105 ( .A1(n6096), .A2(n4307), .ZN(n4822) );
  INV_X1 U6106 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4967) );
  AND2_X1 U6107 ( .A1(n5012), .A2(n5011), .ZN(n4825) );
  INV_X1 U6108 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5002) );
  AND3_X1 U6109 ( .A1(n7068), .A2(n7067), .A3(n7066), .ZN(n9277) );
  AND2_X1 U6110 ( .A1(n8102), .A2(n7665), .ZN(n4827) );
  INV_X1 U6111 ( .A(n8900), .ZN(n6587) );
  INV_X1 U6112 ( .A(n7032), .ZN(n7029) );
  OR2_X1 U6113 ( .A1(n7661), .A2(n7671), .ZN(n4829) );
  INV_X1 U6114 ( .A(n8399), .ZN(n9785) );
  NAND2_X1 U6115 ( .A1(n8870), .A2(n8930), .ZN(n8912) );
  AND2_X1 U6116 ( .A1(n7612), .A2(n7606), .ZN(n7607) );
  NAND2_X1 U6117 ( .A1(n7666), .A2(n4827), .ZN(n7667) );
  AND4_X1 U6118 ( .A1(n5188), .A2(n5634), .A3(n5436), .A4(n5093), .ZN(n4869)
         );
  NAND2_X1 U6119 ( .A1(n7524), .A2(n7523), .ZN(n7525) );
  INV_X1 U6120 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5439) );
  NOR2_X1 U6121 ( .A1(n6090), .A2(n9856), .ZN(n6091) );
  INV_X1 U6122 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5187) );
  AND2_X1 U6123 ( .A1(n8554), .A2(n8556), .ZN(n7298) );
  INV_X1 U6124 ( .A(n8912), .ZN(n7204) );
  INV_X1 U6125 ( .A(n7428), .ZN(n7427) );
  INV_X1 U6126 ( .A(n6981), .ZN(n6983) );
  INV_X1 U6127 ( .A(n7378), .ZN(n7375) );
  INV_X1 U6128 ( .A(n6820), .ZN(n6819) );
  INV_X1 U6129 ( .A(n7449), .ZN(n7663) );
  INV_X1 U6130 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8286) );
  INV_X1 U6131 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5774) );
  OR2_X1 U6132 ( .A1(n7296), .A2(n8609), .ZN(n7301) );
  OR2_X1 U6133 ( .A1(n5425), .A2(n5101), .ZN(n5105) );
  INV_X1 U6134 ( .A(n6713), .ZN(n6600) );
  INV_X1 U6135 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4893) );
  NOR2_X1 U6136 ( .A1(n7029), .A2(n7028), .ZN(n7030) );
  OR2_X1 U6137 ( .A1(n7453), .A2(n7920), .ZN(n7480) );
  OR2_X1 U6138 ( .A1(n7411), .A2(n8299), .ZN(n7420) );
  OR3_X1 U6139 ( .A1(n6566), .A2(n6565), .A3(n6564), .ZN(n6820) );
  OR2_X1 U6140 ( .A1(n6335), .A2(n6339), .ZN(n6336) );
  INV_X1 U6141 ( .A(n5750), .ZN(n5749) );
  OR2_X1 U6142 ( .A1(n6245), .A2(n9873), .ZN(n6356) );
  AND2_X1 U6143 ( .A1(n6405), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U6144 ( .A1(n5295), .A2(n5294), .ZN(n5411) );
  NAND2_X1 U6145 ( .A1(n8702), .A2(n7286), .ZN(n5230) );
  INV_X1 U6146 ( .A(n7280), .ZN(n7281) );
  OR2_X1 U6147 ( .A1(n7065), .A2(n8626), .ZN(n7055) );
  NAND2_X1 U6148 ( .A1(n9325), .A2(n9689), .ZN(n9326) );
  NOR2_X2 U6149 ( .A1(n4852), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n4942) );
  NAND2_X1 U6150 ( .A1(n5183), .A2(n5182), .ZN(n5261) );
  AND2_X1 U6151 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  INV_X1 U6152 ( .A(n7885), .ZN(n7922) );
  AND2_X1 U6153 ( .A1(n7480), .A2(n7454), .ZN(n8092) );
  AOI21_X1 U6154 ( .B1(n5378), .B2(P2_REG2_REG_5__SCAN_IN), .A(n5374), .ZN(
        n5348) );
  AOI21_X1 U6155 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n6016), .A(n5679), .ZN(
        n5682) );
  AOI21_X1 U6156 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6449), .A(n6304), .ZN(
        n6307) );
  AOI21_X1 U6157 ( .B1(n7972), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7971), .ZN(
        n7975) );
  INV_X1 U6158 ( .A(n8132), .ZN(n8035) );
  NAND2_X1 U6159 ( .A1(n7563), .A2(n5749), .ZN(n5804) );
  AND2_X1 U6160 ( .A1(n7654), .A2(n8157), .ZN(n8173) );
  INV_X1 U6161 ( .A(n9900), .ZN(n8489) );
  NAND2_X1 U6162 ( .A1(n7256), .A2(n7257), .ZN(n8643) );
  AND2_X1 U6163 ( .A1(n7089), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7091) );
  OR2_X1 U6164 ( .A1(n8683), .A2(n9736), .ZN(n5536) );
  AND2_X1 U6165 ( .A1(n9313), .A2(n8961), .ZN(n7083) );
  AND2_X1 U6166 ( .A1(n8797), .A2(n8788), .ZN(n8902) );
  AND2_X1 U6167 ( .A1(n9594), .A2(n8776), .ZN(n8894) );
  NAND2_X1 U6168 ( .A1(n8718), .A2(n8766), .ZN(n9622) );
  AND2_X1 U6169 ( .A1(n6762), .A2(n6636), .ZN(n6760) );
  AND2_X1 U6170 ( .A1(n5688), .A2(n5627), .ZN(n5686) );
  INV_X1 U6171 ( .A(n7913), .ZN(n7901) );
  INV_X1 U6172 ( .A(n9751), .ZN(n9456) );
  AND2_X1 U6173 ( .A1(n5329), .A2(n5328), .ZN(n9750) );
  NAND2_X1 U6174 ( .A1(n7653), .A2(n7647), .ZN(n8323) );
  INV_X1 U6175 ( .A(n8022), .ZN(n7717) );
  INV_X1 U6176 ( .A(n8384), .ZN(n9769) );
  INV_X1 U6177 ( .A(n8399), .ZN(n9788) );
  INV_X1 U6178 ( .A(n9500), .ZN(n9902) );
  INV_X1 U6179 ( .A(n9907), .ZN(n8494) );
  AND2_X1 U6180 ( .A1(n5468), .A2(n5449), .ZN(n9892) );
  OR2_X1 U6181 ( .A1(n5606), .A2(n5575), .ZN(n5985) );
  AND2_X1 U6182 ( .A1(n5483), .A2(n5056), .ZN(n9804) );
  AND4_X1 U6183 ( .A1(n7171), .A2(n7170), .A3(n7169), .A4(n7168), .ZN(n9136)
         );
  AND2_X1 U6184 ( .A1(n7061), .A2(n7060), .ZN(n9256) );
  AND4_X1 U6185 ( .A1(n6597), .A2(n6596), .A3(n6595), .A4(n6594), .ZN(n6687)
         );
  OR2_X1 U6186 ( .A1(n5425), .A2(n8997), .ZN(n5416) );
  INV_X1 U6187 ( .A(n9293), .ZN(n9649) );
  INV_X1 U6188 ( .A(n9660), .ZN(n9641) );
  AND2_X1 U6189 ( .A1(n5879), .A2(n5199), .ZN(n9396) );
  XNOR2_X1 U6190 ( .A(n6911), .B(n6910), .ZN(n7436) );
  BUF_X1 U6191 ( .A(n5193), .Z(n5195) );
  XNOR2_X1 U6192 ( .A(n5029), .B(SI_6_), .ZN(n5027) );
  AND2_X1 U6193 ( .A1(n5069), .A2(n5068), .ZN(n9755) );
  INV_X1 U6194 ( .A(n7905), .ZN(n7893) );
  NAND2_X1 U6195 ( .A1(n5587), .A2(n5579), .ZN(n7913) );
  NAND2_X1 U6196 ( .A1(n7470), .A2(n7469), .ZN(n8057) );
  INV_X1 U6197 ( .A(n9750), .ZN(n9449) );
  OR2_X1 U6198 ( .A1(n9793), .A2(n9902), .ZN(n8014) );
  NAND2_X1 U6199 ( .A1(n9785), .A2(n5997), .ZN(n9795) );
  OR2_X1 U6200 ( .A1(n5985), .A2(n5505), .ZN(n9925) );
  OR2_X1 U6201 ( .A1(n5985), .A2(n5599), .ZN(n9908) );
  INV_X1 U6202 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n8288) );
  INV_X1 U6203 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6008) );
  INV_X1 U6204 ( .A(n9690), .ZN(n5901) );
  OR2_X1 U6205 ( .A1(n5237), .A2(n9689), .ZN(n8645) );
  INV_X1 U6206 ( .A(n9161), .ZN(n9142) );
  INV_X1 U6207 ( .A(n9660), .ZN(n9644) );
  INV_X1 U6208 ( .A(n9748), .ZN(n9745) );
  INV_X1 U6209 ( .A(n9729), .ZN(n9727) );
  INV_X1 U6210 ( .A(n9671), .ZN(n9672) );
  INV_X1 U6211 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5082) );
  NOR2_X1 U6212 ( .A1(n9957), .A2(n9956), .ZN(n9955) );
  NOR2_X2 U6213 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4832) );
  NOR2_X2 U6214 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4831) );
  AND4_X2 U6215 ( .A1(n4832), .A2(n4831), .A3(n4830), .A4(n4893), .ZN(n4836)
         );
  AND4_X2 U6216 ( .A1(n8199), .A2(n4911), .A3(n4833), .A4(n4891), .ZN(n4835)
         );
  NOR2_X1 U6217 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4834) );
  NOR2_X2 U6218 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4918) );
  AND2_X2 U6219 ( .A1(n4834), .A2(n4918), .ZN(n4915) );
  INV_X1 U6220 ( .A(n4852), .ZN(n4841) );
  NOR2_X1 U6221 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4839) );
  NOR2_X1 U6222 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4838) );
  NOR2_X1 U6223 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4837) );
  INV_X1 U6224 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U6225 ( .A1(n4848), .A2(n4847), .ZN(n4842) );
  INV_X1 U6226 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4843) );
  XNOR2_X1 U6227 ( .A(n4848), .B(n4847), .ZN(n6907) );
  OR3_X4 U6228 ( .A1(n7333), .A2(n6764), .A3(n6907), .ZN(n5231) );
  NAND2_X1 U6229 ( .A1(n4849), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4850) );
  MUX2_X1 U6230 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4850), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n4851) );
  NAND2_X1 U6231 ( .A1(n4851), .A2(n4309), .ZN(n5015) );
  INV_X1 U6232 ( .A(n5015), .ZN(n6661) );
  NOR2_X1 U6233 ( .A1(n5231), .A2(n6661), .ZN(n4946) );
  INV_X1 U6234 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5640) );
  INV_X1 U6235 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5948) );
  INV_X1 U6236 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5691) );
  INV_X1 U6237 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4853) );
  AND3_X1 U6238 ( .A1(n5948), .A2(n5691), .A3(n4853), .ZN(n4854) );
  AND2_X1 U6239 ( .A1(n5640), .A2(n4854), .ZN(n4855) );
  NAND2_X1 U6240 ( .A1(n4942), .A2(n4855), .ZN(n5196) );
  OAI21_X2 U6241 ( .B1(n5196), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5193) );
  INV_X1 U6242 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6243 ( .A1(n5193), .A2(n5194), .ZN(n4856) );
  NAND2_X1 U6244 ( .A1(n4856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4859) );
  INV_X1 U6245 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U6246 ( .A1(n4859), .A2(n4858), .ZN(n4860) );
  XNOR2_X2 U6247 ( .A(n4857), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8952) );
  OR2_X1 U6248 ( .A1(n4859), .A2(n4858), .ZN(n4861) );
  NAND2_X2 U6249 ( .A1(n8952), .A2(n8917), .ZN(n5219) );
  NAND2_X1 U6250 ( .A1(n5219), .A2(n5231), .ZN(n4862) );
  NAND2_X1 U6251 ( .A1(n4862), .A2(n5015), .ZN(n4960) );
  INV_X1 U6252 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U6253 ( .A1(n4960), .A2(n5846), .ZN(n4866) );
  NAND2_X1 U6254 ( .A1(n4866), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X1 U6255 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4868) );
  NOR2_X1 U6256 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4867) );
  NOR2_X1 U6257 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n4871) );
  NOR2_X1 U6258 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4870) );
  NAND4_X1 U6259 ( .A1(n4871), .A2(n4870), .A3(n4887), .A4(n8286), .ZN(n4872)
         );
  NOR2_X1 U6260 ( .A1(n4873), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6261 ( .A1(n5057), .A2(n8286), .ZN(n4878) );
  INV_X1 U6262 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U6263 ( .A1(n4879), .A2(n4887), .ZN(n4874) );
  NOR2_X1 U6264 ( .A1(n4878), .A2(n4874), .ZN(n4881) );
  INV_X1 U6265 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U6266 ( .A1(n4881), .A2(n4875), .ZN(n4884) );
  NAND2_X1 U6267 ( .A1(n4884), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4876) );
  MUX2_X1 U6268 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4876), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n4877) );
  AND2_X1 U6269 ( .A1(n5064), .A2(n4877), .ZN(n5502) );
  NAND2_X1 U6270 ( .A1(n4878), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U6271 ( .A1(n4888), .A2(n4887), .ZN(n4890) );
  NAND2_X1 U6272 ( .A1(n4890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4880) );
  XNOR2_X1 U6273 ( .A(n4880), .B(n4879), .ZN(n6811) );
  INV_X1 U6274 ( .A(n6811), .ZN(n5499) );
  INV_X1 U6275 ( .A(n4881), .ZN(n4882) );
  NAND2_X1 U6276 ( .A1(n4882), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4883) );
  MUX2_X1 U6277 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4883), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n4885) );
  NAND2_X1 U6278 ( .A1(n4885), .A2(n4884), .ZN(n6906) );
  INV_X1 U6279 ( .A(n6906), .ZN(n4886) );
  NAND3_X1 U6280 ( .A1(n5502), .A2(n5499), .A3(n4886), .ZN(n5483) );
  OR2_X1 U6281 ( .A1(n4888), .A2(n4887), .ZN(n4889) );
  NAND2_X1 U6282 ( .A1(n4890), .A2(n4889), .ZN(n5482) );
  NAND2_X1 U6283 ( .A1(n5482), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9840) );
  NOR2_X2 U6284 ( .A1(n5483), .A2(n9840), .ZN(P2_U3966) );
  NAND2_X1 U6285 ( .A1(n4915), .A2(n4916), .ZN(n4910) );
  NAND2_X1 U6286 ( .A1(n4911), .A2(n4891), .ZN(n4892) );
  NOR2_X1 U6287 ( .A1(n4910), .A2(n4892), .ZN(n4934) );
  NAND2_X1 U6288 ( .A1(n4934), .A2(n4893), .ZN(n4904) );
  OAI21_X1 U6289 ( .B1(n4899), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4897) );
  INV_X1 U6290 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U6291 ( .A1(n4897), .A2(n4894), .ZN(n4895) );
  NAND2_X1 U6292 ( .A1(n4895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4896) );
  XNOR2_X1 U6293 ( .A(n4896), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6707) );
  XNOR2_X1 U6294 ( .A(n4897), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U6295 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6590), .ZN(n4898) );
  OAI21_X1 U6296 ( .B1(n6590), .B2(P1_REG2_REG_12__SCAN_IN), .A(n4898), .ZN(
        n5706) );
  NAND2_X1 U6297 ( .A1(n4899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4900) );
  XNOR2_X1 U6298 ( .A(n4900), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9578) );
  NOR2_X1 U6299 ( .A1(n9578), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4901) );
  AOI21_X1 U6300 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9578), .A(n4901), .ZN(
        n9582) );
  NAND2_X1 U6301 ( .A1(n4902), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4903) );
  XNOR2_X1 U6302 ( .A(n4903), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U6303 ( .A1(n4904), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4909) );
  INV_X1 U6304 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U6305 ( .A1(n4909), .A2(n4905), .ZN(n4906) );
  NAND2_X1 U6306 ( .A1(n4906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4907) );
  XNOR2_X1 U6307 ( .A(n4907), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U6308 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6385), .ZN(n4908) );
  OAI21_X1 U6309 ( .B1(n6385), .B2(P1_REG2_REG_9__SCAN_IN), .A(n4908), .ZN(
        n5246) );
  XNOR2_X1 U6310 ( .A(n4909), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U6311 ( .A1(n4910), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U6312 ( .A1(n4914), .A2(n4911), .ZN(n4912) );
  NAND2_X1 U6313 ( .A1(n4912), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4913) );
  XNOR2_X1 U6314 ( .A(n4913), .B(P1_IR_REG_6__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U6315 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n5847), .ZN(n4932) );
  XNOR2_X1 U6316 ( .A(n4914), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9563) );
  NOR2_X1 U6317 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9563), .ZN(n4929) );
  INV_X1 U6318 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n8220) );
  OR2_X1 U6319 ( .A1(n4915), .A2(n4933), .ZN(n4917) );
  XNOR2_X1 U6320 ( .A(n4917), .B(n4916), .ZN(n9017) );
  OR2_X1 U6321 ( .A1(n4918), .A2(n4933), .ZN(n4923) );
  INV_X1 U6322 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U6323 ( .A1(n4923), .A2(n4922), .ZN(n4921) );
  NAND2_X1 U6324 ( .A1(n4921), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4920) );
  INV_X1 U6325 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4919) );
  XNOR2_X1 U6326 ( .A(n4920), .B(n4919), .ZN(n9421) );
  INV_X1 U6327 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5424) );
  INV_X1 U6328 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8999) );
  INV_X1 U6329 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9645) );
  INV_X1 U6330 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4925) );
  NAND2_X1 U6331 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9558), .ZN(n4924) );
  MUX2_X1 U6332 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9645), .S(n8977), .Z(n4926)
         );
  INV_X1 U6333 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5100) );
  INV_X1 U6334 ( .A(n9558), .ZN(n8993) );
  NOR2_X1 U6335 ( .A1(n8977), .A2(n9645), .ZN(n9000) );
  MUX2_X1 U6336 ( .A(n8999), .B(P1_REG2_REG_2__SCAN_IN), .S(n9006), .Z(n4927)
         );
  MUX2_X1 U6337 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n5424), .S(n9421), .Z(n4928)
         );
  INV_X1 U6338 ( .A(n4928), .ZN(n9425) );
  OAI21_X1 U6339 ( .B1(n9421), .B2(n5424), .A(n9424), .ZN(n9022) );
  MUX2_X1 U6340 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n8220), .S(n9017), .Z(n9021)
         );
  NOR2_X1 U6341 ( .A1(n9022), .A2(n9021), .ZN(n9020) );
  INV_X1 U6342 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5662) );
  MUX2_X1 U6343 ( .A(n5662), .B(P1_REG2_REG_5__SCAN_IN), .S(n9563), .Z(n9569)
         );
  INV_X1 U6344 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n4930) );
  MUX2_X1 U6345 ( .A(n4930), .B(P1_REG2_REG_6__SCAN_IN), .S(n5847), .Z(n4931)
         );
  INV_X1 U6346 ( .A(n4931), .ZN(n5133) );
  NAND2_X1 U6347 ( .A1(n4932), .A2(n5132), .ZN(n5167) );
  OR2_X1 U6348 ( .A1(n4934), .A2(n4933), .ZN(n4935) );
  XNOR2_X1 U6349 ( .A(n4935), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6053) );
  INV_X1 U6350 ( .A(n6053), .ZN(n5162) );
  INV_X1 U6351 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5855) );
  NOR2_X1 U6352 ( .A1(n5162), .A2(n5855), .ZN(n5165) );
  OR2_X1 U6353 ( .A1(n6053), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5160) );
  OAI21_X1 U6354 ( .B1(n5167), .B2(n5165), .A(n5160), .ZN(n5159) );
  INV_X1 U6355 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6079) );
  MUX2_X1 U6356 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6079), .S(n6281), .Z(n5152)
         );
  INV_X1 U6357 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6438) );
  MUX2_X1 U6358 ( .A(n6438), .B(P1_REG2_REG_10__SCAN_IN), .S(n9037), .Z(n9033)
         );
  NOR2_X1 U6359 ( .A1(n9034), .A2(n9033), .ZN(n9032) );
  AOI21_X1 U6360 ( .B1(n9037), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9032), .ZN(
        n9581) );
  INV_X1 U6361 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n4936) );
  MUX2_X1 U6362 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n4936), .S(n6707), .Z(n4937)
         );
  INV_X1 U6363 ( .A(n4937), .ZN(n5936) );
  NOR2_X1 U6364 ( .A1(n5937), .A2(n5936), .ZN(n5935) );
  AOI21_X1 U6365 ( .B1(n6707), .B2(P1_REG2_REG_13__SCAN_IN), .A(n5935), .ZN(
        n4940) );
  NAND2_X1 U6366 ( .A1(n4938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4939) );
  XNOR2_X1 U6367 ( .A(n4939), .B(P1_IR_REG_14__SCAN_IN), .ZN(n6768) );
  INV_X1 U6368 ( .A(n6768), .ZN(n5278) );
  NAND2_X1 U6369 ( .A1(n4940), .A2(n5278), .ZN(n4941) );
  XNOR2_X1 U6370 ( .A(n6768), .B(n4940), .ZN(n6159) );
  INV_X1 U6371 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U6372 ( .A1(n6159), .A2(n6158), .ZN(n6157) );
  NAND2_X1 U6373 ( .A1(n4941), .A2(n6157), .ZN(n9042) );
  INV_X1 U6374 ( .A(n5641), .ZN(n4943) );
  NAND2_X1 U6375 ( .A1(n4943), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4944) );
  XNOR2_X1 U6376 ( .A(n4944), .B(n5640), .ZN(n9048) );
  INV_X1 U6377 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8200) );
  NOR2_X1 U6378 ( .A1(n8991), .A2(P1_U3084), .ZN(n6944) );
  NAND2_X1 U6379 ( .A1(n4960), .A2(n6944), .ZN(n9094) );
  NOR2_X1 U6380 ( .A1(n9094), .A2(n4283), .ZN(n9588) );
  INV_X1 U6381 ( .A(n9588), .ZN(n9571) );
  AOI211_X1 U6382 ( .C1(n4945), .C2(n8200), .A(n9043), .B(n9571), .ZN(n4965)
         );
  OR2_X1 U6383 ( .A1(P1_U3083), .A2(n4946), .ZN(n9593) );
  INV_X1 U6384 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n4947) );
  NOR2_X1 U6385 ( .A1(n9593), .A2(n4947), .ZN(n4964) );
  INV_X1 U6386 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9522) );
  NOR2_X1 U6387 ( .A1(n5278), .A2(n9522), .ZN(n4948) );
  AOI21_X1 U6388 ( .B1(n9522), .B2(n5278), .A(n4948), .ZN(n6161) );
  INV_X1 U6389 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6602) );
  MUX2_X1 U6390 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6602), .S(n6707), .Z(n5934)
         );
  INV_X1 U6391 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6593) );
  MUX2_X1 U6392 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6593), .S(n6590), .Z(n5700)
         );
  INV_X1 U6393 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9543) );
  INV_X1 U6394 ( .A(n9578), .ZN(n5142) );
  AOI22_X1 U6395 ( .A1(n9578), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n9543), .B2(
        n5142), .ZN(n9585) );
  NOR2_X1 U6396 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n9037), .ZN(n4949) );
  AOI21_X1 U6397 ( .B1(n9037), .B2(P1_REG1_REG_10__SCAN_IN), .A(n4949), .ZN(
        n9030) );
  NOR2_X1 U6398 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6385), .ZN(n4950) );
  AOI21_X1 U6399 ( .B1(n6385), .B2(P1_REG1_REG_9__SCAN_IN), .A(n4950), .ZN(
        n5241) );
  NOR2_X1 U6400 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n5847), .ZN(n4957) );
  INV_X1 U6401 ( .A(n5847), .ZN(n5036) );
  INV_X1 U6402 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9739) );
  AOI22_X1 U6403 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n5036), .B1(n5847), .B2(
        n9739), .ZN(n5128) );
  NAND2_X1 U6404 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9563), .ZN(n4956) );
  INV_X1 U6405 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9736) );
  INV_X1 U6406 ( .A(n9421), .ZN(n4954) );
  INV_X1 U6407 ( .A(n9006), .ZN(n4953) );
  INV_X1 U6408 ( .A(n8977), .ZN(n8973) );
  XOR2_X1 U6409 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n8977), .Z(n8981) );
  INV_X1 U6410 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9730) );
  NOR3_X1 U6411 ( .A1(n8981), .A2(n8993), .A3(n9730), .ZN(n8982) );
  INV_X1 U6412 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9732) );
  MUX2_X1 U6413 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9732), .S(n9006), .Z(n4951)
         );
  INV_X1 U6414 ( .A(n9008), .ZN(n4952) );
  INV_X1 U6415 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9734) );
  MUX2_X1 U6416 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9734), .S(n9421), .Z(n9429)
         );
  NOR2_X1 U6417 ( .A1(n9430), .A2(n9429), .ZN(n9428) );
  AOI21_X1 U6418 ( .B1(n4954), .B2(P1_REG1_REG_3__SCAN_IN), .A(n9428), .ZN(
        n9016) );
  MUX2_X1 U6419 ( .A(n9736), .B(P1_REG1_REG_4__SCAN_IN), .S(n9017), .Z(n9015)
         );
  NAND2_X1 U6420 ( .A1(n9016), .A2(n9015), .ZN(n9014) );
  INV_X1 U6421 ( .A(n9014), .ZN(n4955) );
  AOI21_X1 U6422 ( .B1(n9736), .B2(n9017), .A(n4955), .ZN(n9567) );
  INV_X1 U6423 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5664) );
  MUX2_X1 U6424 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5664), .S(n9563), .Z(n9566)
         );
  NAND2_X1 U6425 ( .A1(n9567), .A2(n9566), .ZN(n9565) );
  NAND2_X1 U6426 ( .A1(n4956), .A2(n9565), .ZN(n5127) );
  NOR2_X1 U6427 ( .A1(n4957), .A2(n5126), .ZN(n5169) );
  INV_X1 U6428 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9741) );
  NOR2_X1 U6429 ( .A1(n5162), .A2(n9741), .ZN(n5168) );
  NOR2_X1 U6430 ( .A1(n6281), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4958) );
  AOI21_X1 U6431 ( .B1(n6281), .B2(P1_REG1_REG_8__SCAN_IN), .A(n4958), .ZN(
        n5149) );
  NAND2_X1 U6432 ( .A1(n5163), .A2(n5149), .ZN(n5148) );
  OAI21_X1 U6433 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6281), .A(n5148), .ZN(
        n5242) );
  NAND2_X1 U6434 ( .A1(n9030), .A2(n9031), .ZN(n9029) );
  OAI21_X1 U6435 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9037), .A(n9029), .ZN(
        n9584) );
  NAND2_X1 U6436 ( .A1(n5700), .A2(n5701), .ZN(n5699) );
  OAI21_X1 U6437 ( .B1(n6590), .B2(P1_REG1_REG_12__SCAN_IN), .A(n5699), .ZN(
        n5933) );
  NAND2_X1 U6438 ( .A1(n5934), .A2(n5933), .ZN(n5932) );
  OAI21_X1 U6439 ( .B1(n6707), .B2(P1_REG1_REG_13__SCAN_IN), .A(n5932), .ZN(
        n6162) );
  NAND2_X1 U6440 ( .A1(n6161), .A2(n6162), .ZN(n6160) );
  OAI21_X1 U6441 ( .B1(n6768), .B2(P1_REG1_REG_14__SCAN_IN), .A(n6160), .ZN(
        n9047) );
  XNOR2_X1 U6442 ( .A(n9048), .B(n9047), .ZN(n4961) );
  INV_X1 U6443 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9516) );
  NOR2_X1 U6444 ( .A1(n9516), .A2(n4961), .ZN(n9049) );
  AND2_X1 U6445 ( .A1(n5846), .A2(P1_STATE_REG_SCAN_IN), .ZN(n4959) );
  AND2_X1 U6446 ( .A1(n4960), .A2(n4959), .ZN(n9560) );
  AND2_X1 U6447 ( .A1(n9560), .A2(n8991), .ZN(n9587) );
  INV_X1 U6448 ( .A(n9587), .ZN(n9427) );
  AOI211_X1 U6449 ( .C1(n4961), .C2(n9516), .A(n9049), .B(n9427), .ZN(n4963)
         );
  INV_X1 U6450 ( .A(n9094), .ZN(n5166) );
  AND2_X1 U6451 ( .A1(n5166), .A2(n4283), .ZN(n9579) );
  INV_X1 U6452 ( .A(n9579), .ZN(n9422) );
  NAND2_X1 U6453 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8663) );
  OAI21_X1 U6454 ( .B1(n9422), .B2(n9048), .A(n8663), .ZN(n4962) );
  OR4_X1 U6455 ( .A1(n4965), .A2(n4964), .A3(n4963), .A4(n4962), .ZN(P1_U3256)
         );
  INV_X1 U6456 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4966) );
  INV_X1 U6457 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6458 ( .A1(n7532), .A2(P1_U3084), .ZN(n7364) );
  AND2_X1 U6459 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4969) );
  NAND2_X1 U6460 ( .A1(n4986), .A2(n4969), .ZN(n5216) );
  INV_X1 U6461 ( .A(SI_1_), .ZN(n4970) );
  MUX2_X1 U6462 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4986), .Z(n4971) );
  XNOR2_X1 U6463 ( .A(n4972), .B(n4971), .ZN(n5456) );
  OAI222_X1 U6464 ( .A1(n7361), .A2(n5284), .B1(n7364), .B2(n5456), .C1(
        P1_U3084), .C2(n8977), .ZN(P1_U3352) );
  INV_X1 U6465 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6466 ( .A1(n4972), .A2(n4971), .ZN(n4975) );
  NAND2_X1 U6467 ( .A1(n4973), .A2(SI_1_), .ZN(n4974) );
  INV_X1 U6468 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5555) );
  MUX2_X1 U6469 ( .A(n5555), .B(n5418), .S(n4986), .Z(n4983) );
  XNOR2_X1 U6470 ( .A(n4981), .B(n4982), .ZN(n5556) );
  OAI222_X1 U6471 ( .A1(n7361), .A2(n5418), .B1(n7364), .B2(n5556), .C1(
        P1_U3084), .C2(n9006), .ZN(P1_U3351) );
  AND2_X1 U6472 ( .A1(n7532), .A2(P2_U3152), .ZN(n8525) );
  INV_X1 U6473 ( .A(n8525), .ZN(n7817) );
  INV_X1 U6474 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5457) );
  MUX2_X1 U6475 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4976), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n4979) );
  INV_X1 U6476 ( .A(n4977), .ZN(n4978) );
  NAND2_X1 U6477 ( .A1(n4979), .A2(n4978), .ZN(n5314) );
  OAI222_X1 U6478 ( .A1(n7817), .A2(n5457), .B1(n7800), .B2(n5456), .C1(n5314), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  NAND2_X1 U6479 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4320), .ZN(n4980) );
  INV_X1 U6480 ( .A(n5365), .ZN(n5574) );
  INV_X1 U6481 ( .A(n4983), .ZN(n4984) );
  NAND2_X1 U6482 ( .A1(n4984), .A2(SI_2_), .ZN(n4985) );
  INV_X1 U6483 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5572) );
  INV_X1 U6484 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5514) );
  MUX2_X1 U6485 ( .A(n5572), .B(n5514), .S(n4986), .Z(n4992) );
  XNOR2_X1 U6486 ( .A(n4992), .B(SI_3_), .ZN(n4990) );
  XNOR2_X1 U6487 ( .A(n4991), .B(n4990), .ZN(n5571) );
  OAI222_X1 U6488 ( .A1(n5574), .A2(P2_U3152), .B1(n7800), .B2(n5571), .C1(
        n5572), .C2(n7817), .ZN(P2_U3355) );
  OR2_X1 U6489 ( .A1(n4977), .A2(n8522), .ZN(n4988) );
  INV_X1 U6490 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4987) );
  OAI222_X1 U6491 ( .A1(n7817), .A2(n5555), .B1(n7800), .B2(n5556), .C1(n5559), 
        .C2(P2_U3152), .ZN(P2_U3356) );
  NAND2_X1 U6492 ( .A1(n5005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4989) );
  XNOR2_X1 U6493 ( .A(n4989), .B(P2_IR_REG_4__SCAN_IN), .ZN(n5721) );
  INV_X1 U6494 ( .A(n5721), .ZN(n4995) );
  INV_X1 U6495 ( .A(n4992), .ZN(n4993) );
  NAND2_X1 U6496 ( .A1(n4993), .A2(SI_3_), .ZN(n4994) );
  INV_X1 U6497 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5719) );
  INV_X1 U6498 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5645) );
  MUX2_X1 U6499 ( .A(n5719), .B(n5645), .S(n4986), .Z(n5000) );
  XNOR2_X1 U6500 ( .A(n5000), .B(SI_4_), .ZN(n4998) );
  XNOR2_X1 U6501 ( .A(n4999), .B(n4998), .ZN(n5717) );
  OAI222_X1 U6502 ( .A1(n4995), .A2(P2_U3152), .B1(n7800), .B2(n5717), .C1(
        n5719), .C2(n7817), .ZN(P2_U3354) );
  OR2_X1 U6503 ( .A1(n5005), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U6504 ( .A1(n4996), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4997) );
  XNOR2_X1 U6505 ( .A(n4997), .B(P2_IR_REG_5__SCAN_IN), .ZN(n5378) );
  INV_X1 U6506 ( .A(n5378), .ZN(n5819) );
  NAND2_X1 U6507 ( .A1(n4999), .A2(n4998), .ZN(n5014) );
  INV_X1 U6508 ( .A(n5000), .ZN(n5001) );
  NAND2_X1 U6509 ( .A1(n5001), .A2(SI_4_), .ZN(n5009) );
  NAND2_X1 U6510 ( .A1(n5014), .A2(n5009), .ZN(n5003) );
  INV_X1 U6511 ( .A(SI_5_), .ZN(n8293) );
  XNOR2_X1 U6512 ( .A(n5003), .B(n5010), .ZN(n5817) );
  OAI222_X1 U6513 ( .A1(n5819), .A2(P2_U3152), .B1(n7800), .B2(n5817), .C1(
        n5002), .C2(n7817), .ZN(P2_U3353) );
  NOR2_X1 U6514 ( .A1(n5005), .A2(n5004), .ZN(n5006) );
  OR2_X1 U6515 ( .A1(n5006), .A2(n8522), .ZN(n5007) );
  XNOR2_X1 U6516 ( .A(n5007), .B(P2_IR_REG_6__SCAN_IN), .ZN(n5404) );
  INV_X1 U6517 ( .A(n5404), .ZN(n6010) );
  NAND2_X1 U6518 ( .A1(n5008), .A2(SI_5_), .ZN(n5012) );
  AND2_X1 U6519 ( .A1(n5009), .A2(n5012), .ZN(n5013) );
  INV_X1 U6520 ( .A(n5010), .ZN(n5011) );
  INV_X1 U6521 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5037) );
  MUX2_X1 U6522 ( .A(n6008), .B(n5037), .S(n7532), .Z(n5029) );
  OAI222_X1 U6523 ( .A1(n6010), .A2(P2_U3152), .B1(n7800), .B2(n6007), .C1(
        n6008), .C2(n7817), .ZN(P2_U3352) );
  NAND2_X1 U6524 ( .A1(n5231), .A2(n5015), .ZN(n5523) );
  INV_X1 U6525 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8224) );
  NAND3_X1 U6526 ( .A1(n6907), .A2(P1_B_REG_SCAN_IN), .A3(n6764), .ZN(n5019)
         );
  INV_X1 U6527 ( .A(n6764), .ZN(n5017) );
  INV_X1 U6528 ( .A(P1_B_REG_SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6529 ( .A1(n5017), .A2(n5016), .ZN(n5018) );
  NAND2_X1 U6530 ( .A1(n5019), .A2(n5018), .ZN(n5020) );
  OR2_X1 U6531 ( .A1(n9664), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U6532 ( .A1(n7333), .A2(n6907), .ZN(n5021) );
  NAND2_X1 U6533 ( .A1(n9665), .A2(n9393), .ZN(n5023) );
  OAI21_X1 U6534 ( .B1(n9665), .B2(n8224), .A(n5023), .ZN(P1_U3441) );
  INV_X1 U6535 ( .A(n9665), .ZN(n5220) );
  OR2_X1 U6536 ( .A1(n9664), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6537 ( .A1(n7333), .A2(n6764), .ZN(n5024) );
  NAND2_X1 U6538 ( .A1(n5025), .A2(n5024), .ZN(n5875) );
  NAND2_X1 U6539 ( .A1(n5220), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5026) );
  OAI21_X1 U6540 ( .B1(n5220), .B2(n5875), .A(n5026), .ZN(P1_U3440) );
  NAND2_X1 U6541 ( .A1(n5028), .A2(n5027), .ZN(n5032) );
  INV_X1 U6542 ( .A(n5029), .ZN(n5030) );
  NAND2_X1 U6543 ( .A1(n5030), .A2(SI_6_), .ZN(n5031) );
  MUX2_X1 U6544 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7532), .Z(n5043) );
  XNOR2_X1 U6545 ( .A(n5042), .B(n5040), .ZN(n6052) );
  INV_X1 U6546 ( .A(n6052), .ZN(n5038) );
  OR2_X1 U6547 ( .A1(n5033), .A2(n8522), .ZN(n5034) );
  XNOR2_X1 U6548 ( .A(n5034), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6016) );
  AOI22_X1 U6549 ( .A1(n6016), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8525), .ZN(n5035) );
  OAI21_X1 U6550 ( .B1(n5038), .B2(n7800), .A(n5035), .ZN(P2_U3351) );
  INV_X1 U6551 ( .A(n7364), .ZN(n6660) );
  INV_X1 U6552 ( .A(n6660), .ZN(n9417) );
  OAI222_X1 U6553 ( .A1(n7361), .A2(n5514), .B1(n9417), .B2(n5571), .C1(
        P1_U3084), .C2(n9421), .ZN(P1_U3350) );
  INV_X1 U6554 ( .A(n9563), .ZN(n5766) );
  OAI222_X1 U6555 ( .A1(n7361), .A2(n4508), .B1(n9417), .B2(n5817), .C1(
        P1_U3084), .C2(n5766), .ZN(P1_U3348) );
  OAI222_X1 U6556 ( .A1(n7361), .A2(n5037), .B1(n9417), .B2(n6007), .C1(
        P1_U3084), .C2(n5036), .ZN(P1_U3347) );
  OAI222_X1 U6557 ( .A1(n7361), .A2(n5645), .B1(n9417), .B2(n5717), .C1(
        P1_U3084), .C2(n9017), .ZN(P1_U3349) );
  INV_X1 U6558 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5039) );
  OAI222_X1 U6559 ( .A1(n7361), .A2(n5039), .B1(n7364), .B2(n5038), .C1(
        P1_U3084), .C2(n5162), .ZN(P1_U3346) );
  NAND2_X1 U6560 ( .A1(n5042), .A2(n5041), .ZN(n5045) );
  NAND2_X1 U6561 ( .A1(n5043), .A2(SI_7_), .ZN(n5044) );
  NAND2_X1 U6562 ( .A1(n5045), .A2(n5044), .ZN(n5071) );
  INV_X1 U6563 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5046) );
  MUX2_X1 U6564 ( .A(n5046), .B(n5055), .S(n7532), .Z(n5048) );
  INV_X1 U6565 ( .A(SI_8_), .ZN(n5047) );
  INV_X1 U6566 ( .A(n5048), .ZN(n5049) );
  NAND2_X1 U6567 ( .A1(n5049), .A2(SI_8_), .ZN(n5050) );
  XNOR2_X1 U6568 ( .A(n5071), .B(n5070), .ZN(n6280) );
  INV_X1 U6569 ( .A(n6280), .ZN(n5054) );
  NAND2_X1 U6570 ( .A1(n5051), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5052) );
  XNOR2_X1 U6571 ( .A(n5052), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6134) );
  AOI22_X1 U6572 ( .A1(n6134), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n8525), .ZN(n5053) );
  OAI21_X1 U6573 ( .B1(n5054), .B2(n7800), .A(n5053), .ZN(P2_U3350) );
  INV_X1 U6574 ( .A(n6281), .ZN(n5154) );
  OAI222_X1 U6575 ( .A1(n7361), .A2(n5055), .B1(n9417), .B2(n5054), .C1(
        P1_U3084), .C2(n5154), .ZN(P1_U3345) );
  INV_X1 U6576 ( .A(n9840), .ZN(n5056) );
  INV_X1 U6577 ( .A(n9804), .ZN(n5588) );
  NOR2_X1 U6578 ( .A1(n5482), .A2(P2_U3152), .ZN(n7733) );
  INV_X1 U6579 ( .A(n7733), .ZN(n7737) );
  NAND2_X1 U6580 ( .A1(n5588), .A2(n7737), .ZN(n5069) );
  INV_X1 U6581 ( .A(n5057), .ZN(n5058) );
  NAND2_X1 U6582 ( .A1(n5058), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6583 ( .A1(n4873), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5061) );
  INV_X1 U6584 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5060) );
  XNOR2_X1 U6585 ( .A(n5061), .B(n5060), .ZN(n7727) );
  INV_X1 U6586 ( .A(n7727), .ZN(n7550) );
  NAND2_X1 U6587 ( .A1(n7738), .A2(n7550), .ZN(n5578) );
  INV_X1 U6588 ( .A(n5578), .ZN(n5485) );
  NAND2_X1 U6589 ( .A1(n9804), .A2(n5485), .ZN(n5067) );
  INV_X1 U6590 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U6591 ( .A1(n5067), .A2(n5466), .ZN(n5068) );
  NOR2_X1 U6592 ( .A1(n9755), .A2(P2_U3966), .ZN(P2_U3151) );
  OR2_X2 U6593 ( .A1(n5071), .A2(n5070), .ZN(n5073) );
  INV_X1 U6594 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5074) );
  MUX2_X1 U6595 ( .A(n5074), .B(n5082), .S(n7532), .Z(n5075) );
  INV_X1 U6596 ( .A(SI_9_), .ZN(n8256) );
  INV_X1 U6597 ( .A(n5075), .ZN(n5076) );
  NAND2_X1 U6598 ( .A1(n5076), .A2(SI_9_), .ZN(n5077) );
  INV_X1 U6599 ( .A(n6384), .ZN(n5083) );
  NAND2_X1 U6600 ( .A1(n5079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5080) );
  XNOR2_X1 U6601 ( .A(n5080), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6332) );
  AOI22_X1 U6602 ( .A1(n6332), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8525), .ZN(n5081) );
  OAI21_X1 U6603 ( .B1(n5083), .B2(n7800), .A(n5081), .ZN(P2_U3349) );
  INV_X1 U6604 ( .A(n6385), .ZN(n5244) );
  OAI222_X1 U6605 ( .A1(n7364), .A2(n5083), .B1(n5244), .B2(P1_U3084), .C1(
        n5082), .C2(n7361), .ZN(P1_U3344) );
  NAND2_X1 U6606 ( .A1(n5084), .A2(n4828), .ZN(n5086) );
  NAND2_X1 U6607 ( .A1(n5086), .A2(n5085), .ZN(n5138) );
  INV_X1 U6608 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5088) );
  INV_X1 U6609 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5087) );
  MUX2_X1 U6610 ( .A(n5088), .B(n5087), .S(n7532), .Z(n5090) );
  INV_X1 U6611 ( .A(SI_10_), .ZN(n5089) );
  INV_X1 U6612 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U6613 ( .A1(n5091), .A2(SI_10_), .ZN(n5092) );
  XNOR2_X1 U6614 ( .A(n5138), .B(n4826), .ZN(n6448) );
  INV_X1 U6615 ( .A(n6448), .ZN(n5096) );
  XNOR2_X1 U6616 ( .A(n5143), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6449) );
  AOI22_X1 U6617 ( .A1(n6449), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8525), .ZN(n5094) );
  OAI21_X1 U6618 ( .B1(n5096), .B2(n7800), .A(n5094), .ZN(P2_U3348) );
  INV_X1 U6619 ( .A(n7361), .ZN(n6945) );
  AOI22_X1 U6620 ( .A1(n9037), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n6945), .ZN(n5095) );
  OAI21_X1 U6621 ( .B1(n5096), .B2(n9417), .A(n5095), .ZN(P1_U3343) );
  INV_X1 U6622 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5111) );
  INV_X1 U6623 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9413) );
  INV_X1 U6624 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5101) );
  OR2_X1 U6625 ( .A1(n5300), .A2(n9730), .ZN(n5104) );
  AND2_X1 U6626 ( .A1(n5105), .A2(n5104), .ZN(n5108) );
  INV_X1 U6627 ( .A(n5299), .ZN(n5528) );
  INV_X1 U6628 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5106) );
  OR2_X1 U6629 ( .A1(n4286), .A2(n5106), .ZN(n5107) );
  NAND2_X1 U6630 ( .A1(n8702), .A2(P1_U4006), .ZN(n5110) );
  OAI21_X1 U6631 ( .B1(P1_U4006), .B2(n5111), .A(n5110), .ZN(P1_U3555) );
  INV_X1 U6632 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6633 ( .A1(n5115), .A2(n5116), .ZN(n8523) );
  INV_X1 U6634 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5113) );
  XNOR2_X2 U6635 ( .A(n5114), .B(n5113), .ZN(n7797) );
  XNOR2_X2 U6636 ( .A(n5117), .B(n5116), .ZN(n5451) );
  AND2_X2 U6637 ( .A1(n7797), .A2(n5451), .ZN(n6027) );
  NAND2_X1 U6638 ( .A1(n7517), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5123) );
  INV_X1 U6639 ( .A(n5451), .ZN(n5118) );
  INV_X1 U6640 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5119) );
  OR2_X1 U6641 ( .A1(n7522), .A2(n5119), .ZN(n5122) );
  INV_X1 U6642 ( .A(n7797), .ZN(n5120) );
  INV_X1 U6643 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8007) );
  OR2_X1 U6644 ( .A1(n4278), .A2(n8007), .ZN(n5121) );
  AND3_X1 U6645 ( .A1(n5123), .A2(n5122), .A3(n5121), .ZN(n7540) );
  INV_X1 U6646 ( .A(n7540), .ZN(n8011) );
  NAND2_X1 U6647 ( .A1(n8011), .A2(P2_U3966), .ZN(n5124) );
  OAI21_X1 U6648 ( .B1(P2_U3966), .B2(n5125), .A(n5124), .ZN(P2_U3583) );
  AOI21_X1 U6649 ( .B1(n5128), .B2(n5127), .A(n5126), .ZN(n5137) );
  NAND2_X1 U6650 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3084), .ZN(n5862) );
  INV_X1 U6651 ( .A(n5862), .ZN(n5131) );
  INV_X1 U6652 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n5129) );
  NOR2_X1 U6653 ( .A1(n9593), .A2(n5129), .ZN(n5130) );
  AOI211_X1 U6654 ( .C1(n9579), .C2(n5847), .A(n5131), .B(n5130), .ZN(n5136)
         );
  OAI211_X1 U6655 ( .C1(n5134), .C2(n5133), .A(n9588), .B(n5132), .ZN(n5135)
         );
  OAI211_X1 U6656 ( .C1(n5137), .C2(n9427), .A(n5136), .B(n5135), .ZN(P1_U3247) );
  NAND2_X1 U6657 ( .A1(n5138), .A2(n4826), .ZN(n5140) );
  INV_X1 U6658 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5146) );
  INV_X1 U6659 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5141) );
  MUX2_X1 U6660 ( .A(n5146), .B(n5141), .S(n7532), .Z(n5178) );
  XNOR2_X1 U6661 ( .A(n5181), .B(n5177), .ZN(n6584) );
  INV_X1 U6662 ( .A(n6584), .ZN(n5147) );
  OAI222_X1 U6663 ( .A1(n7364), .A2(n5147), .B1(n5142), .B2(P1_U3084), .C1(
        n5141), .C2(n7361), .ZN(P1_U3342) );
  NAND2_X1 U6664 ( .A1(n5143), .A2(n5188), .ZN(n5144) );
  NAND2_X1 U6665 ( .A1(n5144), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5145) );
  XNOR2_X1 U6666 ( .A(n5145), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6496) );
  INV_X1 U6667 ( .A(n6496), .ZN(n6315) );
  OAI222_X1 U6668 ( .A1(P2_U3152), .A2(n6315), .B1(n7800), .B2(n5147), .C1(
        n5146), .C2(n7817), .ZN(P2_U3347) );
  OAI21_X1 U6669 ( .B1(n5149), .B2(n5163), .A(n5148), .ZN(n5150) );
  NAND2_X1 U6670 ( .A1(n5150), .A2(n9587), .ZN(n5158) );
  OAI21_X1 U6671 ( .B1(n5152), .B2(n5159), .A(n5151), .ZN(n5156) );
  NAND2_X1 U6672 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3084), .ZN(n6325) );
  INV_X1 U6673 ( .A(n9593), .ZN(n9564) );
  NAND2_X1 U6674 ( .A1(n9564), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n5153) );
  OAI211_X1 U6675 ( .C1(n9422), .C2(n5154), .A(n6325), .B(n5153), .ZN(n5155)
         );
  AOI21_X1 U6676 ( .B1(n5156), .B2(n9588), .A(n5155), .ZN(n5157) );
  NAND2_X1 U6677 ( .A1(n5158), .A2(n5157), .ZN(P1_U3249) );
  OAI211_X1 U6678 ( .C1(n5167), .C2(n5160), .A(n5159), .B(n9588), .ZN(n5161)
         );
  OAI21_X1 U6679 ( .B1(n9422), .B2(n5162), .A(n5161), .ZN(n5175) );
  NAND2_X1 U6680 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n5173) );
  NAND2_X1 U6681 ( .A1(n5162), .A2(n9741), .ZN(n5164) );
  OAI211_X1 U6682 ( .C1(n5169), .C2(n5164), .A(n5163), .B(n9587), .ZN(n5172)
         );
  NAND3_X1 U6683 ( .A1(n5167), .A2(n5166), .A3(n5165), .ZN(n5171) );
  NAND3_X1 U6684 ( .A1(n9587), .A2(n5169), .A3(n5168), .ZN(n5170) );
  NAND4_X1 U6685 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n5174)
         );
  AOI211_X1 U6686 ( .C1(n9564), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n5175), .B(
        n5174), .ZN(n5176) );
  INV_X1 U6687 ( .A(n5176), .ZN(P1_U3248) );
  INV_X1 U6688 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5186) );
  INV_X1 U6689 ( .A(n5178), .ZN(n5179) );
  INV_X1 U6690 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5192) );
  MUX2_X1 U6691 ( .A(n5192), .B(n5186), .S(n7532), .Z(n5183) );
  INV_X1 U6692 ( .A(SI_12_), .ZN(n5182) );
  INV_X1 U6693 ( .A(n5183), .ZN(n5184) );
  NAND2_X1 U6694 ( .A1(n5184), .A2(SI_12_), .ZN(n5185) );
  XNOR2_X1 U6695 ( .A(n5263), .B(n5262), .ZN(n6589) );
  INV_X1 U6696 ( .A(n6589), .ZN(n5191) );
  INV_X1 U6697 ( .A(n6590), .ZN(n5704) );
  OAI222_X1 U6698 ( .A1(n7361), .A2(n5186), .B1(n7364), .B2(n5191), .C1(
        P1_U3084), .C2(n5704), .ZN(P1_U3341) );
  NAND2_X1 U6699 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  OR2_X1 U6700 ( .A1(n5272), .A2(n8522), .ZN(n5190) );
  XNOR2_X1 U6701 ( .A(n5190), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6557) );
  INV_X1 U6702 ( .A(n6557), .ZN(n6507) );
  OAI222_X1 U6703 ( .A1(n7817), .A2(n5192), .B1(n7800), .B2(n5191), .C1(n6507), 
        .C2(P2_U3152), .ZN(P2_U3346) );
  XNOR2_X1 U6704 ( .A(n5195), .B(n5194), .ZN(n6260) );
  NAND2_X1 U6705 ( .A1(n5196), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5198) );
  INV_X1 U6706 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5197) );
  XNOR2_X1 U6707 ( .A(n5198), .B(n5197), .ZN(n9188) );
  AND2_X1 U6708 ( .A1(n6260), .A2(n9188), .ZN(n8948) );
  OR2_X1 U6709 ( .A1(n5219), .A2(n8948), .ZN(n5525) );
  INV_X1 U6710 ( .A(n6260), .ZN(n8946) );
  OR2_X1 U6711 ( .A1(n9693), .A2(n8917), .ZN(n5199) );
  NOR4_X1 U6712 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n8309) );
  NOR2_X1 U6713 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n5202) );
  NOR4_X1 U6714 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5201) );
  NOR4_X1 U6715 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5200) );
  NAND4_X1 U6716 ( .A1(n8309), .A2(n5202), .A3(n5201), .A4(n5200), .ZN(n5208)
         );
  NOR4_X1 U6717 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5206) );
  NOR4_X1 U6718 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5205) );
  NOR4_X1 U6719 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n5204) );
  NOR4_X1 U6720 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5203) );
  NAND4_X1 U6721 ( .A1(n5206), .A2(n5205), .A3(n5204), .A4(n5203), .ZN(n5207)
         );
  NOR2_X1 U6722 ( .A1(n5208), .A2(n5207), .ZN(n5209) );
  NOR2_X1 U6723 ( .A1(n9664), .A2(n5209), .ZN(n5874) );
  OR2_X1 U6724 ( .A1(n5874), .A2(n5875), .ZN(n5392) );
  INV_X1 U6725 ( .A(n5392), .ZN(n5210) );
  NAND2_X1 U6726 ( .A1(n5210), .A2(n9393), .ZN(n5221) );
  AND2_X1 U6727 ( .A1(n9396), .A2(n5221), .ZN(n5527) );
  INV_X1 U6728 ( .A(n5527), .ZN(n5211) );
  AND2_X1 U6729 ( .A1(n5211), .A2(n5879), .ZN(n5432) );
  INV_X1 U6730 ( .A(n8917), .ZN(n8934) );
  OR2_X1 U6731 ( .A1(n9652), .A2(n6260), .ZN(n5895) );
  OR2_X1 U6732 ( .A1(n9652), .A2(n9188), .ZN(n5213) );
  NAND2_X1 U6733 ( .A1(n5895), .A2(n5213), .ZN(n9689) );
  INV_X1 U6734 ( .A(n8671), .ZN(n8656) );
  NAND2_X1 U6735 ( .A1(n7532), .A2(SI_0_), .ZN(n5215) );
  INV_X1 U6736 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6737 ( .A1(n5215), .A2(n5214), .ZN(n5217) );
  AND2_X1 U6738 ( .A1(n5217), .A2(n5216), .ZN(n9419) );
  MUX2_X1 U6739 ( .A(n9558), .B(n9419), .S(n5846), .Z(n9654) );
  INV_X1 U6740 ( .A(n5432), .ZN(n8590) );
  INV_X1 U6741 ( .A(n8948), .ZN(n5218) );
  NOR2_X1 U6742 ( .A1(n9646), .A2(n5220), .ZN(n8950) );
  INV_X1 U6743 ( .A(n5221), .ZN(n5236) );
  AND2_X1 U6744 ( .A1(n8950), .A2(n5236), .ZN(n5301) );
  INV_X1 U6745 ( .A(n5301), .ZN(n5222) );
  INV_X1 U6746 ( .A(n4283), .ZN(n8949) );
  INV_X1 U6747 ( .A(n8664), .ZN(n8653) );
  NAND2_X1 U6748 ( .A1(n4284), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5227) );
  INV_X1 U6749 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8975) );
  OR2_X1 U6750 ( .A1(n5425), .A2(n8975), .ZN(n5226) );
  NAND2_X1 U6751 ( .A1(n5299), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5225) );
  INV_X1 U6752 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5223) );
  AOI22_X1 U6753 ( .A1(n8590), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n8653), .B2(
        n5380), .ZN(n5239) );
  NOR2_X1 U6754 ( .A1(n5231), .A2(n8993), .ZN(n5228) );
  AOI21_X1 U6755 ( .B1(n9654), .B2(n7290), .A(n5228), .ZN(n5229) );
  NOR2_X1 U6756 ( .A1(n5231), .A2(n9730), .ZN(n5232) );
  AOI21_X1 U6757 ( .B1(n9654), .B2(n4282), .A(n5232), .ZN(n5233) );
  NAND2_X1 U6758 ( .A1(n5234), .A2(n5233), .ZN(n5279) );
  NAND2_X1 U6759 ( .A1(n5235), .A2(n5279), .ZN(n5283) );
  OAI21_X1 U6760 ( .B1(n5235), .B2(n5279), .A(n5283), .ZN(n8989) );
  NAND3_X1 U6761 ( .A1(n5236), .A2(n9665), .A3(n5219), .ZN(n5237) );
  INV_X1 U6762 ( .A(n8645), .ZN(n8657) );
  NAND2_X1 U6763 ( .A1(n8989), .A2(n8657), .ZN(n5238) );
  OAI211_X1 U6764 ( .C1(n8656), .C2(n8701), .A(n5239), .B(n5238), .ZN(P1_U3230) );
  OAI21_X1 U6765 ( .B1(n5242), .B2(n5241), .A(n5240), .ZN(n5250) );
  NAND2_X1 U6766 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n6411) );
  NAND2_X1 U6767 ( .A1(n9564), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n5243) );
  OAI211_X1 U6768 ( .C1(n9422), .C2(n5244), .A(n6411), .B(n5243), .ZN(n5249)
         );
  AOI211_X1 U6769 ( .C1(n5247), .C2(n5246), .A(n5245), .B(n9571), .ZN(n5248)
         );
  AOI211_X1 U6770 ( .C1(n9587), .C2(n5250), .A(n5249), .B(n5248), .ZN(n5251)
         );
  INV_X1 U6771 ( .A(n5251), .ZN(P1_U3250) );
  INV_X1 U6772 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6603) );
  INV_X1 U6773 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6604) );
  INV_X1 U6774 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8208) );
  INV_X1 U6775 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6880) );
  INV_X1 U6776 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7069) );
  INV_X1 U6777 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8626) );
  INV_X1 U6778 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6779 ( .A1(n7055), .A2(n5252), .ZN(n5253) );
  AND2_X1 U6780 ( .A1(n7103), .A2(n5253), .ZN(n9232) );
  INV_X1 U6781 ( .A(n7167), .ZN(n5254) );
  INV_X1 U6782 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5258) );
  BUF_X4 U6783 ( .A(n5299), .Z(n8678) );
  NAND2_X1 U6784 ( .A1(n8678), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6785 ( .A1(n4284), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5256) );
  OAI211_X1 U6786 ( .C1(n5258), .C2(n8683), .A(n5257), .B(n5256), .ZN(n5259)
         );
  INV_X1 U6787 ( .A(P1_U4006), .ZN(n8972) );
  NAND2_X1 U6788 ( .A1(n8972), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5260) );
  OAI21_X1 U6789 ( .B1(n9242), .B2(n8972), .A(n5260), .ZN(P1_U3576) );
  INV_X1 U6790 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5265) );
  INV_X1 U6791 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5264) );
  MUX2_X1 U6792 ( .A(n5265), .B(n5264), .S(n7532), .Z(n5267) );
  INV_X1 U6793 ( .A(SI_13_), .ZN(n5266) );
  NAND2_X1 U6794 ( .A1(n5267), .A2(n5266), .ZN(n5276) );
  INV_X1 U6795 ( .A(n5267), .ZN(n5268) );
  NAND2_X1 U6796 ( .A1(n5268), .A2(SI_13_), .ZN(n5269) );
  XNOR2_X1 U6797 ( .A(n5275), .B(n4820), .ZN(n6812) );
  INV_X1 U6798 ( .A(n6812), .ZN(n5274) );
  AOI22_X1 U6799 ( .A1(n6707), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6945), .ZN(n5270) );
  OAI21_X1 U6800 ( .B1(n5274), .B2(n9417), .A(n5270), .ZN(P1_U3340) );
  OR2_X1 U6801 ( .A1(n5438), .A2(n8522), .ZN(n5307) );
  XNOR2_X1 U6802 ( .A(n5307), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6849) );
  AOI22_X1 U6803 ( .A1(n6849), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8525), .ZN(n5273) );
  OAI21_X1 U6804 ( .B1(n5274), .B2(n7800), .A(n5273), .ZN(P2_U3345) );
  INV_X1 U6805 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5277) );
  MUX2_X1 U6806 ( .A(n8288), .B(n5277), .S(n7532), .Z(n5615) );
  XNOR2_X1 U6807 ( .A(n5614), .B(n5612), .ZN(n6816) );
  INV_X1 U6808 ( .A(n6816), .ZN(n5309) );
  OAI222_X1 U6809 ( .A1(n9417), .A2(n5309), .B1(n5278), .B2(P1_U3084), .C1(
        n5277), .C2(n7361), .ZN(P1_U3339) );
  AND2_X4 U6810 ( .A1(n9323), .A2(n5281), .ZN(n5653) );
  NAND2_X1 U6811 ( .A1(n5283), .A2(n5282), .ZN(n5295) );
  NAND2_X1 U6812 ( .A1(n5380), .A2(n7290), .ZN(n5290) );
  NAND2_X1 U6813 ( .A1(n5285), .A2(n4968), .ZN(n5513) );
  OR2_X1 U6814 ( .A1(n5513), .A2(n5284), .ZN(n5288) );
  OR2_X1 U6815 ( .A1(n6051), .A2(n5456), .ZN(n5287) );
  OR2_X1 U6816 ( .A1(n5285), .A2(n8977), .ZN(n5286) );
  OR2_X1 U6817 ( .A1(n5382), .A2(n7319), .ZN(n5289) );
  NAND2_X1 U6818 ( .A1(n5290), .A2(n5289), .ZN(n5291) );
  NAND2_X1 U6819 ( .A1(n5412), .A2(n5411), .ZN(n5298) );
  NAND2_X1 U6820 ( .A1(n5380), .A2(n7286), .ZN(n5297) );
  OR2_X1 U6821 ( .A1(n5382), .A2(n7318), .ZN(n5296) );
  NAND2_X1 U6822 ( .A1(n5297), .A2(n5296), .ZN(n5410) );
  XNOR2_X1 U6823 ( .A(n5298), .B(n5410), .ZN(n5305) );
  NAND2_X1 U6824 ( .A1(n8671), .A2(n9634), .ZN(n5303) );
  INV_X1 U6825 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U6826 ( .A1(n8678), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5417) );
  OR2_X1 U6827 ( .A1(n5300), .A2(n9732), .ZN(n5414) );
  NAND4_X1 U6828 ( .A1(n5415), .A2(n5416), .A3(n5417), .A4(n5414), .ZN(n8971)
         );
  AOI22_X1 U6829 ( .A1(n8653), .A2(n8971), .B1(n8666), .B2(n8702), .ZN(n5302)
         );
  OAI211_X1 U6830 ( .C1(n5432), .C2(n8975), .A(n5303), .B(n5302), .ZN(n5304)
         );
  AOI21_X1 U6831 ( .B1(n5305), .B2(n8657), .A(n5304), .ZN(n5306) );
  INV_X1 U6832 ( .A(n5306), .ZN(P1_U3220) );
  NAND2_X1 U6833 ( .A1(n5307), .A2(n5436), .ZN(n5308) );
  NAND2_X1 U6834 ( .A1(n5308), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5635) );
  XNOR2_X1 U6835 ( .A(n5635), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6959) );
  INV_X1 U6836 ( .A(n6959), .ZN(n6854) );
  OAI222_X1 U6837 ( .A1(P2_U3152), .A2(n6854), .B1(n7800), .B2(n5309), .C1(
        n8288), .C2(n7817), .ZN(P2_U3344) );
  OR2_X1 U6838 ( .A1(n5310), .A2(P2_U3152), .ZN(n6952) );
  NAND2_X1 U6839 ( .A1(n9804), .A2(n5578), .ZN(n5311) );
  OAI211_X1 U6840 ( .C1(n5483), .C2(n6952), .A(n5311), .B(n7737), .ZN(n5322)
         );
  NAND2_X1 U6841 ( .A1(n5322), .A2(n5466), .ZN(n5312) );
  INV_X2 U6842 ( .A(P2_U3966), .ZN(n7941) );
  NAND2_X1 U6843 ( .A1(n5312), .A2(n7941), .ZN(n5329) );
  NAND2_X1 U6844 ( .A1(n5329), .A2(n5310), .ZN(n9751) );
  INV_X1 U6845 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5313) );
  MUX2_X1 U6846 ( .A(n5313), .B(P2_REG1_REG_4__SCAN_IN), .S(n5721), .Z(n5317)
         );
  INV_X1 U6847 ( .A(n5559), .ZN(n9455) );
  INV_X1 U6848 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9758) );
  INV_X1 U6849 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9911) );
  NOR3_X1 U6850 ( .A1(n9758), .A2(n9911), .A3(n9436), .ZN(n9435) );
  AOI21_X1 U6851 ( .B1(n9443), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9435), .ZN(
        n9448) );
  XOR2_X1 U6852 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5559), .Z(n9447) );
  NOR2_X1 U6853 ( .A1(n9448), .A2(n9447), .ZN(n9446) );
  OR2_X1 U6854 ( .A1(n5365), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6855 ( .A1(n5365), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6856 ( .A1(n5316), .A2(n5315), .ZN(n5352) );
  NOR2_X1 U6857 ( .A1(n5353), .A2(n5352), .ZN(n5354) );
  NAND2_X1 U6858 ( .A1(n5317), .A2(n5318), .ZN(n5320) );
  NOR2_X1 U6859 ( .A1(n5318), .A2(n5317), .ZN(n5336) );
  INV_X1 U6860 ( .A(n5336), .ZN(n5319) );
  NAND2_X1 U6861 ( .A1(n5320), .A2(n5319), .ZN(n5325) );
  AND2_X1 U6862 ( .A1(n5466), .A2(n8009), .ZN(n5321) );
  NAND2_X1 U6863 ( .A1(n5322), .A2(n5321), .ZN(n9753) );
  NAND2_X1 U6864 ( .A1(n9755), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6865 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n5323) );
  OAI211_X1 U6866 ( .C1(n5325), .C2(n9753), .A(n5324), .B(n5323), .ZN(n5333)
         );
  INV_X1 U6867 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U6868 ( .A1(n9443), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5326) );
  INV_X1 U6869 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6870 ( .A1(n5365), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5327) );
  OAI21_X1 U6871 ( .B1(n5365), .B2(P2_REG2_REG_3__SCAN_IN), .A(n5327), .ZN(
        n5361) );
  NOR2_X1 U6872 ( .A1(n5362), .A2(n5361), .ZN(n5360) );
  MUX2_X1 U6873 ( .A(n8206), .B(P2_REG2_REG_4__SCAN_IN), .S(n5721), .Z(n5330)
         );
  NOR2_X1 U6874 ( .A1(n5310), .A2(n8009), .ZN(n5328) );
  AOI211_X1 U6875 ( .C1(n5331), .C2(n5330), .A(n5344), .B(n9449), .ZN(n5332)
         );
  AOI211_X1 U6876 ( .C1(n9456), .C2(n5721), .A(n5333), .B(n5332), .ZN(n5334)
         );
  INV_X1 U6877 ( .A(n5334), .ZN(P2_U3249) );
  OR2_X1 U6878 ( .A1(n5404), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6879 ( .A1(n5404), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6880 ( .A1(n5335), .A2(n5397), .ZN(n5339) );
  AOI21_X1 U6881 ( .B1(n5721), .B2(P2_REG1_REG_4__SCAN_IN), .A(n5336), .ZN(
        n5367) );
  OR2_X1 U6882 ( .A1(n5378), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6883 ( .A1(n5378), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6884 ( .A1(n5338), .A2(n5337), .ZN(n5368) );
  NOR2_X1 U6885 ( .A1(n5367), .A2(n5368), .ZN(n5369) );
  NAND2_X1 U6886 ( .A1(n5339), .A2(n5340), .ZN(n5341) );
  NAND2_X1 U6887 ( .A1(n5341), .A2(n5396), .ZN(n5343) );
  NAND2_X1 U6888 ( .A1(n9755), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6889 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7906) );
  OAI211_X1 U6890 ( .C1(n9753), .C2(n5343), .A(n5342), .B(n7906), .ZN(n5350)
         );
  NAND2_X1 U6891 ( .A1(n5378), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5345) );
  OAI21_X1 U6892 ( .B1(n5378), .B2(P2_REG2_REG_5__SCAN_IN), .A(n5345), .ZN(
        n5375) );
  NAND2_X1 U6893 ( .A1(n5404), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5346) );
  OAI21_X1 U6894 ( .B1(n5404), .B2(P2_REG2_REG_6__SCAN_IN), .A(n5346), .ZN(
        n5347) );
  NOR2_X1 U6895 ( .A1(n5348), .A2(n5347), .ZN(n5403) );
  AOI211_X1 U6896 ( .C1(n5348), .C2(n5347), .A(n5403), .B(n9449), .ZN(n5349)
         );
  AOI211_X1 U6897 ( .C1(n9456), .C2(n5404), .A(n5350), .B(n5349), .ZN(n5351)
         );
  INV_X1 U6898 ( .A(n5351), .ZN(P2_U3251) );
  NAND2_X1 U6899 ( .A1(n5353), .A2(n5352), .ZN(n5356) );
  INV_X1 U6900 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U6901 ( .A1(n5356), .A2(n5355), .ZN(n5359) );
  NAND2_X1 U6902 ( .A1(n9755), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6903 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n5357) );
  OAI211_X1 U6904 ( .C1(n5359), .C2(n9753), .A(n5358), .B(n5357), .ZN(n5364)
         );
  AOI211_X1 U6905 ( .C1(n5362), .C2(n5361), .A(n5360), .B(n9449), .ZN(n5363)
         );
  AOI211_X1 U6906 ( .C1(n9456), .C2(n5365), .A(n5364), .B(n5363), .ZN(n5366)
         );
  INV_X1 U6907 ( .A(n5366), .ZN(P2_U3248) );
  NAND2_X1 U6908 ( .A1(n5368), .A2(n5367), .ZN(n5371) );
  INV_X1 U6909 ( .A(n5369), .ZN(n5370) );
  NAND2_X1 U6910 ( .A1(n5371), .A2(n5370), .ZN(n5373) );
  NAND2_X1 U6911 ( .A1(n9755), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6912 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5831) );
  OAI211_X1 U6913 ( .C1(n5373), .C2(n9753), .A(n5372), .B(n5831), .ZN(n5377)
         );
  AOI211_X1 U6914 ( .C1(n4373), .C2(n5375), .A(n5374), .B(n9449), .ZN(n5376)
         );
  AOI211_X1 U6915 ( .C1(n9456), .C2(n5378), .A(n5377), .B(n5376), .ZN(n5379)
         );
  INV_X1 U6916 ( .A(n5379), .ZN(P2_U3250) );
  INV_X1 U6917 ( .A(n9693), .ZN(n9720) );
  NAND2_X1 U6918 ( .A1(n5381), .A2(n5383), .ZN(n5869) );
  OAI21_X1 U6919 ( .B1(n5383), .B2(n5381), .A(n5869), .ZN(n5390) );
  INV_X1 U6920 ( .A(n5390), .ZN(n9640) );
  OR2_X1 U6921 ( .A1(n9652), .A2(n8946), .ZN(n9295) );
  OAI211_X1 U6922 ( .C1(n8701), .C2(n5382), .A(n9625), .B(n5922), .ZN(n9637)
         );
  OAI21_X1 U6923 ( .B1(n5382), .B2(n9723), .A(n9637), .ZN(n5391) );
  INV_X1 U6924 ( .A(n5383), .ZN(n8887) );
  XNOR2_X1 U6925 ( .A(n8887), .B(n8886), .ZN(n5386) );
  NAND2_X1 U6926 ( .A1(n8952), .A2(n9638), .ZN(n5385) );
  NAND2_X1 U6927 ( .A1(n8917), .A2(n8946), .ZN(n5384) );
  INV_X1 U6928 ( .A(n9289), .ZN(n9617) );
  NAND2_X1 U6929 ( .A1(n5386), .A2(n9617), .ZN(n5389) );
  OR2_X1 U6930 ( .A1(n5219), .A2(n8949), .ZN(n9293) );
  INV_X1 U6931 ( .A(n5219), .ZN(n5387) );
  AOI22_X1 U6932 ( .A1(n8971), .A2(n9649), .B1(n9614), .B2(n8702), .ZN(n5388)
         );
  OAI211_X1 U6933 ( .C1(n5390), .C2(n9323), .A(n5389), .B(n5388), .ZN(n9632)
         );
  AOI211_X1 U6934 ( .C1(n9720), .C2(n9640), .A(n5391), .B(n9632), .ZN(n9674)
         );
  NOR2_X1 U6935 ( .A1(n5392), .A2(n9393), .ZN(n5393) );
  AND2_X2 U6936 ( .A1(n9396), .A2(n5393), .ZN(n9748) );
  NAND2_X1 U6937 ( .A1(n9745), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5394) );
  OAI21_X1 U6938 ( .B1(n9674), .B2(n9745), .A(n5394), .ZN(P1_U3524) );
  INV_X1 U6939 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5395) );
  XNOR2_X1 U6940 ( .A(n6016), .B(n5395), .ZN(n5399) );
  NAND2_X1 U6941 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  NAND2_X1 U6942 ( .A1(n5399), .A2(n5398), .ZN(n5674) );
  OAI21_X1 U6943 ( .B1(n5399), .B2(n5398), .A(n5674), .ZN(n5402) );
  NAND2_X1 U6944 ( .A1(n9755), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6945 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n5400) );
  OAI211_X1 U6946 ( .C1(n5402), .C2(n9753), .A(n5401), .B(n5400), .ZN(n5408)
         );
  AOI21_X1 U6947 ( .B1(n5404), .B2(P2_REG2_REG_6__SCAN_IN), .A(n5403), .ZN(
        n5406) );
  XNOR2_X1 U6948 ( .A(n6016), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n5405) );
  NOR2_X1 U6949 ( .A1(n5405), .A2(n5406), .ZN(n5679) );
  AOI211_X1 U6950 ( .C1(n5406), .C2(n5405), .A(n5679), .B(n9449), .ZN(n5407)
         );
  AOI211_X1 U6951 ( .C1(n9456), .C2(n6016), .A(n5408), .B(n5407), .ZN(n5409)
         );
  INV_X1 U6952 ( .A(n5409), .ZN(P2_U3252) );
  NAND2_X1 U6953 ( .A1(n5411), .A2(n5410), .ZN(n5413) );
  AND2_X2 U6954 ( .A1(n5413), .A2(n5412), .ZN(n5508) );
  AND4_X2 U6955 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n6121)
         );
  OR2_X1 U6956 ( .A1(n5513), .A2(n5418), .ZN(n5419) );
  OAI211_X2 U6957 ( .C1(n5846), .C2(n9006), .A(n5420), .B(n5419), .ZN(n5923)
         );
  OAI22_X1 U6958 ( .A1(n6121), .A2(n7318), .B1(n9677), .B2(n7319), .ZN(n5421)
         );
  XNOR2_X1 U6959 ( .A(n5421), .B(n5653), .ZN(n5511) );
  NAND2_X1 U6960 ( .A1(n5923), .A2(n4285), .ZN(n5422) );
  NAND2_X1 U6961 ( .A1(n5423), .A2(n5422), .ZN(n5509) );
  XNOR2_X1 U6962 ( .A(n5511), .B(n5509), .ZN(n5507) );
  XNOR2_X1 U6963 ( .A(n5508), .B(n5507), .ZN(n5434) );
  NAND2_X1 U6964 ( .A1(n8671), .A2(n5923), .ZN(n5431) );
  NAND2_X1 U6965 ( .A1(n8678), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5429) );
  OR2_X1 U6966 ( .A1(n4280), .A2(n5424), .ZN(n5428) );
  OR2_X1 U6967 ( .A1(n5425), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5426) );
  AOI22_X1 U6968 ( .A1(n8653), .A2(n8970), .B1(n8666), .B2(n5380), .ZN(n5430)
         );
  OAI211_X1 U6969 ( .C1(n5432), .C2(n8997), .A(n5431), .B(n5430), .ZN(n5433)
         );
  AOI21_X1 U6970 ( .B1(n5434), .B2(n8657), .A(n5433), .ZN(n5435) );
  INV_X1 U6971 ( .A(n5435), .ZN(P1_U3235) );
  AND3_X1 U6972 ( .A1(n5634), .A2(n5436), .A3(n5637), .ZN(n5437) );
  INV_X1 U6973 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5440) );
  INV_X1 U6974 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5442) );
  INV_X1 U6975 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5445) );
  INV_X1 U6976 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6977 ( .A1(n5468), .A2(n7550), .ZN(n5986) );
  XNOR2_X1 U6978 ( .A(n5986), .B(n7738), .ZN(n8336) );
  NAND2_X1 U6979 ( .A1(n8336), .A2(n8375), .ZN(n9781) );
  NOR2_X1 U6980 ( .A1(n8375), .A2(n7738), .ZN(n5449) );
  INV_X1 U6981 ( .A(n9892), .ZN(n8500) );
  NAND2_X1 U6982 ( .A1(n9781), .A2(n8500), .ZN(n9907) );
  INV_X1 U6983 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6265) );
  OR2_X1 U6984 ( .A1(n4278), .A2(n6265), .ZN(n5454) );
  OR2_X2 U6985 ( .A1(n7797), .A2(n5451), .ZN(n5580) );
  INV_X1 U6986 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6262) );
  OR2_X2 U6987 ( .A1(n4279), .A2(n6262), .ZN(n5453) );
  NAND2_X1 U6988 ( .A1(n6027), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5452) );
  NAND4_X4 U6989 ( .A1(n5455), .A2(n5454), .A3(n5453), .A4(n5452), .ZN(n5545)
         );
  NAND2_X1 U6990 ( .A1(n6027), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5464) );
  OR2_X1 U6991 ( .A1(n4277), .A2(n6151), .ZN(n5463) );
  INV_X1 U6992 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5460) );
  OR2_X1 U6993 ( .A1(n4279), .A2(n5460), .ZN(n5462) );
  NAND2_X1 U6994 ( .A1(n4968), .A2(SI_0_), .ZN(n5465) );
  XNOR2_X1 U6995 ( .A(n5465), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8527) );
  MUX2_X1 U6996 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8527), .S(n5466), .Z(n6150) );
  INV_X1 U6997 ( .A(n6150), .ZN(n9843) );
  NAND2_X1 U6998 ( .A1(n5470), .A2(n5467), .ZN(n5746) );
  OAI21_X1 U6999 ( .B1(n5470), .B2(n5467), .A(n5746), .ZN(n6270) );
  OAI21_X1 U7000 ( .B1(n9843), .B2(n6266), .A(n6525), .ZN(n6267) );
  NAND2_X1 U7001 ( .A1(n6642), .A2(n7727), .ZN(n9844) );
  INV_X1 U7002 ( .A(n9844), .ZN(n5469) );
  NAND2_X1 U7003 ( .A1(n5544), .A2(n5469), .ZN(n9900) );
  OAI22_X1 U7004 ( .A1(n6267), .A2(n9902), .B1(n9900), .B2(n6266), .ZN(n5481)
         );
  NAND2_X1 U7005 ( .A1(n5786), .A2(n6150), .ZN(n6149) );
  XNOR2_X1 U7006 ( .A(n5470), .B(n6149), .ZN(n5471) );
  OR2_X1 U7007 ( .A1(n5468), .A2(n7727), .ZN(n7543) );
  INV_X1 U7008 ( .A(n5542), .ZN(n7547) );
  NAND2_X1 U7009 ( .A1(n5471), .A2(n9776), .ZN(n5480) );
  INV_X1 U7010 ( .A(n5786), .ZN(n7942) );
  INV_X1 U7011 ( .A(n5310), .ZN(n5472) );
  AND2_X2 U7012 ( .A1(n5485), .A2(n5472), .ZN(n9772) );
  OR2_X1 U7013 ( .A1(n5472), .A2(n5578), .ZN(n8384) );
  NAND2_X1 U7014 ( .A1(n6027), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5478) );
  OR2_X1 U7015 ( .A1(n4278), .A2(n5473), .ZN(n5477) );
  INV_X1 U7016 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5474) );
  OR2_X1 U7017 ( .A1(n4279), .A2(n5474), .ZN(n5476) );
  INV_X1 U7018 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9913) );
  OR2_X1 U7019 ( .A1(n6985), .A2(n9913), .ZN(n5475) );
  AOI22_X1 U7020 ( .A1(n7942), .A2(n9772), .B1(n9769), .B2(n7940), .ZN(n5479)
         );
  NAND2_X1 U7021 ( .A1(n5480), .A2(n5479), .ZN(n6261) );
  AOI211_X1 U7022 ( .C1(n9907), .C2(n6270), .A(n5481), .B(n6261), .ZN(n5600)
         );
  NAND2_X1 U7023 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  AOI21_X1 U7024 ( .B1(n5544), .B2(n5485), .A(n5484), .ZN(n5592) );
  NAND2_X1 U7025 ( .A1(n5592), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5606) );
  NOR4_X1 U7026 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5494) );
  INV_X1 U7027 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9833) );
  INV_X1 U7028 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9806) );
  INV_X1 U7029 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9822) );
  INV_X1 U7030 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9836) );
  NAND4_X1 U7031 ( .A1(n9833), .A2(n9806), .A3(n9822), .A4(n9836), .ZN(n5491)
         );
  NOR4_X1 U7032 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5489) );
  NOR4_X1 U7033 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5488) );
  NOR4_X1 U7034 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5487) );
  NOR4_X1 U7035 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5486) );
  NAND4_X1 U7036 ( .A1(n5489), .A2(n5488), .A3(n5487), .A4(n5486), .ZN(n5490)
         );
  NOR4_X1 U7037 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        n5491), .A4(n5490), .ZN(n5493) );
  NOR4_X1 U7038 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5492) );
  NAND3_X1 U7039 ( .A1(n5494), .A2(n5493), .A3(n5492), .ZN(n5497) );
  XNOR2_X1 U7040 ( .A(n6811), .B(P2_B_REG_SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7041 ( .A1(n6906), .A2(n5495), .ZN(n5496) );
  AND2_X1 U7042 ( .A1(n5497), .A2(n9803), .ZN(n5575) );
  NAND2_X1 U7043 ( .A1(n9892), .A2(n7727), .ZN(n5598) );
  INV_X1 U7044 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7045 ( .A1(n9803), .A2(n5498), .ZN(n5500) );
  OR2_X1 U7046 ( .A1(n5502), .A2(n5499), .ZN(n9837) );
  NAND2_X1 U7047 ( .A1(n5500), .A2(n9837), .ZN(n5982) );
  INV_X1 U7048 ( .A(n5982), .ZN(n5504) );
  INV_X1 U7049 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7050 ( .A1(n9803), .A2(n5501), .ZN(n5503) );
  INV_X1 U7051 ( .A(n5502), .ZN(n6920) );
  NAND2_X1 U7052 ( .A1(n6920), .A2(n6906), .ZN(n9839) );
  NAND2_X1 U7053 ( .A1(n5503), .A2(n9839), .ZN(n5981) );
  NAND3_X1 U7054 ( .A1(n5598), .A2(n5504), .A3(n5981), .ZN(n5505) );
  NAND2_X1 U7055 ( .A1(n9925), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5506) );
  OAI21_X1 U7056 ( .B1(n5600), .B2(n9925), .A(n5506), .ZN(P2_U3521) );
  INV_X1 U7057 ( .A(n5509), .ZN(n5510) );
  NAND2_X1 U7058 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  NAND2_X1 U7059 ( .A1(n8970), .A2(n7290), .ZN(n5519) );
  OR2_X1 U7060 ( .A1(n6051), .A2(n5571), .ZN(n5517) );
  OR2_X1 U7061 ( .A1(n5513), .A2(n5514), .ZN(n5516) );
  OR2_X1 U7062 ( .A1(n5846), .A2(n9421), .ZN(n5515) );
  OR2_X1 U7063 ( .A1(n9683), .A2(n7319), .ZN(n5518) );
  NAND2_X1 U7064 ( .A1(n5519), .A2(n5518), .ZN(n5520) );
  XNOR2_X1 U7065 ( .A(n5520), .B(n5653), .ZN(n5652) );
  NAND2_X1 U7066 ( .A1(n8970), .A2(n7286), .ZN(n5522) );
  OR2_X1 U7067 ( .A1(n9683), .A2(n7318), .ZN(n5521) );
  NAND2_X1 U7068 ( .A1(n5522), .A2(n5521), .ZN(n5650) );
  XNOR2_X1 U7069 ( .A(n5652), .B(n5650), .ZN(n5648) );
  XOR2_X1 U7070 ( .A(n5648), .B(n5649), .Z(n5541) );
  INV_X1 U7071 ( .A(n9683), .ZN(n6116) );
  INV_X1 U7072 ( .A(n8666), .ZN(n8650) );
  INV_X1 U7073 ( .A(n5523), .ZN(n5524) );
  AOI21_X1 U7074 ( .B1(n5525), .B2(n5524), .A(P1_U3084), .ZN(n5526) );
  INV_X1 U7075 ( .A(n4275), .ZN(n8576) );
  INV_X1 U7076 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9420) );
  NAND2_X1 U7077 ( .A1(n8576), .A2(n9420), .ZN(n5538) );
  INV_X1 U7078 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5529) );
  OR2_X1 U7079 ( .A1(n5528), .A2(n5529), .ZN(n5535) );
  INV_X1 U7080 ( .A(n5663), .ZN(n5532) );
  INV_X1 U7081 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7082 ( .A1(n9420), .A2(n5530), .ZN(n5531) );
  NAND2_X1 U7083 ( .A1(n5532), .A2(n5531), .ZN(n5896) );
  OR2_X1 U7084 ( .A1(n7167), .A2(n5896), .ZN(n5534) );
  OR2_X1 U7085 ( .A1(n4280), .A2(n8220), .ZN(n5533) );
  INV_X1 U7086 ( .A(n6120), .ZN(n8969) );
  AOI22_X1 U7087 ( .A1(n8653), .A2(n8969), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3084), .ZN(n5537) );
  OAI211_X1 U7088 ( .C1(n6121), .C2(n8650), .A(n5538), .B(n5537), .ZN(n5539)
         );
  AOI21_X1 U7089 ( .B1(n8671), .B2(n6116), .A(n5539), .ZN(n5540) );
  OAI21_X1 U7090 ( .B1(n5541), .B2(n8645), .A(n5540), .ZN(P1_U3216) );
  NAND3_X1 U7091 ( .A1(n5542), .A2(n7727), .A3(n9844), .ZN(n5543) );
  NAND2_X1 U7092 ( .A1(n5560), .A2(n5545), .ZN(n5547) );
  NAND2_X1 U7093 ( .A1(n5546), .A2(n5547), .ZN(n5552) );
  INV_X1 U7094 ( .A(n5546), .ZN(n5549) );
  INV_X1 U7095 ( .A(n5547), .ZN(n5548) );
  NAND2_X1 U7096 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U7097 ( .A1(n5552), .A2(n5550), .ZN(n5604) );
  NOR2_X1 U7098 ( .A1(n5725), .A2(n5786), .ZN(n5551) );
  MUX2_X1 U7099 ( .A(n6486), .B(n5551), .S(n6150), .Z(n5605) );
  INV_X1 U7100 ( .A(n5552), .ZN(n5553) );
  NOR2_X1 U7101 ( .A1(n5603), .A2(n5553), .ZN(n5793) );
  OR2_X1 U7102 ( .A1(n5718), .A2(n5555), .ZN(n5558) );
  XNOR2_X1 U7103 ( .A(n5554), .B(n6526), .ZN(n5562) );
  NAND2_X1 U7104 ( .A1(n5560), .A2(n7940), .ZN(n5561) );
  XNOR2_X1 U7105 ( .A(n5562), .B(n5561), .ZN(n5792) );
  INV_X1 U7106 ( .A(n5561), .ZN(n5563) );
  AOI22_X1 U7107 ( .A1(n5793), .A2(n5792), .B1(n5563), .B2(n5562), .ZN(n5716)
         );
  NAND2_X1 U7108 ( .A1(n5450), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5570) );
  INV_X1 U7109 ( .A(n6027), .ZN(n7392) );
  INV_X1 U7110 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5564) );
  OR2_X1 U7111 ( .A1(n7392), .A2(n5564), .ZN(n5569) );
  OR2_X1 U7112 ( .A1(n4279), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5568) );
  INV_X1 U7113 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5565) );
  OR2_X1 U7114 ( .A1(n4277), .A2(n5565), .ZN(n5567) );
  NAND4_X1 U7115 ( .A1(n5570), .A2(n5569), .A3(n5568), .A4(n5567), .ZN(n7939)
         );
  NAND2_X1 U7116 ( .A1(n5560), .A2(n7939), .ZN(n5713) );
  OR2_X1 U7117 ( .A1(n6015), .A2(n5571), .ZN(n5573) );
  XNOR2_X1 U7118 ( .A(n5554), .B(n5798), .ZN(n5712) );
  XOR2_X1 U7119 ( .A(n5713), .B(n5712), .Z(n5715) );
  XNOR2_X1 U7120 ( .A(n5716), .B(n5715), .ZN(n5597) );
  NOR2_X1 U7121 ( .A1(n5982), .A2(n5981), .ZN(n5577) );
  INV_X1 U7122 ( .A(n5575), .ZN(n5576) );
  AND2_X1 U7123 ( .A1(n5577), .A2(n5576), .ZN(n5590) );
  AND2_X1 U7124 ( .A1(n9900), .A2(n5578), .ZN(n5579) );
  INV_X1 U7125 ( .A(n5544), .ZN(n7735) );
  NAND2_X1 U7126 ( .A1(n5587), .A2(n7735), .ZN(n7792) );
  INV_X1 U7127 ( .A(n7792), .ZN(n7924) );
  NAND2_X1 U7128 ( .A1(n6027), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7129 ( .A1(n5450), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5583) );
  OAI21_X1 U7130 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5734), .ZN(n5741) );
  OR2_X1 U7131 ( .A1(n4279), .A2(n5741), .ZN(n5582) );
  OR2_X1 U7132 ( .A1(n4277), .A2(n8206), .ZN(n5581) );
  NAND4_X1 U7133 ( .A1(n5584), .A2(n5583), .A3(n5582), .A4(n5581), .ZN(n7938)
         );
  INV_X1 U7134 ( .A(n7938), .ZN(n5586) );
  INV_X1 U7135 ( .A(n7940), .ZN(n5585) );
  INV_X1 U7136 ( .A(n9772), .ZN(n8386) );
  OAI22_X1 U7137 ( .A1(n5586), .A2(n8384), .B1(n5585), .B2(n8386), .ZN(n5753)
         );
  AOI22_X1 U7138 ( .A1(n7924), .A2(n5753), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n5596) );
  NOR2_X1 U7139 ( .A1(n5468), .A2(n9844), .ZN(n5997) );
  NAND2_X1 U7140 ( .A1(n5587), .A2(n5997), .ZN(n5589) );
  INV_X1 U7141 ( .A(n5590), .ZN(n5591) );
  NAND2_X1 U7142 ( .A1(n5598), .A2(n5591), .ZN(n5607) );
  NAND2_X1 U7143 ( .A1(n5607), .A2(n5592), .ZN(n5593) );
  INV_X1 U7144 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5594) );
  AOI22_X1 U7145 ( .A1(n5798), .A2(n7903), .B1(n7885), .B2(n5594), .ZN(n5595)
         );
  OAI211_X1 U7146 ( .C1(n5597), .C2(n7913), .A(n5596), .B(n5595), .ZN(P2_U3220) );
  NAND3_X1 U7147 ( .A1(n5598), .A2(n5982), .A3(n5981), .ZN(n5599) );
  INV_X2 U7148 ( .A(n9908), .ZN(n9910) );
  INV_X1 U7149 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5602) );
  OR2_X1 U7150 ( .A1(n5600), .A2(n9908), .ZN(n5601) );
  OAI21_X1 U7151 ( .B1(n9910), .B2(n5602), .A(n5601), .ZN(P2_U3454) );
  AOI21_X1 U7152 ( .B1(n5605), .B2(n5604), .A(n5603), .ZN(n5611) );
  INV_X1 U7153 ( .A(n5606), .ZN(n5608) );
  NAND2_X1 U7154 ( .A1(n5608), .A2(n5607), .ZN(n5794) );
  AOI22_X1 U7155 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n5794), .B1(n7903), .B2(
        n5459), .ZN(n5610) );
  NAND2_X1 U7156 ( .A1(n7924), .A2(n9772), .ZN(n7892) );
  INV_X1 U7157 ( .A(n7892), .ZN(n7909) );
  NOR2_X1 U7158 ( .A1(n7792), .A2(n8384), .ZN(n7905) );
  AOI22_X1 U7159 ( .A1(n7909), .A2(n7942), .B1(n7905), .B2(n7940), .ZN(n5609)
         );
  OAI211_X1 U7160 ( .C1(n5611), .C2(n7913), .A(n5610), .B(n5609), .ZN(P2_U3224) );
  INV_X1 U7161 ( .A(n5612), .ZN(n5613) );
  INV_X1 U7162 ( .A(n5615), .ZN(n5616) );
  NAND2_X1 U7163 ( .A1(n5616), .A2(SI_14_), .ZN(n5617) );
  INV_X1 U7164 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6969) );
  INV_X1 U7165 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5633) );
  MUX2_X1 U7166 ( .A(n6969), .B(n5633), .S(n7532), .Z(n5619) );
  INV_X1 U7167 ( .A(SI_15_), .ZN(n5618) );
  INV_X1 U7168 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U7169 ( .A1(n5620), .A2(SI_15_), .ZN(n5621) );
  INV_X1 U7170 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5623) );
  INV_X1 U7171 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5643) );
  MUX2_X1 U7172 ( .A(n5623), .B(n5643), .S(n7532), .Z(n5625) );
  INV_X1 U7173 ( .A(SI_16_), .ZN(n5624) );
  NAND2_X1 U7174 ( .A1(n5625), .A2(n5624), .ZN(n5688) );
  INV_X1 U7175 ( .A(n5625), .ZN(n5626) );
  NAND2_X1 U7176 ( .A1(n5626), .A2(SI_16_), .ZN(n5627) );
  XNOR2_X1 U7177 ( .A(n5687), .B(n5686), .ZN(n7080) );
  INV_X1 U7178 ( .A(n7080), .ZN(n5644) );
  OR2_X1 U7179 ( .A1(n5628), .A2(n8522), .ZN(n5629) );
  XNOR2_X1 U7180 ( .A(n5629), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7972) );
  AOI22_X1 U7181 ( .A1(n7972), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8525), .ZN(n5630) );
  OAI21_X1 U7182 ( .B1(n5644), .B2(n7800), .A(n5630), .ZN(P2_U3342) );
  XNOR2_X1 U7183 ( .A(n5632), .B(n5631), .ZN(n6968) );
  INV_X1 U7184 ( .A(n6968), .ZN(n5639) );
  OAI222_X1 U7185 ( .A1(n7361), .A2(n5633), .B1(n7364), .B2(n5639), .C1(
        P1_U3084), .C2(n9048), .ZN(P1_U3338) );
  NAND2_X1 U7186 ( .A1(n5635), .A2(n5634), .ZN(n5636) );
  NAND2_X1 U7187 ( .A1(n5636), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5638) );
  XNOR2_X1 U7188 ( .A(n5638), .B(n5637), .ZN(n7953) );
  OAI222_X1 U7189 ( .A1(n7817), .A2(n6969), .B1(n7800), .B2(n5639), .C1(n7953), 
        .C2(P2_U3152), .ZN(P2_U3343) );
  NAND2_X1 U7190 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  NAND2_X1 U7191 ( .A1(n5642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5692) );
  XNOR2_X1 U7192 ( .A(n5692), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9064) );
  INV_X1 U7193 ( .A(n9064), .ZN(n9056) );
  OAI222_X1 U7194 ( .A1(n9417), .A2(n5644), .B1(n9056), .B2(P1_U3084), .C1(
        n5643), .C2(n7361), .ZN(P1_U3337) );
  OR2_X1 U7195 ( .A1(n5513), .A2(n5645), .ZN(n5647) );
  OR2_X1 U7196 ( .A1(n6051), .A2(n5717), .ZN(n5646) );
  OAI211_X1 U7197 ( .C1(n5846), .C2(n9017), .A(n5647), .B(n5646), .ZN(n9690)
         );
  INV_X1 U7198 ( .A(n5650), .ZN(n5651) );
  OAI22_X1 U7199 ( .A1(n6120), .A2(n7318), .B1(n5901), .B2(n7319), .ZN(n5654)
         );
  XNOR2_X1 U7200 ( .A(n5654), .B(n7320), .ZN(n5763) );
  OR2_X1 U7201 ( .A1(n6120), .A2(n7322), .ZN(n5656) );
  NAND2_X1 U7202 ( .A1(n9690), .A2(n4285), .ZN(n5655) );
  NAND2_X1 U7203 ( .A1(n5656), .A2(n5655), .ZN(n5762) );
  XNOR2_X1 U7204 ( .A(n5763), .B(n5762), .ZN(n5658) );
  AOI21_X1 U7205 ( .B1(n5657), .B2(n5658), .A(n8645), .ZN(n5661) );
  INV_X1 U7206 ( .A(n5657), .ZN(n5660) );
  NAND2_X1 U7207 ( .A1(n5660), .A2(n5659), .ZN(n5840) );
  NAND2_X1 U7208 ( .A1(n5661), .A2(n5840), .ZN(n5672) );
  NAND2_X1 U7209 ( .A1(n8678), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5668) );
  OR2_X1 U7210 ( .A1(n4280), .A2(n5662), .ZN(n5667) );
  OAI21_X1 U7211 ( .B1(n5663), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5775), .ZN(
        n5911) );
  OR2_X1 U7212 ( .A1(n7167), .A2(n5911), .ZN(n5666) );
  OR2_X1 U7213 ( .A1(n8683), .A2(n5664), .ZN(n5665) );
  NAND4_X1 U7214 ( .A1(n5668), .A2(n5667), .A3(n5666), .A4(n5665), .ZN(n8968)
         );
  INV_X1 U7215 ( .A(n8968), .ZN(n6214) );
  NAND2_X1 U7216 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n9023) );
  OAI21_X1 U7217 ( .B1(n8664), .B2(n6214), .A(n9023), .ZN(n5670) );
  NOR2_X1 U7218 ( .A1(n4275), .A2(n5896), .ZN(n5669) );
  AOI211_X1 U7219 ( .C1(n8666), .C2(n8970), .A(n5670), .B(n5669), .ZN(n5671)
         );
  OAI211_X1 U7220 ( .C1(n5901), .C2(n8656), .A(n5672), .B(n5671), .ZN(P1_U3228) );
  INV_X1 U7221 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9918) );
  MUX2_X1 U7222 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9918), .S(n6134), .Z(n5676)
         );
  NAND2_X1 U7223 ( .A1(n6016), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7224 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  NAND2_X1 U7225 ( .A1(n5675), .A2(n5676), .ZN(n5967) );
  OAI21_X1 U7226 ( .B1(n5676), .B2(n5675), .A(n5967), .ZN(n5678) );
  NAND2_X1 U7227 ( .A1(n9755), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7228 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6144) );
  OAI211_X1 U7229 ( .C1(n9753), .C2(n5678), .A(n5677), .B(n6144), .ZN(n5684)
         );
  NAND2_X1 U7230 ( .A1(n6134), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5680) );
  OAI21_X1 U7231 ( .B1(n6134), .B2(P2_REG2_REG_8__SCAN_IN), .A(n5680), .ZN(
        n5681) );
  NOR2_X1 U7232 ( .A1(n5682), .A2(n5681), .ZN(n5973) );
  AOI211_X1 U7233 ( .C1(n5682), .C2(n5681), .A(n5973), .B(n9449), .ZN(n5683)
         );
  AOI211_X1 U7234 ( .C1(n9456), .C2(n6134), .A(n5684), .B(n5683), .ZN(n5685)
         );
  INV_X1 U7235 ( .A(n5685), .ZN(P2_U3253) );
  INV_X1 U7236 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5690) );
  INV_X1 U7237 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5689) );
  MUX2_X1 U7238 ( .A(n5690), .B(n5689), .S(n7532), .Z(n5945) );
  XNOR2_X1 U7239 ( .A(n5945), .B(SI_17_), .ZN(n5944) );
  XNOR2_X1 U7240 ( .A(n5947), .B(n5944), .ZN(n7076) );
  INV_X1 U7241 ( .A(n7076), .ZN(n5698) );
  NAND2_X1 U7242 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  NAND2_X1 U7243 ( .A1(n5693), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U7244 ( .A(n5949), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9077) );
  AOI22_X1 U7245 ( .A1(n9077), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6945), .ZN(n5694) );
  OAI21_X1 U7246 ( .B1(n5698), .B2(n9417), .A(n5694), .ZN(P1_U3336) );
  NAND2_X1 U7247 ( .A1(n5695), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5696) );
  XNOR2_X1 U7248 ( .A(n5696), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7985) );
  AOI22_X1 U7249 ( .A1(n7985), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8525), .ZN(n5697) );
  OAI21_X1 U7250 ( .B1(n5698), .B2(n7800), .A(n5697), .ZN(P2_U3341) );
  OAI21_X1 U7251 ( .B1(n5701), .B2(n5700), .A(n5699), .ZN(n5710) );
  NAND2_X1 U7252 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n5703) );
  NAND2_X1 U7253 ( .A1(n9564), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n5702) );
  OAI211_X1 U7254 ( .C1(n9422), .C2(n5704), .A(n5703), .B(n5702), .ZN(n5709)
         );
  AOI211_X1 U7255 ( .C1(n5707), .C2(n5706), .A(n5705), .B(n9571), .ZN(n5708)
         );
  AOI211_X1 U7256 ( .C1(n9587), .C2(n5710), .A(n5709), .B(n5708), .ZN(n5711)
         );
  INV_X1 U7257 ( .A(n5711), .ZN(P1_U3253) );
  INV_X1 U7258 ( .A(n5712), .ZN(n5714) );
  OAI22_X1 U7259 ( .A1(n5716), .A2(n5715), .B1(n5714), .B2(n5713), .ZN(n5729)
         );
  OR2_X1 U7260 ( .A1(n6015), .A2(n5717), .ZN(n5724) );
  OR2_X1 U7261 ( .A1(n4287), .A2(n5719), .ZN(n5723) );
  NAND2_X1 U7262 ( .A1(n5720), .A2(n5721), .ZN(n5722) );
  XNOR2_X1 U7263 ( .A(n5554), .B(n5801), .ZN(n5727) );
  NAND2_X1 U7264 ( .A1(n5560), .A2(n7938), .ZN(n5726) );
  NAND2_X1 U7265 ( .A1(n5727), .A2(n5726), .ZN(n5814) );
  OAI21_X1 U7266 ( .B1(n5727), .B2(n5726), .A(n5814), .ZN(n5728) );
  AOI21_X1 U7267 ( .B1(n5729), .B2(n5728), .A(n5816), .ZN(n5744) );
  NAND2_X1 U7268 ( .A1(n6027), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5740) );
  INV_X1 U7269 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5730) );
  OR2_X1 U7270 ( .A1(n4278), .A2(n5730), .ZN(n5739) );
  INV_X1 U7271 ( .A(n5734), .ZN(n5732) );
  NAND2_X1 U7272 ( .A1(n5732), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5822) );
  INV_X1 U7273 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7274 ( .A1(n5734), .A2(n5733), .ZN(n5735) );
  NAND2_X1 U7275 ( .A1(n5822), .A2(n5735), .ZN(n5995) );
  INV_X1 U7276 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5736) );
  OR2_X1 U7277 ( .A1(n6985), .A2(n5736), .ZN(n5737) );
  OAI22_X1 U7278 ( .A1(n4632), .A2(n8384), .B1(n4401), .B2(n8386), .ZN(n5806)
         );
  AOI22_X1 U7279 ( .A1(n7924), .A2(n5806), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n5743) );
  INV_X1 U7280 ( .A(n5741), .ZN(n6196) );
  AOI22_X1 U7281 ( .A1(n6198), .A2(n7903), .B1(n7885), .B2(n6196), .ZN(n5742)
         );
  OAI211_X1 U7282 ( .C1(n5744), .C2(n7913), .A(n5743), .B(n5742), .ZN(P2_U3232) );
  OR2_X1 U7283 ( .A1(n5545), .A2(n5459), .ZN(n5745) );
  NAND2_X1 U7284 ( .A1(n5746), .A2(n5745), .ZN(n6522) );
  OR2_X1 U7285 ( .A1(n7940), .A2(n9850), .ZN(n7557) );
  NAND2_X1 U7286 ( .A1(n6522), .A2(n6527), .ZN(n6523) );
  OR2_X1 U7287 ( .A1(n7940), .A2(n6526), .ZN(n5747) );
  NAND2_X1 U7288 ( .A1(n6523), .A2(n5747), .ZN(n5748) );
  NAND2_X1 U7289 ( .A1(n7939), .A2(n9796), .ZN(n7573) );
  NAND2_X1 U7290 ( .A1(n5748), .A2(n7700), .ZN(n5800) );
  OAI21_X1 U7291 ( .B1(n5748), .B2(n7700), .A(n5800), .ZN(n5754) );
  INV_X1 U7292 ( .A(n5754), .ZN(n9797) );
  INV_X1 U7293 ( .A(n9781), .ZN(n5755) );
  INV_X1 U7294 ( .A(n7700), .ZN(n7563) );
  NAND2_X1 U7295 ( .A1(n6149), .A2(n7556), .ZN(n7551) );
  NAND2_X1 U7296 ( .A1(n7551), .A2(n7554), .ZN(n6530) );
  NAND2_X1 U7297 ( .A1(n6530), .A2(n7557), .ZN(n6528) );
  NAND2_X1 U7298 ( .A1(n6528), .A2(n7698), .ZN(n5750) );
  NAND2_X1 U7299 ( .A1(n5750), .A2(n7700), .ZN(n5751) );
  AOI21_X1 U7300 ( .B1(n5804), .B2(n5751), .A(n8371), .ZN(n5752) );
  AOI211_X1 U7301 ( .C1(n5755), .C2(n5754), .A(n5753), .B(n5752), .ZN(n9802)
         );
  INV_X1 U7302 ( .A(n6524), .ZN(n5756) );
  AOI211_X1 U7303 ( .C1(n5798), .C2(n5756), .A(n9902), .B(n4428), .ZN(n9791)
         );
  AOI21_X1 U7304 ( .B1(n8489), .B2(n5798), .A(n9791), .ZN(n5757) );
  OAI211_X1 U7305 ( .C1(n9797), .C2(n8500), .A(n9802), .B(n5757), .ZN(n5759)
         );
  NAND2_X1 U7306 ( .A1(n5759), .A2(n9910), .ZN(n5758) );
  OAI21_X1 U7307 ( .B1(n9910), .B2(n5564), .A(n5758), .ZN(P2_U3460) );
  INV_X2 U7308 ( .A(n9925), .ZN(n9927) );
  INV_X1 U7309 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7310 ( .A1(n5759), .A2(n9927), .ZN(n5760) );
  OAI21_X1 U7311 ( .B1(n9927), .B2(n5761), .A(n5760), .ZN(P2_U3523) );
  NAND2_X1 U7312 ( .A1(n5763), .A2(n5762), .ZN(n5838) );
  NAND2_X1 U7313 ( .A1(n5840), .A2(n5838), .ZN(n5773) );
  NAND2_X1 U7314 ( .A1(n8968), .A2(n4285), .ZN(n5768) );
  OR2_X1 U7315 ( .A1(n5817), .A2(n6051), .ZN(n5765) );
  OR2_X1 U7316 ( .A1(n5513), .A2(n4508), .ZN(n5764) );
  OAI211_X1 U7317 ( .C1(n5846), .C2(n5766), .A(n5765), .B(n5764), .ZN(n6213)
         );
  NAND2_X1 U7318 ( .A1(n6213), .A2(n7289), .ZN(n5767) );
  NAND2_X1 U7319 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  XNOR2_X1 U7320 ( .A(n5769), .B(n7320), .ZN(n5841) );
  NAND2_X1 U7321 ( .A1(n8968), .A2(n7286), .ZN(n5771) );
  NAND2_X1 U7322 ( .A1(n6213), .A2(n4285), .ZN(n5770) );
  NAND2_X1 U7323 ( .A1(n5771), .A2(n5770), .ZN(n5836) );
  INV_X1 U7324 ( .A(n5836), .ZN(n5842) );
  XNOR2_X1 U7325 ( .A(n5841), .B(n5842), .ZN(n5772) );
  XNOR2_X1 U7326 ( .A(n5773), .B(n5772), .ZN(n5785) );
  NAND2_X1 U7327 ( .A1(n8678), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5780) );
  OR2_X1 U7328 ( .A1(n4280), .A2(n4930), .ZN(n5779) );
  AND2_X1 U7329 ( .A1(n5775), .A2(n5774), .ZN(n5776) );
  OR2_X1 U7330 ( .A1(n5776), .A2(n5856), .ZN(n6209) );
  OR2_X1 U7331 ( .A1(n7167), .A2(n6209), .ZN(n5778) );
  OR2_X1 U7332 ( .A1(n8683), .A2(n9739), .ZN(n5777) );
  NAND2_X1 U7333 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n9575) );
  OAI21_X1 U7334 ( .B1(n8664), .B2(n6274), .A(n9575), .ZN(n5781) );
  AOI21_X1 U7335 ( .B1(n8666), .B2(n8969), .A(n5781), .ZN(n5782) );
  OAI21_X1 U7336 ( .B1(n4275), .B2(n5911), .A(n5782), .ZN(n5783) );
  AOI21_X1 U7337 ( .B1(n8671), .B2(n6213), .A(n5783), .ZN(n5784) );
  OAI21_X1 U7338 ( .B1(n5785), .B2(n8645), .A(n5784), .ZN(P1_U3225) );
  AOI22_X1 U7339 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n5794), .B1(n7903), .B2(
        n6150), .ZN(n5791) );
  INV_X1 U7340 ( .A(n6149), .ZN(n5789) );
  OR2_X1 U7341 ( .A1(n5786), .A2(n6150), .ZN(n7555) );
  INV_X1 U7342 ( .A(n7555), .ZN(n5787) );
  MUX2_X1 U7343 ( .A(n6150), .B(n5787), .S(n5560), .Z(n5788) );
  OAI21_X1 U7344 ( .B1(n5789), .B2(n5788), .A(n7901), .ZN(n5790) );
  OAI211_X1 U7345 ( .C1(n7893), .C2(n5458), .A(n5791), .B(n5790), .ZN(P2_U3234) );
  XNOR2_X1 U7346 ( .A(n5793), .B(n5792), .ZN(n5797) );
  AOI22_X1 U7347 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(n5794), .B1(n7903), .B2(
        n6526), .ZN(n5796) );
  AOI22_X1 U7348 ( .A1(n7909), .A2(n5545), .B1(n7905), .B2(n7939), .ZN(n5795)
         );
  OAI211_X1 U7349 ( .C1(n5797), .C2(n7913), .A(n5796), .B(n5795), .ZN(P2_U3239) );
  OR2_X1 U7350 ( .A1(n7939), .A2(n5798), .ZN(n5799) );
  NAND2_X1 U7351 ( .A1(n5800), .A2(n5799), .ZN(n5802) );
  OR2_X1 U7352 ( .A1(n7938), .A2(n5801), .ZN(n7567) );
  NAND2_X1 U7353 ( .A1(n7938), .A2(n5801), .ZN(n7574) );
  NAND2_X1 U7354 ( .A1(n7567), .A2(n7574), .ZN(n5805) );
  NAND2_X1 U7355 ( .A1(n5802), .A2(n5805), .ZN(n5980) );
  OAI21_X1 U7356 ( .B1(n5802), .B2(n5805), .A(n5980), .ZN(n6202) );
  INV_X1 U7357 ( .A(n6202), .ZN(n5809) );
  INV_X1 U7358 ( .A(n5993), .ZN(n5994) );
  AOI211_X1 U7359 ( .C1(n6198), .C2(n5803), .A(n9902), .B(n5994), .ZN(n6197)
         );
  AOI21_X1 U7360 ( .B1(n8489), .B2(n6198), .A(n6197), .ZN(n5808) );
  NAND2_X1 U7361 ( .A1(n5804), .A2(n7566), .ZN(n5988) );
  INV_X1 U7362 ( .A(n5805), .ZN(n7702) );
  XNOR2_X1 U7363 ( .A(n5988), .B(n7702), .ZN(n5807) );
  AOI21_X1 U7364 ( .B1(n5807), .B2(n9776), .A(n5806), .ZN(n6204) );
  OAI211_X1 U7365 ( .C1(n5809), .C2(n8494), .A(n5808), .B(n6204), .ZN(n5811)
         );
  NAND2_X1 U7366 ( .A1(n5811), .A2(n9927), .ZN(n5810) );
  OAI21_X1 U7367 ( .B1(n9927), .B2(n5313), .A(n5810), .ZN(P2_U3524) );
  INV_X1 U7368 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7369 ( .A1(n5811), .A2(n9910), .ZN(n5812) );
  OAI21_X1 U7370 ( .B1(n9910), .B2(n5813), .A(n5812), .ZN(P2_U3463) );
  INV_X1 U7371 ( .A(n5814), .ZN(n5815) );
  OR2_X1 U7372 ( .A1(n4287), .A2(n5002), .ZN(n5818) );
  XNOR2_X1 U7373 ( .A(n5554), .B(n5998), .ZN(n6004) );
  NAND2_X1 U7374 ( .A1(n5560), .A2(n7937), .ZN(n6002) );
  XNOR2_X1 U7375 ( .A(n6004), .B(n6002), .ZN(n6005) );
  XNOR2_X1 U7376 ( .A(n6006), .B(n6005), .ZN(n5835) );
  NAND2_X1 U7377 ( .A1(n7938), .A2(n9772), .ZN(n5830) );
  NAND2_X1 U7378 ( .A1(n6027), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5828) );
  INV_X1 U7379 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6102) );
  OR2_X1 U7380 ( .A1(n4278), .A2(n6102), .ZN(n5827) );
  INV_X1 U7381 ( .A(n5822), .ZN(n5820) );
  NAND2_X1 U7382 ( .A1(n5820), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6021) );
  INV_X1 U7383 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7384 ( .A1(n5822), .A2(n5821), .ZN(n5823) );
  NAND2_X1 U7385 ( .A1(n6021), .A2(n5823), .ZN(n7907) );
  INV_X1 U7386 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5824) );
  OR2_X1 U7387 ( .A1(n6985), .A2(n5824), .ZN(n5825) );
  NAND2_X1 U7388 ( .A1(n7936), .A2(n9769), .ZN(n5829) );
  NAND2_X1 U7389 ( .A1(n5830), .A2(n5829), .ZN(n5990) );
  INV_X1 U7390 ( .A(n5831), .ZN(n5833) );
  INV_X1 U7391 ( .A(n7903), .ZN(n7927) );
  OAI22_X1 U7392 ( .A1(n9856), .A2(n7927), .B1(n7922), .B2(n5995), .ZN(n5832)
         );
  AOI211_X1 U7393 ( .C1(n7924), .C2(n5990), .A(n5833), .B(n5832), .ZN(n5834)
         );
  OAI21_X1 U7394 ( .B1(n5835), .B2(n7913), .A(n5834), .ZN(P2_U3229) );
  NAND2_X1 U7395 ( .A1(n5841), .A2(n5836), .ZN(n5837) );
  AND2_X1 U7396 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  NAND2_X1 U7397 ( .A1(n5840), .A2(n5839), .ZN(n5845) );
  INV_X1 U7398 ( .A(n5841), .ZN(n5843) );
  NAND2_X1 U7399 ( .A1(n5843), .A2(n5842), .ZN(n5844) );
  OR2_X1 U7400 ( .A1(n6007), .A2(n6051), .ZN(n5849) );
  AOI22_X1 U7401 ( .A1(n7086), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7085), .B2(
        n5847), .ZN(n5848) );
  NAND2_X1 U7402 ( .A1(n5849), .A2(n5848), .ZN(n6211) );
  NAND2_X1 U7403 ( .A1(n6211), .A2(n7289), .ZN(n5850) );
  OAI21_X1 U7404 ( .B1(n6274), .B2(n7283), .A(n5850), .ZN(n5851) );
  XNOR2_X1 U7405 ( .A(n5851), .B(n5653), .ZN(n6066) );
  INV_X1 U7406 ( .A(n6066), .ZN(n6069) );
  OR2_X1 U7407 ( .A1(n6274), .A2(n7322), .ZN(n5853) );
  NAND2_X1 U7408 ( .A1(n6211), .A2(n4285), .ZN(n5852) );
  NAND2_X1 U7409 ( .A1(n5853), .A2(n5852), .ZN(n6067) );
  XNOR2_X1 U7410 ( .A(n6069), .B(n6067), .ZN(n5854) );
  XNOR2_X1 U7411 ( .A(n6068), .B(n5854), .ZN(n5867) );
  NAND2_X1 U7412 ( .A1(n8678), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5861) );
  OR2_X1 U7413 ( .A1(n4280), .A2(n5855), .ZN(n5860) );
  OR2_X1 U7414 ( .A1(n5856), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7415 ( .A1(n6077), .A2(n5857), .ZN(n9618) );
  OR2_X1 U7416 ( .A1(n7167), .A2(n9618), .ZN(n5859) );
  OR2_X1 U7417 ( .A1(n8683), .A2(n9741), .ZN(n5858) );
  OAI21_X1 U7418 ( .B1(n8664), .B2(n6277), .A(n5862), .ZN(n5863) );
  AOI21_X1 U7419 ( .B1(n8666), .B2(n8968), .A(n5863), .ZN(n5864) );
  OAI21_X1 U7420 ( .B1(n4275), .B2(n6209), .A(n5864), .ZN(n5865) );
  AOI21_X1 U7421 ( .B1(n8671), .B2(n6211), .A(n5865), .ZN(n5866) );
  OAI21_X1 U7422 ( .B1(n5867), .B2(n8645), .A(n5866), .ZN(P1_U3237) );
  NAND2_X1 U7423 ( .A1(n6120), .A2(n9690), .ZN(n8711) );
  NAND2_X1 U7424 ( .A1(n5380), .A2(n9634), .ZN(n5868) );
  NAND2_X1 U7425 ( .A1(n5869), .A2(n5868), .ZN(n5920) );
  INV_X1 U7426 ( .A(n5920), .ZN(n5870) );
  NAND2_X1 U7427 ( .A1(n8971), .A2(n9677), .ZN(n8706) );
  NAND2_X1 U7428 ( .A1(n5886), .A2(n8706), .ZN(n5885) );
  NAND2_X1 U7429 ( .A1(n5870), .A2(n5885), .ZN(n5919) );
  NAND2_X1 U7430 ( .A1(n6121), .A2(n9677), .ZN(n5871) );
  NAND2_X1 U7431 ( .A1(n5919), .A2(n5871), .ZN(n6113) );
  NAND2_X1 U7432 ( .A1(n6113), .A2(n8889), .ZN(n5873) );
  INV_X1 U7433 ( .A(n8970), .ZN(n5888) );
  NAND2_X1 U7434 ( .A1(n5888), .A2(n9683), .ZN(n5872) );
  NAND2_X1 U7435 ( .A1(n5873), .A2(n5872), .ZN(n5900) );
  XNOR2_X1 U7436 ( .A(n8890), .B(n5900), .ZN(n5892) );
  INV_X1 U7437 ( .A(n5892), .ZN(n9694) );
  INV_X1 U7438 ( .A(n5874), .ZN(n5876) );
  NAND2_X1 U7439 ( .A1(n5876), .A2(n5875), .ZN(n9394) );
  INV_X1 U7440 ( .A(n9393), .ZN(n5877) );
  NOR2_X1 U7441 ( .A1(n9394), .A2(n5877), .ZN(n5878) );
  NAND2_X1 U7442 ( .A1(n5879), .A2(n5878), .ZN(n5894) );
  NAND2_X1 U7443 ( .A1(n9665), .A2(n8934), .ZN(n5880) );
  NAND2_X1 U7444 ( .A1(n5881), .A2(n9638), .ZN(n5907) );
  INV_X1 U7445 ( .A(n5907), .ZN(n5882) );
  AND2_X1 U7446 ( .A1(n9641), .A2(n5882), .ZN(n9639) );
  INV_X1 U7447 ( .A(n9639), .ZN(n6659) );
  INV_X1 U7448 ( .A(n9323), .ZN(n6890) );
  NAND2_X1 U7449 ( .A1(n8887), .A2(n8886), .ZN(n5884) );
  INV_X1 U7450 ( .A(n5380), .ZN(n8704) );
  NAND2_X1 U7451 ( .A1(n8704), .A2(n9634), .ZN(n5883) );
  NAND2_X1 U7452 ( .A1(n5884), .A2(n5883), .ZN(n5925) );
  NAND2_X1 U7453 ( .A1(n5925), .A2(n8888), .ZN(n5887) );
  NAND2_X1 U7454 ( .A1(n5887), .A2(n5886), .ZN(n6118) );
  INV_X1 U7455 ( .A(n8889), .ZN(n6119) );
  NAND2_X1 U7456 ( .A1(n5888), .A2(n6116), .ZN(n8708) );
  XNOR2_X1 U7457 ( .A(n8755), .B(n8890), .ZN(n5890) );
  AOI22_X1 U7458 ( .A1(n9614), .A2(n8970), .B1(n8968), .B2(n9649), .ZN(n5889)
         );
  OAI21_X1 U7459 ( .B1(n5890), .B2(n9289), .A(n5889), .ZN(n5891) );
  AOI21_X1 U7460 ( .B1(n6890), .B2(n5892), .A(n5891), .ZN(n9692) );
  MUX2_X1 U7461 ( .A(n8220), .B(n9692), .S(n9641), .Z(n5899) );
  NAND2_X1 U7462 ( .A1(n6115), .A2(n9683), .ZN(n6114) );
  OR2_X1 U7463 ( .A1(n6114), .A2(n9690), .ZN(n5908) );
  INV_X1 U7464 ( .A(n5908), .ZN(n5893) );
  AOI211_X1 U7465 ( .C1(n9690), .C2(n6114), .A(n9295), .B(n5893), .ZN(n9688)
         );
  NOR2_X2 U7466 ( .A1(n5894), .A2(n9638), .ZN(n9628) );
  INV_X1 U7467 ( .A(n5895), .ZN(n9633) );
  NAND2_X1 U7468 ( .A1(n9644), .A2(n9633), .ZN(n9263) );
  OAI22_X1 U7469 ( .A1(n9263), .A2(n5901), .B1(n5896), .B2(n9306), .ZN(n5897)
         );
  AOI21_X1 U7470 ( .B1(n9688), .B2(n9628), .A(n5897), .ZN(n5898) );
  OAI211_X1 U7471 ( .C1(n9694), .C2(n6659), .A(n5899), .B(n5898), .ZN(P1_U3287) );
  NAND2_X1 U7472 ( .A1(n5900), .A2(n8890), .ZN(n5903) );
  NAND2_X1 U7473 ( .A1(n6120), .A2(n5901), .ZN(n5902) );
  NAND2_X1 U7474 ( .A1(n5903), .A2(n5902), .ZN(n5905) );
  INV_X1 U7475 ( .A(n5905), .ZN(n5904) );
  XNOR2_X1 U7476 ( .A(n8968), .B(n6213), .ZN(n8893) );
  INV_X1 U7477 ( .A(n8893), .ZN(n5912) );
  NAND2_X1 U7478 ( .A1(n5904), .A2(n5912), .ZN(n6206) );
  NAND2_X1 U7479 ( .A1(n5905), .A2(n8893), .ZN(n5906) );
  AND2_X1 U7480 ( .A1(n6206), .A2(n5906), .ZN(n9699) );
  NAND2_X1 U7481 ( .A1(n9323), .A2(n5907), .ZN(n6416) );
  NOR2_X1 U7482 ( .A1(n5908), .A2(n6213), .ZN(n6208) );
  NAND2_X1 U7483 ( .A1(n5908), .A2(n6213), .ZN(n5909) );
  NAND2_X1 U7484 ( .A1(n5909), .A2(n9625), .ZN(n5910) );
  OR2_X1 U7485 ( .A1(n6208), .A2(n5910), .ZN(n9696) );
  OAI22_X1 U7486 ( .A1(n9696), .A2(n9638), .B1(n9306), .B2(n5911), .ZN(n5916)
         );
  NAND2_X1 U7487 ( .A1(n8757), .A2(n8754), .ZN(n6215) );
  XNOR2_X1 U7488 ( .A(n6215), .B(n5912), .ZN(n5914) );
  INV_X1 U7489 ( .A(n9614), .ZN(n9291) );
  OAI22_X1 U7490 ( .A1(n6274), .A2(n9293), .B1(n6120), .B2(n9291), .ZN(n5913)
         );
  AOI21_X1 U7491 ( .B1(n5914), .B2(n9617), .A(n5913), .ZN(n9700) );
  INV_X1 U7492 ( .A(n9700), .ZN(n5915) );
  AOI211_X1 U7493 ( .C1(n9699), .C2(n6416), .A(n5916), .B(n5915), .ZN(n5918)
         );
  AOI22_X1 U7494 ( .A1(n9620), .A2(n6213), .B1(n9660), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n5917) );
  OAI21_X1 U7495 ( .B1(n5918), .B2(n9660), .A(n5917), .ZN(P1_U3286) );
  NAND2_X1 U7496 ( .A1(n5920), .A2(n8888), .ZN(n5921) );
  NAND2_X1 U7497 ( .A1(n5919), .A2(n5921), .ZN(n9680) );
  AOI211_X1 U7498 ( .C1(n5923), .C2(n5922), .A(n9295), .B(n6115), .ZN(n9675)
         );
  INV_X1 U7499 ( .A(n9306), .ZN(n9661) );
  AOI22_X1 U7500 ( .A1(n9675), .A2(n9628), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9661), .ZN(n5924) );
  OAI21_X1 U7501 ( .B1(n9677), .B2(n9263), .A(n5924), .ZN(n5930) );
  XNOR2_X1 U7502 ( .A(n5885), .B(n5925), .ZN(n5928) );
  NAND2_X1 U7503 ( .A1(n9680), .A2(n6890), .ZN(n5927) );
  AOI22_X1 U7504 ( .A1(n9614), .A2(n5380), .B1(n8970), .B2(n9649), .ZN(n5926)
         );
  OAI211_X1 U7505 ( .C1(n5928), .C2(n9289), .A(n5927), .B(n5926), .ZN(n9678)
         );
  MUX2_X1 U7506 ( .A(n9678), .B(P1_REG2_REG_2__SCAN_IN), .S(n9660), .Z(n5929)
         );
  AOI211_X1 U7507 ( .C1(n9639), .C2(n9680), .A(n5930), .B(n5929), .ZN(n5931)
         );
  INV_X1 U7508 ( .A(n5931), .ZN(P1_U3289) );
  INV_X1 U7509 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n5943) );
  OAI21_X1 U7510 ( .B1(n5934), .B2(n5933), .A(n5932), .ZN(n5939) );
  AOI211_X1 U7511 ( .C1(n5937), .C2(n5936), .A(n5935), .B(n9571), .ZN(n5938)
         );
  AOI21_X1 U7512 ( .B1(n9587), .B2(n5939), .A(n5938), .ZN(n5942) );
  NAND2_X1 U7513 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3084), .ZN(n6753) );
  INV_X1 U7514 ( .A(n6753), .ZN(n5940) );
  AOI21_X1 U7515 ( .B1(n9579), .B2(n6707), .A(n5940), .ZN(n5941) );
  OAI211_X1 U7516 ( .C1(n9593), .C2(n5943), .A(n5942), .B(n5941), .ZN(P1_U3254) );
  INV_X1 U7517 ( .A(n5945), .ZN(n5946) );
  MUX2_X1 U7518 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7532), .Z(n6043) );
  XNOR2_X1 U7519 ( .A(n6043), .B(SI_18_), .ZN(n6040) );
  XNOR2_X1 U7520 ( .A(n6042), .B(n6040), .ZN(n7366) );
  INV_X1 U7521 ( .A(n7366), .ZN(n5955) );
  NAND2_X1 U7522 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  NAND2_X1 U7523 ( .A1(n5950), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U7524 ( .A(n5951), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9091) );
  AOI22_X1 U7525 ( .A1(n9091), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n6945), .ZN(n5952) );
  OAI21_X1 U7526 ( .B1(n5955), .B2(n9417), .A(n5952), .ZN(P1_U3335) );
  XNOR2_X1 U7527 ( .A(n5953), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7995) );
  AOI22_X1 U7528 ( .A1(n7995), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8525), .ZN(n5954) );
  OAI21_X1 U7529 ( .B1(n5955), .B2(n7800), .A(n5954), .ZN(P2_U3340) );
  NAND2_X1 U7530 ( .A1(n5255), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5964) );
  INV_X1 U7531 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5956) );
  OR2_X1 U7532 ( .A1(n5528), .A2(n5956), .ZN(n5963) );
  INV_X1 U7533 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U7534 ( .A1(n7113), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7114) );
  INV_X1 U7535 ( .A(n7145), .ZN(n5958) );
  NAND2_X1 U7536 ( .A1(n5958), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7156) );
  INV_X1 U7537 ( .A(n7156), .ZN(n5959) );
  NAND2_X1 U7538 ( .A1(n5959), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n7165) );
  INV_X1 U7539 ( .A(n7165), .ZN(n5960) );
  NAND2_X1 U7540 ( .A1(n5960), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7193) );
  OR2_X1 U7541 ( .A1(n7167), .A2(n7193), .ZN(n5962) );
  INV_X1 U7542 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7194) );
  OR2_X1 U7543 ( .A1(n4280), .A2(n7194), .ZN(n5961) );
  NAND2_X1 U7544 ( .A1(n8972), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5965) );
  OAI21_X1 U7545 ( .B1(n9115), .B2(n8972), .A(n5965), .ZN(P1_U3584) );
  INV_X1 U7546 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9920) );
  MUX2_X1 U7547 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9920), .S(n6332), .Z(n5969)
         );
  NAND2_X1 U7548 ( .A1(n6134), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7549 ( .A1(n5967), .A2(n5966), .ZN(n5968) );
  NAND2_X1 U7550 ( .A1(n5968), .A2(n5969), .ZN(n6170) );
  OAI21_X1 U7551 ( .B1(n5969), .B2(n5968), .A(n6170), .ZN(n5972) );
  NAND2_X1 U7552 ( .A1(n9755), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7553 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n5970) );
  OAI211_X1 U7554 ( .C1(n5972), .C2(n9753), .A(n5971), .B(n5970), .ZN(n5977)
         );
  XNOR2_X1 U7555 ( .A(n6332), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n5974) );
  AOI211_X1 U7556 ( .C1(n5975), .C2(n5974), .A(n6176), .B(n9449), .ZN(n5976)
         );
  AOI211_X1 U7557 ( .C1(n9456), .C2(n6332), .A(n5977), .B(n5976), .ZN(n5978)
         );
  INV_X1 U7558 ( .A(n5978), .ZN(P2_U3254) );
  OR2_X1 U7559 ( .A1(n7938), .A2(n6198), .ZN(n5979) );
  NAND2_X1 U7560 ( .A1(n7937), .A2(n9856), .ZN(n7575) );
  NAND2_X1 U7561 ( .A1(n7568), .A2(n7575), .ZN(n7705) );
  NAND2_X1 U7562 ( .A1(n6090), .A2(n7705), .ZN(n6089) );
  OAI21_X1 U7563 ( .B1(n6090), .B2(n7705), .A(n6089), .ZN(n9859) );
  INV_X1 U7564 ( .A(n9859), .ZN(n6001) );
  INV_X1 U7565 ( .A(n5981), .ZN(n5983) );
  NAND2_X1 U7566 ( .A1(n5983), .A2(n5982), .ZN(n5984) );
  OR2_X1 U7567 ( .A1(n5986), .A2(n8375), .ZN(n6236) );
  NAND2_X1 U7568 ( .A1(n9781), .A2(n6236), .ZN(n5987) );
  NAND2_X1 U7569 ( .A1(n9785), .A2(n5987), .ZN(n8362) );
  XNOR2_X1 U7570 ( .A(n6097), .B(n7705), .ZN(n5989) );
  NAND2_X1 U7571 ( .A1(n5989), .A2(n9776), .ZN(n5992) );
  INV_X1 U7572 ( .A(n5990), .ZN(n5991) );
  NAND2_X1 U7573 ( .A1(n5992), .A2(n5991), .ZN(n9857) );
  OAI211_X1 U7574 ( .C1(n5994), .C2(n9856), .A(n9500), .B(n6105), .ZN(n9855)
         );
  INV_X1 U7575 ( .A(n8375), .ZN(n7370) );
  OAI22_X1 U7576 ( .A1(n9855), .A2(n7370), .B1(n9792), .B2(n5995), .ZN(n5996)
         );
  OAI21_X1 U7577 ( .B1(n9857), .B2(n5996), .A(n9785), .ZN(n6000) );
  AOI22_X1 U7578 ( .A1(n8380), .A2(n5998), .B1(n8399), .B2(
        P2_REG2_REG_5__SCAN_IN), .ZN(n5999) );
  OAI211_X1 U7579 ( .C1(n6001), .C2(n8362), .A(n6000), .B(n5999), .ZN(P2_U3291) );
  INV_X1 U7580 ( .A(n6002), .ZN(n6003) );
  AND2_X1 U7581 ( .A1(n5560), .A2(n7936), .ZN(n6012) );
  OR2_X1 U7582 ( .A1(n4288), .A2(n6008), .ZN(n6009) );
  XNOR2_X1 U7583 ( .A(n5554), .B(n7904), .ZN(n6011) );
  NOR2_X1 U7584 ( .A1(n6011), .A2(n6012), .ZN(n6013) );
  AOI21_X1 U7585 ( .B1(n6012), .B2(n6011), .A(n6013), .ZN(n7900) );
  INV_X1 U7586 ( .A(n6013), .ZN(n6014) );
  NAND2_X1 U7587 ( .A1(n7898), .A2(n6014), .ZN(n6132) );
  INV_X2 U7588 ( .A(n6015), .ZN(n6133) );
  NAND2_X1 U7589 ( .A1(n6052), .A2(n6133), .ZN(n6018) );
  AOI22_X1 U7590 ( .A1(n7473), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5720), .B2(
        n6016), .ZN(n6017) );
  AND2_X2 U7591 ( .A1(n6018), .A2(n6017), .ZN(n9869) );
  XNOR2_X1 U7592 ( .A(n5554), .B(n9869), .ZN(n6130) );
  NAND2_X1 U7593 ( .A1(n5450), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6026) );
  INV_X1 U7594 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6019) );
  OR2_X1 U7595 ( .A1(n7392), .A2(n6019), .ZN(n6025) );
  INV_X1 U7596 ( .A(n6021), .ZN(n6020) );
  NAND2_X1 U7597 ( .A1(n6020), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6029) );
  INV_X1 U7598 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7599 ( .A1(n6021), .A2(n6035), .ZN(n6022) );
  NAND2_X1 U7600 ( .A1(n6029), .A2(n6022), .ZN(n6187) );
  OR2_X1 U7601 ( .A1(n4279), .A2(n6187), .ZN(n6024) );
  INV_X1 U7602 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6188) );
  OR2_X1 U7603 ( .A1(n4277), .A2(n6188), .ZN(n6023) );
  NAND2_X1 U7604 ( .A1(n5560), .A2(n7935), .ZN(n6129) );
  XNOR2_X1 U7605 ( .A(n6130), .B(n6129), .ZN(n6131) );
  XNOR2_X1 U7606 ( .A(n6132), .B(n6131), .ZN(n6039) );
  NAND2_X1 U7607 ( .A1(n6027), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6034) );
  OR2_X1 U7608 ( .A1(n6985), .A2(n9918), .ZN(n6033) );
  INV_X1 U7609 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7610 ( .A1(n6029), .A2(n6028), .ZN(n6030) );
  NAND2_X1 U7611 ( .A1(n6138), .A2(n6030), .ZN(n6243) );
  OR2_X1 U7612 ( .A1(n4279), .A2(n6243), .ZN(n6032) );
  INV_X1 U7613 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6244) );
  OR2_X1 U7614 ( .A1(n4277), .A2(n6244), .ZN(n6031) );
  NAND4_X1 U7615 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n7934)
         );
  AOI22_X1 U7616 ( .A1(n7909), .A2(n7936), .B1(n7905), .B2(n7934), .ZN(n6038)
         );
  INV_X1 U7617 ( .A(n9869), .ZN(n6222) );
  OAI22_X1 U7618 ( .A1(n7922), .A2(n6187), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6035), .ZN(n6036) );
  AOI21_X1 U7619 ( .B1(n6222), .B2(n7903), .A(n6036), .ZN(n6037) );
  OAI211_X1 U7620 ( .C1(n6039), .C2(n7913), .A(n6038), .B(n6037), .ZN(P2_U3215) );
  INV_X1 U7621 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6050) );
  INV_X1 U7622 ( .A(n6040), .ZN(n6041) );
  NAND2_X1 U7623 ( .A1(n6042), .A2(n6041), .ZN(n6045) );
  NAND2_X1 U7624 ( .A1(n6043), .A2(SI_18_), .ZN(n6044) );
  INV_X1 U7625 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6183) );
  MUX2_X1 U7626 ( .A(n6183), .B(n6050), .S(n7532), .Z(n6047) );
  INV_X1 U7627 ( .A(SI_19_), .ZN(n6046) );
  NAND2_X1 U7628 ( .A1(n6047), .A2(n6046), .ZN(n6251) );
  INV_X1 U7629 ( .A(n6047), .ZN(n6048) );
  NAND2_X1 U7630 ( .A1(n6048), .A2(SI_19_), .ZN(n6049) );
  NAND2_X1 U7631 ( .A1(n6251), .A2(n6049), .ZN(n6252) );
  XNOR2_X1 U7632 ( .A(n6253), .B(n6252), .ZN(n7369) );
  INV_X1 U7633 ( .A(n7369), .ZN(n6184) );
  OAI222_X1 U7634 ( .A1(n7361), .A2(n6050), .B1(n7364), .B2(n6184), .C1(
        P1_U3084), .C2(n9188), .ZN(P1_U3334) );
  INV_X2 U7635 ( .A(n6051), .ZN(n6383) );
  NAND2_X1 U7636 ( .A1(n6052), .A2(n6383), .ZN(n6055) );
  AOI22_X1 U7637 ( .A1(n7086), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7085), .B2(
        n6053), .ZN(n6054) );
  NAND2_X1 U7638 ( .A1(n6055), .A2(n6054), .ZN(n9621) );
  NAND2_X1 U7639 ( .A1(n9621), .A2(n7289), .ZN(n6057) );
  OR2_X1 U7640 ( .A1(n6277), .A2(n7283), .ZN(n6056) );
  NAND2_X1 U7641 ( .A1(n6057), .A2(n6056), .ZN(n6058) );
  XNOR2_X1 U7642 ( .A(n6058), .B(n5653), .ZN(n6061) );
  NAND2_X1 U7643 ( .A1(n9621), .A2(n4285), .ZN(n6060) );
  OR2_X1 U7644 ( .A1(n6277), .A2(n7322), .ZN(n6059) );
  AND2_X1 U7645 ( .A1(n6060), .A2(n6059), .ZN(n6062) );
  NAND2_X1 U7646 ( .A1(n6061), .A2(n6062), .ZN(n6319) );
  INV_X1 U7647 ( .A(n6061), .ZN(n6064) );
  INV_X1 U7648 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7649 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  NAND2_X1 U7650 ( .A1(n6319), .A2(n6065), .ZN(n6074) );
  INV_X1 U7651 ( .A(n6074), .ZN(n6070) );
  INV_X1 U7652 ( .A(n6320), .ZN(n6072) );
  AOI21_X1 U7653 ( .B1(n6074), .B2(n6073), .A(n6072), .ZN(n6088) );
  INV_X1 U7654 ( .A(n6274), .ZN(n9615) );
  NAND2_X1 U7655 ( .A1(n5255), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6083) );
  INV_X1 U7656 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6075) );
  OR2_X1 U7657 ( .A1(n5528), .A2(n6075), .ZN(n6082) );
  NAND2_X1 U7658 ( .A1(n6077), .A2(n6076), .ZN(n6078) );
  NAND2_X1 U7659 ( .A1(n6290), .A2(n6078), .ZN(n6328) );
  OR2_X1 U7660 ( .A1(n7167), .A2(n6328), .ZN(n6081) );
  OR2_X1 U7661 ( .A1(n4280), .A2(n6079), .ZN(n6080) );
  INV_X1 U7662 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8226) );
  OAI22_X1 U7663 ( .A1(n8664), .A2(n6403), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8226), .ZN(n6084) );
  AOI21_X1 U7664 ( .B1(n8666), .B2(n9615), .A(n6084), .ZN(n6085) );
  OAI21_X1 U7665 ( .B1(n4275), .B2(n9618), .A(n6085), .ZN(n6086) );
  AOI21_X1 U7666 ( .B1(n8671), .B2(n9621), .A(n6086), .ZN(n6087) );
  OAI21_X1 U7667 ( .B1(n6088), .B2(n8645), .A(n6087), .ZN(P1_U3211) );
  OR2_X1 U7668 ( .A1(n7936), .A2(n7904), .ZN(n6227) );
  INV_X1 U7669 ( .A(n6227), .ZN(n6095) );
  NAND2_X1 U7670 ( .A1(n6089), .A2(n7937), .ZN(n6093) );
  INV_X1 U7671 ( .A(n6091), .ZN(n6092) );
  AND2_X1 U7672 ( .A1(n7936), .A2(n7904), .ZN(n6224) );
  OR2_X1 U7673 ( .A1(n6337), .A2(n6224), .ZN(n6192) );
  INV_X1 U7674 ( .A(n6224), .ZN(n6094) );
  OAI22_X1 U7675 ( .A1(n6095), .A2(n6192), .B1(n4799), .B2(n4307), .ZN(n9865)
         );
  INV_X1 U7676 ( .A(n9865), .ZN(n6112) );
  INV_X1 U7677 ( .A(n7935), .ZN(n6101) );
  INV_X1 U7678 ( .A(n7575), .ZN(n6096) );
  OR2_X1 U7679 ( .A1(n6097), .A2(n6096), .ZN(n6098) );
  NAND3_X1 U7680 ( .A1(n6098), .A2(n4307), .A3(n7568), .ZN(n6099) );
  AND2_X1 U7681 ( .A1(n6185), .A2(n6099), .ZN(n6100) );
  OAI222_X1 U7682 ( .A1(n8384), .A2(n6101), .B1(n8386), .B2(n4632), .C1(n8371), 
        .C2(n6100), .ZN(n9863) );
  NAND2_X1 U7683 ( .A1(n9863), .A2(n9788), .ZN(n6111) );
  OAI22_X1 U7684 ( .A1(n9788), .A2(n6102), .B1(n7907), .B2(n9792), .ZN(n6109)
         );
  INV_X1 U7685 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7686 ( .A1(n6104), .A2(n8375), .ZN(n9793) );
  INV_X1 U7687 ( .A(n6189), .ZN(n6107) );
  NAND2_X1 U7688 ( .A1(n6105), .A2(n7904), .ZN(n6106) );
  NAND2_X1 U7689 ( .A1(n6107), .A2(n6106), .ZN(n9862) );
  NOR2_X1 U7690 ( .A1(n8014), .A2(n9862), .ZN(n6108) );
  AOI211_X1 U7691 ( .C1(n8380), .C2(n7904), .A(n6109), .B(n6108), .ZN(n6110)
         );
  OAI211_X1 U7692 ( .C1(n6112), .C2(n8362), .A(n6111), .B(n6110), .ZN(P2_U3290) );
  XNOR2_X1 U7693 ( .A(n6113), .B(n6119), .ZN(n6125) );
  INV_X1 U7694 ( .A(n6125), .ZN(n9686) );
  INV_X1 U7695 ( .A(n9628), .ZN(n9310) );
  OAI211_X1 U7696 ( .C1(n6115), .C2(n9683), .A(n6114), .B(n9625), .ZN(n9682)
         );
  AOI22_X1 U7697 ( .A1(n9620), .A2(n6116), .B1(n9661), .B2(n9420), .ZN(n6117)
         );
  OAI21_X1 U7698 ( .B1(n9310), .B2(n9682), .A(n6117), .ZN(n6127) );
  XNOR2_X1 U7699 ( .A(n6118), .B(n6119), .ZN(n6123) );
  OAI22_X1 U7700 ( .A1(n6121), .A2(n9291), .B1(n6120), .B2(n9293), .ZN(n6122)
         );
  AOI21_X1 U7701 ( .B1(n6123), .B2(n9617), .A(n6122), .ZN(n6124) );
  OAI21_X1 U7702 ( .B1(n6125), .B2(n9323), .A(n6124), .ZN(n9684) );
  MUX2_X1 U7703 ( .A(n9684), .B(P1_REG2_REG_3__SCAN_IN), .S(n9660), .Z(n6126)
         );
  AOI211_X1 U7704 ( .C1(n9686), .C2(n9639), .A(n6127), .B(n6126), .ZN(n6128)
         );
  INV_X1 U7705 ( .A(n6128), .ZN(P1_U3288) );
  NAND2_X1 U7706 ( .A1(n6280), .A2(n6133), .ZN(n6136) );
  AOI22_X1 U7707 ( .A1(n7473), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5720), .B2(
        n6134), .ZN(n6135) );
  NAND2_X1 U7708 ( .A1(n6136), .A2(n6135), .ZN(n9873) );
  XNOR2_X1 U7709 ( .A(n5554), .B(n9873), .ZN(n6367) );
  NAND2_X1 U7710 ( .A1(n5560), .A2(n7934), .ZN(n6366) );
  XNOR2_X1 U7711 ( .A(n6367), .B(n6366), .ZN(n6369) );
  XNOR2_X1 U7712 ( .A(n6370), .B(n6369), .ZN(n6148) );
  NAND2_X1 U7713 ( .A1(n6027), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6143) );
  INV_X1 U7714 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6355) );
  OR2_X1 U7715 ( .A1(n4278), .A2(n6355), .ZN(n6142) );
  INV_X1 U7716 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U7717 ( .A1(n6138), .A2(n6377), .ZN(n6139) );
  NAND2_X1 U7718 ( .A1(n6342), .A2(n6139), .ZN(n6376) );
  OR2_X1 U7719 ( .A1(n4279), .A2(n6376), .ZN(n6141) );
  OR2_X1 U7720 ( .A1(n7522), .A2(n9920), .ZN(n6140) );
  NAND4_X1 U7721 ( .A1(n6143), .A2(n6142), .A3(n6141), .A4(n6140), .ZN(n9771)
         );
  AOI22_X1 U7722 ( .A1(n7909), .A2(n7935), .B1(n7905), .B2(n9771), .ZN(n6145)
         );
  OAI211_X1 U7723 ( .C1(n6243), .C2(n7922), .A(n6145), .B(n6144), .ZN(n6146)
         );
  AOI21_X1 U7724 ( .B1(n9873), .B2(n7903), .A(n6146), .ZN(n6147) );
  OAI21_X1 U7725 ( .B1(n6148), .B2(n7913), .A(n6147), .ZN(P2_U3223) );
  NAND2_X1 U7726 ( .A1(n7555), .A2(n6149), .ZN(n9846) );
  INV_X1 U7727 ( .A(n9846), .ZN(n6156) );
  OAI21_X1 U7728 ( .B1(n9767), .B2(n8380), .A(n6150), .ZN(n6155) );
  AOI22_X1 U7729 ( .A1(n9776), .A2(n9846), .B1(n9769), .B2(n5545), .ZN(n9842)
         );
  OAI21_X1 U7730 ( .B1(n5460), .B2(n9792), .A(n9842), .ZN(n6153) );
  NOR2_X1 U7731 ( .A1(n9785), .A2(n6151), .ZN(n6152) );
  AOI21_X1 U7732 ( .B1(n9788), .B2(n6153), .A(n6152), .ZN(n6154) );
  OAI211_X1 U7733 ( .C1(n6156), .C2(n8362), .A(n6155), .B(n6154), .ZN(P2_U3296) );
  INV_X1 U7734 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n6168) );
  OAI21_X1 U7735 ( .B1(n6159), .B2(n6158), .A(n6157), .ZN(n6164) );
  OAI21_X1 U7736 ( .B1(n6162), .B2(n6161), .A(n6160), .ZN(n6163) );
  AOI22_X1 U7737 ( .A1(n9588), .A2(n6164), .B1(n9587), .B2(n6163), .ZN(n6167)
         );
  NAND2_X1 U7738 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n8543) );
  INV_X1 U7739 ( .A(n8543), .ZN(n6165) );
  AOI21_X1 U7740 ( .B1(n9579), .B2(n6768), .A(n6165), .ZN(n6166) );
  OAI211_X1 U7741 ( .C1(n9593), .C2(n6168), .A(n6167), .B(n6166), .ZN(P1_U3255) );
  NAND2_X1 U7742 ( .A1(n6332), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7743 ( .A1(n6170), .A2(n6169), .ZN(n6172) );
  INV_X1 U7744 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9922) );
  MUX2_X1 U7745 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9922), .S(n6449), .Z(n6171)
         );
  AND2_X1 U7746 ( .A1(n6172), .A2(n6171), .ZN(n6309) );
  NOR2_X1 U7747 ( .A1(n6172), .A2(n6171), .ZN(n6173) );
  OR2_X1 U7748 ( .A1(n6309), .A2(n6173), .ZN(n6175) );
  NAND2_X1 U7749 ( .A1(n9755), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7750 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n6487) );
  OAI211_X1 U7751 ( .C1(n9753), .C2(n6175), .A(n6174), .B(n6487), .ZN(n6181)
         );
  NAND2_X1 U7752 ( .A1(n6449), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6177) );
  OAI21_X1 U7753 ( .B1(n6449), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6177), .ZN(
        n6178) );
  AOI211_X1 U7754 ( .C1(n6179), .C2(n6178), .A(n9449), .B(n6304), .ZN(n6180)
         );
  AOI211_X1 U7755 ( .C1(n9456), .C2(n6449), .A(n6181), .B(n6180), .ZN(n6182)
         );
  INV_X1 U7756 ( .A(n6182), .ZN(P2_U3255) );
  OAI222_X1 U7757 ( .A1(P2_U3152), .A2(n8375), .B1(n7800), .B2(n6184), .C1(
        n6183), .C2(n7817), .ZN(P2_U3339) );
  INV_X1 U7758 ( .A(n7904), .ZN(n9861) );
  OR2_X1 U7759 ( .A1(n7936), .A2(n9861), .ZN(n7582) );
  OR2_X1 U7760 ( .A1(n7935), .A2(n9869), .ZN(n7583) );
  NAND2_X1 U7761 ( .A1(n7935), .A2(n9869), .ZN(n7584) );
  INV_X1 U7762 ( .A(n7706), .ZN(n7581) );
  XNOR2_X1 U7763 ( .A(n6349), .B(n7581), .ZN(n6186) );
  AOI222_X1 U7764 ( .A1(n7936), .A2(n9772), .B1(n7934), .B2(n9769), .C1(n9776), 
        .C2(n6186), .ZN(n9868) );
  OAI22_X1 U7765 ( .A1(n9788), .A2(n6188), .B1(n6187), .B2(n9792), .ZN(n6191)
         );
  NAND2_X1 U7766 ( .A1(n6189), .A2(n9869), .ZN(n6245) );
  OAI211_X1 U7767 ( .C1(n6189), .C2(n9869), .A(n6245), .B(n9500), .ZN(n9867)
         );
  NOR2_X1 U7768 ( .A1(n9867), .A2(n9793), .ZN(n6190) );
  AOI211_X1 U7769 ( .C1(n8380), .C2(n6222), .A(n6191), .B(n6190), .ZN(n6195)
         );
  NAND2_X1 U7770 ( .A1(n6192), .A2(n6227), .ZN(n6193) );
  XNOR2_X1 U7771 ( .A(n6193), .B(n7706), .ZN(n9871) );
  INV_X1 U7772 ( .A(n8362), .ZN(n8143) );
  NAND2_X1 U7773 ( .A1(n9871), .A2(n8143), .ZN(n6194) );
  OAI211_X1 U7774 ( .C1(n9868), .C2(n8399), .A(n6195), .B(n6194), .ZN(P2_U3289) );
  INV_X1 U7775 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8206) );
  INV_X1 U7776 ( .A(n9793), .ZN(n6534) );
  INV_X1 U7777 ( .A(n9792), .ZN(n8397) );
  AOI22_X1 U7778 ( .A1(n6197), .A2(n6534), .B1(n6196), .B2(n8397), .ZN(n6200)
         );
  NAND2_X1 U7779 ( .A1(n8380), .A2(n6198), .ZN(n6199) );
  OAI211_X1 U7780 ( .C1(n8206), .C2(n9788), .A(n6200), .B(n6199), .ZN(n6201)
         );
  AOI21_X1 U7781 ( .B1(n8143), .B2(n6202), .A(n6201), .ZN(n6203) );
  OAI21_X1 U7782 ( .B1(n8399), .B2(n6204), .A(n6203), .ZN(P2_U3292) );
  NAND2_X1 U7783 ( .A1(n8968), .A2(n6213), .ZN(n6205) );
  NAND2_X1 U7784 ( .A1(n6274), .A2(n6211), .ZN(n8714) );
  NAND2_X1 U7785 ( .A1(n9704), .A2(n9615), .ZN(n8715) );
  NAND2_X1 U7786 ( .A1(n8714), .A2(n8715), .ZN(n8891) );
  OAI21_X1 U7787 ( .B1(n4371), .B2(n8891), .A(n6276), .ZN(n9707) );
  INV_X1 U7788 ( .A(n9626), .ZN(n6207) );
  OAI211_X1 U7789 ( .C1(n9704), .C2(n6208), .A(n6207), .B(n9625), .ZN(n9703)
         );
  INV_X1 U7790 ( .A(n6209), .ZN(n6210) );
  AOI22_X1 U7791 ( .A1(n9620), .A2(n6211), .B1(n6210), .B2(n9661), .ZN(n6212)
         );
  OAI21_X1 U7792 ( .B1(n9703), .B2(n9310), .A(n6212), .ZN(n6220) );
  INV_X1 U7793 ( .A(n6213), .ZN(n9697) );
  AND2_X1 U7794 ( .A1(n8968), .A2(n9697), .ZN(n8713) );
  NAND2_X1 U7795 ( .A1(n6214), .A2(n6213), .ZN(n8710) );
  XNOR2_X1 U7796 ( .A(n6286), .B(n8891), .ZN(n6218) );
  NAND2_X1 U7797 ( .A1(n9707), .A2(n6890), .ZN(n6217) );
  INV_X1 U7798 ( .A(n6277), .ZN(n8967) );
  AOI22_X1 U7799 ( .A1(n8967), .A2(n9649), .B1(n9614), .B2(n8968), .ZN(n6216)
         );
  OAI211_X1 U7800 ( .C1(n9289), .C2(n6218), .A(n6217), .B(n6216), .ZN(n9705)
         );
  MUX2_X1 U7801 ( .A(n9705), .B(P1_REG2_REG_6__SCAN_IN), .S(n9660), .Z(n6219)
         );
  AOI211_X1 U7802 ( .C1(n9639), .C2(n9707), .A(n6220), .B(n6219), .ZN(n6221)
         );
  INV_X1 U7803 ( .A(n6221), .ZN(P1_U3285) );
  INV_X1 U7804 ( .A(n6226), .ZN(n6223) );
  NOR2_X1 U7805 ( .A1(n6223), .A2(n7706), .ZN(n6229) );
  OR2_X1 U7806 ( .A1(n6224), .A2(n6229), .ZN(n6335) );
  OR2_X1 U7807 ( .A1(n6337), .A2(n6335), .ZN(n6232) );
  INV_X1 U7808 ( .A(n7934), .ZN(n6225) );
  OR2_X1 U7809 ( .A1(n6225), .A2(n9873), .ZN(n7588) );
  NAND2_X1 U7810 ( .A1(n6225), .A2(n9873), .ZN(n7589) );
  INV_X1 U7811 ( .A(n7709), .ZN(n6230) );
  AND2_X1 U7812 ( .A1(n6227), .A2(n6226), .ZN(n6228) );
  OR2_X1 U7813 ( .A1(n6229), .A2(n6228), .ZN(n6231) );
  AND2_X1 U7814 ( .A1(n6230), .A2(n6231), .ZN(n6338) );
  NAND2_X1 U7815 ( .A1(n6232), .A2(n6338), .ZN(n6235) );
  NAND2_X1 U7816 ( .A1(n6232), .A2(n6231), .ZN(n6233) );
  NAND2_X1 U7817 ( .A1(n6233), .A2(n7709), .ZN(n6234) );
  NAND2_X1 U7818 ( .A1(n6235), .A2(n6234), .ZN(n9872) );
  OR2_X1 U7819 ( .A1(n8399), .A2(n6236), .ZN(n9798) );
  AOI22_X1 U7820 ( .A1(n9772), .A2(n7935), .B1(n9771), .B2(n9769), .ZN(n6242)
         );
  OR2_X1 U7821 ( .A1(n6349), .A2(n7706), .ZN(n6237) );
  AND2_X1 U7822 ( .A1(n6237), .A2(n7584), .ZN(n6239) );
  AND2_X1 U7823 ( .A1(n7709), .A2(n7584), .ZN(n6350) );
  NAND2_X1 U7824 ( .A1(n6237), .A2(n6350), .ZN(n6238) );
  OAI21_X1 U7825 ( .B1(n7709), .B2(n6239), .A(n6238), .ZN(n6240) );
  NAND2_X1 U7826 ( .A1(n6240), .A2(n9776), .ZN(n6241) );
  OAI211_X1 U7827 ( .C1(n9872), .C2(n9781), .A(n6242), .B(n6241), .ZN(n9876)
         );
  NAND2_X1 U7828 ( .A1(n9876), .A2(n9788), .ZN(n6250) );
  OAI22_X1 U7829 ( .A1(n9785), .A2(n6244), .B1(n6243), .B2(n9792), .ZN(n6248)
         );
  NAND2_X1 U7830 ( .A1(n6245), .A2(n9873), .ZN(n6246) );
  NAND2_X1 U7831 ( .A1(n6356), .A2(n6246), .ZN(n9875) );
  NOR2_X1 U7832 ( .A1(n9875), .A2(n8014), .ZN(n6247) );
  AOI211_X1 U7833 ( .C1(n8380), .C2(n9873), .A(n6248), .B(n6247), .ZN(n6249)
         );
  OAI211_X1 U7834 ( .C1(n9872), .C2(n9798), .A(n6250), .B(n6249), .ZN(P2_U3288) );
  INV_X1 U7835 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7051) );
  INV_X1 U7836 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6364) );
  MUX2_X1 U7837 ( .A(n6364), .B(n7051), .S(n7532), .Z(n6255) );
  INV_X1 U7838 ( .A(SI_20_), .ZN(n6254) );
  NAND2_X1 U7839 ( .A1(n6255), .A2(n6254), .ZN(n6272) );
  INV_X1 U7840 ( .A(n6255), .ZN(n6256) );
  NAND2_X1 U7841 ( .A1(n6256), .A2(SI_20_), .ZN(n6257) );
  OAI21_X1 U7842 ( .B1(n6259), .B2(n6258), .A(n6273), .ZN(n7385) );
  INV_X1 U7843 ( .A(n7385), .ZN(n6365) );
  OAI222_X1 U7844 ( .A1(n7361), .A2(n7051), .B1(n7364), .B2(n6365), .C1(
        P1_U3084), .C2(n6260), .ZN(P1_U3333) );
  NAND2_X1 U7845 ( .A1(n9785), .A2(n6261), .ZN(n6264) );
  OR2_X1 U7846 ( .A1(n9792), .A2(n6262), .ZN(n6263) );
  OAI211_X1 U7847 ( .C1(n9788), .C2(n6265), .A(n6264), .B(n6263), .ZN(n6269)
         );
  OAI22_X1 U7848 ( .A1(n8014), .A2(n6267), .B1(n6266), .B2(n9795), .ZN(n6268)
         );
  AOI211_X1 U7849 ( .C1(n8143), .C2(n6270), .A(n6269), .B(n6268), .ZN(n6271)
         );
  INV_X1 U7850 ( .A(n6271), .ZN(P2_U3295) );
  INV_X1 U7851 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6362) );
  INV_X1 U7852 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7097) );
  MUX2_X1 U7853 ( .A(n6362), .B(n7097), .S(n7532), .Z(n6624) );
  XNOR2_X1 U7854 ( .A(n6624), .B(SI_21_), .ZN(n6623) );
  INV_X1 U7855 ( .A(n7398), .ZN(n6363) );
  OAI222_X1 U7856 ( .A1(n7364), .A2(n6363), .B1(n8934), .B2(P1_U3084), .C1(
        n7097), .C2(n7361), .ZN(P1_U3332) );
  NAND2_X1 U7857 ( .A1(n6274), .A2(n9704), .ZN(n6275) );
  OR2_X1 U7858 ( .A1(n9621), .A2(n6277), .ZN(n8718) );
  NAND2_X1 U7859 ( .A1(n9621), .A2(n6277), .ZN(n8766) );
  OR2_X1 U7860 ( .A1(n9621), .A2(n8967), .ZN(n6278) );
  NAND2_X1 U7861 ( .A1(n6279), .A2(n6278), .ZN(n6421) );
  NAND2_X1 U7862 ( .A1(n6280), .A2(n6383), .ZN(n6283) );
  AOI22_X1 U7863 ( .A1(n7086), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7085), .B2(
        n6281), .ZN(n6282) );
  NAND2_X1 U7864 ( .A1(n6283), .A2(n6282), .ZN(n6417) );
  OR2_X1 U7865 ( .A1(n6417), .A2(n6403), .ZN(n9594) );
  NAND2_X1 U7866 ( .A1(n6417), .A2(n6403), .ZN(n8776) );
  OR2_X1 U7867 ( .A1(n6421), .A2(n8894), .ZN(n9603) );
  NAND2_X1 U7868 ( .A1(n6421), .A2(n8894), .ZN(n6284) );
  NAND2_X1 U7869 ( .A1(n9603), .A2(n6284), .ZN(n9715) );
  INV_X1 U7870 ( .A(n8714), .ZN(n6285) );
  OAI21_X1 U7871 ( .B1(n6286), .B2(n6285), .A(n8715), .ZN(n9612) );
  INV_X1 U7872 ( .A(n9612), .ZN(n6287) );
  INV_X1 U7873 ( .A(n8718), .ZN(n8765) );
  XOR2_X1 U7874 ( .A(n8894), .B(n4370), .Z(n6288) );
  NAND2_X1 U7875 ( .A1(n6288), .A2(n9617), .ZN(n6298) );
  NAND2_X1 U7876 ( .A1(n5255), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6296) );
  AND2_X1 U7877 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  OR2_X1 U7878 ( .A1(n6291), .A2(n6405), .ZN(n9599) );
  OR2_X1 U7879 ( .A1(n7167), .A2(n9599), .ZN(n6295) );
  OR2_X1 U7880 ( .A1(n5528), .A2(n9728), .ZN(n6294) );
  INV_X1 U7881 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6292) );
  OR2_X1 U7882 ( .A1(n4280), .A2(n6292), .ZN(n6293) );
  NAND4_X1 U7883 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(n8966)
         );
  AOI22_X1 U7884 ( .A1(n8967), .A2(n9614), .B1(n9649), .B2(n8966), .ZN(n6297)
         );
  OAI211_X1 U7885 ( .C1(n9323), .C2(n9715), .A(n6298), .B(n6297), .ZN(n9717)
         );
  NAND2_X1 U7886 ( .A1(n9717), .A2(n9641), .ZN(n6303) );
  OAI22_X1 U7887 ( .A1(n9641), .A2(n6079), .B1(n6328), .B2(n9306), .ZN(n6301)
         );
  INV_X1 U7888 ( .A(n9621), .ZN(n9711) );
  INV_X1 U7889 ( .A(n9624), .ZN(n6299) );
  OAI211_X1 U7890 ( .C1(n6299), .C2(n4446), .A(n9625), .B(n9606), .ZN(n9716)
         );
  NOR2_X1 U7891 ( .A1(n9716), .A2(n9310), .ZN(n6300) );
  AOI211_X1 U7892 ( .C1(n9620), .C2(n6417), .A(n6301), .B(n6300), .ZN(n6302)
         );
  OAI211_X1 U7893 ( .C1(n9715), .C2(n6659), .A(n6303), .B(n6302), .ZN(P1_U3283) );
  NOR2_X1 U7894 ( .A1(n6496), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6305) );
  AOI21_X1 U7895 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n6496), .A(n6305), .ZN(
        n6306) );
  NAND2_X1 U7896 ( .A1(n6307), .A2(n6306), .ZN(n6494) );
  OAI21_X1 U7897 ( .B1(n6307), .B2(n6306), .A(n6494), .ZN(n6308) );
  NAND2_X1 U7898 ( .A1(n6308), .A2(n9750), .ZN(n6314) );
  AND2_X1 U7899 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7880) );
  INV_X1 U7900 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6455) );
  MUX2_X1 U7901 ( .A(n6455), .B(P2_REG1_REG_11__SCAN_IN), .S(n6496), .Z(n6310)
         );
  NOR2_X1 U7902 ( .A1(n6311), .A2(n6310), .ZN(n6495) );
  AOI211_X1 U7903 ( .C1(n6311), .C2(n6310), .A(n6495), .B(n9753), .ZN(n6312)
         );
  AOI211_X1 U7904 ( .C1(n9755), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7880), .B(
        n6312), .ZN(n6313) );
  OAI211_X1 U7905 ( .C1(n9751), .C2(n6315), .A(n6314), .B(n6313), .ZN(P2_U3256) );
  NAND2_X1 U7906 ( .A1(n6417), .A2(n7289), .ZN(n6317) );
  OR2_X1 U7907 ( .A1(n6403), .A2(n7283), .ZN(n6316) );
  NAND2_X1 U7908 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  XNOR2_X1 U7909 ( .A(n6318), .B(n7320), .ZN(n6397) );
  NOR2_X1 U7910 ( .A1(n6403), .A2(n7322), .ZN(n6321) );
  AOI21_X1 U7911 ( .B1(n6417), .B2(n4285), .A(n6321), .ZN(n6323) );
  INV_X1 U7912 ( .A(n6323), .ZN(n6322) );
  NAND2_X1 U7913 ( .A1(n6399), .A2(n6398), .ZN(n6324) );
  XOR2_X1 U7914 ( .A(n6397), .B(n6324), .Z(n6331) );
  INV_X1 U7915 ( .A(n8966), .ZN(n6424) );
  OAI21_X1 U7916 ( .B1(n8664), .B2(n6424), .A(n6325), .ZN(n6326) );
  AOI21_X1 U7917 ( .B1(n8666), .B2(n8967), .A(n6326), .ZN(n6327) );
  OAI21_X1 U7918 ( .B1(n4275), .B2(n6328), .A(n6327), .ZN(n6329) );
  AOI21_X1 U7919 ( .B1(n8671), .B2(n6417), .A(n6329), .ZN(n6330) );
  OAI21_X1 U7920 ( .B1(n6331), .B2(n8645), .A(n6330), .ZN(P1_U3219) );
  NAND2_X1 U7921 ( .A1(n6384), .A2(n6133), .ZN(n6334) );
  AOI22_X1 U7922 ( .A1(n7473), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5720), .B2(
        n6332), .ZN(n6333) );
  INV_X1 U7923 ( .A(n9771), .ZN(n6488) );
  OR2_X1 U7924 ( .A1(n6471), .A2(n6488), .ZN(n7596) );
  NAND2_X1 U7925 ( .A1(n6471), .A2(n6488), .ZN(n7592) );
  AND2_X1 U7926 ( .A1(n9873), .A2(n7934), .ZN(n6339) );
  XOR2_X1 U7927 ( .A(n7708), .B(n6473), .Z(n9880) );
  NAND2_X1 U7928 ( .A1(n5450), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U7929 ( .A1(n7517), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6346) );
  INV_X1 U7930 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U7931 ( .A1(n6342), .A2(n6341), .ZN(n6343) );
  NAND2_X1 U7932 ( .A1(n6458), .A2(n6343), .ZN(n9783) );
  OR2_X1 U7933 ( .A1(n4279), .A2(n9783), .ZN(n6345) );
  INV_X1 U7934 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9784) );
  OR2_X1 U7935 ( .A1(n4277), .A2(n9784), .ZN(n6344) );
  NAND4_X1 U7936 ( .A1(n6347), .A2(n6346), .A3(n6345), .A4(n6344), .ZN(n7933)
         );
  AOI22_X1 U7937 ( .A1(n9769), .A2(n7933), .B1(n7934), .B2(n9772), .ZN(n6378)
         );
  INV_X1 U7938 ( .A(n7589), .ZN(n6351) );
  OR2_X1 U7939 ( .A1(n7706), .A2(n6351), .ZN(n6348) );
  OR2_X1 U7940 ( .A1(n6349), .A2(n6348), .ZN(n6446) );
  OR2_X1 U7941 ( .A1(n6351), .A2(n6350), .ZN(n6444) );
  AND2_X1 U7942 ( .A1(n6446), .A2(n6444), .ZN(n6352) );
  XNOR2_X1 U7943 ( .A(n6352), .B(n7708), .ZN(n6353) );
  NAND2_X1 U7944 ( .A1(n6353), .A2(n9776), .ZN(n6354) );
  OAI211_X1 U7945 ( .C1(n9880), .C2(n9781), .A(n6378), .B(n6354), .ZN(n9883)
         );
  NAND2_X1 U7946 ( .A1(n9883), .A2(n9788), .ZN(n6361) );
  OAI22_X1 U7947 ( .A1(n9785), .A2(n6355), .B1(n6376), .B2(n9792), .ZN(n6359)
         );
  AND2_X1 U7948 ( .A1(n6356), .A2(n6471), .ZN(n6357) );
  OR2_X1 U7949 ( .A1(n6357), .A2(n9765), .ZN(n9882) );
  NOR2_X1 U7950 ( .A1(n9882), .A2(n8014), .ZN(n6358) );
  AOI211_X1 U7951 ( .C1(n8380), .C2(n6471), .A(n6359), .B(n6358), .ZN(n6360)
         );
  OAI211_X1 U7952 ( .C1(n9880), .C2(n9798), .A(n6361), .B(n6360), .ZN(P2_U3287) );
  OAI222_X1 U7953 ( .A1(P2_U3152), .A2(n7727), .B1(n7800), .B2(n6363), .C1(
        n6362), .C2(n7817), .ZN(P2_U3337) );
  OAI222_X1 U7954 ( .A1(P2_U3152), .A2(n5468), .B1(n7800), .B2(n6365), .C1(
        n6364), .C2(n7817), .ZN(P2_U3338) );
  INV_X1 U7955 ( .A(n6471), .ZN(n9881) );
  INV_X1 U7956 ( .A(n6366), .ZN(n6368) );
  AND2_X1 U7957 ( .A1(n5560), .A2(n9771), .ZN(n6372) );
  XNOR2_X1 U7958 ( .A(n5554), .B(n6471), .ZN(n6371) );
  NOR2_X1 U7959 ( .A1(n6371), .A2(n6372), .ZN(n6484) );
  AOI21_X1 U7960 ( .B1(n6372), .B2(n6371), .A(n6484), .ZN(n6373) );
  OAI21_X1 U7961 ( .B1(n6374), .B2(n6373), .A(n6485), .ZN(n6375) );
  NAND2_X1 U7962 ( .A1(n6375), .A2(n7901), .ZN(n6382) );
  INV_X1 U7963 ( .A(n6376), .ZN(n6380) );
  OAI22_X1 U7964 ( .A1(n7792), .A2(n6378), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6377), .ZN(n6379) );
  AOI21_X1 U7965 ( .B1(n6380), .B2(n7885), .A(n6379), .ZN(n6381) );
  OAI211_X1 U7966 ( .C1(n9881), .C2(n7927), .A(n6382), .B(n6381), .ZN(P2_U3233) );
  NAND2_X1 U7967 ( .A1(n6384), .A2(n6383), .ZN(n6387) );
  AOI22_X1 U7968 ( .A1(n7086), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7085), .B2(
        n6385), .ZN(n6386) );
  NAND2_X1 U7969 ( .A1(n6387), .A2(n6386), .ZN(n9601) );
  NAND2_X1 U7970 ( .A1(n9601), .A2(n7289), .ZN(n6389) );
  NAND2_X1 U7971 ( .A1(n8966), .A2(n4285), .ZN(n6388) );
  NAND2_X1 U7972 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  XNOR2_X1 U7973 ( .A(n6390), .B(n5653), .ZN(n6392) );
  AND2_X1 U7974 ( .A1(n8966), .A2(n7286), .ZN(n6391) );
  AOI21_X1 U7975 ( .B1(n9601), .B2(n4285), .A(n6391), .ZN(n6393) );
  NAND2_X1 U7976 ( .A1(n6392), .A2(n6393), .ZN(n6543) );
  INV_X1 U7977 ( .A(n6392), .ZN(n6395) );
  INV_X1 U7978 ( .A(n6393), .ZN(n6394) );
  NAND2_X1 U7979 ( .A1(n6395), .A2(n6394), .ZN(n6396) );
  AND2_X1 U7980 ( .A1(n6543), .A2(n6396), .ZN(n6401) );
  OAI21_X1 U7981 ( .B1(n6401), .B2(n6400), .A(n6544), .ZN(n6402) );
  NAND2_X1 U7982 ( .A1(n6402), .A2(n8657), .ZN(n6415) );
  INV_X1 U7983 ( .A(n6403), .ZN(n9613) );
  NAND2_X1 U7984 ( .A1(n5255), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6410) );
  INV_X1 U7985 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6404) );
  OR2_X1 U7986 ( .A1(n5528), .A2(n6404), .ZN(n6409) );
  NOR2_X1 U7987 ( .A1(n6405), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6406) );
  OR2_X1 U7988 ( .A1(n6427), .A2(n6406), .ZN(n6550) );
  OR2_X1 U7989 ( .A1(n7167), .A2(n6550), .ZN(n6408) );
  OR2_X1 U7990 ( .A1(n4280), .A2(n6438), .ZN(n6407) );
  OAI21_X1 U7991 ( .B1(n8664), .B2(n6679), .A(n6411), .ZN(n6413) );
  NOR2_X1 U7992 ( .A1(n4275), .A2(n9599), .ZN(n6412) );
  AOI211_X1 U7993 ( .C1(n8666), .C2(n9613), .A(n6413), .B(n6412), .ZN(n6414)
         );
  OAI211_X1 U7994 ( .C1(n4445), .C2(n8656), .A(n6415), .B(n6414), .ZN(P1_U3229) );
  NAND2_X1 U7995 ( .A1(n9644), .A2(n6416), .ZN(n9301) );
  NAND2_X1 U7996 ( .A1(n6417), .A2(n9613), .ZN(n9602) );
  NAND2_X1 U7997 ( .A1(n9601), .A2(n8966), .ZN(n6418) );
  AND2_X1 U7998 ( .A1(n9602), .A2(n6418), .ZN(n6419) );
  OR2_X1 U7999 ( .A1(n4317), .A2(n6419), .ZN(n6420) );
  NAND2_X1 U8000 ( .A1(n6448), .A2(n6383), .ZN(n6423) );
  AOI22_X1 U8001 ( .A1(n7086), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7085), .B2(
        n9037), .ZN(n6422) );
  NAND2_X2 U8002 ( .A1(n6423), .A2(n6422), .ZN(n6582) );
  OR2_X2 U8003 ( .A1(n6582), .A2(n6679), .ZN(n8782) );
  NAND2_X1 U8004 ( .A1(n6582), .A2(n6679), .ZN(n8773) );
  XNOR2_X1 U8005 ( .A(n6583), .B(n8881), .ZN(n9463) );
  INV_X1 U8006 ( .A(n9463), .ZN(n6443) );
  OR2_X1 U8007 ( .A1(n9601), .A2(n6424), .ZN(n8882) );
  AND2_X1 U8008 ( .A1(n8882), .A2(n9594), .ZN(n8777) );
  AND2_X1 U8009 ( .A1(n9601), .A2(n6424), .ZN(n8883) );
  INV_X1 U8010 ( .A(n8782), .ZN(n6425) );
  NOR2_X1 U8011 ( .A1(n6647), .A2(n6425), .ZN(n6435) );
  OAI21_X1 U8012 ( .B1(n6426), .B2(n8881), .A(n9617), .ZN(n6434) );
  NAND2_X1 U8013 ( .A1(n8678), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6432) );
  INV_X1 U8014 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6652) );
  OR2_X1 U8015 ( .A1(n4280), .A2(n6652), .ZN(n6431) );
  OR2_X1 U8016 ( .A1(n6427), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8017 ( .A1(n6605), .A2(n6428), .ZN(n6676) );
  OR2_X1 U8018 ( .A1(n7167), .A2(n6676), .ZN(n6430) );
  OR2_X1 U8019 ( .A1(n8683), .A2(n9543), .ZN(n6429) );
  NAND4_X1 U8020 ( .A1(n6432), .A2(n6431), .A3(n6430), .A4(n6429), .ZN(n8965)
         );
  AOI22_X1 U8021 ( .A1(n9614), .A2(n8966), .B1(n8965), .B2(n9649), .ZN(n6433)
         );
  OAI21_X1 U8022 ( .B1(n6435), .B2(n6434), .A(n6433), .ZN(n9461) );
  INV_X1 U8023 ( .A(n6654), .ZN(n6437) );
  AOI21_X1 U8024 ( .B1(n9607), .B2(n6582), .A(n9295), .ZN(n6436) );
  NAND2_X1 U8025 ( .A1(n6437), .A2(n6436), .ZN(n9459) );
  OAI22_X1 U8026 ( .A1(n9641), .A2(n6438), .B1(n6550), .B2(n9306), .ZN(n6439)
         );
  AOI21_X1 U8027 ( .B1(n6582), .B2(n9620), .A(n6439), .ZN(n6440) );
  OAI21_X1 U8028 ( .B1(n9459), .B2(n9310), .A(n6440), .ZN(n6441) );
  AOI21_X1 U8029 ( .B1(n9461), .B2(n9641), .A(n6441), .ZN(n6442) );
  OAI21_X1 U8030 ( .B1(n9301), .B2(n6443), .A(n6442), .ZN(P1_U3281) );
  AND2_X1 U8031 ( .A1(n6444), .A2(n7596), .ZN(n6445) );
  NAND2_X1 U8032 ( .A1(n6446), .A2(n6445), .ZN(n6447) );
  NAND2_X1 U8033 ( .A1(n6448), .A2(n6133), .ZN(n6451) );
  AOI22_X1 U8034 ( .A1(n7473), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5720), .B2(
        n6449), .ZN(n6450) );
  INV_X1 U8035 ( .A(n7933), .ZN(n6452) );
  OR2_X1 U8036 ( .A1(n6491), .A2(n6452), .ZN(n7599) );
  NAND2_X1 U8037 ( .A1(n6491), .A2(n6452), .ZN(n7595) );
  INV_X1 U8038 ( .A(n9777), .ZN(n9773) );
  NAND2_X1 U8039 ( .A1(n6584), .A2(n6133), .ZN(n6454) );
  AOI22_X1 U8040 ( .A1(n7473), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5720), .B2(
        n6496), .ZN(n6453) );
  NAND2_X2 U8041 ( .A1(n6454), .A2(n6453), .ZN(n7882) );
  NAND2_X1 U8042 ( .A1(n7517), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6463) );
  OR2_X1 U8043 ( .A1(n6985), .A2(n6455), .ZN(n6462) );
  INV_X1 U8044 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U8045 ( .A1(n6458), .A2(n6457), .ZN(n6459) );
  NAND2_X1 U8046 ( .A1(n6566), .A2(n6459), .ZN(n7883) );
  OR2_X1 U8047 ( .A1(n4279), .A2(n7883), .ZN(n6461) );
  INV_X1 U8048 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6479) );
  OR2_X1 U8049 ( .A1(n4278), .A2(n6479), .ZN(n6460) );
  NAND4_X1 U8050 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(n9770)
         );
  INV_X1 U8051 ( .A(n9770), .ZN(n6803) );
  NAND2_X1 U8052 ( .A1(n7882), .A2(n6803), .ZN(n7610) );
  NAND2_X1 U8053 ( .A1(n7606), .A2(n7610), .ZN(n7711) );
  XNOR2_X1 U8054 ( .A(n6561), .B(n7711), .ZN(n6470) );
  NAND2_X1 U8055 ( .A1(n7933), .A2(n9772), .ZN(n6469) );
  NAND2_X1 U8056 ( .A1(n7517), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6467) );
  INV_X1 U8057 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6497) );
  OR2_X1 U8058 ( .A1(n6985), .A2(n6497), .ZN(n6466) );
  INV_X1 U8059 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6565) );
  XNOR2_X1 U8060 ( .A(n6566), .B(n6565), .ZN(n6802) );
  OR2_X1 U8061 ( .A1(n4279), .A2(n6802), .ZN(n6465) );
  INV_X1 U8062 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6576) );
  OR2_X1 U8063 ( .A1(n4278), .A2(n6576), .ZN(n6464) );
  NAND4_X1 U8064 ( .A1(n6467), .A2(n6466), .A3(n6465), .A4(n6464), .ZN(n7932)
         );
  NAND2_X1 U8065 ( .A1(n7932), .A2(n9769), .ZN(n6468) );
  NAND2_X1 U8066 ( .A1(n6469), .A2(n6468), .ZN(n7881) );
  AOI21_X1 U8067 ( .B1(n6470), .B2(n9776), .A(n7881), .ZN(n9895) );
  OR2_X1 U8068 ( .A1(n6471), .A2(n9771), .ZN(n6472) );
  INV_X1 U8069 ( .A(n9761), .ZN(n6474) );
  NAND2_X1 U8070 ( .A1(n6474), .A2(n9773), .ZN(n9760) );
  NAND2_X1 U8071 ( .A1(n6491), .A2(n7933), .ZN(n6475) );
  NAND2_X1 U8072 ( .A1(n9760), .A2(n6475), .ZN(n6476) );
  OAI21_X1 U8073 ( .B1(n6476), .B2(n7711), .A(n6556), .ZN(n6477) );
  INV_X1 U8074 ( .A(n6477), .ZN(n9898) );
  INV_X1 U8075 ( .A(n6491), .ZN(n9887) );
  XNOR2_X1 U8076 ( .A(n9763), .B(n7882), .ZN(n6478) );
  NAND2_X1 U8077 ( .A1(n6478), .A2(n9500), .ZN(n9894) );
  OAI22_X1 U8078 ( .A1(n9788), .A2(n6479), .B1(n7883), .B2(n9792), .ZN(n6480)
         );
  AOI21_X1 U8079 ( .B1(n8380), .B2(n7882), .A(n6480), .ZN(n6481) );
  OAI21_X1 U8080 ( .B1(n9894), .B2(n9793), .A(n6481), .ZN(n6482) );
  AOI21_X1 U8081 ( .B1(n9898), .B2(n8143), .A(n6482), .ZN(n6483) );
  OAI21_X1 U8082 ( .B1(n8399), .B2(n9895), .A(n6483), .ZN(P2_U3285) );
  XNOR2_X1 U8083 ( .A(n6491), .B(n6486), .ZN(n6791) );
  NAND2_X1 U8084 ( .A1(n5560), .A2(n7933), .ZN(n6790) );
  XNOR2_X1 U8085 ( .A(n6791), .B(n6790), .ZN(n6792) );
  XNOR2_X1 U8086 ( .A(n6793), .B(n6792), .ZN(n6493) );
  OAI21_X1 U8087 ( .B1(n7922), .B2(n9783), .A(n6487), .ZN(n6490) );
  OAI22_X1 U8088 ( .A1(n7893), .A2(n6803), .B1(n6488), .B2(n7892), .ZN(n6489)
         );
  AOI211_X1 U8089 ( .C1(n6491), .C2(n7903), .A(n6490), .B(n6489), .ZN(n6492)
         );
  OAI21_X1 U8090 ( .B1(n6493), .B2(n7913), .A(n6492), .ZN(P2_U3219) );
  OAI21_X1 U8091 ( .B1(n6496), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6494), .ZN(
        n6509) );
  XNOR2_X1 U8092 ( .A(n6557), .B(n6576), .ZN(n6508) );
  XOR2_X1 U8093 ( .A(n6509), .B(n6508), .Z(n6506) );
  AOI21_X1 U8094 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n6496), .A(n6495), .ZN(
        n6499) );
  MUX2_X1 U8095 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6497), .S(n6557), .Z(n6498)
         );
  NAND2_X1 U8096 ( .A1(n6498), .A2(n6499), .ZN(n6515) );
  OAI21_X1 U8097 ( .B1(n6499), .B2(n6498), .A(n6515), .ZN(n6500) );
  INV_X1 U8098 ( .A(n6500), .ZN(n6503) );
  NAND2_X1 U8099 ( .A1(n9755), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6502) );
  AND2_X1 U8100 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6805) );
  INV_X1 U8101 ( .A(n6805), .ZN(n6501) );
  OAI211_X1 U8102 ( .C1(n6503), .C2(n9753), .A(n6502), .B(n6501), .ZN(n6504)
         );
  AOI21_X1 U8103 ( .B1(n9456), .B2(n6557), .A(n6504), .ZN(n6505) );
  OAI21_X1 U8104 ( .B1(n6506), .B2(n9449), .A(n6505), .ZN(P2_U3257) );
  AOI22_X1 U8105 ( .A1(n6509), .A2(n6508), .B1(n6507), .B2(n6576), .ZN(n6512)
         );
  INV_X1 U8106 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6510) );
  MUX2_X1 U8107 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n6510), .S(n6849), .Z(n6511)
         );
  OAI21_X1 U8108 ( .B1(n6512), .B2(n6511), .A(n9750), .ZN(n6521) );
  INV_X1 U8109 ( .A(n9755), .ZN(n7989) );
  INV_X1 U8110 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8111 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n6513) );
  OAI21_X1 U8112 ( .B1(n7989), .B2(n6514), .A(n6513), .ZN(n6519) );
  XNOR2_X1 U8113 ( .A(n6849), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n6517) );
  OAI21_X1 U8114 ( .B1(n6557), .B2(P2_REG1_REG_12__SCAN_IN), .A(n6515), .ZN(
        n6516) );
  NOR2_X1 U8115 ( .A1(n6516), .A2(n6517), .ZN(n6843) );
  AOI211_X1 U8116 ( .C1(n6517), .C2(n6516), .A(n6843), .B(n9753), .ZN(n6518)
         );
  AOI211_X1 U8117 ( .C1(n9456), .C2(n6849), .A(n6519), .B(n6518), .ZN(n6520)
         );
  OAI21_X1 U8118 ( .B1(n6521), .B2(n6848), .A(n6520), .ZN(P2_U3258) );
  OAI21_X1 U8119 ( .B1(n6522), .B2(n6527), .A(n6523), .ZN(n9853) );
  INV_X1 U8120 ( .A(n6527), .ZN(n6531) );
  INV_X1 U8121 ( .A(n6528), .ZN(n7703) );
  NAND2_X1 U8122 ( .A1(n7703), .A2(n7698), .ZN(n6529) );
  OAI211_X1 U8123 ( .C1(n6531), .C2(n6530), .A(n6529), .B(n9776), .ZN(n6533)
         );
  AOI22_X1 U8124 ( .A1(n9772), .A2(n5545), .B1(n7939), .B2(n9769), .ZN(n6532)
         );
  NAND2_X1 U8125 ( .A1(n6533), .A2(n6532), .ZN(n9852) );
  AOI22_X1 U8126 ( .A1(n6534), .A2(n9848), .B1(n9788), .B2(n9852), .ZN(n6535)
         );
  OAI21_X1 U8127 ( .B1(n9850), .B2(n9795), .A(n6535), .ZN(n6537) );
  OAI22_X1 U8128 ( .A1(n9792), .A2(n5474), .B1(n5473), .B2(n9788), .ZN(n6536)
         );
  AOI211_X1 U8129 ( .C1(n8143), .C2(n9853), .A(n6537), .B(n6536), .ZN(n6538)
         );
  INV_X1 U8130 ( .A(n6538), .ZN(P2_U3294) );
  INV_X1 U8131 ( .A(n6582), .ZN(n9460) );
  NAND2_X1 U8132 ( .A1(n6582), .A2(n7289), .ZN(n6540) );
  OR2_X1 U8133 ( .A1(n6679), .A2(n7283), .ZN(n6539) );
  NAND2_X1 U8134 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  XNOR2_X1 U8135 ( .A(n6541), .B(n7320), .ZN(n6663) );
  NOR2_X1 U8136 ( .A1(n6679), .A2(n7322), .ZN(n6542) );
  AOI21_X1 U8137 ( .B1(n6582), .B2(n4285), .A(n6542), .ZN(n6664) );
  XNOR2_X1 U8138 ( .A(n6663), .B(n6664), .ZN(n6547) );
  NAND2_X1 U8139 ( .A1(n6546), .A2(n6547), .ZN(n6673) );
  OAI21_X1 U8140 ( .B1(n6547), .B2(n6546), .A(n6545), .ZN(n6548) );
  NAND2_X1 U8141 ( .A1(n6548), .A2(n8657), .ZN(n6554) );
  INV_X1 U8142 ( .A(n8965), .ZN(n6599) );
  INV_X1 U8143 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6549) );
  OAI22_X1 U8144 ( .A1(n8664), .A2(n6599), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6549), .ZN(n6552) );
  NOR2_X1 U8145 ( .A1(n4275), .A2(n6550), .ZN(n6551) );
  AOI211_X1 U8146 ( .C1(n8666), .C2(n8966), .A(n6552), .B(n6551), .ZN(n6553)
         );
  OAI211_X1 U8147 ( .C1(n9460), .C2(n8656), .A(n6554), .B(n6553), .ZN(P1_U3215) );
  NAND2_X1 U8148 ( .A1(n7882), .A2(n9770), .ZN(n6555) );
  NAND2_X1 U8149 ( .A1(n6589), .A2(n6133), .ZN(n6559) );
  AOI22_X1 U8150 ( .A1(n7473), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5720), .B2(
        n6557), .ZN(n6558) );
  INV_X1 U8151 ( .A(n7932), .ZN(n6862) );
  NAND2_X1 U8152 ( .A1(n6836), .A2(n6862), .ZN(n7609) );
  OAI21_X1 U8153 ( .B1(n4372), .B2(n7712), .A(n6838), .ZN(n9906) );
  INV_X1 U8154 ( .A(n9906), .ZN(n6581) );
  INV_X1 U8155 ( .A(n7606), .ZN(n6560) );
  OAI211_X1 U8156 ( .C1(n4281), .C2(n4388), .A(n9776), .B(n6815), .ZN(n6573)
         );
  NAND2_X1 U8157 ( .A1(n7517), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6571) );
  INV_X1 U8158 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6563) );
  OR2_X1 U8159 ( .A1(n7522), .A2(n6563), .ZN(n6570) );
  INV_X1 U8160 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6564) );
  OAI21_X1 U8161 ( .B1(n6566), .B2(n6565), .A(n6564), .ZN(n6567) );
  NAND2_X1 U8162 ( .A1(n6567), .A2(n6820), .ZN(n7353) );
  OR2_X1 U8163 ( .A1(n4279), .A2(n7353), .ZN(n6569) );
  OR2_X1 U8164 ( .A1(n4277), .A2(n6510), .ZN(n6568) );
  NAND4_X1 U8165 ( .A1(n6571), .A2(n6570), .A3(n6569), .A4(n6568), .ZN(n7931)
         );
  AOI22_X1 U8166 ( .A1(n9772), .A2(n9770), .B1(n7931), .B2(n9769), .ZN(n6572)
         );
  NAND2_X1 U8167 ( .A1(n6573), .A2(n6572), .ZN(n9904) );
  INV_X1 U8168 ( .A(n7882), .ZN(n9896) );
  NAND2_X1 U8169 ( .A1(n6574), .A2(n6836), .ZN(n6575) );
  NAND2_X1 U8170 ( .A1(n7354), .A2(n6575), .ZN(n9903) );
  OAI22_X1 U8171 ( .A1(n9788), .A2(n6576), .B1(n6802), .B2(n9792), .ZN(n6577)
         );
  AOI21_X1 U8172 ( .B1(n8380), .B2(n6836), .A(n6577), .ZN(n6578) );
  OAI21_X1 U8173 ( .B1(n9903), .B2(n8014), .A(n6578), .ZN(n6579) );
  AOI21_X1 U8174 ( .B1(n9904), .B2(n9788), .A(n6579), .ZN(n6580) );
  OAI21_X1 U8175 ( .B1(n6581), .B2(n8362), .A(n6580), .ZN(P2_U3284) );
  INV_X1 U8176 ( .A(n6679), .ZN(n9597) );
  NAND2_X1 U8177 ( .A1(n6584), .A2(n6383), .ZN(n6586) );
  AOI22_X1 U8178 ( .A1(n7086), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7085), .B2(
        n9578), .ZN(n6585) );
  XNOR2_X1 U8179 ( .A(n6670), .B(n8965), .ZN(n8900) );
  NAND2_X1 U8180 ( .A1(n6670), .A2(n8965), .ZN(n6588) );
  NAND2_X1 U8181 ( .A1(n6646), .A2(n6588), .ZN(n6704) );
  NAND2_X1 U8182 ( .A1(n6589), .A2(n6383), .ZN(n6592) );
  AOI22_X1 U8183 ( .A1(n7086), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7085), .B2(
        n6590), .ZN(n6591) );
  NAND2_X2 U8184 ( .A1(n6592), .A2(n6591), .ZN(n9530) );
  NAND2_X1 U8185 ( .A1(n8678), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6597) );
  INV_X1 U8186 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6618) );
  OR2_X1 U8187 ( .A1(n4280), .A2(n6618), .ZN(n6596) );
  XNOR2_X1 U8188 ( .A(n6605), .B(n6604), .ZN(n6698) );
  OR2_X1 U8189 ( .A1(n7167), .A2(n6698), .ZN(n6595) );
  OR2_X1 U8190 ( .A1(n8683), .A2(n6593), .ZN(n6594) );
  NAND2_X1 U8191 ( .A1(n9530), .A2(n6687), .ZN(n8774) );
  NAND2_X1 U8192 ( .A1(n8781), .A2(n8774), .ZN(n8899) );
  INV_X1 U8193 ( .A(n8899), .ZN(n6711) );
  XNOR2_X1 U8194 ( .A(n6704), .B(n6711), .ZN(n9534) );
  NAND2_X1 U8195 ( .A1(n9534), .A2(n6890), .ZN(n6616) );
  OR2_X1 U8196 ( .A1(n6670), .A2(n6599), .ZN(n6598) );
  AND2_X1 U8197 ( .A1(n8782), .A2(n6598), .ZN(n6601) );
  NAND2_X1 U8198 ( .A1(n6670), .A2(n6599), .ZN(n6713) );
  XNOR2_X1 U8199 ( .A(n6712), .B(n8899), .ZN(n6614) );
  NAND2_X1 U8200 ( .A1(n8678), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6610) );
  OR2_X1 U8201 ( .A1(n8683), .A2(n6602), .ZN(n6609) );
  OAI21_X1 U8202 ( .B1(n6605), .B2(n6604), .A(n6603), .ZN(n6606) );
  NAND2_X1 U8203 ( .A1(n6606), .A2(n6721), .ZN(n6756) );
  OR2_X1 U8204 ( .A1(n7167), .A2(n6756), .ZN(n6608) );
  OR2_X1 U8205 ( .A1(n4280), .A2(n4936), .ZN(n6607) );
  NAND4_X1 U8206 ( .A1(n6610), .A2(n6609), .A3(n6608), .A4(n6607), .ZN(n8963)
         );
  NAND2_X1 U8207 ( .A1(n8963), .A2(n9649), .ZN(n6612) );
  NAND2_X1 U8208 ( .A1(n8965), .A2(n9614), .ZN(n6611) );
  NAND2_X1 U8209 ( .A1(n6612), .A2(n6611), .ZN(n6613) );
  AOI21_X1 U8210 ( .B1(n6614), .B2(n9617), .A(n6613), .ZN(n6615) );
  AND2_X1 U8211 ( .A1(n6616), .A2(n6615), .ZN(n9536) );
  INV_X1 U8212 ( .A(n6670), .ZN(n9539) );
  NAND2_X1 U8213 ( .A1(n6654), .A2(n9539), .ZN(n6653) );
  AOI21_X1 U8214 ( .B1(n6653), .B2(n9530), .A(n9295), .ZN(n6617) );
  NAND2_X1 U8215 ( .A1(n6617), .A2(n6732), .ZN(n9532) );
  OAI22_X1 U8216 ( .A1(n9641), .A2(n6618), .B1(n6698), .B2(n9306), .ZN(n6619)
         );
  AOI21_X1 U8217 ( .B1(n9530), .B2(n9620), .A(n6619), .ZN(n6620) );
  OAI21_X1 U8218 ( .B1(n9532), .B2(n9310), .A(n6620), .ZN(n6621) );
  AOI21_X1 U8219 ( .B1(n9534), .B2(n9639), .A(n6621), .ZN(n6622) );
  OAI21_X1 U8220 ( .B1(n9536), .B2(n9660), .A(n6622), .ZN(P1_U3279) );
  INV_X1 U8221 ( .A(n6624), .ZN(n6625) );
  INV_X1 U8222 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n6641) );
  INV_X1 U8223 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7100) );
  MUX2_X1 U8224 ( .A(n6641), .B(n7100), .S(n7532), .Z(n6628) );
  INV_X1 U8225 ( .A(SI_22_), .ZN(n6627) );
  NAND2_X1 U8226 ( .A1(n6628), .A2(n6627), .ZN(n6631) );
  INV_X1 U8227 ( .A(n6628), .ZN(n6629) );
  NAND2_X1 U8228 ( .A1(n6629), .A2(SI_22_), .ZN(n6630) );
  NAND2_X1 U8229 ( .A1(n6631), .A2(n6630), .ZN(n6639) );
  INV_X1 U8230 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n6632) );
  INV_X1 U8231 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7110) );
  MUX2_X1 U8232 ( .A(n6632), .B(n7110), .S(n7532), .Z(n6634) );
  INV_X1 U8233 ( .A(SI_23_), .ZN(n6633) );
  NAND2_X1 U8234 ( .A1(n6634), .A2(n6633), .ZN(n6762) );
  INV_X1 U8235 ( .A(n6634), .ZN(n6635) );
  NAND2_X1 U8236 ( .A1(n6635), .A2(SI_23_), .ZN(n6636) );
  XNOR2_X1 U8237 ( .A(n6761), .B(n6760), .ZN(n7417) );
  INV_X1 U8238 ( .A(n7417), .ZN(n6638) );
  AOI21_X1 U8239 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8525), .A(n7733), .ZN(
        n6637) );
  OAI21_X1 U8240 ( .B1(n6638), .B2(n7800), .A(n6637), .ZN(P2_U3335) );
  XNOR2_X1 U8241 ( .A(n6640), .B(n6639), .ZN(n7408) );
  INV_X1 U8242 ( .A(n7408), .ZN(n6643) );
  OAI222_X1 U8243 ( .A1(n6642), .A2(P2_U3152), .B1(n7800), .B2(n6643), .C1(
        n6641), .C2(n7817), .ZN(P2_U3336) );
  OAI222_X1 U8244 ( .A1(n7361), .A2(n7100), .B1(n7364), .B2(n6643), .C1(
        P1_U3084), .C2(n5212), .ZN(P1_U3331) );
  NAND2_X1 U8245 ( .A1(n6644), .A2(n8900), .ZN(n6645) );
  NAND2_X1 U8246 ( .A1(n6646), .A2(n6645), .ZN(n9537) );
  NAND2_X1 U8247 ( .A1(n6647), .A2(n8782), .ZN(n6648) );
  XNOR2_X1 U8248 ( .A(n6648), .B(n6587), .ZN(n6650) );
  OAI22_X1 U8249 ( .A1(n6679), .A2(n9291), .B1(n6687), .B2(n9293), .ZN(n6649)
         );
  AOI21_X1 U8250 ( .B1(n6650), .B2(n9617), .A(n6649), .ZN(n6651) );
  OAI21_X1 U8251 ( .B1(n9537), .B2(n9323), .A(n6651), .ZN(n9540) );
  NAND2_X1 U8252 ( .A1(n9540), .A2(n9641), .ZN(n6658) );
  OAI22_X1 U8253 ( .A1(n9641), .A2(n6652), .B1(n6676), .B2(n9306), .ZN(n6656)
         );
  OAI211_X1 U8254 ( .C1(n6654), .C2(n9539), .A(n6653), .B(n9625), .ZN(n9538)
         );
  NOR2_X1 U8255 ( .A1(n9538), .A2(n9310), .ZN(n6655) );
  AOI211_X1 U8256 ( .C1(n9620), .C2(n6670), .A(n6656), .B(n6655), .ZN(n6657)
         );
  OAI211_X1 U8257 ( .C1(n9537), .C2(n6659), .A(n6658), .B(n6657), .ZN(P1_U3280) );
  NAND2_X1 U8258 ( .A1(n7417), .A2(n6660), .ZN(n6662) );
  NAND2_X1 U8259 ( .A1(n6661), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8954) );
  OAI211_X1 U8260 ( .C1(n7110), .C2(n7361), .A(n6662), .B(n8954), .ZN(P1_U3330) );
  INV_X1 U8261 ( .A(n6663), .ZN(n6665) );
  NAND2_X1 U8262 ( .A1(n6665), .A2(n6664), .ZN(n6671) );
  AND2_X1 U8263 ( .A1(n6545), .A2(n6671), .ZN(n6675) );
  NAND2_X1 U8264 ( .A1(n6670), .A2(n7289), .ZN(n6667) );
  NAND2_X1 U8265 ( .A1(n8965), .A2(n4285), .ZN(n6666) );
  NAND2_X1 U8266 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  XNOR2_X1 U8267 ( .A(n6668), .B(n7320), .ZN(n6691) );
  AND2_X1 U8268 ( .A1(n8965), .A2(n7286), .ZN(n6669) );
  AOI21_X1 U8269 ( .B1(n6670), .B2(n4285), .A(n6669), .ZN(n6689) );
  XNOR2_X1 U8270 ( .A(n6691), .B(n6689), .ZN(n6674) );
  AND2_X1 U8271 ( .A1(n6674), .A2(n6671), .ZN(n6672) );
  OAI211_X1 U8272 ( .C1(n6675), .C2(n6674), .A(n8657), .B(n6695), .ZN(n6683)
         );
  INV_X1 U8273 ( .A(n6676), .ZN(n6681) );
  INV_X1 U8274 ( .A(n6687), .ZN(n8964) );
  INV_X1 U8275 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6677) );
  NOR2_X1 U8276 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6677), .ZN(n9577) );
  AOI21_X1 U8277 ( .B1(n8653), .B2(n8964), .A(n9577), .ZN(n6678) );
  OAI21_X1 U8278 ( .B1(n8650), .B2(n6679), .A(n6678), .ZN(n6680) );
  AOI21_X1 U8279 ( .B1(n6681), .B2(n8576), .A(n6680), .ZN(n6682) );
  OAI211_X1 U8280 ( .C1(n9539), .C2(n8656), .A(n6683), .B(n6682), .ZN(P1_U3234) );
  INV_X1 U8281 ( .A(n9530), .ZN(n6703) );
  NAND2_X1 U8282 ( .A1(n9530), .A2(n7289), .ZN(n6685) );
  OR2_X1 U8283 ( .A1(n6687), .A2(n7283), .ZN(n6684) );
  NAND2_X1 U8284 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  XNOR2_X1 U8285 ( .A(n6686), .B(n7320), .ZN(n6738) );
  NOR2_X1 U8286 ( .A1(n6687), .A2(n7322), .ZN(n6688) );
  AOI21_X1 U8287 ( .B1(n9530), .B2(n4285), .A(n6688), .ZN(n6739) );
  XNOR2_X1 U8288 ( .A(n6738), .B(n6739), .ZN(n6693) );
  INV_X1 U8289 ( .A(n6689), .ZN(n6690) );
  NAND2_X1 U8290 ( .A1(n6691), .A2(n6690), .ZN(n6694) );
  AND2_X1 U8291 ( .A1(n6693), .A2(n6694), .ZN(n6692) );
  INV_X1 U8292 ( .A(n6742), .ZN(n6697) );
  AOI21_X1 U8293 ( .B1(n6695), .B2(n6694), .A(n6693), .ZN(n6696) );
  OAI21_X1 U8294 ( .B1(n6697), .B2(n6696), .A(n8657), .ZN(n6702) );
  INV_X1 U8295 ( .A(n8963), .ZN(n6710) );
  OAI22_X1 U8296 ( .A1(n8664), .A2(n6710), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6604), .ZN(n6700) );
  NOR2_X1 U8297 ( .A1(n4275), .A2(n6698), .ZN(n6699) );
  AOI211_X1 U8298 ( .C1(n8666), .C2(n8965), .A(n6700), .B(n6699), .ZN(n6701)
         );
  OAI211_X1 U8299 ( .C1(n6703), .C2(n8656), .A(n6702), .B(n6701), .ZN(P1_U3222) );
  NAND2_X1 U8300 ( .A1(n6704), .A2(n8899), .ZN(n6706) );
  NAND2_X1 U8301 ( .A1(n9530), .A2(n8964), .ZN(n6705) );
  NAND2_X1 U8302 ( .A1(n6706), .A2(n6705), .ZN(n6767) );
  NAND2_X1 U8303 ( .A1(n6812), .A2(n6383), .ZN(n6709) );
  AOI22_X1 U8304 ( .A1(n7086), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7085), .B2(
        n6707), .ZN(n6708) );
  OR2_X1 U8305 ( .A1(n9523), .A2(n6710), .ZN(n8797) );
  NAND2_X1 U8306 ( .A1(n9523), .A2(n6710), .ZN(n8788) );
  XNOR2_X1 U8307 ( .A(n6767), .B(n8902), .ZN(n9527) );
  NAND2_X1 U8308 ( .A1(n6712), .A2(n6711), .ZN(n6718) );
  OR2_X1 U8309 ( .A1(n8899), .A2(n6587), .ZN(n6714) );
  NAND2_X1 U8310 ( .A1(n8774), .A2(n6713), .ZN(n8699) );
  NAND2_X1 U8311 ( .A1(n8699), .A2(n8781), .ZN(n8789) );
  NAND2_X1 U8312 ( .A1(n6718), .A2(n8786), .ZN(n6716) );
  INV_X1 U8313 ( .A(n8902), .ZN(n6715) );
  NAND2_X1 U8314 ( .A1(n6716), .A2(n6715), .ZN(n6719) );
  AND2_X1 U8315 ( .A1(n8902), .A2(n8786), .ZN(n6717) );
  NAND2_X1 U8316 ( .A1(n6718), .A2(n6717), .ZN(n6772) );
  NAND2_X1 U8317 ( .A1(n6719), .A2(n6772), .ZN(n6720) );
  NAND2_X1 U8318 ( .A1(n6720), .A2(n9617), .ZN(n6729) );
  NAND2_X1 U8319 ( .A1(n8678), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6727) );
  OR2_X1 U8320 ( .A1(n8683), .A2(n9522), .ZN(n6726) );
  INV_X1 U8321 ( .A(n6775), .ZN(n6723) );
  NAND2_X1 U8322 ( .A1(n6721), .A2(n8208), .ZN(n6722) );
  NAND2_X1 U8323 ( .A1(n6723), .A2(n6722), .ZN(n8545) );
  OR2_X1 U8324 ( .A1(n7167), .A2(n8545), .ZN(n6725) );
  OR2_X1 U8325 ( .A1(n4280), .A2(n6158), .ZN(n6724) );
  NAND4_X1 U8326 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .ZN(n8962)
         );
  AOI22_X1 U8327 ( .A1(n8964), .A2(n9614), .B1(n9649), .B2(n8962), .ZN(n6728)
         );
  NAND2_X1 U8328 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  AOI21_X1 U8329 ( .B1(n9527), .B2(n6890), .A(n6730), .ZN(n9529) );
  NAND2_X1 U8330 ( .A1(n6732), .A2(n9523), .ZN(n6731) );
  NAND2_X1 U8331 ( .A1(n6731), .A2(n9625), .ZN(n6733) );
  OR2_X1 U8332 ( .A1(n6733), .A2(n6784), .ZN(n9524) );
  OAI22_X1 U8333 ( .A1(n9641), .A2(n4936), .B1(n6756), .B2(n9306), .ZN(n6734)
         );
  AOI21_X1 U8334 ( .B1(n9523), .B2(n9620), .A(n6734), .ZN(n6735) );
  OAI21_X1 U8335 ( .B1(n9524), .B2(n9310), .A(n6735), .ZN(n6736) );
  AOI21_X1 U8336 ( .B1(n9527), .B2(n9639), .A(n6736), .ZN(n6737) );
  OAI21_X1 U8337 ( .B1(n9529), .B2(n9660), .A(n6737), .ZN(P1_U3278) );
  INV_X1 U8338 ( .A(n6738), .ZN(n6740) );
  NAND2_X1 U8339 ( .A1(n6740), .A2(n6739), .ZN(n6741) );
  NAND2_X1 U8340 ( .A1(n9523), .A2(n7289), .ZN(n6744) );
  NAND2_X1 U8341 ( .A1(n8963), .A2(n4285), .ZN(n6743) );
  NAND2_X1 U8342 ( .A1(n6744), .A2(n6743), .ZN(n6745) );
  XNOR2_X1 U8343 ( .A(n6745), .B(n5653), .ZN(n6747) );
  AND2_X1 U8344 ( .A1(n8963), .A2(n7286), .ZN(n6746) );
  AOI21_X1 U8345 ( .B1(n9523), .B2(n4285), .A(n6746), .ZN(n6748) );
  AND2_X1 U8346 ( .A1(n6747), .A2(n6748), .ZN(n7216) );
  INV_X1 U8347 ( .A(n7216), .ZN(n6751) );
  INV_X1 U8348 ( .A(n6747), .ZN(n6750) );
  INV_X1 U8349 ( .A(n6748), .ZN(n6749) );
  NAND2_X1 U8350 ( .A1(n6750), .A2(n6749), .ZN(n7215) );
  NAND2_X1 U8351 ( .A1(n6751), .A2(n7215), .ZN(n6752) );
  XNOR2_X1 U8352 ( .A(n7217), .B(n6752), .ZN(n6759) );
  INV_X1 U8353 ( .A(n8962), .ZN(n8695) );
  OAI21_X1 U8354 ( .B1(n8664), .B2(n8695), .A(n6753), .ZN(n6754) );
  AOI21_X1 U8355 ( .B1(n8666), .B2(n8964), .A(n6754), .ZN(n6755) );
  OAI21_X1 U8356 ( .B1(n4275), .B2(n6756), .A(n6755), .ZN(n6757) );
  AOI21_X1 U8357 ( .B1(n9523), .B2(n8671), .A(n6757), .ZN(n6758) );
  OAI21_X1 U8358 ( .B1(n6759), .B2(n8645), .A(n6758), .ZN(P1_U3232) );
  NAND2_X1 U8359 ( .A1(n6761), .A2(n6760), .ZN(n6763) );
  INV_X1 U8360 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n6809) );
  INV_X1 U8361 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7122) );
  MUX2_X1 U8362 ( .A(n6809), .B(n7122), .S(n7532), .Z(n6897) );
  XNOR2_X1 U8363 ( .A(n6897), .B(SI_24_), .ZN(n6896) );
  XNOR2_X1 U8364 ( .A(n6901), .B(n6896), .ZN(n7424) );
  INV_X1 U8365 ( .A(n7424), .ZN(n6810) );
  OAI222_X1 U8366 ( .A1(n7364), .A2(n6810), .B1(n6764), .B2(P1_U3084), .C1(
        n7122), .C2(n7361), .ZN(P1_U3329) );
  AND2_X1 U8367 ( .A1(n9523), .A2(n8963), .ZN(n6766) );
  OR2_X1 U8368 ( .A1(n9523), .A2(n8963), .ZN(n6765) );
  NAND2_X1 U8369 ( .A1(n6816), .A2(n6383), .ZN(n6770) );
  AOI22_X1 U8370 ( .A1(n7086), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7085), .B2(
        n6768), .ZN(n6769) );
  XNOR2_X1 U8371 ( .A(n8696), .B(n8695), .ZN(n8904) );
  XNOR2_X1 U8372 ( .A(n6868), .B(n8904), .ZN(n9521) );
  INV_X1 U8373 ( .A(n9521), .ZN(n6789) );
  AND2_X1 U8374 ( .A1(n6772), .A2(n8788), .ZN(n6774) );
  INV_X1 U8375 ( .A(n8904), .ZN(n6773) );
  AND2_X1 U8376 ( .A1(n6773), .A2(n8788), .ZN(n6771) );
  NAND2_X1 U8377 ( .A1(n6772), .A2(n6771), .ZN(n6876) );
  OAI211_X1 U8378 ( .C1(n6774), .C2(n6773), .A(n9617), .B(n6876), .ZN(n6782)
         );
  NAND2_X1 U8379 ( .A1(n8678), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6780) );
  OR2_X1 U8380 ( .A1(n8683), .A2(n9516), .ZN(n6779) );
  OR2_X1 U8381 ( .A1(n6775), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8382 ( .A1(n6881), .A2(n6776), .ZN(n8668) );
  OR2_X1 U8383 ( .A1(n7167), .A2(n8668), .ZN(n6778) );
  OR2_X1 U8384 ( .A1(n4280), .A2(n8200), .ZN(n6777) );
  NAND4_X1 U8385 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n9303)
         );
  AOI22_X1 U8386 ( .A1(n9614), .A2(n8963), .B1(n9303), .B2(n9649), .ZN(n6781)
         );
  NAND2_X1 U8387 ( .A1(n6782), .A2(n6781), .ZN(n9519) );
  INV_X1 U8388 ( .A(n6891), .ZN(n6783) );
  OAI211_X1 U8389 ( .C1(n9518), .C2(n6784), .A(n6783), .B(n9625), .ZN(n9517)
         );
  OAI22_X1 U8390 ( .A1(n9641), .A2(n6158), .B1(n8545), .B2(n9306), .ZN(n6785)
         );
  AOI21_X1 U8391 ( .B1(n8696), .B2(n9620), .A(n6785), .ZN(n6786) );
  OAI21_X1 U8392 ( .B1(n9517), .B2(n9310), .A(n6786), .ZN(n6787) );
  AOI21_X1 U8393 ( .B1(n9519), .B2(n9641), .A(n6787), .ZN(n6788) );
  OAI21_X1 U8394 ( .B1(n6789), .B2(n9301), .A(n6788), .ZN(P1_U3277) );
  INV_X1 U8395 ( .A(n6836), .ZN(n9901) );
  OAI22_X1 U8396 ( .A1(n6793), .A2(n6792), .B1(n6791), .B2(n6790), .ZN(n7877)
         );
  XNOR2_X1 U8397 ( .A(n7882), .B(n5554), .ZN(n6795) );
  NAND2_X1 U8398 ( .A1(n5560), .A2(n9770), .ZN(n6794) );
  XNOR2_X1 U8399 ( .A(n6795), .B(n6794), .ZN(n7878) );
  INV_X1 U8400 ( .A(n6794), .ZN(n6796) );
  AND2_X1 U8401 ( .A1(n5560), .A2(n7932), .ZN(n6798) );
  XNOR2_X1 U8402 ( .A(n6836), .B(n5554), .ZN(n6797) );
  NOR2_X1 U8403 ( .A1(n6797), .A2(n6798), .ZN(n6859) );
  AOI21_X1 U8404 ( .B1(n6798), .B2(n6797), .A(n6859), .ZN(n6799) );
  NAND2_X1 U8405 ( .A1(n6800), .A2(n6799), .ZN(n6861) );
  OAI21_X1 U8406 ( .B1(n6800), .B2(n6799), .A(n6861), .ZN(n6801) );
  NAND2_X1 U8407 ( .A1(n6801), .A2(n7901), .ZN(n6808) );
  INV_X1 U8408 ( .A(n6802), .ZN(n6806) );
  OAI22_X1 U8409 ( .A1(n7893), .A2(n6932), .B1(n6803), .B2(n7892), .ZN(n6804)
         );
  AOI211_X1 U8410 ( .C1(n7885), .C2(n6806), .A(n6805), .B(n6804), .ZN(n6807)
         );
  OAI211_X1 U8411 ( .C1(n9901), .C2(n7927), .A(n6808), .B(n6807), .ZN(P2_U3226) );
  OAI222_X1 U8412 ( .A1(P2_U3152), .A2(n6811), .B1(n7800), .B2(n6810), .C1(
        n6809), .C2(n7817), .ZN(P2_U3334) );
  NAND2_X1 U8413 ( .A1(n6812), .A2(n6133), .ZN(n6814) );
  AOI22_X1 U8414 ( .A1(n7473), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5720), .B2(
        n6849), .ZN(n6813) );
  XNOR2_X1 U8415 ( .A(n8495), .B(n6932), .ZN(n7714) );
  NAND2_X1 U8416 ( .A1(n6816), .A2(n6133), .ZN(n6818) );
  AOI22_X1 U8417 ( .A1(n5720), .A2(n6959), .B1(n7473), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U8418 ( .A1(n6027), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6825) );
  INV_X1 U8419 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6844) );
  OR2_X1 U8420 ( .A1(n6985), .A2(n6844), .ZN(n6824) );
  INV_X1 U8421 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U8422 ( .A1(n6820), .A2(n8259), .ZN(n6821) );
  NAND2_X1 U8423 ( .A1(n6981), .A2(n6821), .ZN(n6931) );
  OR2_X1 U8424 ( .A1(n4279), .A2(n6931), .ZN(n6823) );
  INV_X1 U8425 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6833) );
  OR2_X1 U8426 ( .A1(n4277), .A2(n6833), .ZN(n6822) );
  NAND4_X1 U8427 ( .A1(n6825), .A2(n6824), .A3(n6823), .A4(n6822), .ZN(n7930)
         );
  INV_X1 U8428 ( .A(n7930), .ZN(n7001) );
  XNOR2_X1 U8429 ( .A(n8488), .B(n7001), .ZN(n6840) );
  INV_X1 U8430 ( .A(n6840), .ZN(n7715) );
  OAI211_X1 U8431 ( .C1(n6826), .C2(n7715), .A(n6978), .B(n9776), .ZN(n6832)
         );
  NAND2_X1 U8432 ( .A1(n7517), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6830) );
  INV_X1 U8433 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6960) );
  OR2_X1 U8434 ( .A1(n6985), .A2(n6960), .ZN(n6829) );
  INV_X1 U8435 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6999) );
  XNOR2_X1 U8436 ( .A(n6981), .B(n6999), .ZN(n7000) );
  OR2_X1 U8437 ( .A1(n4279), .A2(n7000), .ZN(n6828) );
  INV_X1 U8438 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8271) );
  OR2_X1 U8439 ( .A1(n4278), .A2(n8271), .ZN(n6827) );
  NAND4_X1 U8440 ( .A1(n6830), .A2(n6829), .A3(n6828), .A4(n6827), .ZN(n8020)
         );
  AOI22_X1 U8441 ( .A1(n9772), .A2(n7931), .B1(n8020), .B2(n9769), .ZN(n6831)
         );
  AND2_X1 U8442 ( .A1(n6832), .A2(n6831), .ZN(n8492) );
  XNOR2_X1 U8443 ( .A(n7355), .B(n8488), .ZN(n8490) );
  INV_X1 U8444 ( .A(n8488), .ZN(n6973) );
  NOR2_X1 U8445 ( .A1(n6973), .A2(n9795), .ZN(n6835) );
  OAI22_X1 U8446 ( .A1(n9788), .A2(n6833), .B1(n6931), .B2(n9792), .ZN(n6834)
         );
  AOI211_X1 U8447 ( .C1(n8490), .C2(n9767), .A(n6835), .B(n6834), .ZN(n6842)
         );
  OR2_X1 U8448 ( .A1(n6836), .A2(n7932), .ZN(n6837) );
  NAND2_X1 U8449 ( .A1(n8495), .A2(n7931), .ZN(n7615) );
  NAND2_X1 U8450 ( .A1(n6839), .A2(n6840), .ZN(n6967) );
  OAI21_X1 U8451 ( .B1(n6839), .B2(n6840), .A(n6967), .ZN(n8487) );
  NAND2_X1 U8452 ( .A1(n8487), .A2(n8143), .ZN(n6841) );
  OAI211_X1 U8453 ( .C1(n8492), .C2(n8399), .A(n6842), .B(n6841), .ZN(P2_U3282) );
  AOI22_X1 U8454 ( .A1(n6959), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n6844), .B2(
        n6854), .ZN(n6845) );
  NAND2_X1 U8455 ( .A1(n6846), .A2(n6845), .ZN(n6958) );
  OAI21_X1 U8456 ( .B1(n6846), .B2(n6845), .A(n6958), .ZN(n6847) );
  INV_X1 U8457 ( .A(n6847), .ZN(n6858) );
  NOR2_X1 U8458 ( .A1(n6959), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6850) );
  AOI21_X1 U8459 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6959), .A(n6850), .ZN(
        n6851) );
  OAI21_X1 U8460 ( .B1(n6852), .B2(n6851), .A(n6953), .ZN(n6856) );
  NOR2_X1 U8461 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8259), .ZN(n6934) );
  AOI21_X1 U8462 ( .B1(n9755), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n6934), .ZN(
        n6853) );
  OAI21_X1 U8463 ( .B1(n9751), .B2(n6854), .A(n6853), .ZN(n6855) );
  AOI21_X1 U8464 ( .B1(n6856), .B2(n9750), .A(n6855), .ZN(n6857) );
  OAI21_X1 U8465 ( .B1(n6858), .B2(n9753), .A(n6857), .ZN(P2_U3259) );
  INV_X1 U8466 ( .A(n6859), .ZN(n6860) );
  XNOR2_X1 U8467 ( .A(n8495), .B(n5554), .ZN(n6925) );
  NAND2_X1 U8468 ( .A1(n5560), .A2(n7931), .ZN(n6923) );
  XNOR2_X1 U8469 ( .A(n6925), .B(n6923), .ZN(n6926) );
  XNOR2_X1 U8470 ( .A(n6927), .B(n6926), .ZN(n6866) );
  OAI22_X1 U8471 ( .A1(n7922), .A2(n7353), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6564), .ZN(n6864) );
  OAI22_X1 U8472 ( .A1(n7893), .A2(n7001), .B1(n6862), .B2(n7892), .ZN(n6863)
         );
  AOI211_X1 U8473 ( .C1(n8495), .C2(n7903), .A(n6864), .B(n6863), .ZN(n6865)
         );
  OAI21_X1 U8474 ( .B1(n6866), .B2(n7913), .A(n6865), .ZN(P2_U3236) );
  NOR2_X1 U8475 ( .A1(n8696), .A2(n8962), .ZN(n6867) );
  NAND2_X1 U8476 ( .A1(n6968), .A2(n6383), .ZN(n6871) );
  INV_X1 U8477 ( .A(n9048), .ZN(n6869) );
  AOI22_X1 U8478 ( .A1(n7086), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7085), .B2(
        n6869), .ZN(n6870) );
  INV_X1 U8479 ( .A(n9303), .ZN(n8544) );
  OR2_X1 U8480 ( .A1(n8672), .A2(n8544), .ZN(n8806) );
  NAND2_X1 U8481 ( .A1(n8672), .A2(n8544), .ZN(n8805) );
  NAND2_X1 U8482 ( .A1(n8806), .A2(n8805), .ZN(n6874) );
  INV_X1 U8483 ( .A(n6874), .ZN(n8903) );
  XNOR2_X1 U8484 ( .A(n7079), .B(n8903), .ZN(n9513) );
  AND2_X1 U8485 ( .A1(n9518), .A2(n8962), .ZN(n8801) );
  INV_X1 U8486 ( .A(n8801), .ZN(n6872) );
  NAND2_X1 U8487 ( .A1(n6876), .A2(n6872), .ZN(n6873) );
  NAND2_X1 U8488 ( .A1(n6873), .A2(n6874), .ZN(n6877) );
  NOR2_X1 U8489 ( .A1(n6874), .A2(n8801), .ZN(n6875) );
  NAND2_X1 U8490 ( .A1(n6877), .A2(n7197), .ZN(n6878) );
  NAND2_X1 U8491 ( .A1(n6878), .A2(n9617), .ZN(n6888) );
  NAND2_X1 U8492 ( .A1(n5255), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6886) );
  INV_X1 U8493 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6879) );
  OR2_X1 U8494 ( .A1(n5528), .A2(n6879), .ZN(n6885) );
  NAND2_X1 U8495 ( .A1(n6881), .A2(n6880), .ZN(n6882) );
  NAND2_X1 U8496 ( .A1(n7070), .A2(n6882), .ZN(n9307) );
  OR2_X1 U8497 ( .A1(n7167), .A2(n9307), .ZN(n6884) );
  INV_X1 U8498 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9308) );
  OR2_X1 U8499 ( .A1(n4280), .A2(n9308), .ZN(n6883) );
  INV_X1 U8500 ( .A(n9290), .ZN(n8961) );
  AOI22_X1 U8501 ( .A1(n8961), .A2(n9649), .B1(n9614), .B2(n8962), .ZN(n6887)
         );
  NAND2_X1 U8502 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  AOI21_X1 U8503 ( .B1(n9513), .B2(n6890), .A(n6889), .ZN(n9515) );
  OAI211_X1 U8504 ( .C1(n6891), .C2(n9511), .A(n9625), .B(n9309), .ZN(n9510)
         );
  OAI22_X1 U8505 ( .A1(n9641), .A2(n8200), .B1(n8668), .B2(n9306), .ZN(n6892)
         );
  AOI21_X1 U8506 ( .B1(n8672), .B2(n9620), .A(n6892), .ZN(n6893) );
  OAI21_X1 U8507 ( .B1(n9510), .B2(n9310), .A(n6893), .ZN(n6894) );
  AOI21_X1 U8508 ( .B1(n9513), .B2(n9639), .A(n6894), .ZN(n6895) );
  OAI21_X1 U8509 ( .B1(n9515), .B2(n9660), .A(n6895), .ZN(P1_U3276) );
  INV_X1 U8510 ( .A(n6896), .ZN(n6900) );
  INV_X1 U8511 ( .A(n6897), .ZN(n6898) );
  NAND2_X1 U8512 ( .A1(n6898), .A2(SI_24_), .ZN(n6899) );
  INV_X1 U8513 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n6905) );
  INV_X1 U8514 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7131) );
  MUX2_X1 U8515 ( .A(n6905), .B(n7131), .S(n7532), .Z(n6902) );
  INV_X1 U8516 ( .A(SI_25_), .ZN(n8221) );
  NAND2_X1 U8517 ( .A1(n6902), .A2(n8221), .ZN(n6909) );
  INV_X1 U8518 ( .A(n6902), .ZN(n6903) );
  NAND2_X1 U8519 ( .A1(n6903), .A2(SI_25_), .ZN(n6904) );
  NAND2_X1 U8520 ( .A1(n6909), .A2(n6904), .ZN(n6910) );
  INV_X1 U8521 ( .A(n7436), .ZN(n6908) );
  OAI222_X1 U8522 ( .A1(n6906), .A2(P2_U3152), .B1(n7800), .B2(n6908), .C1(
        n6905), .C2(n7817), .ZN(P2_U3333) );
  OAI222_X1 U8523 ( .A1(n7361), .A2(n7131), .B1(n9417), .B2(n6908), .C1(
        P1_U3084), .C2(n6907), .ZN(P1_U3328) );
  INV_X1 U8524 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6919) );
  INV_X1 U8525 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7335) );
  MUX2_X1 U8526 ( .A(n6919), .B(n7335), .S(n7532), .Z(n6913) );
  INV_X1 U8527 ( .A(SI_26_), .ZN(n6912) );
  NAND2_X1 U8528 ( .A1(n6913), .A2(n6912), .ZN(n6938) );
  INV_X1 U8529 ( .A(n6913), .ZN(n6914) );
  NAND2_X1 U8530 ( .A1(n6914), .A2(SI_26_), .ZN(n6915) );
  AND2_X1 U8531 ( .A1(n6938), .A2(n6915), .ZN(n6916) );
  OR2_X1 U8532 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  NAND2_X1 U8533 ( .A1(n6939), .A2(n6918), .ZN(n7450) );
  INV_X1 U8534 ( .A(n7450), .ZN(n7334) );
  OAI222_X1 U8535 ( .A1(n6920), .A2(P2_U3152), .B1(n7800), .B2(n7334), .C1(
        n6919), .C2(n7817), .ZN(P2_U3332) );
  AND2_X1 U8536 ( .A1(n5560), .A2(n7930), .ZN(n6922) );
  XNOR2_X1 U8537 ( .A(n8488), .B(n5554), .ZN(n6921) );
  NOR2_X1 U8538 ( .A1(n6921), .A2(n6922), .ZN(n6995) );
  AOI21_X1 U8539 ( .B1(n6922), .B2(n6921), .A(n6995), .ZN(n6929) );
  INV_X1 U8540 ( .A(n6923), .ZN(n6924) );
  OAI21_X1 U8541 ( .B1(n6929), .B2(n6928), .A(n6996), .ZN(n6930) );
  NAND2_X1 U8542 ( .A1(n6930), .A2(n7901), .ZN(n6937) );
  INV_X1 U8543 ( .A(n6931), .ZN(n6935) );
  INV_X1 U8544 ( .A(n8020), .ZN(n8387) );
  OAI22_X1 U8545 ( .A1(n7893), .A2(n8387), .B1(n6932), .B2(n7892), .ZN(n6933)
         );
  AOI211_X1 U8546 ( .C1(n7885), .C2(n6935), .A(n6934), .B(n6933), .ZN(n6936)
         );
  OAI211_X1 U8547 ( .C1(n6973), .C2(n7927), .A(n6937), .B(n6936), .ZN(P2_U3217) );
  INV_X1 U8548 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6947) );
  INV_X1 U8549 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8267) );
  MUX2_X1 U8550 ( .A(n6947), .B(n8267), .S(n7532), .Z(n6941) );
  INV_X1 U8551 ( .A(SI_27_), .ZN(n6940) );
  NAND2_X1 U8552 ( .A1(n6941), .A2(n6940), .ZN(n7184) );
  INV_X1 U8553 ( .A(n6941), .ZN(n6942) );
  NAND2_X1 U8554 ( .A1(n6942), .A2(SI_27_), .ZN(n6943) );
  AND2_X1 U8555 ( .A1(n7184), .A2(n6943), .ZN(n7180) );
  INV_X1 U8556 ( .A(n7462), .ZN(n6948) );
  AOI21_X1 U8557 ( .B1(n6945), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n6944), .ZN(
        n6946) );
  OAI21_X1 U8558 ( .B1(n6948), .B2(n9417), .A(n6946), .ZN(P1_U3326) );
  OAI222_X1 U8559 ( .A1(P2_U3152), .A2(n8009), .B1(n7800), .B2(n6948), .C1(
        n6947), .C2(n7817), .ZN(P2_U3331) );
  INV_X1 U8560 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6949) );
  INV_X1 U8561 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7344) );
  MUX2_X1 U8562 ( .A(n6949), .B(n7344), .S(n7532), .Z(n7177) );
  XNOR2_X1 U8563 ( .A(n7177), .B(SI_28_), .ZN(n7178) );
  INV_X1 U8564 ( .A(n7472), .ZN(n7345) );
  NAND2_X1 U8565 ( .A1(n8525), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6951) );
  OAI211_X1 U8566 ( .C1(n7345), .C2(n7800), .A(n6952), .B(n6951), .ZN(P2_U3330) );
  NAND2_X1 U8567 ( .A1(n6954), .A2(n8271), .ZN(n7954) );
  OAI21_X1 U8568 ( .B1(n6954), .B2(n8271), .A(n7954), .ZN(n6964) );
  INV_X1 U8569 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6957) );
  OR2_X1 U8570 ( .A1(n9751), .A2(n7953), .ZN(n6956) );
  NAND2_X1 U8571 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n6955) );
  OAI211_X1 U8572 ( .C1(n6957), .C2(n7989), .A(n6956), .B(n6955), .ZN(n6963)
         );
  OAI21_X1 U8573 ( .B1(n6959), .B2(P2_REG1_REG_14__SCAN_IN), .A(n6958), .ZN(
        n7943) );
  XNOR2_X1 U8574 ( .A(n7943), .B(n7953), .ZN(n6961) );
  NOR2_X1 U8575 ( .A1(n6960), .A2(n6961), .ZN(n7944) );
  AOI211_X1 U8576 ( .C1(n6961), .C2(n6960), .A(n7944), .B(n9753), .ZN(n6962)
         );
  AOI211_X1 U8577 ( .C1(n9750), .C2(n6964), .A(n6963), .B(n6962), .ZN(n6965)
         );
  INV_X1 U8578 ( .A(n6965), .ZN(P2_U3260) );
  OR2_X1 U8579 ( .A1(n8488), .A2(n7930), .ZN(n6966) );
  NAND2_X1 U8580 ( .A1(n6968), .A2(n6133), .ZN(n6972) );
  OAI22_X1 U8581 ( .A1(n7953), .A2(n5466), .B1(n4288), .B2(n6969), .ZN(n6970)
         );
  INV_X1 U8582 ( .A(n6970), .ZN(n6971) );
  NAND2_X1 U8583 ( .A1(n8482), .A2(n8387), .ZN(n7634) );
  NAND2_X1 U8584 ( .A1(n7630), .A2(n7634), .ZN(n8022) );
  XNOR2_X1 U8585 ( .A(n8023), .B(n7717), .ZN(n8486) );
  INV_X1 U8586 ( .A(n8482), .ZN(n6977) );
  INV_X1 U8587 ( .A(n8393), .ZN(n6974) );
  AOI21_X1 U8588 ( .B1(n8482), .B2(n4369), .A(n6974), .ZN(n8483) );
  INV_X1 U8589 ( .A(n7000), .ZN(n6975) );
  AOI22_X1 U8590 ( .A1(n8399), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n6975), .B2(
        n8397), .ZN(n6976) );
  OAI21_X1 U8591 ( .B1(n6977), .B2(n9795), .A(n6976), .ZN(n6993) );
  NAND2_X1 U8592 ( .A1(n6979), .A2(n7717), .ZN(n7365) );
  OAI211_X1 U8593 ( .C1(n6979), .C2(n7717), .A(n7365), .B(n9776), .ZN(n6991)
         );
  NAND2_X1 U8594 ( .A1(n7490), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6989) );
  INV_X1 U8595 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8283) );
  OR2_X1 U8596 ( .A1(n7392), .A2(n8283), .ZN(n6988) );
  INV_X1 U8597 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6980) );
  OAI21_X1 U8598 ( .B1(n6981), .B2(n6999), .A(n6980), .ZN(n6984) );
  AND2_X1 U8599 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n6982) );
  NAND2_X1 U8600 ( .A1(n6984), .A2(n7018), .ZN(n8396) );
  OR2_X1 U8601 ( .A1(n4279), .A2(n8396), .ZN(n6987) );
  INV_X1 U8602 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7946) );
  OR2_X1 U8603 ( .A1(n6985), .A2(n7946), .ZN(n6986) );
  NAND4_X1 U8604 ( .A1(n6989), .A2(n6988), .A3(n6987), .A4(n6986), .ZN(n7929)
         );
  AOI22_X1 U8605 ( .A1(n9772), .A2(n7930), .B1(n7929), .B2(n9769), .ZN(n6990)
         );
  AND2_X1 U8606 ( .A1(n6991), .A2(n6990), .ZN(n8485) );
  NOR2_X1 U8607 ( .A1(n8485), .A2(n8399), .ZN(n6992) );
  AOI211_X1 U8608 ( .C1(n8483), .C2(n9767), .A(n6993), .B(n6992), .ZN(n6994)
         );
  OAI21_X1 U8609 ( .B1(n8486), .B2(n8362), .A(n6994), .ZN(P2_U3281) );
  XNOR2_X1 U8610 ( .A(n8482), .B(n6486), .ZN(n7034) );
  NOR2_X1 U8611 ( .A1(n7031), .A2(n7034), .ZN(n7008) );
  INV_X1 U8612 ( .A(n7008), .ZN(n6997) );
  NAND2_X1 U8613 ( .A1(n7031), .A2(n7034), .ZN(n7006) );
  NAND2_X1 U8614 ( .A1(n6997), .A2(n7006), .ZN(n6998) );
  NAND2_X1 U8615 ( .A1(n5560), .A2(n8020), .ZN(n7033) );
  XNOR2_X1 U8616 ( .A(n6998), .B(n7033), .ZN(n7005) );
  OAI22_X1 U8617 ( .A1(n7922), .A2(n7000), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6999), .ZN(n7003) );
  INV_X1 U8618 ( .A(n7929), .ZN(n8372) );
  OAI22_X1 U8619 ( .A1(n7893), .A2(n8372), .B1(n7001), .B2(n7892), .ZN(n7002)
         );
  AOI211_X1 U8620 ( .C1(n8482), .C2(n7903), .A(n7003), .B(n7002), .ZN(n7004)
         );
  OAI21_X1 U8621 ( .B1(n7005), .B2(n7913), .A(n7004), .ZN(P2_U3243) );
  INV_X1 U8622 ( .A(n7033), .ZN(n7007) );
  OAI21_X1 U8623 ( .B1(n7008), .B2(n7007), .A(n7006), .ZN(n7016) );
  NAND2_X1 U8624 ( .A1(n7080), .A2(n6133), .ZN(n7010) );
  AOI22_X1 U8625 ( .A1(n7473), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7972), .B2(
        n5720), .ZN(n7009) );
  XNOR2_X1 U8626 ( .A(n8477), .B(n5554), .ZN(n7011) );
  AND2_X1 U8627 ( .A1(n5560), .A2(n7929), .ZN(n7012) );
  NAND2_X1 U8628 ( .A1(n7011), .A2(n7012), .ZN(n7032) );
  INV_X1 U8629 ( .A(n7011), .ZN(n7014) );
  INV_X1 U8630 ( .A(n7012), .ZN(n7013) );
  NAND2_X1 U8631 ( .A1(n7014), .A2(n7013), .ZN(n7036) );
  NAND2_X1 U8632 ( .A1(n7032), .A2(n7036), .ZN(n7015) );
  XNOR2_X1 U8633 ( .A(n7016), .B(n7015), .ZN(n7027) );
  NAND2_X1 U8634 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n7950) );
  OAI21_X1 U8635 ( .B1(n7922), .B2(n8396), .A(n7950), .ZN(n7025) );
  NAND2_X1 U8636 ( .A1(n5450), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7023) );
  INV_X1 U8637 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7017) );
  OR2_X1 U8638 ( .A1(n7392), .A2(n7017), .ZN(n7022) );
  INV_X1 U8639 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7042) );
  NAND2_X1 U8640 ( .A1(n7018), .A2(n7042), .ZN(n7019) );
  NAND2_X1 U8641 ( .A1(n7378), .A2(n7019), .ZN(n8376) );
  OR2_X1 U8642 ( .A1(n4279), .A2(n8376), .ZN(n7021) );
  INV_X1 U8643 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8377) );
  OR2_X1 U8644 ( .A1(n4277), .A2(n8377), .ZN(n7020) );
  NAND4_X1 U8645 ( .A1(n7023), .A2(n7022), .A3(n7021), .A4(n7020), .ZN(n8026)
         );
  INV_X1 U8646 ( .A(n8026), .ZN(n8385) );
  OAI22_X1 U8647 ( .A1(n7893), .A2(n8385), .B1(n8387), .B2(n7892), .ZN(n7024)
         );
  AOI211_X1 U8648 ( .C1(n8477), .C2(n7903), .A(n7025), .B(n7024), .ZN(n7026)
         );
  OAI21_X1 U8649 ( .B1(n7027), .B2(n7913), .A(n7026), .ZN(P2_U3228) );
  NOR2_X1 U8650 ( .A1(n7034), .A2(n7033), .ZN(n7028) );
  NAND2_X1 U8651 ( .A1(n7031), .A2(n7030), .ZN(n7039) );
  NAND2_X1 U8652 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  NAND2_X1 U8653 ( .A1(n7039), .A2(n7038), .ZN(n7745) );
  NAND2_X1 U8654 ( .A1(n5560), .A2(n8026), .ZN(n7742) );
  NAND2_X1 U8655 ( .A1(n7076), .A2(n6133), .ZN(n7041) );
  AOI22_X1 U8656 ( .A1(n7985), .A2(n5720), .B1(n7473), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n7040) );
  XNOR2_X1 U8657 ( .A(n8474), .B(n5554), .ZN(n7741) );
  XOR2_X1 U8658 ( .A(n7742), .B(n7741), .Z(n7744) );
  XNOR2_X1 U8659 ( .A(n7745), .B(n7744), .ZN(n7050) );
  OAI22_X1 U8660 ( .A1(n7922), .A2(n8376), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7042), .ZN(n7048) );
  NAND2_X1 U8661 ( .A1(n6027), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7046) );
  INV_X1 U8662 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7983) );
  OR2_X1 U8663 ( .A1(n7522), .A2(n7983), .ZN(n7045) );
  INV_X1 U8664 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7377) );
  XNOR2_X1 U8665 ( .A(n7378), .B(n7377), .ZN(n8356) );
  OR2_X1 U8666 ( .A1(n4279), .A2(n8356), .ZN(n7044) );
  INV_X1 U8667 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8357) );
  OR2_X1 U8668 ( .A1(n4277), .A2(n8357), .ZN(n7043) );
  NAND4_X1 U8669 ( .A1(n7046), .A2(n7045), .A3(n7044), .A4(n7043), .ZN(n8027)
         );
  INV_X1 U8670 ( .A(n8027), .ZN(n8373) );
  OAI22_X1 U8671 ( .A1(n7893), .A2(n8373), .B1(n8372), .B2(n7892), .ZN(n7047)
         );
  AOI211_X1 U8672 ( .C1(n8474), .C2(n7903), .A(n7048), .B(n7047), .ZN(n7049)
         );
  OAI21_X1 U8673 ( .B1(n7050), .B2(n7913), .A(n7049), .ZN(P2_U3230) );
  NAND2_X1 U8674 ( .A1(n7385), .A2(n6383), .ZN(n7053) );
  OR2_X1 U8675 ( .A1(n8687), .A2(n7051), .ZN(n7052) );
  NAND2_X1 U8676 ( .A1(n7065), .A2(n8626), .ZN(n7054) );
  NAND2_X1 U8677 ( .A1(n7055), .A2(n7054), .ZN(n9245) );
  OR2_X1 U8678 ( .A1(n9245), .A2(n7167), .ZN(n7061) );
  INV_X1 U8679 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U8680 ( .A1(n8678), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7057) );
  NAND2_X1 U8681 ( .A1(n4284), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7056) );
  OAI211_X1 U8682 ( .C1(n7058), .C2(n8683), .A(n7057), .B(n7056), .ZN(n7059)
         );
  INV_X1 U8683 ( .A(n7059), .ZN(n7060) );
  INV_X1 U8684 ( .A(n9256), .ZN(n8958) );
  NAND2_X1 U8685 ( .A1(n7369), .A2(n6383), .ZN(n7063) );
  AOI22_X1 U8686 ( .A1(n7086), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9638), .B2(
        n7085), .ZN(n7062) );
  OR2_X1 U8687 ( .A1(n7091), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7064) );
  AND2_X1 U8688 ( .A1(n7065), .A2(n7064), .ZN(n9260) );
  NAND2_X1 U8689 ( .A1(n9260), .A2(n5254), .ZN(n7068) );
  AOI22_X1 U8690 ( .A1(n5255), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n8678), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n7067) );
  NAND2_X1 U8691 ( .A1(n4284), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7066) );
  INV_X1 U8692 ( .A(n9277), .ZN(n8959) );
  AND2_X1 U8693 ( .A1(n7070), .A2(n7069), .ZN(n7071) );
  OR2_X1 U8694 ( .A1(n7071), .A2(n7089), .ZN(n9296) );
  NAND2_X1 U8695 ( .A1(n8678), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7073) );
  NAND2_X1 U8696 ( .A1(n5255), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7072) );
  AND2_X1 U8697 ( .A1(n7073), .A2(n7072), .ZN(n7075) );
  NAND2_X1 U8698 ( .A1(n4284), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7074) );
  OAI211_X1 U8699 ( .C1(n9296), .C2(n7167), .A(n7075), .B(n7074), .ZN(n9304)
         );
  NAND2_X1 U8700 ( .A1(n7076), .A2(n6383), .ZN(n7078) );
  AOI22_X1 U8701 ( .A1(n7086), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7085), .B2(
        n9077), .ZN(n7077) );
  INV_X1 U8702 ( .A(n9304), .ZN(n9276) );
  NAND2_X1 U8703 ( .A1(n7080), .A2(n6383), .ZN(n7082) );
  AOI22_X1 U8704 ( .A1(n7086), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7085), .B2(
        n9064), .ZN(n7081) );
  NAND2_X1 U8705 ( .A1(n9313), .A2(n9290), .ZN(n8810) );
  NAND2_X1 U8706 ( .A1(n8811), .A2(n8810), .ZN(n8906) );
  OAI21_X1 U8707 ( .B1(n7243), .B2(n9276), .A(n9285), .ZN(n7084) );
  NAND2_X1 U8708 ( .A1(n7366), .A2(n6383), .ZN(n7088) );
  AOI22_X1 U8709 ( .A1(n7086), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7085), .B2(
        n9091), .ZN(n7087) );
  NOR2_X1 U8710 ( .A1(n7089), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7090) );
  OR2_X1 U8711 ( .A1(n7091), .A2(n7090), .ZN(n9268) );
  AOI22_X1 U8712 ( .A1(n5255), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8678), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n7093) );
  INV_X1 U8713 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9269) );
  OR2_X1 U8714 ( .A1(n4280), .A2(n9269), .ZN(n7092) );
  OAI211_X1 U8715 ( .C1(n9268), .C2(n7167), .A(n7093), .B(n7092), .ZN(n8960)
         );
  INV_X1 U8716 ( .A(n8960), .ZN(n9292) );
  OR2_X1 U8717 ( .A1(n9384), .A2(n9292), .ZN(n8816) );
  NAND2_X1 U8718 ( .A1(n9384), .A2(n9292), .ZN(n8751) );
  AOI21_X1 U8719 ( .B1(n9256), .B2(n9249), .A(n9238), .ZN(n7096) );
  AOI21_X2 U8720 ( .B1(n9373), .B2(n8958), .A(n7096), .ZN(n9226) );
  NAND2_X1 U8721 ( .A1(n7398), .A2(n6383), .ZN(n7099) );
  OR2_X1 U8722 ( .A1(n8687), .A2(n7097), .ZN(n7098) );
  NAND2_X1 U8723 ( .A1(n9368), .A2(n9242), .ZN(n8691) );
  INV_X1 U8724 ( .A(n9368), .ZN(n9235) );
  NAND2_X1 U8725 ( .A1(n7408), .A2(n6383), .ZN(n7102) );
  OR2_X1 U8726 ( .A1(n8687), .A2(n7100), .ZN(n7101) );
  AND2_X1 U8727 ( .A1(n7103), .A2(n8635), .ZN(n7104) );
  OR2_X1 U8728 ( .A1(n7104), .A2(n7113), .ZN(n8638) );
  INV_X1 U8729 ( .A(n8638), .ZN(n9219) );
  INV_X1 U8730 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U8731 ( .A1(n5255), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7106) );
  NAND2_X1 U8732 ( .A1(n8678), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7105) );
  OAI211_X1 U8733 ( .C1(n7107), .C2(n4280), .A(n7106), .B(n7105), .ZN(n7108)
         );
  AOI21_X1 U8734 ( .B1(n9219), .B2(n5254), .A(n7108), .ZN(n9230) );
  NOR2_X1 U8735 ( .A1(n9222), .A2(n9230), .ZN(n7109) );
  INV_X1 U8736 ( .A(n9230), .ZN(n9207) );
  NAND2_X1 U8737 ( .A1(n7417), .A2(n6383), .ZN(n7112) );
  OR2_X1 U8738 ( .A1(n8687), .A2(n7110), .ZN(n7111) );
  OR2_X1 U8739 ( .A1(n7113), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7115) );
  AND2_X1 U8740 ( .A1(n7115), .A2(n7114), .ZN(n9198) );
  NAND2_X1 U8741 ( .A1(n9198), .A2(n5254), .ZN(n7121) );
  INV_X1 U8742 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7118) );
  NAND2_X1 U8743 ( .A1(n8678), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7117) );
  NAND2_X1 U8744 ( .A1(n4284), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7116) );
  OAI211_X1 U8745 ( .C1(n7118), .C2(n8683), .A(n7117), .B(n7116), .ZN(n7119)
         );
  INV_X1 U8746 ( .A(n7119), .ZN(n7120) );
  NAND2_X1 U8747 ( .A1(n7121), .A2(n7120), .ZN(n9183) );
  INV_X1 U8748 ( .A(n9357), .ZN(n9200) );
  INV_X1 U8749 ( .A(n9183), .ZN(n9216) );
  NAND2_X1 U8750 ( .A1(n7424), .A2(n6383), .ZN(n7124) );
  OR2_X1 U8751 ( .A1(n5513), .A2(n7122), .ZN(n7123) );
  NAND2_X1 U8752 ( .A1(n5255), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n7130) );
  INV_X1 U8753 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n7125) );
  OR2_X1 U8754 ( .A1(n5528), .A2(n7125), .ZN(n7129) );
  OAI21_X1 U8755 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n7126), .A(n7135), .ZN(
        n9190) );
  OR2_X1 U8756 ( .A1(n7167), .A2(n9190), .ZN(n7128) );
  INV_X1 U8757 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9191) );
  OR2_X1 U8758 ( .A1(n4280), .A2(n9191), .ZN(n7127) );
  NAND2_X1 U8759 ( .A1(n7436), .A2(n6383), .ZN(n7133) );
  OR2_X1 U8760 ( .A1(n8687), .A2(n7131), .ZN(n7132) );
  NAND2_X1 U8761 ( .A1(n8678), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7140) );
  INV_X1 U8762 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7134) );
  OR2_X1 U8763 ( .A1(n8683), .A2(n7134), .ZN(n7139) );
  INV_X1 U8764 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U8765 ( .A1(n8585), .A2(n7135), .ZN(n7136) );
  NAND2_X1 U8766 ( .A1(n7145), .A2(n7136), .ZN(n9169) );
  OR2_X1 U8767 ( .A1(n7167), .A2(n9169), .ZN(n7138) );
  INV_X1 U8768 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9170) );
  OR2_X1 U8769 ( .A1(n4280), .A2(n9170), .ZN(n7137) );
  NAND2_X1 U8770 ( .A1(n9176), .A2(n8957), .ZN(n8848) );
  AOI22_X1 U8771 ( .A1(n9168), .A2(n9167), .B1(n8957), .B2(n9173), .ZN(n9146)
         );
  NAND2_X1 U8772 ( .A1(n7450), .A2(n6383), .ZN(n7142) );
  OR2_X1 U8773 ( .A1(n8687), .A2(n7335), .ZN(n7141) );
  NAND2_X1 U8774 ( .A1(n5255), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7150) );
  INV_X1 U8775 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n7143) );
  OR2_X1 U8776 ( .A1(n5528), .A2(n7143), .ZN(n7149) );
  INV_X1 U8777 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7144) );
  NAND2_X1 U8778 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  NAND2_X1 U8779 ( .A1(n7156), .A2(n7146), .ZN(n9149) );
  OR2_X1 U8780 ( .A1(n7167), .A2(n9149), .ZN(n7148) );
  INV_X1 U8781 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9150) );
  OR2_X1 U8782 ( .A1(n4280), .A2(n9150), .ZN(n7147) );
  NAND2_X1 U8783 ( .A1(n9153), .A2(n9161), .ZN(n7151) );
  NAND2_X1 U8784 ( .A1(n7462), .A2(n6383), .ZN(n7153) );
  OR2_X1 U8785 ( .A1(n8687), .A2(n8267), .ZN(n7152) );
  NAND2_X1 U8786 ( .A1(n8678), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7162) );
  INV_X1 U8787 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7154) );
  OR2_X1 U8788 ( .A1(n8683), .A2(n7154), .ZN(n7161) );
  INV_X1 U8789 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7155) );
  NAND2_X1 U8790 ( .A1(n7156), .A2(n7155), .ZN(n7157) );
  NAND2_X1 U8791 ( .A1(n7165), .A2(n7157), .ZN(n9133) );
  OR2_X1 U8792 ( .A1(n7167), .A2(n9133), .ZN(n7160) );
  INV_X1 U8793 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n7158) );
  OR2_X1 U8794 ( .A1(n4280), .A2(n7158), .ZN(n7159) );
  NAND2_X1 U8795 ( .A1(n9337), .A2(n7327), .ZN(n8859) );
  OR2_X1 U8796 ( .A1(n8687), .A2(n7344), .ZN(n7174) );
  NAND2_X1 U8797 ( .A1(n8678), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7171) );
  INV_X1 U8798 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7163) );
  OR2_X1 U8799 ( .A1(n8683), .A2(n7163), .ZN(n7170) );
  INV_X1 U8800 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U8801 ( .A1(n7165), .A2(n7164), .ZN(n7166) );
  NAND2_X1 U8802 ( .A1(n7193), .A2(n7166), .ZN(n9123) );
  OR2_X1 U8803 ( .A1(n7167), .A2(n9123), .ZN(n7169) );
  INV_X1 U8804 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9124) );
  OR2_X1 U8805 ( .A1(n4280), .A2(n9124), .ZN(n7168) );
  INV_X1 U8806 ( .A(n9136), .ZN(n7172) );
  AND2_X1 U8807 ( .A1(n7174), .A2(n7172), .ZN(n7173) );
  NAND2_X1 U8808 ( .A1(n9114), .A2(n9117), .ZN(n9113) );
  NAND2_X1 U8809 ( .A1(n9332), .A2(n7172), .ZN(n7175) );
  NAND2_X1 U8810 ( .A1(n9113), .A2(n7175), .ZN(n7190) );
  INV_X1 U8811 ( .A(SI_28_), .ZN(n7176) );
  NAND2_X1 U8812 ( .A1(n7177), .A2(n7176), .ZN(n7183) );
  INV_X1 U8813 ( .A(n7183), .ZN(n7179) );
  OR2_X1 U8814 ( .A1(n7179), .A2(n7178), .ZN(n7506) );
  AND2_X1 U8815 ( .A1(n7180), .A2(n7506), .ZN(n7181) );
  INV_X1 U8816 ( .A(n7506), .ZN(n7185) );
  AND2_X1 U8817 ( .A1(n7184), .A2(n7183), .ZN(n7501) );
  OR2_X1 U8818 ( .A1(n7185), .A2(n7501), .ZN(n7498) );
  MUX2_X1 U8819 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7532), .Z(n7504) );
  INV_X1 U8820 ( .A(SI_29_), .ZN(n7505) );
  XNOR2_X1 U8821 ( .A(n7504), .B(n7505), .ZN(n7186) );
  NAND2_X1 U8822 ( .A1(n7489), .A2(n6383), .ZN(n7189) );
  INV_X1 U8823 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7362) );
  OR2_X1 U8824 ( .A1(n8687), .A2(n7362), .ZN(n7188) );
  NAND2_X1 U8825 ( .A1(n9325), .A2(n9115), .ZN(n8930) );
  INV_X1 U8826 ( .A(n9384), .ZN(n9278) );
  INV_X1 U8827 ( .A(n9121), .ZN(n7191) );
  INV_X1 U8828 ( .A(n9325), .ZN(n7192) );
  AOI211_X1 U8829 ( .C1(n9325), .C2(n7191), .A(n9295), .B(n9107), .ZN(n9324)
         );
  NOR2_X1 U8830 ( .A1(n7192), .A2(n9263), .ZN(n7196) );
  OAI22_X1 U8831 ( .A1(n9641), .A2(n7194), .B1(n7193), .B2(n9306), .ZN(n7195)
         );
  AOI211_X1 U8832 ( .C1(n9324), .C2(n9628), .A(n7196), .B(n7195), .ZN(n7214)
         );
  INV_X1 U8833 ( .A(n8810), .ZN(n7198) );
  NAND2_X1 U8834 ( .A1(n9390), .A2(n9276), .ZN(n8809) );
  OR2_X1 U8835 ( .A1(n9390), .A2(n9276), .ZN(n9271) );
  AND2_X1 U8836 ( .A1(n8816), .A2(n9271), .ZN(n8753) );
  INV_X1 U8837 ( .A(n8751), .ZN(n7199) );
  AOI21_X2 U8838 ( .B1(n9272), .B2(n8753), .A(n7199), .ZN(n9254) );
  OR2_X1 U8839 ( .A1(n9378), .A2(n9277), .ZN(n8815) );
  NAND2_X1 U8840 ( .A1(n9378), .A2(n9277), .ZN(n8818) );
  NAND2_X1 U8841 ( .A1(n8815), .A2(n8818), .ZN(n9253) );
  NAND2_X1 U8842 ( .A1(n9373), .A2(n9256), .ZN(n8817) );
  INV_X1 U8843 ( .A(n8691), .ZN(n7200) );
  NAND2_X1 U8844 ( .A1(n9222), .A2(n9207), .ZN(n8836) );
  NAND2_X1 U8845 ( .A1(n9363), .A2(n9230), .ZN(n8692) );
  INV_X1 U8846 ( .A(n8836), .ZN(n7201) );
  NAND2_X1 U8847 ( .A1(n9357), .A2(n9216), .ZN(n8834) );
  NAND2_X1 U8848 ( .A1(n8844), .A2(n8834), .ZN(n9203) );
  INV_X1 U8849 ( .A(n8844), .ZN(n7202) );
  XNOR2_X1 U8850 ( .A(n9352), .B(n9166), .ZN(n9181) );
  NAND2_X1 U8851 ( .A1(n9182), .A2(n9181), .ZN(n9180) );
  NAND2_X1 U8852 ( .A1(n9352), .A2(n9201), .ZN(n8845) );
  NAND2_X1 U8853 ( .A1(n9342), .A2(n9161), .ZN(n8856) );
  NAND2_X1 U8854 ( .A1(n9154), .A2(n8856), .ZN(n9138) );
  NOR2_X1 U8855 ( .A1(n9332), .A2(n9136), .ZN(n7203) );
  NOR2_X1 U8856 ( .A1(n9116), .A2(n7203), .ZN(n7205) );
  XNOR2_X1 U8857 ( .A(n7205), .B(n7204), .ZN(n7206) );
  INV_X1 U8858 ( .A(n8991), .ZN(n9557) );
  AND2_X1 U8859 ( .A1(n9557), .A2(P1_B_REG_SCAN_IN), .ZN(n7207) );
  NOR2_X1 U8860 ( .A1(n9293), .A2(n7207), .ZN(n9103) );
  INV_X1 U8861 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7210) );
  NAND2_X1 U8862 ( .A1(n4284), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U8863 ( .A1(n8678), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7208) );
  OAI211_X1 U8864 ( .C1(n8683), .C2(n7210), .A(n7209), .B(n7208), .ZN(n8956)
         );
  AOI22_X1 U8865 ( .A1(n9103), .A2(n8956), .B1(n7172), .B2(n9614), .ZN(n7211)
         );
  NAND2_X1 U8866 ( .A1(n9329), .A2(n9644), .ZN(n7213) );
  OAI211_X1 U8867 ( .C1(n9330), .C2(n9301), .A(n7214), .B(n7213), .ZN(P1_U3355) );
  NAND2_X1 U8868 ( .A1(n8696), .A2(n7289), .ZN(n7219) );
  NAND2_X1 U8869 ( .A1(n8962), .A2(n4285), .ZN(n7218) );
  NAND2_X1 U8870 ( .A1(n7219), .A2(n7218), .ZN(n7220) );
  XNOR2_X1 U8871 ( .A(n7220), .B(n7320), .ZN(n7224) );
  NAND2_X1 U8872 ( .A1(n8672), .A2(n7289), .ZN(n7222) );
  NAND2_X1 U8873 ( .A1(n9303), .A2(n4285), .ZN(n7221) );
  NAND2_X1 U8874 ( .A1(n7222), .A2(n7221), .ZN(n7223) );
  XNOR2_X1 U8875 ( .A(n7223), .B(n5653), .ZN(n7232) );
  NAND2_X1 U8876 ( .A1(n8696), .A2(n4285), .ZN(n7227) );
  NAND2_X1 U8877 ( .A1(n8962), .A2(n7286), .ZN(n7226) );
  NAND2_X1 U8878 ( .A1(n7227), .A2(n7226), .ZN(n8537) );
  NAND2_X1 U8879 ( .A1(n7228), .A2(n8541), .ZN(n8661) );
  NAND2_X1 U8880 ( .A1(n8672), .A2(n4285), .ZN(n7230) );
  NAND2_X1 U8881 ( .A1(n9303), .A2(n7286), .ZN(n7229) );
  NAND2_X1 U8882 ( .A1(n7230), .A2(n7229), .ZN(n8660) );
  NAND2_X1 U8883 ( .A1(n8541), .A2(n7231), .ZN(n7234) );
  INV_X1 U8884 ( .A(n7232), .ZN(n7233) );
  NAND2_X1 U8885 ( .A1(n9313), .A2(n7289), .ZN(n7236) );
  NAND2_X1 U8886 ( .A1(n8961), .A2(n4285), .ZN(n7235) );
  NAND2_X1 U8887 ( .A1(n7236), .A2(n7235), .ZN(n7237) );
  XNOR2_X1 U8888 ( .A(n7237), .B(n5653), .ZN(n7240) );
  NOR2_X1 U8889 ( .A1(n9290), .A2(n7322), .ZN(n7238) );
  AOI21_X1 U8890 ( .B1(n9313), .B2(n4285), .A(n7238), .ZN(n7239) );
  XNOR2_X1 U8891 ( .A(n7240), .B(n7239), .ZN(n8594) );
  NAND2_X1 U8892 ( .A1(n7240), .A2(n7239), .ZN(n7241) );
  OAI22_X1 U8893 ( .A1(n7243), .A2(n7319), .B1(n9276), .B2(n7283), .ZN(n7242)
         );
  XNOR2_X1 U8894 ( .A(n7242), .B(n5653), .ZN(n7248) );
  OR2_X1 U8895 ( .A1(n7243), .A2(n7283), .ZN(n7245) );
  NAND2_X1 U8896 ( .A1(n9304), .A2(n7286), .ZN(n7244) );
  NAND2_X1 U8897 ( .A1(n7245), .A2(n7244), .ZN(n7246) );
  XNOR2_X1 U8898 ( .A(n7248), .B(n7246), .ZN(n8601) );
  NAND2_X1 U8899 ( .A1(n8600), .A2(n8601), .ZN(n7250) );
  INV_X1 U8900 ( .A(n7246), .ZN(n7247) );
  NAND2_X1 U8901 ( .A1(n7248), .A2(n7247), .ZN(n7249) );
  NAND2_X1 U8902 ( .A1(n9384), .A2(n7289), .ZN(n7252) );
  NAND2_X1 U8903 ( .A1(n8960), .A2(n4285), .ZN(n7251) );
  NAND2_X1 U8904 ( .A1(n7252), .A2(n7251), .ZN(n7253) );
  XNOR2_X1 U8905 ( .A(n7253), .B(n5653), .ZN(n7257) );
  NAND2_X1 U8906 ( .A1(n9384), .A2(n4285), .ZN(n7255) );
  NAND2_X1 U8907 ( .A1(n8960), .A2(n7286), .ZN(n7254) );
  NAND2_X1 U8908 ( .A1(n7255), .A2(n7254), .ZN(n8642) );
  INV_X1 U8909 ( .A(n7256), .ZN(n7259) );
  INV_X1 U8910 ( .A(n7257), .ZN(n7258) );
  OAI22_X1 U8911 ( .A1(n9264), .A2(n7319), .B1(n9277), .B2(n7283), .ZN(n7260)
         );
  XNOR2_X1 U8912 ( .A(n7260), .B(n7320), .ZN(n8565) );
  OAI22_X1 U8913 ( .A1(n9264), .A2(n7283), .B1(n9277), .B2(n7322), .ZN(n8566)
         );
  NAND2_X1 U8914 ( .A1(n8564), .A2(n8565), .ZN(n7261) );
  OAI22_X1 U8915 ( .A1(n9249), .A2(n7319), .B1(n9256), .B2(n7283), .ZN(n7262)
         );
  XNOR2_X1 U8916 ( .A(n7262), .B(n7320), .ZN(n7265) );
  OR2_X1 U8917 ( .A1(n9249), .A2(n7283), .ZN(n7264) );
  NAND2_X1 U8918 ( .A1(n8958), .A2(n7286), .ZN(n7263) );
  NAND2_X1 U8919 ( .A1(n7264), .A2(n7263), .ZN(n7266) );
  AND2_X1 U8920 ( .A1(n7265), .A2(n7266), .ZN(n8621) );
  INV_X1 U8921 ( .A(n7265), .ZN(n7268) );
  INV_X1 U8922 ( .A(n7266), .ZN(n7267) );
  NAND2_X1 U8923 ( .A1(n7268), .A2(n7267), .ZN(n8619) );
  NAND2_X1 U8924 ( .A1(n8624), .A2(n8619), .ZN(n8573) );
  NAND2_X1 U8925 ( .A1(n9368), .A2(n7289), .ZN(n7270) );
  OR2_X1 U8926 ( .A1(n9242), .A2(n7283), .ZN(n7269) );
  NAND2_X1 U8927 ( .A1(n7270), .A2(n7269), .ZN(n7271) );
  XNOR2_X1 U8928 ( .A(n7271), .B(n7320), .ZN(n7273) );
  NOR2_X1 U8929 ( .A1(n9242), .A2(n7322), .ZN(n7272) );
  AOI21_X1 U8930 ( .B1(n9368), .B2(n4285), .A(n7272), .ZN(n7274) );
  XNOR2_X1 U8931 ( .A(n7273), .B(n7274), .ZN(n8574) );
  NAND2_X1 U8932 ( .A1(n8573), .A2(n8574), .ZN(n7277) );
  INV_X1 U8933 ( .A(n7273), .ZN(n7275) );
  NAND2_X1 U8934 ( .A1(n7275), .A2(n7274), .ZN(n7276) );
  NOR2_X1 U8935 ( .A1(n9230), .A2(n7322), .ZN(n7278) );
  AOI21_X1 U8936 ( .B1(n9363), .B2(n4285), .A(n7278), .ZN(n7280) );
  OAI22_X1 U8937 ( .A1(n9222), .A2(n7319), .B1(n9230), .B2(n7283), .ZN(n7279)
         );
  XNOR2_X1 U8938 ( .A(n7279), .B(n7320), .ZN(n8634) );
  OAI22_X1 U8939 ( .A1(n9192), .A2(n7319), .B1(n9201), .B2(n7283), .ZN(n7282)
         );
  XNOR2_X1 U8940 ( .A(n7282), .B(n7320), .ZN(n8610) );
  OR2_X1 U8941 ( .A1(n9192), .A2(n7283), .ZN(n7285) );
  OR2_X1 U8942 ( .A1(n9201), .A2(n7322), .ZN(n7284) );
  NAND2_X1 U8943 ( .A1(n7285), .A2(n7284), .ZN(n8609) );
  NAND2_X1 U8944 ( .A1(n9357), .A2(n4285), .ZN(n7288) );
  NAND2_X1 U8945 ( .A1(n9183), .A2(n7286), .ZN(n7287) );
  NAND2_X1 U8946 ( .A1(n7288), .A2(n7287), .ZN(n7295) );
  NAND2_X1 U8947 ( .A1(n9357), .A2(n7289), .ZN(n7292) );
  NAND2_X1 U8948 ( .A1(n9183), .A2(n4285), .ZN(n7291) );
  NAND2_X1 U8949 ( .A1(n7292), .A2(n7291), .ZN(n7293) );
  XNOR2_X1 U8950 ( .A(n7293), .B(n7320), .ZN(n8552) );
  AOI22_X1 U8951 ( .A1(n8610), .A2(n8609), .B1(n7295), .B2(n8552), .ZN(n7294)
         );
  NAND2_X1 U8952 ( .A1(n8550), .A2(n7294), .ZN(n7303) );
  INV_X1 U8953 ( .A(n8552), .ZN(n8554) );
  INV_X1 U8954 ( .A(n7298), .ZN(n7296) );
  INV_X1 U8955 ( .A(n8609), .ZN(n7299) );
  INV_X1 U8956 ( .A(n8610), .ZN(n7297) );
  OAI21_X1 U8957 ( .B1(n7299), .B2(n7298), .A(n7297), .ZN(n7300) );
  NAND2_X1 U8958 ( .A1(n7303), .A2(n7302), .ZN(n8582) );
  OAI22_X1 U8959 ( .A1(n9173), .A2(n7319), .B1(n8957), .B2(n7283), .ZN(n7304)
         );
  XNOR2_X1 U8960 ( .A(n7304), .B(n7320), .ZN(n7306) );
  NOR2_X1 U8961 ( .A1(n8957), .A2(n7322), .ZN(n7305) );
  AOI21_X1 U8962 ( .B1(n9176), .B2(n4285), .A(n7305), .ZN(n7307) );
  XNOR2_X1 U8963 ( .A(n7306), .B(n7307), .ZN(n8583) );
  INV_X1 U8964 ( .A(n7306), .ZN(n7308) );
  OAI22_X1 U8965 ( .A1(n9153), .A2(n7283), .B1(n9161), .B2(n7322), .ZN(n7311)
         );
  OAI22_X1 U8966 ( .A1(n9153), .A2(n7319), .B1(n9161), .B2(n7283), .ZN(n7309)
         );
  XNOR2_X1 U8967 ( .A(n7309), .B(n7320), .ZN(n7310) );
  XOR2_X1 U8968 ( .A(n7311), .B(n7310), .Z(n7337) );
  NAND2_X1 U8969 ( .A1(n7336), .A2(n7312), .ZN(n8528) );
  OAI22_X1 U8970 ( .A1(n4491), .A2(n7319), .B1(n7327), .B2(n7283), .ZN(n7313)
         );
  XOR2_X1 U8971 ( .A(n7320), .B(n7313), .Z(n8530) );
  NOR2_X1 U8972 ( .A1(n7327), .A2(n7322), .ZN(n7314) );
  AOI21_X1 U8973 ( .B1(n9337), .B2(n4285), .A(n7314), .ZN(n7315) );
  NAND2_X1 U8974 ( .A1(n8530), .A2(n7315), .ZN(n7317) );
  INV_X1 U8975 ( .A(n7315), .ZN(n8529) );
  OAI22_X1 U8976 ( .A1(n9122), .A2(n7319), .B1(n9136), .B2(n7283), .ZN(n7321)
         );
  XNOR2_X1 U8977 ( .A(n7321), .B(n7320), .ZN(n7324) );
  OAI22_X1 U8978 ( .A1(n9122), .A2(n7283), .B1(n9136), .B2(n7322), .ZN(n7323)
         );
  XNOR2_X1 U8979 ( .A(n7324), .B(n7323), .ZN(n7325) );
  XNOR2_X1 U8980 ( .A(n7326), .B(n7325), .ZN(n7332) );
  NOR2_X1 U8981 ( .A1(n4275), .A2(n9123), .ZN(n7330) );
  AOI22_X1 U8982 ( .A1(n8666), .A2(n4490), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7328) );
  OAI21_X1 U8983 ( .B1(n9115), .B2(n8664), .A(n7328), .ZN(n7329) );
  AOI211_X1 U8984 ( .C1(n9332), .C2(n8671), .A(n7330), .B(n7329), .ZN(n7331)
         );
  OAI21_X1 U8985 ( .B1(n7332), .B2(n8645), .A(n7331), .ZN(P1_U3218) );
  OAI222_X1 U8986 ( .A1(n7361), .A2(n7335), .B1(n7364), .B2(n7334), .C1(
        P1_U3084), .C2(n7333), .ZN(P1_U3327) );
  OAI211_X1 U8987 ( .C1(n7338), .C2(n7337), .A(n7336), .B(n8657), .ZN(n7343)
         );
  INV_X1 U8988 ( .A(n9149), .ZN(n7341) );
  AOI22_X1 U8989 ( .A1(n8653), .A2(n4490), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n7339) );
  OAI21_X1 U8990 ( .B1(n8957), .B2(n8650), .A(n7339), .ZN(n7340) );
  AOI21_X1 U8991 ( .B1(n7341), .B2(n8576), .A(n7340), .ZN(n7342) );
  OAI211_X1 U8992 ( .C1(n9153), .C2(n8656), .A(n7343), .B(n7342), .ZN(P1_U3238) );
  OAI222_X1 U8993 ( .A1(n7364), .A2(n7345), .B1(n4283), .B2(P1_U3084), .C1(
        n7344), .C2(n7361), .ZN(P1_U3325) );
  OAI21_X1 U8994 ( .B1(n7347), .B2(n7714), .A(n7346), .ZN(n8501) );
  AOI22_X1 U8995 ( .A1(n9772), .A2(n7932), .B1(n7930), .B2(n9769), .ZN(n7352)
         );
  AND2_X1 U8996 ( .A1(n7348), .A2(n7714), .ZN(n7349) );
  OAI21_X1 U8997 ( .B1(n7350), .B2(n7349), .A(n9776), .ZN(n7351) );
  OAI211_X1 U8998 ( .C1(n8501), .C2(n9781), .A(n7352), .B(n7351), .ZN(n8503)
         );
  NAND2_X1 U8999 ( .A1(n8503), .A2(n9788), .ZN(n7360) );
  OAI22_X1 U9000 ( .A1(n9788), .A2(n6510), .B1(n7353), .B2(n9792), .ZN(n7358)
         );
  AND2_X1 U9001 ( .A1(n7354), .A2(n8495), .ZN(n7356) );
  OR2_X1 U9002 ( .A1(n7356), .A2(n7355), .ZN(n8497) );
  NOR2_X1 U9003 ( .A1(n8497), .A2(n8014), .ZN(n7357) );
  AOI211_X1 U9004 ( .C1(n8380), .C2(n8495), .A(n7358), .B(n7357), .ZN(n7359)
         );
  OAI211_X1 U9005 ( .C1(n8501), .C2(n9798), .A(n7360), .B(n7359), .ZN(P2_U3283) );
  INV_X1 U9006 ( .A(n7489), .ZN(n7819) );
  OAI222_X1 U9007 ( .A1(n7364), .A2(n7819), .B1(n7363), .B2(P1_U3084), .C1(
        n7362), .C2(n7361), .ZN(P1_U3324) );
  NAND2_X1 U9008 ( .A1(n7365), .A2(n7630), .ZN(n8383) );
  NAND2_X1 U9009 ( .A1(n8477), .A2(n8372), .ZN(n7633) );
  NOR2_X1 U9010 ( .A1(n8477), .A2(n8372), .ZN(n7621) );
  AOI21_X1 U9011 ( .B1(n8383), .B2(n7633), .A(n7621), .ZN(n8369) );
  NAND2_X1 U9012 ( .A1(n8474), .A2(n8385), .ZN(n7638) );
  NAND2_X1 U9013 ( .A1(n7366), .A2(n6133), .ZN(n7368) );
  AOI22_X1 U9014 ( .A1(n7995), .A2(n5720), .B1(n7473), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n7367) );
  OR2_X1 U9015 ( .A1(n8467), .A2(n8373), .ZN(n7642) );
  NAND2_X1 U9016 ( .A1(n8467), .A2(n8373), .ZN(n7645) );
  NAND2_X1 U9017 ( .A1(n7642), .A2(n7645), .ZN(n8351) );
  NAND2_X1 U9018 ( .A1(n7369), .A2(n6133), .ZN(n7372) );
  AOI22_X1 U9019 ( .A1(n7370), .A2(n5720), .B1(n7473), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n7371) );
  NAND2_X1 U9020 ( .A1(n7517), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7383) );
  INV_X1 U9021 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7373) );
  OR2_X1 U9022 ( .A1(n7522), .A2(n7373), .ZN(n7382) );
  AND2_X1 U9023 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n7374) );
  INV_X1 U9024 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7376) );
  OAI21_X1 U9025 ( .B1(n7378), .B2(n7377), .A(n7376), .ZN(n7379) );
  NAND2_X1 U9026 ( .A1(n7388), .A2(n7379), .ZN(n8341) );
  OR2_X1 U9027 ( .A1(n4279), .A2(n8341), .ZN(n7381) );
  INV_X1 U9028 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8342) );
  OR2_X1 U9029 ( .A1(n4278), .A2(n8342), .ZN(n7380) );
  NAND4_X1 U9030 ( .A1(n7383), .A2(n7382), .A3(n7381), .A4(n7380), .ZN(n8327)
         );
  INV_X1 U9031 ( .A(n8327), .ZN(n8353) );
  NAND2_X1 U9032 ( .A1(n8344), .A2(n8353), .ZN(n7384) );
  INV_X1 U9033 ( .A(n7384), .ZN(n8322) );
  NAND2_X1 U9034 ( .A1(n7385), .A2(n6133), .ZN(n7387) );
  NAND2_X1 U9035 ( .A1(n7473), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7386) );
  INV_X1 U9036 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U9037 ( .A1(n7388), .A2(n7864), .ZN(n7389) );
  NAND2_X1 U9038 ( .A1(n7402), .A2(n7389), .ZN(n8318) );
  OR2_X1 U9039 ( .A1(n8318), .A2(n4279), .ZN(n7397) );
  INV_X1 U9040 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7390) );
  OR2_X1 U9041 ( .A1(n7522), .A2(n7390), .ZN(n7396) );
  INV_X1 U9042 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n7391) );
  OR2_X1 U9043 ( .A1(n7392), .A2(n7391), .ZN(n7395) );
  INV_X1 U9044 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n7393) );
  OR2_X1 U9045 ( .A1(n4277), .A2(n7393), .ZN(n7394) );
  NAND4_X1 U9046 ( .A1(n7397), .A2(n7396), .A3(n7395), .A4(n7394), .ZN(n8174)
         );
  INV_X1 U9047 ( .A(n8174), .ZN(n8335) );
  NAND2_X1 U9048 ( .A1(n8457), .A2(n8335), .ZN(n7647) );
  NAND2_X1 U9049 ( .A1(n7398), .A2(n6133), .ZN(n7400) );
  NAND2_X1 U9050 ( .A1(n7473), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7399) );
  INV_X1 U9051 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U9052 ( .A1(n7402), .A2(n7837), .ZN(n7403) );
  NAND2_X1 U9053 ( .A1(n7411), .A2(n7403), .ZN(n8167) );
  OR2_X1 U9054 ( .A1(n8167), .A2(n4279), .ZN(n7407) );
  NAND2_X1 U9055 ( .A1(n7517), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7406) );
  INV_X1 U9056 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8237) );
  OR2_X1 U9057 ( .A1(n7522), .A2(n8237), .ZN(n7405) );
  NAND2_X1 U9058 ( .A1(n7490), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7404) );
  NAND4_X1 U9059 ( .A1(n7407), .A2(n7406), .A3(n7405), .A4(n7404), .ZN(n8326)
         );
  INV_X1 U9060 ( .A(n8326), .ZN(n8030) );
  OR2_X1 U9061 ( .A1(n8452), .A2(n8030), .ZN(n7654) );
  NAND2_X1 U9062 ( .A1(n8452), .A2(n8030), .ZN(n8157) );
  NAND2_X1 U9063 ( .A1(n7408), .A2(n6133), .ZN(n7410) );
  NAND2_X1 U9064 ( .A1(n7473), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7409) );
  INV_X1 U9065 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n7415) );
  INV_X1 U9066 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U9067 ( .A1(n7411), .A2(n8299), .ZN(n7412) );
  NAND2_X1 U9068 ( .A1(n7420), .A2(n7412), .ZN(n8150) );
  OR2_X1 U9069 ( .A1(n8150), .A2(n4279), .ZN(n7414) );
  AOI22_X1 U9070 ( .A1(n7490), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n7517), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n7413) );
  OAI211_X1 U9071 ( .C1(n7522), .C2(n7415), .A(n7414), .B(n7413), .ZN(n8175)
         );
  INV_X1 U9072 ( .A(n8175), .ZN(n8032) );
  NAND2_X1 U9073 ( .A1(n8447), .A2(n8032), .ZN(n7657) );
  NAND2_X1 U9074 ( .A1(n8128), .A2(n7657), .ZN(n8033) );
  NAND2_X1 U9075 ( .A1(n7417), .A2(n6133), .ZN(n7419) );
  NAND2_X1 U9076 ( .A1(n7473), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7418) );
  INV_X1 U9077 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U9078 ( .A1(n7420), .A2(n7824), .ZN(n7421) );
  NAND2_X1 U9079 ( .A1(n7428), .A2(n7421), .ZN(n8136) );
  AOI22_X1 U9080 ( .A1(n5450), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n6027), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9081 ( .A1(n7490), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7422) );
  OAI211_X1 U9082 ( .C1(n8136), .C2(n4279), .A(n7423), .B(n7422), .ZN(n8154)
         );
  INV_X1 U9083 ( .A(n8154), .ZN(n8034) );
  OR2_X1 U9084 ( .A1(n8440), .A2(n8034), .ZN(n7659) );
  NAND2_X1 U9085 ( .A1(n8440), .A2(n8034), .ZN(n8118) );
  NAND2_X1 U9086 ( .A1(n7424), .A2(n6133), .ZN(n7426) );
  NAND2_X1 U9087 ( .A1(n7473), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7425) );
  INV_X1 U9088 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U9089 ( .A1(n7428), .A2(n7854), .ZN(n7429) );
  NAND2_X1 U9090 ( .A1(n7441), .A2(n7429), .ZN(n8115) );
  OR2_X1 U9091 ( .A1(n8115), .A2(n4279), .ZN(n7434) );
  INV_X1 U9092 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U9093 ( .A1(n7517), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7431) );
  NAND2_X1 U9094 ( .A1(n7490), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7430) );
  OAI211_X1 U9095 ( .C1(n7522), .C2(n8223), .A(n7431), .B(n7430), .ZN(n7432)
         );
  INV_X1 U9096 ( .A(n7432), .ZN(n7433) );
  NAND2_X1 U9097 ( .A1(n7434), .A2(n7433), .ZN(n8132) );
  NAND2_X1 U9098 ( .A1(n8435), .A2(n8035), .ZN(n7660) );
  NAND2_X1 U9099 ( .A1(n7436), .A2(n6133), .ZN(n7438) );
  NAND2_X1 U9100 ( .A1(n7473), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7437) );
  INV_X1 U9101 ( .A(n7441), .ZN(n7439) );
  NAND2_X1 U9102 ( .A1(n7439), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7453) );
  INV_X1 U9103 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U9104 ( .A1(n7441), .A2(n7440), .ZN(n7442) );
  NAND2_X1 U9105 ( .A1(n7453), .A2(n7442), .ZN(n8098) );
  OR2_X1 U9106 ( .A1(n8098), .A2(n4279), .ZN(n7448) );
  INV_X1 U9107 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n7445) );
  NAND2_X1 U9108 ( .A1(n7490), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7444) );
  NAND2_X1 U9109 ( .A1(n7517), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7443) );
  OAI211_X1 U9110 ( .C1(n7522), .C2(n7445), .A(n7444), .B(n7443), .ZN(n7446)
         );
  INV_X1 U9111 ( .A(n7446), .ZN(n7447) );
  NAND2_X1 U9112 ( .A1(n7448), .A2(n7447), .ZN(n8122) );
  INV_X1 U9113 ( .A(n8122), .ZN(n7855) );
  NAND2_X1 U9114 ( .A1(n8432), .A2(n7855), .ZN(n7669) );
  NAND2_X1 U9115 ( .A1(n7450), .A2(n6133), .ZN(n7452) );
  NAND2_X1 U9116 ( .A1(n7473), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7451) );
  INV_X1 U9117 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U9118 ( .A1(n7453), .A2(n7920), .ZN(n7454) );
  NAND2_X1 U9119 ( .A1(n8092), .A2(n5731), .ZN(n7460) );
  INV_X1 U9120 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7457) );
  NAND2_X1 U9121 ( .A1(n7490), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7456) );
  NAND2_X1 U9122 ( .A1(n7517), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7455) );
  OAI211_X1 U9123 ( .C1(n7522), .C2(n7457), .A(n7456), .B(n7455), .ZN(n7458)
         );
  INV_X1 U9124 ( .A(n7458), .ZN(n7459) );
  NAND2_X1 U9125 ( .A1(n7460), .A2(n7459), .ZN(n7928) );
  NAND2_X1 U9126 ( .A1(n8426), .A2(n8036), .ZN(n7695) );
  INV_X1 U9127 ( .A(n7695), .ZN(n7461) );
  NAND2_X1 U9128 ( .A1(n7462), .A2(n6133), .ZN(n7464) );
  NAND2_X1 U9129 ( .A1(n7473), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7463) );
  XNOR2_X1 U9130 ( .A(n7480), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U9131 ( .A1(n8080), .A2(n5731), .ZN(n7470) );
  INV_X1 U9132 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7467) );
  NAND2_X1 U9133 ( .A1(n7490), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7466) );
  NAND2_X1 U9134 ( .A1(n7517), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7465) );
  OAI211_X1 U9135 ( .C1(n7522), .C2(n7467), .A(n7466), .B(n7465), .ZN(n7468)
         );
  INV_X1 U9136 ( .A(n7468), .ZN(n7469) );
  NAND2_X1 U9137 ( .A1(n8074), .A2(n8057), .ZN(n7471) );
  NAND2_X1 U9138 ( .A1(n8075), .A2(n7471), .ZN(n8056) );
  NAND2_X1 U9139 ( .A1(n7472), .A2(n6133), .ZN(n7475) );
  NAND2_X1 U9140 ( .A1(n7473), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7474) );
  INV_X1 U9141 ( .A(n7480), .ZN(n7477) );
  AND2_X1 U9142 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n7476) );
  NAND2_X1 U9143 ( .A1(n7477), .A2(n7476), .ZN(n8046) );
  INV_X1 U9144 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7479) );
  INV_X1 U9145 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7478) );
  OAI21_X1 U9146 ( .B1(n7480), .B2(n7479), .A(n7478), .ZN(n7481) );
  NAND2_X1 U9147 ( .A1(n8046), .A2(n7481), .ZN(n7804) );
  OR2_X1 U9148 ( .A1(n7804), .A2(n4279), .ZN(n7487) );
  INV_X1 U9149 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U9150 ( .A1(n7490), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U9151 ( .A1(n7517), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7482) );
  OAI211_X1 U9152 ( .C1(n7522), .C2(n7484), .A(n7483), .B(n7482), .ZN(n7485)
         );
  INV_X1 U9153 ( .A(n7485), .ZN(n7486) );
  NAND2_X1 U9154 ( .A1(n7487), .A2(n7486), .ZN(n8042) );
  INV_X1 U9155 ( .A(n8042), .ZN(n8037) );
  NAND2_X1 U9156 ( .A1(n8415), .A2(n8037), .ZN(n7693) );
  INV_X1 U9157 ( .A(n7694), .ZN(n7676) );
  INV_X1 U9158 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7818) );
  NOR2_X1 U9159 ( .A1(n4287), .A2(n7818), .ZN(n7488) );
  OR2_X1 U9160 ( .A1(n8046), .A2(n4279), .ZN(n7496) );
  INV_X1 U9161 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7493) );
  NAND2_X1 U9162 ( .A1(n7517), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U9163 ( .A1(n7490), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7491) );
  OAI211_X1 U9164 ( .C1(n7522), .C2(n7493), .A(n7492), .B(n7491), .ZN(n7494)
         );
  INV_X1 U9165 ( .A(n7494), .ZN(n7495) );
  NAND2_X1 U9166 ( .A1(n7496), .A2(n7495), .ZN(n8058) );
  INV_X1 U9167 ( .A(n7678), .ZN(n7497) );
  AND2_X1 U9168 ( .A1(n7498), .A2(SI_29_), .ZN(n7499) );
  NAND2_X1 U9169 ( .A1(n7500), .A2(n7499), .ZN(n7511) );
  AND2_X1 U9170 ( .A1(n7501), .A2(n7504), .ZN(n7502) );
  NAND2_X1 U9171 ( .A1(n7503), .A2(n7502), .ZN(n7510) );
  INV_X1 U9172 ( .A(n7504), .ZN(n7508) );
  AND2_X1 U9173 ( .A1(n7506), .A2(n7505), .ZN(n7507) );
  OR2_X1 U9174 ( .A1(n7508), .A2(n7507), .ZN(n7509) );
  NAND3_X1 U9175 ( .A1(n7511), .A2(n7510), .A3(n7509), .ZN(n7529) );
  MUX2_X1 U9176 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7532), .Z(n7528) );
  NAND2_X1 U9177 ( .A1(n8685), .A2(n6133), .ZN(n7513) );
  INV_X1 U9178 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7798) );
  OR2_X1 U9179 ( .A1(n4288), .A2(n7798), .ZN(n7512) );
  NAND2_X1 U9180 ( .A1(n7540), .A2(n7550), .ZN(n7523) );
  NOR2_X1 U9181 ( .A1(n8410), .A2(n8058), .ZN(n7677) );
  INV_X1 U9182 ( .A(n7677), .ZN(n7514) );
  OAI21_X1 U9183 ( .B1(n9498), .B2(n7523), .A(n7514), .ZN(n7515) );
  INV_X1 U9184 ( .A(n7515), .ZN(n7516) );
  INV_X1 U9185 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n7521) );
  NAND2_X1 U9186 ( .A1(n7517), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7520) );
  INV_X1 U9187 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n7518) );
  OR2_X1 U9188 ( .A1(n4277), .A2(n7518), .ZN(n7519) );
  OAI211_X1 U9189 ( .C1(n7522), .C2(n7521), .A(n7520), .B(n7519), .ZN(n8040)
         );
  INV_X1 U9190 ( .A(n8040), .ZN(n7539) );
  INV_X1 U9191 ( .A(n7683), .ZN(n7524) );
  INV_X1 U9192 ( .A(n7526), .ZN(n7527) );
  NAND2_X1 U9193 ( .A1(n7527), .A2(SI_30_), .ZN(n7531) );
  NAND2_X1 U9194 ( .A1(n7529), .A2(n7528), .ZN(n7530) );
  NAND2_X1 U9195 ( .A1(n7531), .A2(n7530), .ZN(n7535) );
  MUX2_X1 U9196 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7532), .Z(n7533) );
  XNOR2_X1 U9197 ( .A(n7533), .B(SI_31_), .ZN(n7534) );
  NAND2_X1 U9198 ( .A1(n8676), .A2(n6133), .ZN(n7538) );
  INV_X1 U9199 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7536) );
  OR2_X1 U9200 ( .A1(n4287), .A2(n7536), .ZN(n7537) );
  OR2_X1 U9201 ( .A1(n8405), .A2(n7540), .ZN(n7687) );
  NAND2_X1 U9202 ( .A1(n8016), .A2(n7539), .ZN(n7685) );
  AOI21_X1 U9203 ( .B1(n7541), .B2(n7680), .A(n7682), .ZN(n7542) );
  XNOR2_X1 U9204 ( .A(n7542), .B(n8375), .ZN(n7545) );
  NAND2_X1 U9205 ( .A1(n5560), .A2(n7543), .ZN(n7544) );
  NAND2_X1 U9206 ( .A1(n7545), .A2(n7544), .ZN(n7732) );
  OAI21_X1 U9207 ( .B1(n7729), .B2(n7738), .A(n5544), .ZN(n7546) );
  OR2_X1 U9208 ( .A1(n7738), .A2(n7727), .ZN(n7548) );
  AND2_X1 U9209 ( .A1(n7555), .A2(n7550), .ZN(n7552) );
  OAI211_X1 U9210 ( .C1(n7552), .C2(n7551), .A(n7698), .B(n7554), .ZN(n7553)
         );
  NAND2_X1 U9211 ( .A1(n7553), .A2(n7557), .ZN(n7560) );
  NAND2_X1 U9212 ( .A1(n7555), .A2(n7554), .ZN(n7701) );
  NAND3_X1 U9213 ( .A1(n7701), .A2(n7557), .A3(n7556), .ZN(n7558) );
  NAND2_X1 U9214 ( .A1(n7558), .A2(n7698), .ZN(n7559) );
  MUX2_X1 U9215 ( .A(n7560), .B(n7559), .S(n7671), .Z(n7565) );
  NAND2_X1 U9216 ( .A1(n7567), .A2(n7568), .ZN(n7562) );
  NAND2_X1 U9217 ( .A1(n7574), .A2(n7575), .ZN(n7561) );
  MUX2_X1 U9218 ( .A(n7562), .B(n7561), .S(n7690), .Z(n7577) );
  INV_X1 U9219 ( .A(n7577), .ZN(n7564) );
  NAND3_X1 U9220 ( .A1(n7565), .A2(n7564), .A3(n7563), .ZN(n7572) );
  AND2_X1 U9221 ( .A1(n7567), .A2(n7566), .ZN(n7569) );
  OAI211_X1 U9222 ( .C1(n7577), .C2(n7569), .A(n7568), .B(n7582), .ZN(n7570)
         );
  NAND2_X1 U9223 ( .A1(n7570), .A2(n7690), .ZN(n7571) );
  NAND2_X1 U9224 ( .A1(n7572), .A2(n7571), .ZN(n7580) );
  NAND2_X1 U9225 ( .A1(n7936), .A2(n9861), .ZN(n7579) );
  AND2_X1 U9226 ( .A1(n7574), .A2(n7573), .ZN(n7576) );
  OAI211_X1 U9227 ( .C1(n7577), .C2(n7576), .A(n7575), .B(n7579), .ZN(n7578)
         );
  AOI22_X1 U9228 ( .A1(n7580), .A2(n7579), .B1(n7671), .B2(n7578), .ZN(n7587)
         );
  OAI21_X1 U9229 ( .B1(n7690), .B2(n7582), .A(n7581), .ZN(n7586) );
  MUX2_X1 U9230 ( .A(n7584), .B(n7583), .S(n7690), .Z(n7585) );
  OAI211_X1 U9231 ( .C1(n7587), .C2(n7586), .A(n7709), .B(n7585), .ZN(n7591)
         );
  MUX2_X1 U9232 ( .A(n7589), .B(n7588), .S(n7690), .Z(n7590) );
  NAND3_X1 U9233 ( .A1(n7591), .A2(n7592), .A3(n7590), .ZN(n7594) );
  NAND2_X1 U9234 ( .A1(n7595), .A2(n7592), .ZN(n7593) );
  NAND2_X1 U9235 ( .A1(n7593), .A2(n7690), .ZN(n7598) );
  NAND4_X1 U9236 ( .A1(n7594), .A2(n7598), .A3(n7596), .A4(n7599), .ZN(n7605)
         );
  NAND2_X1 U9237 ( .A1(n7610), .A2(n7595), .ZN(n7602) );
  INV_X1 U9238 ( .A(n7596), .ZN(n7597) );
  NAND2_X1 U9239 ( .A1(n7598), .A2(n7597), .ZN(n7600) );
  NAND3_X1 U9240 ( .A1(n7600), .A2(n7606), .A3(n7599), .ZN(n7601) );
  INV_X1 U9241 ( .A(n7603), .ZN(n7604) );
  NAND2_X1 U9242 ( .A1(n7605), .A2(n7604), .ZN(n7611) );
  NAND2_X1 U9243 ( .A1(n7611), .A2(n7607), .ZN(n7608) );
  NAND3_X1 U9244 ( .A1(n7611), .A2(n7610), .A3(n7609), .ZN(n7613) );
  INV_X1 U9245 ( .A(n7714), .ZN(n7614) );
  MUX2_X1 U9246 ( .A(n7931), .B(n8495), .S(n7671), .Z(n7616) );
  NAND2_X1 U9247 ( .A1(n7616), .A2(n7615), .ZN(n7617) );
  MUX2_X1 U9248 ( .A(n7930), .B(n8488), .S(n7671), .Z(n7618) );
  NAND2_X1 U9249 ( .A1(n7619), .A2(n7618), .ZN(n7629) );
  NAND2_X1 U9250 ( .A1(n7629), .A2(n8488), .ZN(n7620) );
  NAND3_X1 U9251 ( .A1(n7620), .A2(n7634), .A3(n7631), .ZN(n7623) );
  INV_X1 U9252 ( .A(n7621), .ZN(n7622) );
  NAND3_X1 U9253 ( .A1(n7623), .A2(n7622), .A3(n7630), .ZN(n7626) );
  MUX2_X1 U9254 ( .A(n7929), .B(n8477), .S(n7690), .Z(n7624) );
  NAND2_X1 U9255 ( .A1(n8477), .A2(n7929), .ZN(n8024) );
  AND2_X1 U9256 ( .A1(n7624), .A2(n8024), .ZN(n7625) );
  NOR2_X1 U9257 ( .A1(n8368), .A2(n7625), .ZN(n7636) );
  NAND2_X1 U9258 ( .A1(n7626), .A2(n7636), .ZN(n7628) );
  NAND3_X1 U9259 ( .A1(n7628), .A2(n7627), .A3(n7642), .ZN(n7641) );
  NAND2_X1 U9260 ( .A1(n7629), .A2(n7930), .ZN(n7632) );
  NAND3_X1 U9261 ( .A1(n7632), .A2(n7631), .A3(n7630), .ZN(n7635) );
  NAND3_X1 U9262 ( .A1(n7635), .A2(n7634), .A3(n7633), .ZN(n7637) );
  NAND2_X1 U9263 ( .A1(n7637), .A2(n7636), .ZN(n7639) );
  NAND3_X1 U9264 ( .A1(n7639), .A2(n7645), .A3(n7638), .ZN(n7640) );
  AOI21_X1 U9265 ( .B1(n7646), .B2(n7642), .A(n8322), .ZN(n7644) );
  NAND2_X1 U9266 ( .A1(n7653), .A2(n7649), .ZN(n7643) );
  OAI211_X1 U9267 ( .C1(n7644), .C2(n7643), .A(n7647), .B(n8157), .ZN(n7652)
         );
  NAND2_X1 U9268 ( .A1(n7646), .A2(n7645), .ZN(n7650) );
  INV_X1 U9269 ( .A(n7647), .ZN(n7648) );
  AOI211_X1 U9270 ( .C1(n7650), .C2(n7649), .A(n7648), .B(n8322), .ZN(n7651)
         );
  AOI21_X1 U9271 ( .B1(n7654), .B2(n7653), .A(n7671), .ZN(n7656) );
  MUX2_X1 U9272 ( .A(n7654), .B(n8157), .S(n7690), .Z(n7655) );
  MUX2_X1 U9273 ( .A(n7657), .B(n8128), .S(n7690), .Z(n7658) );
  AND2_X1 U9274 ( .A1(n7660), .A2(n8118), .ZN(n7661) );
  INV_X1 U9275 ( .A(n7696), .ZN(n7664) );
  AOI211_X1 U9276 ( .C1(n7666), .C2(n8102), .A(n7664), .B(n7663), .ZN(n7668)
         );
  NAND2_X1 U9277 ( .A1(n7695), .A2(n7669), .ZN(n7670) );
  OAI21_X1 U9278 ( .B1(n7671), .B2(n7696), .A(n8076), .ZN(n7673) );
  NAND3_X1 U9279 ( .A1(n8074), .A2(n7671), .A3(n8057), .ZN(n7672) );
  OAI21_X1 U9280 ( .B1(n8074), .B2(n8057), .A(n7693), .ZN(n7675) );
  MUX2_X1 U9281 ( .A(n7678), .B(n7677), .S(n7690), .Z(n7679) );
  INV_X1 U9282 ( .A(n7680), .ZN(n7725) );
  AOI21_X1 U9283 ( .B1(n7686), .B2(n7683), .A(n7725), .ZN(n7681) );
  NOR2_X1 U9284 ( .A1(n7681), .A2(n7682), .ZN(n7692) );
  INV_X1 U9285 ( .A(n7682), .ZN(n7684) );
  NAND2_X1 U9286 ( .A1(n7684), .A2(n7683), .ZN(n7724) );
  AOI21_X1 U9287 ( .B1(n7686), .B2(n7685), .A(n7724), .ZN(n7689) );
  INV_X1 U9288 ( .A(n7687), .ZN(n7688) );
  NOR2_X1 U9289 ( .A1(n7689), .A2(n7688), .ZN(n7691) );
  NAND2_X1 U9290 ( .A1(n7694), .A2(n7693), .ZN(n8055) );
  INV_X1 U9291 ( .A(n8055), .ZN(n8053) );
  OR2_X1 U9292 ( .A1(n8477), .A2(n7929), .ZN(n7697) );
  INV_X1 U9293 ( .A(n8388), .ZN(n7718) );
  INV_X1 U9294 ( .A(n7698), .ZN(n7699) );
  NOR4_X1 U9295 ( .A1(n7701), .A2(n7700), .A3(n7699), .A4(n5468), .ZN(n7704)
         );
  NAND3_X1 U9296 ( .A1(n7704), .A2(n7703), .A3(n7702), .ZN(n7707) );
  NOR4_X1 U9297 ( .A1(n7707), .A2(n4307), .A3(n7706), .A4(n7705), .ZN(n7710)
         );
  NAND4_X1 U9298 ( .A1(n7710), .A2(n7709), .A3(n9777), .A4(n7708), .ZN(n7713)
         );
  NOR4_X1 U9299 ( .A1(n7714), .A2(n7713), .A3(n7712), .A4(n7711), .ZN(n7716)
         );
  NAND4_X1 U9300 ( .A1(n7718), .A2(n7717), .A3(n7716), .A4(n7715), .ZN(n7719)
         );
  NOR4_X1 U9301 ( .A1(n8323), .A2(n8368), .A3(n8351), .A4(n7719), .ZN(n7720)
         );
  NAND4_X1 U9302 ( .A1(n8156), .A2(n8173), .A3(n8028), .A4(n7720), .ZN(n7721)
         );
  NOR4_X1 U9303 ( .A1(n8088), .A2(n4605), .A3(n8141), .A4(n7721), .ZN(n7722)
         );
  NAND4_X1 U9304 ( .A1(n8053), .A2(n8102), .A3(n7722), .A4(n8076), .ZN(n7723)
         );
  NOR4_X1 U9305 ( .A1(n7725), .A2(n7724), .A3(n4290), .A4(n7723), .ZN(n7726)
         );
  XNOR2_X1 U9306 ( .A(n7726), .B(n8375), .ZN(n7728) );
  OAI211_X1 U9307 ( .C1(n7730), .C2(n7729), .A(n7728), .B(n7727), .ZN(n7731)
         );
  INV_X1 U9308 ( .A(n8009), .ZN(n7734) );
  NAND4_X1 U9309 ( .A1(n7735), .A2(n9804), .A3(n7734), .A4(n9772), .ZN(n7736)
         );
  OAI211_X1 U9310 ( .C1(n7738), .C2(n7737), .A(n7736), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7739) );
  NAND2_X1 U9311 ( .A1(n7740), .A2(n7739), .ZN(P2_U3244) );
  INV_X1 U9312 ( .A(n7741), .ZN(n7743) );
  XNOR2_X1 U9313 ( .A(n8467), .B(n5554), .ZN(n7747) );
  NAND2_X1 U9314 ( .A1(n5560), .A2(n8027), .ZN(n7746) );
  XNOR2_X1 U9315 ( .A(n7747), .B(n7746), .ZN(n7890) );
  INV_X1 U9316 ( .A(n7746), .ZN(n7748) );
  AND2_X1 U9317 ( .A1(n5560), .A2(n8327), .ZN(n7750) );
  XNOR2_X1 U9318 ( .A(n8344), .B(n5554), .ZN(n7749) );
  NOR2_X1 U9319 ( .A1(n7749), .A2(n7750), .ZN(n7756) );
  AOI21_X1 U9320 ( .B1(n7750), .B2(n7749), .A(n7756), .ZN(n7829) );
  XNOR2_X1 U9321 ( .A(n8457), .B(n6486), .ZN(n7755) );
  INV_X1 U9322 ( .A(n7755), .ZN(n7752) );
  NAND2_X1 U9323 ( .A1(n5560), .A2(n8174), .ZN(n7754) );
  INV_X1 U9324 ( .A(n7754), .ZN(n7751) );
  NAND2_X1 U9325 ( .A1(n7752), .A2(n7751), .ZN(n7753) );
  AND2_X1 U9326 ( .A1(n7829), .A2(n7753), .ZN(n7760) );
  INV_X1 U9327 ( .A(n7753), .ZN(n7759) );
  XNOR2_X1 U9328 ( .A(n7755), .B(n7754), .ZN(n7862) );
  INV_X1 U9329 ( .A(n7862), .ZN(n7757) );
  INV_X1 U9330 ( .A(n7756), .ZN(n7860) );
  AND2_X1 U9331 ( .A1(n7757), .A2(n7860), .ZN(n7758) );
  XNOR2_X1 U9332 ( .A(n8452), .B(n5554), .ZN(n7761) );
  NAND2_X1 U9333 ( .A1(n5560), .A2(n8326), .ZN(n7762) );
  XNOR2_X1 U9334 ( .A(n7761), .B(n7762), .ZN(n7836) );
  INV_X1 U9335 ( .A(n7761), .ZN(n7763) );
  XNOR2_X1 U9336 ( .A(n8447), .B(n5554), .ZN(n7764) );
  XNOR2_X1 U9337 ( .A(n7766), .B(n7764), .ZN(n7871) );
  NAND2_X1 U9338 ( .A1(n5560), .A2(n8175), .ZN(n7870) );
  INV_X1 U9339 ( .A(n7764), .ZN(n7765) );
  NAND2_X1 U9340 ( .A1(n7766), .A2(n7765), .ZN(n7767) );
  XOR2_X1 U9341 ( .A(n5554), .B(n8440), .Z(n7768) );
  NAND2_X1 U9342 ( .A1(n8154), .A2(n5560), .ZN(n7822) );
  NAND2_X1 U9343 ( .A1(n7820), .A2(n7822), .ZN(n7770) );
  NAND2_X1 U9344 ( .A1(n7769), .A2(n7768), .ZN(n7821) );
  NAND2_X1 U9345 ( .A1(n7770), .A2(n7821), .ZN(n7771) );
  XNOR2_X1 U9346 ( .A(n8435), .B(n5554), .ZN(n7772) );
  XNOR2_X1 U9347 ( .A(n7771), .B(n7772), .ZN(n7852) );
  AND2_X1 U9348 ( .A1(n8132), .A2(n5560), .ZN(n7853) );
  NAND2_X1 U9349 ( .A1(n7852), .A2(n7853), .ZN(n7775) );
  INV_X1 U9350 ( .A(n7771), .ZN(n7773) );
  NAND2_X1 U9351 ( .A1(n7773), .A2(n7772), .ZN(n7774) );
  XNOR2_X1 U9352 ( .A(n8432), .B(n5554), .ZN(n7843) );
  NAND2_X1 U9353 ( .A1(n8122), .A2(n5560), .ZN(n7842) );
  INV_X1 U9354 ( .A(n7915), .ZN(n7779) );
  XNOR2_X1 U9355 ( .A(n8426), .B(n5554), .ZN(n7777) );
  AND2_X1 U9356 ( .A1(n7928), .A2(n5560), .ZN(n7776) );
  NAND2_X1 U9357 ( .A1(n7777), .A2(n7776), .ZN(n7784) );
  OAI21_X1 U9358 ( .B1(n7777), .B2(n7776), .A(n7784), .ZN(n7914) );
  INV_X1 U9359 ( .A(n7914), .ZN(n7778) );
  NAND2_X1 U9360 ( .A1(n7779), .A2(n7778), .ZN(n7916) );
  NAND2_X1 U9361 ( .A1(n7916), .A2(n7784), .ZN(n7790) );
  XNOR2_X1 U9362 ( .A(n8420), .B(n5554), .ZN(n7781) );
  INV_X1 U9363 ( .A(n7781), .ZN(n7783) );
  AND2_X1 U9364 ( .A1(n8057), .A2(n5560), .ZN(n7780) );
  INV_X1 U9365 ( .A(n7780), .ZN(n7782) );
  AOI21_X1 U9366 ( .B1(n7783), .B2(n7782), .A(n7808), .ZN(n7789) );
  INV_X1 U9367 ( .A(n7789), .ZN(n7785) );
  OR2_X1 U9368 ( .A1(n7914), .A2(n7785), .ZN(n7787) );
  INV_X1 U9369 ( .A(n7788), .ZN(n7816) );
  OAI211_X1 U9370 ( .C1(n7790), .C2(n7789), .A(n7816), .B(n7901), .ZN(n7795)
         );
  AOI22_X1 U9371 ( .A1(n8042), .A2(n9769), .B1(n9772), .B2(n7928), .ZN(n8078)
         );
  AOI22_X1 U9372 ( .A1(n8080), .A2(n7885), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n7791) );
  OAI21_X1 U9373 ( .B1(n8078), .B2(n7792), .A(n7791), .ZN(n7793) );
  AOI21_X1 U9374 ( .B1(n8420), .B2(n7903), .A(n7793), .ZN(n7794) );
  NAND2_X1 U9375 ( .A1(n7795), .A2(n7794), .ZN(P2_U3216) );
  INV_X1 U9376 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8686) );
  INV_X1 U9377 ( .A(n8685), .ZN(n7799) );
  OAI222_X1 U9378 ( .A1(n7361), .A2(n8686), .B1(n9417), .B2(n7799), .C1(
        P1_U3084), .C2(n7796), .ZN(P1_U3323) );
  OAI222_X1 U9379 ( .A1(n7797), .A2(P2_U3152), .B1(n7800), .B2(n7799), .C1(
        n7798), .C2(n7817), .ZN(P2_U3328) );
  NAND2_X1 U9380 ( .A1(n8042), .A2(n5560), .ZN(n7801) );
  XNOR2_X1 U9381 ( .A(n7801), .B(n6486), .ZN(n7802) );
  XNOR2_X1 U9382 ( .A(n8415), .B(n7802), .ZN(n7807) );
  NAND2_X1 U9383 ( .A1(n7807), .A2(n7901), .ZN(n7815) );
  NOR3_X1 U9384 ( .A1(n7807), .A2(n7808), .A3(n7913), .ZN(n7803) );
  NAND2_X1 U9385 ( .A1(n7816), .A2(n7803), .ZN(n7814) );
  INV_X1 U9386 ( .A(n7804), .ZN(n8064) );
  AOI22_X1 U9387 ( .A1(n8064), .A2(n7885), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n7806) );
  NAND2_X1 U9388 ( .A1(n7905), .A2(n8058), .ZN(n7805) );
  OAI211_X1 U9389 ( .C1(n4787), .C2(n7892), .A(n7806), .B(n7805), .ZN(n7812)
         );
  INV_X1 U9390 ( .A(n7807), .ZN(n7810) );
  INV_X1 U9391 ( .A(n7808), .ZN(n7809) );
  NOR3_X1 U9392 ( .A1(n7810), .A2(n7809), .A3(n7913), .ZN(n7811) );
  AOI211_X1 U9393 ( .C1(n8415), .C2(n7903), .A(n7812), .B(n7811), .ZN(n7813)
         );
  OAI211_X1 U9394 ( .C1(n7816), .C2(n7815), .A(n7814), .B(n7813), .ZN(P2_U3222) );
  OAI222_X1 U9395 ( .A1(P2_U3152), .A2(n5451), .B1(n7800), .B2(n7819), .C1(
        n7818), .C2(n7817), .ZN(P2_U3329) );
  NAND2_X1 U9396 ( .A1(n7820), .A2(n7821), .ZN(n7823) );
  XNOR2_X1 U9397 ( .A(n7823), .B(n7822), .ZN(n7828) );
  OAI22_X1 U9398 ( .A1(n7922), .A2(n8136), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7824), .ZN(n7826) );
  OAI22_X1 U9399 ( .A1(n7893), .A2(n8035), .B1(n8032), .B2(n7892), .ZN(n7825)
         );
  AOI211_X1 U9400 ( .C1(n8440), .C2(n7903), .A(n7826), .B(n7825), .ZN(n7827)
         );
  OAI21_X1 U9401 ( .B1(n7828), .B2(n7913), .A(n7827), .ZN(P2_U3218) );
  INV_X1 U9402 ( .A(n8344), .ZN(n8465) );
  NAND2_X1 U9403 ( .A1(n7830), .A2(n7829), .ZN(n7861) );
  OAI21_X1 U9404 ( .B1(n7830), .B2(n7829), .A(n7861), .ZN(n7831) );
  NAND2_X1 U9405 ( .A1(n7831), .A2(n7901), .ZN(n7835) );
  INV_X1 U9406 ( .A(n8341), .ZN(n7833) );
  AND2_X1 U9407 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8006) );
  OAI22_X1 U9408 ( .A1(n7893), .A2(n8335), .B1(n8373), .B2(n7892), .ZN(n7832)
         );
  AOI211_X1 U9409 ( .C1(n7885), .C2(n7833), .A(n8006), .B(n7832), .ZN(n7834)
         );
  OAI211_X1 U9410 ( .C1(n8465), .C2(n7927), .A(n7835), .B(n7834), .ZN(P2_U3221) );
  XNOR2_X1 U9411 ( .A(n4357), .B(n7836), .ZN(n7841) );
  OAI22_X1 U9412 ( .A1(n7922), .A2(n8167), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7837), .ZN(n7839) );
  OAI22_X1 U9413 ( .A1(n7893), .A2(n8032), .B1(n8335), .B2(n7892), .ZN(n7838)
         );
  AOI211_X1 U9414 ( .C1(n8452), .C2(n7903), .A(n7839), .B(n7838), .ZN(n7840)
         );
  OAI21_X1 U9415 ( .B1(n7841), .B2(n7913), .A(n7840), .ZN(P2_U3225) );
  XNOR2_X1 U9416 ( .A(n7843), .B(n7842), .ZN(n7844) );
  XNOR2_X1 U9417 ( .A(n7845), .B(n7844), .ZN(n7851) );
  NAND2_X1 U9418 ( .A1(n7928), .A2(n9769), .ZN(n7847) );
  NAND2_X1 U9419 ( .A1(n8132), .A2(n9772), .ZN(n7846) );
  NAND2_X1 U9420 ( .A1(n7847), .A2(n7846), .ZN(n8104) );
  AOI22_X1 U9421 ( .A1(n8104), .A2(n7924), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n7848) );
  OAI21_X1 U9422 ( .B1(n8098), .B2(n7922), .A(n7848), .ZN(n7849) );
  AOI21_X1 U9423 ( .B1(n8432), .B2(n7903), .A(n7849), .ZN(n7850) );
  OAI21_X1 U9424 ( .B1(n7851), .B2(n7913), .A(n7850), .ZN(P2_U3227) );
  XNOR2_X1 U9425 ( .A(n7852), .B(n7853), .ZN(n7859) );
  OAI22_X1 U9426 ( .A1(n7922), .A2(n8115), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7854), .ZN(n7857) );
  OAI22_X1 U9427 ( .A1(n7893), .A2(n7855), .B1(n8034), .B2(n7892), .ZN(n7856)
         );
  AOI211_X1 U9428 ( .C1(n8435), .C2(n7903), .A(n7857), .B(n7856), .ZN(n7858)
         );
  OAI21_X1 U9429 ( .B1(n7859), .B2(n7913), .A(n7858), .ZN(P2_U3231) );
  NAND2_X1 U9430 ( .A1(n7861), .A2(n7860), .ZN(n7863) );
  XNOR2_X1 U9431 ( .A(n7863), .B(n7862), .ZN(n7868) );
  OAI22_X1 U9432 ( .A1(n7922), .A2(n8318), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7864), .ZN(n7866) );
  OAI22_X1 U9433 ( .A1(n7893), .A2(n8030), .B1(n8353), .B2(n7892), .ZN(n7865)
         );
  AOI211_X1 U9434 ( .C1(n8457), .C2(n7903), .A(n7866), .B(n7865), .ZN(n7867)
         );
  OAI21_X1 U9435 ( .B1(n7868), .B2(n7913), .A(n7867), .ZN(P2_U3235) );
  OAI21_X1 U9436 ( .B1(n7871), .B2(n7870), .A(n7869), .ZN(n7872) );
  NAND2_X1 U9437 ( .A1(n7872), .A2(n7901), .ZN(n7876) );
  OAI22_X1 U9438 ( .A1(n7922), .A2(n8150), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8299), .ZN(n7874) );
  OAI22_X1 U9439 ( .A1(n7893), .A2(n8034), .B1(n8030), .B2(n7892), .ZN(n7873)
         );
  AOI211_X1 U9440 ( .C1(n8447), .C2(n7903), .A(n7874), .B(n7873), .ZN(n7875)
         );
  NAND2_X1 U9441 ( .A1(n7876), .A2(n7875), .ZN(P2_U3237) );
  XOR2_X1 U9442 ( .A(n7878), .B(n7877), .Z(n7879) );
  NAND2_X1 U9443 ( .A1(n7879), .A2(n7901), .ZN(n7889) );
  AOI21_X1 U9444 ( .B1(n7924), .B2(n7881), .A(n7880), .ZN(n7888) );
  NAND2_X1 U9445 ( .A1(n7903), .A2(n7882), .ZN(n7887) );
  INV_X1 U9446 ( .A(n7883), .ZN(n7884) );
  NAND2_X1 U9447 ( .A1(n7885), .A2(n7884), .ZN(n7886) );
  NAND4_X1 U9448 ( .A1(n7889), .A2(n7888), .A3(n7887), .A4(n7886), .ZN(
        P2_U3238) );
  XNOR2_X1 U9449 ( .A(n7891), .B(n7890), .ZN(n7897) );
  NAND2_X1 U9450 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7988) );
  OAI21_X1 U9451 ( .B1(n7922), .B2(n8356), .A(n7988), .ZN(n7895) );
  OAI22_X1 U9452 ( .A1(n7893), .A2(n8353), .B1(n8385), .B2(n7892), .ZN(n7894)
         );
  AOI211_X1 U9453 ( .C1(n8467), .C2(n7903), .A(n7895), .B(n7894), .ZN(n7896)
         );
  OAI21_X1 U9454 ( .B1(n7897), .B2(n7913), .A(n7896), .ZN(P2_U3240) );
  OAI21_X1 U9455 ( .B1(n7900), .B2(n7899), .A(n7898), .ZN(n7902) );
  NAND2_X1 U9456 ( .A1(n7902), .A2(n7901), .ZN(n7912) );
  AOI22_X1 U9457 ( .A1(n7905), .A2(n7935), .B1(n7904), .B2(n7903), .ZN(n7911)
         );
  OAI21_X1 U9458 ( .B1(n7922), .B2(n7907), .A(n7906), .ZN(n7908) );
  AOI21_X1 U9459 ( .B1(n7909), .B2(n7937), .A(n7908), .ZN(n7910) );
  NAND3_X1 U9460 ( .A1(n7912), .A2(n7911), .A3(n7910), .ZN(P2_U3241) );
  INV_X1 U9461 ( .A(n8426), .ZN(n8086) );
  AOI21_X1 U9462 ( .B1(n7915), .B2(n7914), .A(n7913), .ZN(n7917) );
  NAND2_X1 U9463 ( .A1(n7917), .A2(n7916), .ZN(n7926) );
  NAND2_X1 U9464 ( .A1(n8057), .A2(n9769), .ZN(n7919) );
  NAND2_X1 U9465 ( .A1(n8122), .A2(n9772), .ZN(n7918) );
  NAND2_X1 U9466 ( .A1(n7919), .A2(n7918), .ZN(n8089) );
  INV_X1 U9467 ( .A(n8092), .ZN(n7921) );
  OAI22_X1 U9468 ( .A1(n7922), .A2(n7921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7920), .ZN(n7923) );
  AOI21_X1 U9469 ( .B1(n8089), .B2(n7924), .A(n7923), .ZN(n7925) );
  OAI211_X1 U9470 ( .C1(n8086), .C2(n7927), .A(n7926), .B(n7925), .ZN(P2_U3242) );
  MUX2_X1 U9471 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8040), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9472 ( .A(n8058), .B(P2_DATAO_REG_29__SCAN_IN), .S(n7941), .Z(
        P2_U3581) );
  MUX2_X1 U9473 ( .A(n8042), .B(P2_DATAO_REG_28__SCAN_IN), .S(n7941), .Z(
        P2_U3580) );
  MUX2_X1 U9474 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8057), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9475 ( .A(n7928), .B(P2_DATAO_REG_26__SCAN_IN), .S(n7941), .Z(
        P2_U3578) );
  MUX2_X1 U9476 ( .A(n8122), .B(P2_DATAO_REG_25__SCAN_IN), .S(n7941), .Z(
        P2_U3577) );
  MUX2_X1 U9477 ( .A(n8132), .B(P2_DATAO_REG_24__SCAN_IN), .S(n7941), .Z(
        P2_U3576) );
  MUX2_X1 U9478 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8154), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9479 ( .A(n8175), .B(P2_DATAO_REG_22__SCAN_IN), .S(n7941), .Z(
        P2_U3574) );
  MUX2_X1 U9480 ( .A(n8326), .B(P2_DATAO_REG_21__SCAN_IN), .S(n7941), .Z(
        P2_U3573) );
  MUX2_X1 U9481 ( .A(n8174), .B(P2_DATAO_REG_20__SCAN_IN), .S(n7941), .Z(
        P2_U3572) );
  MUX2_X1 U9482 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8327), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9483 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8027), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9484 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8026), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9485 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n7929), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9486 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8020), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9487 ( .A(n7930), .B(P2_DATAO_REG_14__SCAN_IN), .S(n7941), .Z(
        P2_U3566) );
  MUX2_X1 U9488 ( .A(n7931), .B(P2_DATAO_REG_13__SCAN_IN), .S(n7941), .Z(
        P2_U3565) );
  MUX2_X1 U9489 ( .A(n7932), .B(P2_DATAO_REG_12__SCAN_IN), .S(n7941), .Z(
        P2_U3564) );
  MUX2_X1 U9490 ( .A(n9770), .B(P2_DATAO_REG_11__SCAN_IN), .S(n7941), .Z(
        P2_U3563) );
  MUX2_X1 U9491 ( .A(n7933), .B(P2_DATAO_REG_10__SCAN_IN), .S(n7941), .Z(
        P2_U3562) );
  MUX2_X1 U9492 ( .A(n9771), .B(P2_DATAO_REG_9__SCAN_IN), .S(n7941), .Z(
        P2_U3561) );
  MUX2_X1 U9493 ( .A(n7934), .B(P2_DATAO_REG_8__SCAN_IN), .S(n7941), .Z(
        P2_U3560) );
  MUX2_X1 U9494 ( .A(n7935), .B(P2_DATAO_REG_7__SCAN_IN), .S(n7941), .Z(
        P2_U3559) );
  MUX2_X1 U9495 ( .A(n7936), .B(P2_DATAO_REG_6__SCAN_IN), .S(n7941), .Z(
        P2_U3558) );
  MUX2_X1 U9496 ( .A(n7937), .B(P2_DATAO_REG_5__SCAN_IN), .S(n7941), .Z(
        P2_U3557) );
  MUX2_X1 U9497 ( .A(n7938), .B(P2_DATAO_REG_4__SCAN_IN), .S(n7941), .Z(
        P2_U3556) );
  MUX2_X1 U9498 ( .A(n7939), .B(P2_DATAO_REG_3__SCAN_IN), .S(n7941), .Z(
        P2_U3555) );
  MUX2_X1 U9499 ( .A(n7940), .B(P2_DATAO_REG_2__SCAN_IN), .S(n7941), .Z(
        P2_U3554) );
  MUX2_X1 U9500 ( .A(n5545), .B(P2_DATAO_REG_1__SCAN_IN), .S(n7941), .Z(
        P2_U3553) );
  MUX2_X1 U9501 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n7942), .S(P2_U3966), .Z(
        P2_U3552) );
  NOR2_X1 U9502 ( .A1(n7953), .A2(n7943), .ZN(n7945) );
  XNOR2_X1 U9503 ( .A(n7972), .B(n7946), .ZN(n7947) );
  OAI21_X1 U9504 ( .B1(n7948), .B2(n7947), .A(n7963), .ZN(n7949) );
  INV_X1 U9505 ( .A(n7949), .ZN(n7962) );
  INV_X1 U9506 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7951) );
  OAI21_X1 U9507 ( .B1(n7989), .B2(n7951), .A(n7950), .ZN(n7960) );
  NAND2_X1 U9508 ( .A1(n7953), .A2(n7952), .ZN(n7955) );
  NAND2_X1 U9509 ( .A1(n7955), .A2(n7954), .ZN(n7958) );
  NAND2_X1 U9510 ( .A1(n7972), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7956) );
  OAI21_X1 U9511 ( .B1(n7972), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7956), .ZN(
        n7957) );
  NOR2_X1 U9512 ( .A1(n7957), .A2(n7958), .ZN(n7971) );
  AOI211_X1 U9513 ( .C1(n7958), .C2(n7957), .A(n7971), .B(n9449), .ZN(n7959)
         );
  AOI211_X1 U9514 ( .C1(n9456), .C2(n7972), .A(n7960), .B(n7959), .ZN(n7961)
         );
  OAI21_X1 U9515 ( .B1(n7962), .B2(n9753), .A(n7961), .ZN(P2_U3261) );
  XNOR2_X1 U9516 ( .A(n7985), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7965) );
  OAI21_X1 U9517 ( .B1(n7972), .B2(P2_REG1_REG_16__SCAN_IN), .A(n7963), .ZN(
        n7964) );
  NAND2_X1 U9518 ( .A1(n7965), .A2(n7964), .ZN(n7967) );
  NOR2_X1 U9519 ( .A1(n7965), .A2(n7964), .ZN(n7984) );
  INV_X1 U9520 ( .A(n7984), .ZN(n7966) );
  NAND2_X1 U9521 ( .A1(n7967), .A2(n7966), .ZN(n7970) );
  NAND2_X1 U9522 ( .A1(n9755), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U9523 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n7968) );
  OAI211_X1 U9524 ( .C1(n7970), .C2(n9753), .A(n7969), .B(n7968), .ZN(n7977)
         );
  NAND2_X1 U9525 ( .A1(n7985), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7973) );
  OAI21_X1 U9526 ( .B1(n7985), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7973), .ZN(
        n7974) );
  NOR2_X1 U9527 ( .A1(n7975), .A2(n7974), .ZN(n7979) );
  AOI211_X1 U9528 ( .C1(n7975), .C2(n7974), .A(n7979), .B(n9449), .ZN(n7976)
         );
  AOI211_X1 U9529 ( .C1(n9456), .C2(n7985), .A(n7977), .B(n7976), .ZN(n7978)
         );
  INV_X1 U9530 ( .A(n7978), .ZN(P2_U3262) );
  INV_X1 U9531 ( .A(n7995), .ZN(n7994) );
  INV_X1 U9532 ( .A(n7980), .ZN(n7982) );
  NOR2_X1 U9533 ( .A1(n7980), .A2(n8357), .ZN(n8000) );
  INV_X1 U9534 ( .A(n8000), .ZN(n7981) );
  OAI211_X1 U9535 ( .C1(n7982), .C2(P2_REG2_REG_18__SCAN_IN), .A(n7981), .B(
        n9750), .ZN(n7993) );
  INV_X1 U9536 ( .A(n9753), .ZN(n9749) );
  XNOR2_X1 U9537 ( .A(n7995), .B(n7983), .ZN(n7987) );
  AOI21_X1 U9538 ( .B1(n7985), .B2(P2_REG1_REG_17__SCAN_IN), .A(n7984), .ZN(
        n7986) );
  NAND2_X1 U9539 ( .A1(n7987), .A2(n7986), .ZN(n7997) );
  OAI21_X1 U9540 ( .B1(n7987), .B2(n7986), .A(n7997), .ZN(n7991) );
  INV_X1 U9541 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9969) );
  OAI21_X1 U9542 ( .B1(n7989), .B2(n9969), .A(n7988), .ZN(n7990) );
  AOI21_X1 U9543 ( .B1(n9749), .B2(n7991), .A(n7990), .ZN(n7992) );
  OAI211_X1 U9544 ( .C1(n9751), .C2(n7994), .A(n7993), .B(n7992), .ZN(P2_U3263) );
  OR2_X1 U9545 ( .A1(n7995), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U9546 ( .A1(n7997), .A2(n7996), .ZN(n7998) );
  XNOR2_X1 U9547 ( .A(n7998), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8003) );
  OR2_X1 U9548 ( .A1(n8000), .A2(n7999), .ZN(n8001) );
  XNOR2_X1 U9549 ( .A(n8001), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U9550 ( .A1(n8005), .A2(n9750), .ZN(n8002) );
  INV_X1 U9551 ( .A(n8003), .ZN(n8004) );
  NAND2_X1 U9552 ( .A1(n8354), .A2(n8465), .ZN(n8317) );
  NOR2_X2 U9553 ( .A1(n8315), .A2(n8452), .ZN(n8166) );
  INV_X1 U9554 ( .A(n8447), .ZN(n8153) );
  NAND2_X1 U9555 ( .A1(n8074), .A2(n8091), .ZN(n8070) );
  NOR2_X1 U9556 ( .A1(n9785), .A2(n8007), .ZN(n8012) );
  INV_X1 U9557 ( .A(P2_B_REG_SCAN_IN), .ZN(n8008) );
  NOR2_X1 U9558 ( .A1(n8009), .A2(n8008), .ZN(n8010) );
  NOR2_X1 U9559 ( .A1(n8384), .A2(n8010), .ZN(n8041) );
  NAND2_X1 U9560 ( .A1(n8011), .A2(n8041), .ZN(n9497) );
  NOR2_X1 U9561 ( .A1(n8399), .A2(n9497), .ZN(n8017) );
  AOI211_X1 U9562 ( .C1(n8405), .C2(n8380), .A(n8012), .B(n8017), .ZN(n8013)
         );
  OAI21_X1 U9563 ( .B1(n8407), .B2(n8014), .A(n8013), .ZN(P2_U3265) );
  AOI21_X1 U9564 ( .B1(n8016), .B2(n8045), .A(n8015), .ZN(n9501) );
  NAND2_X1 U9565 ( .A1(n9501), .A2(n9767), .ZN(n8019) );
  AOI21_X1 U9566 ( .B1(n8399), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8017), .ZN(
        n8018) );
  OAI211_X1 U9567 ( .C1(n9498), .C2(n9795), .A(n8019), .B(n8018), .ZN(P2_U3266) );
  INV_X1 U9568 ( .A(n8467), .ZN(n8355) );
  NOR2_X1 U9569 ( .A1(n8482), .A2(n8020), .ZN(n8021) );
  INV_X1 U9570 ( .A(n8024), .ZN(n8025) );
  AOI21_X2 U9571 ( .B1(n8389), .B2(n8388), .A(n8025), .ZN(n8366) );
  INV_X1 U9572 ( .A(n8452), .ZN(n8170) );
  NAND2_X1 U9573 ( .A1(n8165), .A2(n4823), .ZN(n8031) );
  INV_X1 U9574 ( .A(n8440), .ZN(n8139) );
  INV_X1 U9575 ( .A(n8415), .ZN(n8066) );
  XNOR2_X1 U9576 ( .A(n8038), .B(n4290), .ZN(n8408) );
  INV_X1 U9577 ( .A(n8408), .ZN(n8052) );
  XNOR2_X1 U9578 ( .A(n8039), .B(n4290), .ZN(n8044) );
  AOI22_X1 U9579 ( .A1(n8042), .A2(n9772), .B1(n8041), .B2(n8040), .ZN(n8043)
         );
  OAI21_X1 U9580 ( .B1(n8044), .B2(n8371), .A(n8043), .ZN(n8412) );
  OAI211_X1 U9581 ( .C1(n8063), .C2(n8410), .A(n9500), .B(n8045), .ZN(n8409)
         );
  NOR2_X1 U9582 ( .A1(n8409), .A2(n9793), .ZN(n8050) );
  INV_X1 U9583 ( .A(n8046), .ZN(n8047) );
  AOI22_X1 U9584 ( .A1(n8399), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8047), .B2(
        n8397), .ZN(n8048) );
  OAI21_X1 U9585 ( .B1(n8410), .B2(n9795), .A(n8048), .ZN(n8049) );
  AOI211_X1 U9586 ( .C1(n8412), .C2(n9788), .A(n8050), .B(n8049), .ZN(n8051)
         );
  OAI21_X1 U9587 ( .B1(n8052), .B2(n8362), .A(n8051), .ZN(P2_U3267) );
  XNOR2_X1 U9588 ( .A(n8054), .B(n8053), .ZN(n8419) );
  NAND2_X1 U9589 ( .A1(n8057), .A2(n9772), .ZN(n8060) );
  NAND2_X1 U9590 ( .A1(n8058), .A2(n9769), .ZN(n8059) );
  OR2_X1 U9591 ( .A1(n8418), .A2(n8399), .ZN(n8069) );
  AOI21_X1 U9592 ( .B1(n8415), .B2(n8070), .A(n8063), .ZN(n8416) );
  AOI22_X1 U9593 ( .A1(n8399), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8064), .B2(
        n8397), .ZN(n8065) );
  OAI21_X1 U9594 ( .B1(n8066), .B2(n9795), .A(n8065), .ZN(n8067) );
  AOI21_X1 U9595 ( .B1(n8416), .B2(n9767), .A(n8067), .ZN(n8068) );
  OAI211_X1 U9596 ( .C1(n8419), .C2(n8362), .A(n8069), .B(n8068), .ZN(P2_U3268) );
  INV_X1 U9597 ( .A(n8091), .ZN(n8072) );
  INV_X1 U9598 ( .A(n8070), .ZN(n8071) );
  AOI21_X1 U9599 ( .B1(n8420), .B2(n8072), .A(n8071), .ZN(n8421) );
  INV_X1 U9600 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8073) );
  OAI22_X1 U9601 ( .A1(n8074), .A2(n9795), .B1(n9788), .B2(n8073), .ZN(n8083)
         );
  OAI211_X1 U9602 ( .C1(n8077), .C2(n8076), .A(n8075), .B(n9776), .ZN(n8079)
         );
  AND2_X1 U9603 ( .A1(n8079), .A2(n8078), .ZN(n8423) );
  NAND2_X1 U9604 ( .A1(n8080), .A2(n8397), .ZN(n8081) );
  AOI21_X1 U9605 ( .B1(n8423), .B2(n8081), .A(n8399), .ZN(n8082) );
  AOI211_X1 U9606 ( .C1(n9767), .C2(n8421), .A(n8083), .B(n8082), .ZN(n8084)
         );
  OAI21_X1 U9607 ( .B1(n8424), .B2(n8362), .A(n8084), .ZN(P2_U3269) );
  XOR2_X1 U9608 ( .A(n8088), .B(n8085), .Z(n8429) );
  NOR2_X1 U9609 ( .A1(n8086), .A2(n9795), .ZN(n8095) );
  XOR2_X1 U9610 ( .A(n8088), .B(n8087), .Z(n8090) );
  AOI211_X1 U9611 ( .C1(n8426), .C2(n8100), .A(n9902), .B(n8091), .ZN(n8425)
         );
  AOI22_X1 U9612 ( .A1(n8425), .A2(n8375), .B1(n8397), .B2(n8092), .ZN(n8093)
         );
  AOI21_X1 U9613 ( .B1(n8428), .B2(n8093), .A(n8399), .ZN(n8094) );
  AOI211_X1 U9614 ( .C1(n8399), .C2(P2_REG2_REG_26__SCAN_IN), .A(n8095), .B(
        n8094), .ZN(n8096) );
  OAI21_X1 U9615 ( .B1(n8429), .B2(n8362), .A(n8096), .ZN(P2_U3270) );
  XOR2_X1 U9616 ( .A(n8102), .B(n8097), .Z(n8434) );
  INV_X1 U9617 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8099) );
  OAI22_X1 U9618 ( .A1(n9788), .A2(n8099), .B1(n8098), .B2(n9792), .ZN(n8110)
         );
  INV_X1 U9619 ( .A(n8100), .ZN(n8101) );
  AOI211_X1 U9620 ( .C1(n8432), .C2(n4413), .A(n9902), .B(n8101), .ZN(n8431)
         );
  OAI21_X1 U9621 ( .B1(n8103), .B2(n8102), .A(n9776), .ZN(n8107) );
  INV_X1 U9622 ( .A(n8104), .ZN(n8105) );
  OAI21_X1 U9623 ( .B1(n8107), .B2(n8106), .A(n8105), .ZN(n8430) );
  AOI21_X1 U9624 ( .B1(n8431), .B2(n8375), .A(n8430), .ZN(n8108) );
  NOR2_X1 U9625 ( .A1(n8108), .A2(n8399), .ZN(n8109) );
  AOI211_X1 U9626 ( .C1(n8380), .C2(n8432), .A(n8110), .B(n8109), .ZN(n8111)
         );
  OAI21_X1 U9627 ( .B1(n8434), .B2(n8362), .A(n8111), .ZN(P2_U3271) );
  AOI21_X1 U9628 ( .B1(n8120), .B2(n8113), .A(n8112), .ZN(n8439) );
  AOI21_X1 U9629 ( .B1(n8435), .B2(n8134), .A(n8114), .ZN(n8436) );
  INV_X1 U9630 ( .A(n8115), .ZN(n8116) );
  AOI22_X1 U9631 ( .A1(n8399), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8116), .B2(
        n8397), .ZN(n8117) );
  OAI21_X1 U9632 ( .B1(n4411), .B2(n9795), .A(n8117), .ZN(n8126) );
  AND2_X1 U9633 ( .A1(n8129), .A2(n8118), .ZN(n8121) );
  OAI211_X1 U9634 ( .C1(n8121), .C2(n8120), .A(n9776), .B(n8119), .ZN(n8124)
         );
  AOI22_X1 U9635 ( .A1(n8122), .A2(n9769), .B1(n9772), .B2(n8154), .ZN(n8123)
         );
  AND2_X1 U9636 ( .A1(n8124), .A2(n8123), .ZN(n8438) );
  NOR2_X1 U9637 ( .A1(n8438), .A2(n8399), .ZN(n8125) );
  AOI211_X1 U9638 ( .C1(n8436), .C2(n9767), .A(n8126), .B(n8125), .ZN(n8127)
         );
  OAI21_X1 U9639 ( .B1(n8439), .B2(n8362), .A(n8127), .ZN(P2_U3272) );
  AND2_X1 U9640 ( .A1(n8155), .A2(n8128), .ZN(n8131) );
  OAI21_X1 U9641 ( .B1(n8131), .B2(n8130), .A(n8129), .ZN(n8133) );
  AOI222_X1 U9642 ( .A1(n9776), .A2(n8133), .B1(n8132), .B2(n9769), .C1(n8175), 
        .C2(n9772), .ZN(n8446) );
  INV_X1 U9643 ( .A(n8134), .ZN(n8135) );
  AOI21_X1 U9644 ( .B1(n8440), .B2(n8147), .A(n8135), .ZN(n8441) );
  INV_X1 U9645 ( .A(n8136), .ZN(n8137) );
  AOI22_X1 U9646 ( .A1(n8399), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8137), .B2(
        n8397), .ZN(n8138) );
  OAI21_X1 U9647 ( .B1(n8139), .B2(n9795), .A(n8138), .ZN(n8140) );
  AOI21_X1 U9648 ( .B1(n8441), .B2(n9767), .A(n8140), .ZN(n8145) );
  OR2_X1 U9649 ( .A1(n8142), .A2(n8141), .ZN(n8443) );
  NAND3_X1 U9650 ( .A1(n8443), .A2(n8442), .A3(n8143), .ZN(n8144) );
  OAI211_X1 U9651 ( .C1(n8446), .C2(n8399), .A(n8145), .B(n8144), .ZN(P2_U3273) );
  XNOR2_X1 U9652 ( .A(n8146), .B(n8156), .ZN(n8451) );
  INV_X1 U9653 ( .A(n8166), .ZN(n8149) );
  INV_X1 U9654 ( .A(n8147), .ZN(n8148) );
  AOI21_X1 U9655 ( .B1(n8447), .B2(n8149), .A(n8148), .ZN(n8448) );
  INV_X1 U9656 ( .A(n8150), .ZN(n8151) );
  AOI22_X1 U9657 ( .A1(n8399), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8151), .B2(
        n8397), .ZN(n8152) );
  OAI21_X1 U9658 ( .B1(n8153), .B2(n9795), .A(n8152), .ZN(n8163) );
  AND2_X1 U9659 ( .A1(n8154), .A2(n9769), .ZN(n8161) );
  INV_X1 U9660 ( .A(n8155), .ZN(n8159) );
  AOI21_X1 U9661 ( .B1(n8171), .B2(n8157), .A(n8156), .ZN(n8158) );
  NOR3_X1 U9662 ( .A1(n8159), .A2(n8158), .A3(n8371), .ZN(n8160) );
  AOI211_X1 U9663 ( .C1(n9772), .C2(n8326), .A(n8161), .B(n8160), .ZN(n8450)
         );
  NOR2_X1 U9664 ( .A1(n8450), .A2(n8399), .ZN(n8162) );
  AOI211_X1 U9665 ( .C1(n8448), .C2(n9767), .A(n8163), .B(n8162), .ZN(n8164)
         );
  OAI21_X1 U9666 ( .B1(n8451), .B2(n8362), .A(n8164), .ZN(P2_U3274) );
  XNOR2_X1 U9667 ( .A(n8165), .B(n8173), .ZN(n8456) );
  AOI21_X1 U9668 ( .B1(n8452), .B2(n8315), .A(n8166), .ZN(n8453) );
  INV_X1 U9669 ( .A(n8167), .ZN(n8168) );
  AOI22_X1 U9670 ( .A1(n8399), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8168), .B2(
        n8397), .ZN(n8169) );
  OAI21_X1 U9671 ( .B1(n8170), .B2(n9795), .A(n8169), .ZN(n8178) );
  OAI21_X1 U9672 ( .B1(n8173), .B2(n8172), .A(n8171), .ZN(n8176) );
  AOI222_X1 U9673 ( .A1(n9776), .A2(n8176), .B1(n8175), .B2(n9769), .C1(n8174), 
        .C2(n9772), .ZN(n8455) );
  NOR2_X1 U9674 ( .A1(n8455), .A2(n8399), .ZN(n8177) );
  AOI211_X1 U9675 ( .C1(n8453), .C2(n9767), .A(n8178), .B(n8177), .ZN(n8179)
         );
  OAI21_X1 U9676 ( .B1(n8362), .B2(n8456), .A(n8179), .ZN(n8313) );
  AOI22_X1 U9677 ( .A1(n9833), .A2(keyinput55), .B1(n4775), .B2(keyinput1), 
        .ZN(n8180) );
  OAI221_X1 U9678 ( .B1(n9833), .B2(keyinput55), .C1(n4775), .C2(keyinput1), 
        .A(n8180), .ZN(n8188) );
  INV_X1 U9679 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9502) );
  INV_X1 U9680 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9669) );
  AOI22_X1 U9681 ( .A1(n9502), .A2(keyinput37), .B1(n9669), .B2(keyinput27), 
        .ZN(n8181) );
  OAI221_X1 U9682 ( .B1(n9502), .B2(keyinput37), .C1(n9669), .C2(keyinput27), 
        .A(n8181), .ZN(n8187) );
  INV_X1 U9683 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U9684 ( .A1(n9899), .A2(keyinput15), .B1(n4879), .B2(keyinput7), 
        .ZN(n8182) );
  OAI221_X1 U9685 ( .B1(n9899), .B2(keyinput15), .C1(n4879), .C2(keyinput7), 
        .A(n8182), .ZN(n8186) );
  INV_X1 U9686 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8184) );
  AOI22_X1 U9687 ( .A1(n8283), .A2(keyinput34), .B1(n8184), .B2(keyinput50), 
        .ZN(n8183) );
  OAI221_X1 U9688 ( .B1(n8283), .B2(keyinput34), .C1(n8184), .C2(keyinput50), 
        .A(n8183), .ZN(n8185) );
  OR4_X1 U9689 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), .ZN(n8194) );
  AOI22_X1 U9690 ( .A1(n5474), .A2(keyinput36), .B1(n8288), .B2(keyinput21), 
        .ZN(n8189) );
  OAI221_X1 U9691 ( .B1(n5474), .B2(keyinput36), .C1(n8288), .C2(keyinput21), 
        .A(n8189), .ZN(n8193) );
  INV_X1 U9692 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9932) );
  INV_X1 U9693 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8279) );
  AOI22_X1 U9694 ( .A1(n9932), .A2(keyinput33), .B1(n8279), .B2(keyinput16), 
        .ZN(n8190) );
  OAI221_X1 U9695 ( .B1(n9932), .B2(keyinput33), .C1(n8279), .C2(keyinput16), 
        .A(n8190), .ZN(n8192) );
  INV_X1 U9696 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9667) );
  XNOR2_X1 U9697 ( .A(n9667), .B(keyinput6), .ZN(n8191) );
  NOR4_X1 U9698 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n8218)
         );
  XOR2_X1 U9699 ( .A(keyinput25), .B(n9822), .Z(n8217) );
  XOR2_X1 U9700 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput11), .Z(n8204) );
  XNOR2_X1 U9701 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput61), .ZN(n8198) );
  XNOR2_X1 U9702 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput4), .ZN(n8197) );
  XNOR2_X1 U9703 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput39), .ZN(n8196) );
  XNOR2_X1 U9704 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput40), .ZN(n8195) );
  NAND4_X1 U9705 ( .A1(n8198), .A2(n8197), .A3(n8196), .A4(n8195), .ZN(n8203)
         );
  XNOR2_X1 U9706 ( .A(n8199), .B(keyinput10), .ZN(n8202) );
  XNOR2_X1 U9707 ( .A(keyinput60), .B(n8200), .ZN(n8201) );
  NOR4_X1 U9708 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(n8216)
         );
  AOI22_X1 U9709 ( .A1(n8206), .A2(keyinput17), .B1(keyinput3), .B2(n8686), 
        .ZN(n8205) );
  OAI221_X1 U9710 ( .B1(n8206), .B2(keyinput17), .C1(n8686), .C2(keyinput3), 
        .A(n8205), .ZN(n8214) );
  AOI22_X1 U9711 ( .A1(n6593), .A2(keyinput44), .B1(n8208), .B2(keyinput0), 
        .ZN(n8207) );
  OAI221_X1 U9712 ( .B1(n6593), .B2(keyinput44), .C1(n8208), .C2(keyinput0), 
        .A(n8207), .ZN(n8213) );
  AOI22_X1 U9713 ( .A1(n9806), .A2(keyinput8), .B1(P1_U3084), .B2(keyinput2), 
        .ZN(n8209) );
  OAI221_X1 U9714 ( .B1(n9806), .B2(keyinput8), .C1(P1_U3084), .C2(keyinput2), 
        .A(n8209), .ZN(n8212) );
  INV_X1 U9715 ( .A(P1_WR_REG_SCAN_IN), .ZN(n8210) );
  XNOR2_X1 U9716 ( .A(n8210), .B(keyinput28), .ZN(n8211) );
  NOR4_X1 U9717 ( .A1(n8214), .A2(n8213), .A3(n8212), .A4(n8211), .ZN(n8215)
         );
  NAND4_X1 U9718 ( .A1(n8218), .A2(n8217), .A3(n8216), .A4(n8215), .ZN(n8253)
         );
  AOI22_X1 U9719 ( .A1(n8221), .A2(keyinput45), .B1(keyinput5), .B2(n8220), 
        .ZN(n8219) );
  OAI221_X1 U9720 ( .B1(n8221), .B2(keyinput45), .C1(n8220), .C2(keyinput5), 
        .A(n8219), .ZN(n8229) );
  AOI22_X1 U9721 ( .A1(n8224), .A2(keyinput13), .B1(keyinput38), .B2(n8223), 
        .ZN(n8222) );
  OAI221_X1 U9722 ( .B1(n8224), .B2(keyinput13), .C1(n8223), .C2(keyinput38), 
        .A(n8222), .ZN(n8228) );
  AOI22_X1 U9723 ( .A1(n8293), .A2(keyinput14), .B1(keyinput24), .B2(n8226), 
        .ZN(n8225) );
  OAI221_X1 U9724 ( .B1(n8293), .B2(keyinput14), .C1(n8226), .C2(keyinput24), 
        .A(n8225), .ZN(n8227) );
  NOR3_X1 U9725 ( .A1(n8229), .A2(n8228), .A3(n8227), .ZN(n8251) );
  AOI22_X1 U9726 ( .A1(n4911), .A2(keyinput46), .B1(keyinput30), .B2(n7376), 
        .ZN(n8230) );
  OAI221_X1 U9727 ( .B1(n4911), .B2(keyinput46), .C1(n7376), .C2(keyinput30), 
        .A(n8230), .ZN(n8234) );
  INV_X1 U9728 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8232) );
  INV_X1 U9729 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9668) );
  AOI22_X1 U9730 ( .A1(n8232), .A2(keyinput18), .B1(n9668), .B2(keyinput23), 
        .ZN(n8231) );
  OAI221_X1 U9731 ( .B1(n8232), .B2(keyinput18), .C1(n9668), .C2(keyinput23), 
        .A(n8231), .ZN(n8233) );
  NOR2_X1 U9732 ( .A1(n8234), .A2(n8233), .ZN(n8250) );
  INV_X1 U9733 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9549) );
  AOI22_X1 U9734 ( .A1(n6602), .A2(keyinput20), .B1(keyinput59), .B2(n9549), 
        .ZN(n8235) );
  OAI221_X1 U9735 ( .B1(n6602), .B2(keyinput20), .C1(n9549), .C2(keyinput59), 
        .A(n8235), .ZN(n8243) );
  INV_X1 U9736 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8238) );
  AOI22_X1 U9737 ( .A1(n8238), .A2(keyinput52), .B1(n8237), .B2(keyinput63), 
        .ZN(n8236) );
  OAI221_X1 U9738 ( .B1(n8238), .B2(keyinput52), .C1(n8237), .C2(keyinput63), 
        .A(n8236), .ZN(n8242) );
  XNOR2_X1 U9739 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput31), .ZN(n8240) );
  XNOR2_X1 U9740 ( .A(keyinput53), .B(P1_REG0_REG_10__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U9741 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  NOR3_X1 U9742 ( .A1(n8243), .A2(n8242), .A3(n8241), .ZN(n8249) );
  INV_X1 U9743 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U9744 ( .A1(n8357), .A2(keyinput12), .B1(keyinput56), .B2(n9879), 
        .ZN(n8244) );
  OAI221_X1 U9745 ( .B1(n8357), .B2(keyinput12), .C1(n9879), .C2(keyinput56), 
        .A(n8244), .ZN(n8247) );
  INV_X1 U9746 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9670) );
  AOI22_X1 U9747 ( .A1(n9670), .A2(keyinput62), .B1(keyinput48), .B2(n6438), 
        .ZN(n8245) );
  OAI221_X1 U9748 ( .B1(n9670), .B2(keyinput62), .C1(n6438), .C2(keyinput48), 
        .A(n8245), .ZN(n8246) );
  NOR2_X1 U9749 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  NAND4_X1 U9750 ( .A1(n8251), .A2(n8250), .A3(n8249), .A4(n8248), .ZN(n8252)
         );
  NOR2_X1 U9751 ( .A1(n8253), .A2(n8252), .ZN(n8278) );
  INV_X1 U9752 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9973) );
  INV_X1 U9753 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9728) );
  AOI22_X1 U9754 ( .A1(n9973), .A2(keyinput51), .B1(n9728), .B2(keyinput26), 
        .ZN(n8254) );
  OAI221_X1 U9755 ( .B1(n9973), .B2(keyinput51), .C1(n9728), .C2(keyinput26), 
        .A(n8254), .ZN(n8265) );
  AOI22_X1 U9756 ( .A1(n9913), .A2(keyinput42), .B1(n8256), .B2(keyinput22), 
        .ZN(n8255) );
  OAI221_X1 U9757 ( .B1(n9913), .B2(keyinput42), .C1(n8256), .C2(keyinput22), 
        .A(n8255), .ZN(n8264) );
  INV_X1 U9758 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n8258) );
  AOI22_X1 U9759 ( .A1(n8259), .A2(keyinput57), .B1(keyinput35), .B2(n8258), 
        .ZN(n8257) );
  OAI221_X1 U9760 ( .B1(n8259), .B2(keyinput57), .C1(n8258), .C2(keyinput35), 
        .A(n8257), .ZN(n8263) );
  INV_X1 U9761 ( .A(SI_18_), .ZN(n8261) );
  AOI22_X1 U9762 ( .A1(n7107), .A2(keyinput47), .B1(n8261), .B2(keyinput29), 
        .ZN(n8260) );
  OAI221_X1 U9763 ( .B1(n7107), .B2(keyinput47), .C1(n8261), .C2(keyinput29), 
        .A(n8260), .ZN(n8262) );
  NOR4_X1 U9764 ( .A1(n8265), .A2(n8264), .A3(n8263), .A4(n8262), .ZN(n8277)
         );
  AOI22_X1 U9765 ( .A1(n5948), .A2(keyinput43), .B1(keyinput32), .B2(n8267), 
        .ZN(n8266) );
  OAI221_X1 U9766 ( .B1(n5948), .B2(keyinput43), .C1(n8267), .C2(keyinput32), 
        .A(n8266), .ZN(n8275) );
  AOI22_X1 U9767 ( .A1(n6079), .A2(keyinput54), .B1(n8585), .B2(keyinput49), 
        .ZN(n8268) );
  OAI221_X1 U9768 ( .B1(n6079), .B2(keyinput54), .C1(n8585), .C2(keyinput49), 
        .A(n8268), .ZN(n8274) );
  INV_X1 U9769 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9666) );
  AOI22_X1 U9770 ( .A1(n9666), .A2(keyinput58), .B1(keyinput19), .B2(n8299), 
        .ZN(n8269) );
  OAI221_X1 U9771 ( .B1(n9666), .B2(keyinput58), .C1(n8299), .C2(keyinput19), 
        .A(n8269), .ZN(n8273) );
  AOI22_X1 U9772 ( .A1(n9918), .A2(keyinput41), .B1(keyinput9), .B2(n8271), 
        .ZN(n8270) );
  OAI221_X1 U9773 ( .B1(n9918), .B2(keyinput41), .C1(n8271), .C2(keyinput9), 
        .A(n8270), .ZN(n8272) );
  NOR4_X1 U9774 ( .A1(n8275), .A2(n8274), .A3(n8273), .A4(n8272), .ZN(n8276)
         );
  NAND3_X1 U9775 ( .A1(n8278), .A2(n8277), .A3(n8276), .ZN(n8311) );
  NOR4_X1 U9776 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n9913), .A3(n5474), .A4(
        n8279), .ZN(n8308) );
  NAND4_X1 U9777 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P2_DATAO_REG_27__SCAN_IN), 
        .A3(SI_25_), .A4(P1_U3084), .ZN(n8282) );
  NAND4_X1 U9778 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .A3(P1_REG3_REG_7__SCAN_IN), .A4(P2_DATAO_REG_30__SCAN_IN), .ZN(n8281)
         );
  NAND4_X1 U9779 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_REG2_REG_10__SCAN_IN), .A4(P2_REG0_REG_30__SCAN_IN), .ZN(n8280) );
  OR3_X1 U9780 ( .A1(n8282), .A2(n8281), .A3(n8280), .ZN(n8306) );
  NOR3_X1 U9781 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(P2_REG2_REG_15__SCAN_IN), 
        .A3(n9879), .ZN(n8298) );
  NAND4_X1 U9782 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_REG1_REG_21__SCAN_IN), .A4(P2_REG2_REG_21__SCAN_IN), .ZN(n8285) );
  NAND4_X1 U9783 ( .A1(n9932), .A2(n8283), .A3(P2_REG0_REG_11__SCAN_IN), .A4(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n8284) );
  NOR2_X1 U9784 ( .A1(n8285), .A2(n8284), .ZN(n8297) );
  INV_X1 U9785 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8287) );
  NAND4_X1 U9786 ( .A1(n8287), .A2(n8286), .A3(P2_IR_REG_1__SCAN_IN), .A4(
        P2_REG3_REG_14__SCAN_IN), .ZN(n8295) );
  NAND4_X1 U9787 ( .A1(SI_18_), .A2(SI_9_), .A3(P2_REG3_REG_19__SCAN_IN), .A4(
        n8288), .ZN(n8289) );
  NOR2_X1 U9788 ( .A1(n8289), .A2(n8357), .ZN(n8291) );
  NOR4_X1 U9789 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG2_REG_22__SCAN_IN), 
        .A3(P1_REG1_REG_13__SCAN_IN), .A4(P1_REG2_REG_15__SCAN_IN), .ZN(n8290)
         );
  AND2_X1 U9790 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  NAND4_X1 U9791 ( .A1(n8293), .A2(P2_DATAO_REG_2__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .A4(n8292), .ZN(n8294) );
  NOR2_X1 U9792 ( .A1(n8295), .A2(n8294), .ZN(n8296) );
  NAND4_X1 U9793 ( .A1(n8298), .A2(n8297), .A3(n9973), .A4(n8296), .ZN(n8305)
         );
  NOR4_X1 U9794 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .A3(
        n9822), .A4(n8299), .ZN(n8303) );
  NOR4_X1 U9795 ( .A1(P1_D_REG_1__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .A3(
        P2_REG1_REG_24__SCAN_IN), .A4(P1_WR_REG_SCAN_IN), .ZN(n8302) );
  NOR4_X1 U9796 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(P1_REG0_REG_9__SCAN_IN), 
        .A3(P1_REG1_REG_1__SCAN_IN), .A4(P2_REG1_REG_23__SCAN_IN), .ZN(n8301)
         );
  NOR4_X1 U9797 ( .A1(P1_REG0_REG_13__SCAN_IN), .A2(P1_REG1_REG_12__SCAN_IN), 
        .A3(P1_REG2_REG_8__SCAN_IN), .A4(P1_REG2_REG_4__SCAN_IN), .ZN(n8300)
         );
  NAND4_X1 U9798 ( .A1(n8303), .A2(n8302), .A3(n8301), .A4(n8300), .ZN(n8304)
         );
  NOR3_X1 U9799 ( .A1(n8306), .A2(n8305), .A3(n8304), .ZN(n8307) );
  NAND3_X1 U9800 ( .A1(n8309), .A2(n8308), .A3(n8307), .ZN(n8310) );
  XNOR2_X1 U9801 ( .A(n8311), .B(n8310), .ZN(n8312) );
  XNOR2_X1 U9802 ( .A(n8313), .B(n8312), .ZN(P2_U3275) );
  XNOR2_X1 U9803 ( .A(n8314), .B(n8323), .ZN(n8461) );
  INV_X1 U9804 ( .A(n8315), .ZN(n8316) );
  AOI21_X1 U9805 ( .B1(n8457), .B2(n8317), .A(n8316), .ZN(n8458) );
  INV_X1 U9806 ( .A(n8457), .ZN(n8321) );
  INV_X1 U9807 ( .A(n8318), .ZN(n8319) );
  AOI22_X1 U9808 ( .A1(n8399), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8319), .B2(
        n8397), .ZN(n8320) );
  OAI21_X1 U9809 ( .B1(n8321), .B2(n9795), .A(n8320), .ZN(n8329) );
  NOR2_X1 U9810 ( .A1(n4308), .A2(n8322), .ZN(n8324) );
  XNOR2_X1 U9811 ( .A(n8324), .B(n8323), .ZN(n8325) );
  AOI222_X1 U9812 ( .A1(n8327), .A2(n9772), .B1(n8326), .B2(n9769), .C1(n9776), 
        .C2(n8325), .ZN(n8460) );
  NOR2_X1 U9813 ( .A1(n8460), .A2(n8399), .ZN(n8328) );
  AOI211_X1 U9814 ( .C1(n8458), .C2(n9767), .A(n8329), .B(n8328), .ZN(n8330)
         );
  OAI21_X1 U9815 ( .B1(n8362), .B2(n8461), .A(n8330), .ZN(P2_U3276) );
  XNOR2_X1 U9816 ( .A(n8331), .B(n8332), .ZN(n8462) );
  INV_X1 U9817 ( .A(n8462), .ZN(n8347) );
  AOI21_X1 U9818 ( .B1(n8333), .B2(n8332), .A(n4308), .ZN(n8334) );
  OAI222_X1 U9819 ( .A1(n8384), .A2(n8335), .B1(n8386), .B2(n8373), .C1(n8371), 
        .C2(n8334), .ZN(n8340) );
  INV_X1 U9820 ( .A(n8336), .ZN(n8338) );
  XNOR2_X1 U9821 ( .A(n8354), .B(n8344), .ZN(n8337) );
  AOI21_X1 U9822 ( .B1(n9500), .B2(n8337), .A(n8340), .ZN(n8464) );
  OAI21_X1 U9823 ( .B1(n8338), .B2(n8347), .A(n8464), .ZN(n8339) );
  OAI211_X1 U9824 ( .C1(n8375), .C2(n8340), .A(n8339), .B(n9785), .ZN(n8346)
         );
  OAI22_X1 U9825 ( .A1(n9785), .A2(n8342), .B1(n8341), .B2(n9792), .ZN(n8343)
         );
  AOI21_X1 U9826 ( .B1(n8344), .B2(n8380), .A(n8343), .ZN(n8345) );
  OAI211_X1 U9827 ( .C1(n8347), .C2(n9798), .A(n8346), .B(n8345), .ZN(P2_U3277) );
  XOR2_X1 U9828 ( .A(n8351), .B(n8348), .Z(n8471) );
  AOI21_X1 U9829 ( .B1(n8351), .B2(n8350), .A(n8349), .ZN(n8352) );
  OAI222_X1 U9830 ( .A1(n8384), .A2(n8353), .B1(n8386), .B2(n8385), .C1(n8371), 
        .C2(n8352), .ZN(n8466) );
  NAND2_X1 U9831 ( .A1(n8466), .A2(n9788), .ZN(n8361) );
  AOI21_X1 U9832 ( .B1(n8467), .B2(n8363), .A(n8354), .ZN(n8468) );
  NOR2_X1 U9833 ( .A1(n8355), .A2(n9795), .ZN(n8359) );
  OAI22_X1 U9834 ( .A1(n9788), .A2(n8357), .B1(n8356), .B2(n9792), .ZN(n8358)
         );
  AOI211_X1 U9835 ( .C1(n8468), .C2(n9767), .A(n8359), .B(n8358), .ZN(n8360)
         );
  OAI211_X1 U9836 ( .C1(n8471), .C2(n8362), .A(n8361), .B(n8360), .ZN(P2_U3278) );
  INV_X1 U9837 ( .A(n8363), .ZN(n8364) );
  AOI211_X1 U9838 ( .C1(n8474), .C2(n8395), .A(n9902), .B(n8364), .ZN(n8473)
         );
  OAI21_X1 U9839 ( .B1(n8366), .B2(n8368), .A(n8365), .ZN(n8367) );
  INV_X1 U9840 ( .A(n8367), .ZN(n8476) );
  NOR2_X1 U9841 ( .A1(n8476), .A2(n9781), .ZN(n8374) );
  XNOR2_X1 U9842 ( .A(n8369), .B(n8368), .ZN(n8370) );
  OAI222_X1 U9843 ( .A1(n8384), .A2(n8373), .B1(n8386), .B2(n8372), .C1(n8371), 
        .C2(n8370), .ZN(n8472) );
  AOI211_X1 U9844 ( .C1(n8473), .C2(n8375), .A(n8374), .B(n8472), .ZN(n8382)
         );
  OAI22_X1 U9845 ( .A1(n9785), .A2(n8377), .B1(n8376), .B2(n9792), .ZN(n8379)
         );
  NOR2_X1 U9846 ( .A1(n8476), .A2(n9798), .ZN(n8378) );
  AOI211_X1 U9847 ( .C1(n8380), .C2(n8474), .A(n8379), .B(n8378), .ZN(n8381)
         );
  OAI21_X1 U9848 ( .B1(n8382), .B2(n8399), .A(n8381), .ZN(P2_U3279) );
  XNOR2_X1 U9849 ( .A(n8383), .B(n8388), .ZN(n8392) );
  OAI22_X1 U9850 ( .A1(n8387), .A2(n8386), .B1(n8385), .B2(n8384), .ZN(n8391)
         );
  XNOR2_X1 U9851 ( .A(n8389), .B(n8388), .ZN(n8481) );
  NOR2_X1 U9852 ( .A1(n8481), .A2(n9781), .ZN(n8390) );
  AOI211_X1 U9853 ( .C1(n8392), .C2(n9776), .A(n8391), .B(n8390), .ZN(n8480)
         );
  NAND2_X1 U9854 ( .A1(n8393), .A2(n8477), .ZN(n8394) );
  AND2_X1 U9855 ( .A1(n8395), .A2(n8394), .ZN(n8478) );
  INV_X1 U9856 ( .A(n8477), .ZN(n8401) );
  INV_X1 U9857 ( .A(n8396), .ZN(n8398) );
  AOI22_X1 U9858 ( .A1(n8399), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8398), .B2(
        n8397), .ZN(n8400) );
  OAI21_X1 U9859 ( .B1(n8401), .B2(n9795), .A(n8400), .ZN(n8403) );
  NOR2_X1 U9860 ( .A1(n8481), .A2(n9798), .ZN(n8402) );
  AOI211_X1 U9861 ( .C1(n8478), .C2(n9767), .A(n8403), .B(n8402), .ZN(n8404)
         );
  OAI21_X1 U9862 ( .B1(n8480), .B2(n8399), .A(n8404), .ZN(P2_U3280) );
  NAND2_X1 U9863 ( .A1(n8405), .A2(n8489), .ZN(n8406) );
  OAI211_X1 U9864 ( .C1(n8407), .C2(n9902), .A(n9497), .B(n8406), .ZN(n8504)
         );
  MUX2_X1 U9865 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8504), .S(n9927), .Z(
        P2_U3551) );
  NAND2_X1 U9866 ( .A1(n8408), .A2(n9907), .ZN(n8414) );
  OAI21_X1 U9867 ( .B1(n8410), .B2(n9900), .A(n8409), .ZN(n8411) );
  NOR2_X1 U9868 ( .A1(n8412), .A2(n8411), .ZN(n8413) );
  NAND2_X1 U9869 ( .A1(n8414), .A2(n8413), .ZN(n8505) );
  MUX2_X1 U9870 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8505), .S(n9927), .Z(
        P2_U3549) );
  AOI22_X1 U9871 ( .A1(n8416), .A2(n9500), .B1(n8489), .B2(n8415), .ZN(n8417)
         );
  OAI211_X1 U9872 ( .C1(n8419), .C2(n8494), .A(n8418), .B(n8417), .ZN(n8506)
         );
  MUX2_X1 U9873 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8506), .S(n9927), .Z(
        P2_U3548) );
  AOI22_X1 U9874 ( .A1(n8421), .A2(n9500), .B1(n8489), .B2(n8420), .ZN(n8422)
         );
  OAI211_X1 U9875 ( .C1(n8424), .C2(n8494), .A(n8423), .B(n8422), .ZN(n8507)
         );
  MUX2_X1 U9876 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8507), .S(n9927), .Z(
        P2_U3547) );
  AOI21_X1 U9877 ( .B1(n8489), .B2(n8426), .A(n8425), .ZN(n8427) );
  OAI211_X1 U9878 ( .C1(n8429), .C2(n8494), .A(n8428), .B(n8427), .ZN(n8508)
         );
  MUX2_X1 U9879 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8508), .S(n9927), .Z(
        P2_U3546) );
  AOI211_X1 U9880 ( .C1(n8489), .C2(n8432), .A(n8431), .B(n8430), .ZN(n8433)
         );
  OAI21_X1 U9881 ( .B1(n8434), .B2(n8494), .A(n8433), .ZN(n8509) );
  MUX2_X1 U9882 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8509), .S(n9927), .Z(
        P2_U3545) );
  AOI22_X1 U9883 ( .A1(n8436), .A2(n9500), .B1(n8489), .B2(n8435), .ZN(n8437)
         );
  OAI211_X1 U9884 ( .C1(n8439), .C2(n8494), .A(n8438), .B(n8437), .ZN(n8510)
         );
  MUX2_X1 U9885 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8510), .S(n9927), .Z(
        P2_U3544) );
  AOI22_X1 U9886 ( .A1(n8441), .A2(n9500), .B1(n8489), .B2(n8440), .ZN(n8445)
         );
  NAND3_X1 U9887 ( .A1(n8443), .A2(n8442), .A3(n9907), .ZN(n8444) );
  NAND3_X1 U9888 ( .A1(n8446), .A2(n8445), .A3(n8444), .ZN(n8511) );
  MUX2_X1 U9889 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8511), .S(n9927), .Z(
        P2_U3543) );
  AOI22_X1 U9890 ( .A1(n8448), .A2(n9500), .B1(n8489), .B2(n8447), .ZN(n8449)
         );
  OAI211_X1 U9891 ( .C1(n8494), .C2(n8451), .A(n8450), .B(n8449), .ZN(n8512)
         );
  MUX2_X1 U9892 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8512), .S(n9927), .Z(
        P2_U3542) );
  AOI22_X1 U9893 ( .A1(n8453), .A2(n9500), .B1(n8489), .B2(n8452), .ZN(n8454)
         );
  OAI211_X1 U9894 ( .C1(n8494), .C2(n8456), .A(n8455), .B(n8454), .ZN(n8513)
         );
  MUX2_X1 U9895 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8513), .S(n9927), .Z(
        P2_U3541) );
  AOI22_X1 U9896 ( .A1(n8458), .A2(n9500), .B1(n8489), .B2(n8457), .ZN(n8459)
         );
  OAI211_X1 U9897 ( .C1(n8494), .C2(n8461), .A(n8460), .B(n8459), .ZN(n8514)
         );
  MUX2_X1 U9898 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8514), .S(n9927), .Z(
        P2_U3540) );
  NAND2_X1 U9899 ( .A1(n8462), .A2(n9907), .ZN(n8463) );
  OAI211_X1 U9900 ( .C1(n8465), .C2(n9900), .A(n8464), .B(n8463), .ZN(n8515)
         );
  MUX2_X1 U9901 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8515), .S(n9927), .Z(
        P2_U3539) );
  INV_X1 U9902 ( .A(n8466), .ZN(n8470) );
  AOI22_X1 U9903 ( .A1(n8468), .A2(n9500), .B1(n8489), .B2(n8467), .ZN(n8469)
         );
  OAI211_X1 U9904 ( .C1(n8494), .C2(n8471), .A(n8470), .B(n8469), .ZN(n8516)
         );
  MUX2_X1 U9905 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8516), .S(n9927), .Z(
        P2_U3538) );
  AOI211_X1 U9906 ( .C1(n8489), .C2(n8474), .A(n8473), .B(n8472), .ZN(n8475)
         );
  OAI21_X1 U9907 ( .B1(n8494), .B2(n8476), .A(n8475), .ZN(n8517) );
  MUX2_X1 U9908 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8517), .S(n9927), .Z(
        P2_U3537) );
  AOI22_X1 U9909 ( .A1(n8478), .A2(n9500), .B1(n8489), .B2(n8477), .ZN(n8479)
         );
  OAI211_X1 U9910 ( .C1(n8500), .C2(n8481), .A(n8480), .B(n8479), .ZN(n8518)
         );
  MUX2_X1 U9911 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8518), .S(n9927), .Z(
        P2_U3536) );
  AOI22_X1 U9912 ( .A1(n8483), .A2(n9500), .B1(n8489), .B2(n8482), .ZN(n8484)
         );
  OAI211_X1 U9913 ( .C1(n8494), .C2(n8486), .A(n8485), .B(n8484), .ZN(n8519)
         );
  MUX2_X1 U9914 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8519), .S(n9927), .Z(
        P2_U3535) );
  INV_X1 U9915 ( .A(n8487), .ZN(n8493) );
  AOI22_X1 U9916 ( .A1(n8490), .A2(n9500), .B1(n8489), .B2(n8488), .ZN(n8491)
         );
  OAI211_X1 U9917 ( .C1(n8494), .C2(n8493), .A(n8492), .B(n8491), .ZN(n8520)
         );
  MUX2_X1 U9918 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8520), .S(n9927), .Z(
        P2_U3534) );
  INV_X1 U9919 ( .A(n8495), .ZN(n8496) );
  OAI22_X1 U9920 ( .A1(n8497), .A2(n9902), .B1(n8496), .B2(n9900), .ZN(n8498)
         );
  INV_X1 U9921 ( .A(n8498), .ZN(n8499) );
  OAI21_X1 U9922 ( .B1(n8501), .B2(n8500), .A(n8499), .ZN(n8502) );
  OR2_X1 U9923 ( .A1(n8503), .A2(n8502), .ZN(n8521) );
  MUX2_X1 U9924 ( .A(n8521), .B(P2_REG1_REG_13__SCAN_IN), .S(n9925), .Z(
        P2_U3533) );
  MUX2_X1 U9925 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8504), .S(n9910), .Z(
        P2_U3519) );
  MUX2_X1 U9926 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8505), .S(n9910), .Z(
        P2_U3517) );
  MUX2_X1 U9927 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8506), .S(n9910), .Z(
        P2_U3516) );
  MUX2_X1 U9928 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8507), .S(n9910), .Z(
        P2_U3515) );
  MUX2_X1 U9929 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8508), .S(n9910), .Z(
        P2_U3514) );
  MUX2_X1 U9930 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8509), .S(n9910), .Z(
        P2_U3513) );
  MUX2_X1 U9931 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8510), .S(n9910), .Z(
        P2_U3512) );
  MUX2_X1 U9932 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8511), .S(n9910), .Z(
        P2_U3511) );
  MUX2_X1 U9933 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8512), .S(n9910), .Z(
        P2_U3510) );
  MUX2_X1 U9934 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8513), .S(n9910), .Z(
        P2_U3509) );
  MUX2_X1 U9935 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8514), .S(n9910), .Z(
        P2_U3508) );
  MUX2_X1 U9936 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8515), .S(n9910), .Z(
        P2_U3507) );
  MUX2_X1 U9937 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8516), .S(n9910), .Z(
        P2_U3505) );
  MUX2_X1 U9938 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8517), .S(n9910), .Z(
        P2_U3502) );
  MUX2_X1 U9939 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8518), .S(n9910), .Z(
        P2_U3499) );
  MUX2_X1 U9940 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8519), .S(n9910), .Z(
        P2_U3496) );
  MUX2_X1 U9941 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8520), .S(n9910), .Z(
        P2_U3493) );
  MUX2_X1 U9942 ( .A(n8521), .B(P2_REG0_REG_13__SCAN_IN), .S(n9908), .Z(
        P2_U3490) );
  INV_X1 U9943 ( .A(n8676), .ZN(n9418) );
  NOR4_X1 U9944 ( .A1(n8523), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n8522), .ZN(n8524) );
  AOI21_X1 U9945 ( .B1(n8525), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8524), .ZN(
        n8526) );
  OAI21_X1 U9946 ( .B1(n9418), .B2(n7800), .A(n8526), .ZN(P2_U3327) );
  MUX2_X1 U9947 ( .A(n8527), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U9948 ( .A(n8530), .B(n8529), .ZN(n8531) );
  XNOR2_X1 U9949 ( .A(n8528), .B(n8531), .ZN(n8536) );
  NOR2_X1 U9950 ( .A1(n4275), .A2(n9133), .ZN(n8534) );
  AOI22_X1 U9951 ( .A1(n8666), .A2(n9142), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8532) );
  OAI21_X1 U9952 ( .B1(n9136), .B2(n8664), .A(n8532), .ZN(n8533) );
  AOI211_X1 U9953 ( .C1(n9337), .C2(n8671), .A(n8534), .B(n8533), .ZN(n8535)
         );
  OAI21_X1 U9954 ( .B1(n8536), .B2(n8645), .A(n8535), .ZN(P1_U3212) );
  INV_X1 U9955 ( .A(n7231), .ZN(n8542) );
  AOI21_X1 U9956 ( .B1(n8538), .B2(n7231), .A(n8537), .ZN(n8539) );
  NOR2_X1 U9957 ( .A1(n8539), .A2(n8645), .ZN(n8540) );
  OAI21_X1 U9958 ( .B1(n8542), .B2(n8541), .A(n8540), .ZN(n8549) );
  OAI21_X1 U9959 ( .B1(n8664), .B2(n8544), .A(n8543), .ZN(n8547) );
  NOR2_X1 U9960 ( .A1(n4275), .A2(n8545), .ZN(n8546) );
  AOI211_X1 U9961 ( .C1(n8666), .C2(n8963), .A(n8547), .B(n8546), .ZN(n8548)
         );
  OAI211_X1 U9962 ( .C1(n9518), .C2(n8656), .A(n8549), .B(n8548), .ZN(P1_U3213) );
  INV_X1 U9964 ( .A(n8551), .ZN(n8553) );
  NAND2_X1 U9965 ( .A1(n8553), .A2(n8552), .ZN(n8557) );
  NAND2_X1 U9966 ( .A1(n8557), .A2(n8556), .ZN(n8608) );
  NAND2_X1 U9967 ( .A1(n8551), .A2(n8554), .ZN(n8607) );
  INV_X1 U9968 ( .A(n8607), .ZN(n8555) );
  NOR2_X1 U9969 ( .A1(n8608), .A2(n8555), .ZN(n8559) );
  AOI21_X1 U9970 ( .B1(n8557), .B2(n8607), .A(n8556), .ZN(n8558) );
  OAI21_X1 U9971 ( .B1(n8559), .B2(n8558), .A(n8657), .ZN(n8563) );
  AOI22_X1 U9972 ( .A1(n8653), .A2(n9166), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8560) );
  OAI21_X1 U9973 ( .B1(n9230), .B2(n8650), .A(n8560), .ZN(n8561) );
  AOI21_X1 U9974 ( .B1(n9198), .B2(n8576), .A(n8561), .ZN(n8562) );
  OAI211_X1 U9975 ( .C1(n9200), .C2(n8656), .A(n8563), .B(n8562), .ZN(P1_U3214) );
  XOR2_X1 U9976 ( .A(n8566), .B(n8565), .Z(n8567) );
  XNOR2_X1 U9977 ( .A(n8564), .B(n8567), .ZN(n8572) );
  NAND2_X1 U9978 ( .A1(n8666), .A2(n8960), .ZN(n8568) );
  NAND2_X1 U9979 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9098) );
  OAI211_X1 U9980 ( .C1(n9256), .C2(n8664), .A(n8568), .B(n9098), .ZN(n8570)
         );
  NOR2_X1 U9981 ( .A1(n9264), .A2(n8656), .ZN(n8569) );
  AOI211_X1 U9982 ( .C1(n9260), .C2(n8576), .A(n8570), .B(n8569), .ZN(n8571)
         );
  OAI21_X1 U9983 ( .B1(n8572), .B2(n8645), .A(n8571), .ZN(P1_U3217) );
  XOR2_X1 U9984 ( .A(n8574), .B(n8573), .Z(n8581) );
  AOI22_X1 U9985 ( .A1(n8958), .A2(n8666), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8578) );
  NAND2_X1 U9986 ( .A1(n8576), .A2(n9232), .ZN(n8577) );
  OAI211_X1 U9987 ( .C1(n9230), .C2(n8664), .A(n8578), .B(n8577), .ZN(n8579)
         );
  AOI21_X1 U9988 ( .B1(n9368), .B2(n8671), .A(n8579), .ZN(n8580) );
  OAI21_X1 U9989 ( .B1(n8581), .B2(n8645), .A(n8580), .ZN(P1_U3221) );
  NAND2_X1 U9990 ( .A1(n9176), .A2(n9689), .ZN(n9348) );
  XNOR2_X1 U9991 ( .A(n8582), .B(n8583), .ZN(n8584) );
  NAND2_X1 U9992 ( .A1(n8584), .A2(n8657), .ZN(n8589) );
  OAI22_X1 U9993 ( .A1(n8664), .A2(n9161), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8585), .ZN(n8587) );
  NOR2_X1 U9994 ( .A1(n4275), .A2(n9169), .ZN(n8586) );
  AOI211_X1 U9995 ( .C1(n8666), .C2(n9166), .A(n8587), .B(n8586), .ZN(n8588)
         );
  OAI211_X1 U9996 ( .C1(n8590), .C2(n9348), .A(n8589), .B(n8588), .ZN(P1_U3223) );
  INV_X1 U9997 ( .A(n8591), .ZN(n8592) );
  AOI21_X1 U9998 ( .B1(n8594), .B2(n8593), .A(n8592), .ZN(n8599) );
  NAND2_X1 U9999 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9055) );
  OAI21_X1 U10000 ( .B1(n8664), .B2(n9276), .A(n9055), .ZN(n8595) );
  AOI21_X1 U10001 ( .B1(n8666), .B2(n9303), .A(n8595), .ZN(n8596) );
  OAI21_X1 U10002 ( .B1(n4275), .B2(n9307), .A(n8596), .ZN(n8597) );
  AOI21_X1 U10003 ( .B1(n9313), .B2(n8671), .A(n8597), .ZN(n8598) );
  OAI21_X1 U10004 ( .B1(n8599), .B2(n8645), .A(n8598), .ZN(P1_U3224) );
  XOR2_X1 U10005 ( .A(n8600), .B(n8601), .Z(n8606) );
  NAND2_X1 U10006 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9068) );
  OAI21_X1 U10007 ( .B1(n8650), .B2(n9290), .A(n9068), .ZN(n8602) );
  AOI21_X1 U10008 ( .B1(n8653), .B2(n8960), .A(n8602), .ZN(n8603) );
  OAI21_X1 U10009 ( .B1(n4275), .B2(n9296), .A(n8603), .ZN(n8604) );
  AOI21_X1 U10010 ( .B1(n9390), .B2(n8671), .A(n8604), .ZN(n8605) );
  OAI21_X1 U10011 ( .B1(n8606), .B2(n8645), .A(n8605), .ZN(P1_U3226) );
  NAND2_X1 U10012 ( .A1(n8608), .A2(n8607), .ZN(n8612) );
  XNOR2_X1 U10013 ( .A(n8610), .B(n8609), .ZN(n8611) );
  XNOR2_X1 U10014 ( .A(n8612), .B(n8611), .ZN(n8618) );
  INV_X1 U10015 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8613) );
  OAI22_X1 U10016 ( .A1(n8664), .A2(n8957), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8613), .ZN(n8614) );
  AOI21_X1 U10017 ( .B1(n9183), .B2(n8666), .A(n8614), .ZN(n8615) );
  OAI21_X1 U10018 ( .B1(n4275), .B2(n9190), .A(n8615), .ZN(n8616) );
  AOI21_X1 U10019 ( .B1(n9352), .B2(n8671), .A(n8616), .ZN(n8617) );
  OAI21_X1 U10020 ( .B1(n8618), .B2(n8645), .A(n8617), .ZN(P1_U3227) );
  INV_X1 U10021 ( .A(n8619), .ZN(n8623) );
  OAI21_X1 U10022 ( .B1(n8621), .B2(n8623), .A(n8620), .ZN(n8622) );
  OAI21_X1 U10023 ( .B1(n8624), .B2(n8623), .A(n8622), .ZN(n8625) );
  NAND2_X1 U10024 ( .A1(n8625), .A2(n8657), .ZN(n8630) );
  NOR2_X1 U10025 ( .A1(n4275), .A2(n9245), .ZN(n8628) );
  OAI22_X1 U10026 ( .A1(n9242), .A2(n8664), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8626), .ZN(n8627) );
  AOI211_X1 U10027 ( .C1(n8666), .C2(n8959), .A(n8628), .B(n8627), .ZN(n8629)
         );
  OAI211_X1 U10028 ( .C1(n9249), .C2(n8656), .A(n8630), .B(n8629), .ZN(
        P1_U3231) );
  NAND2_X1 U10029 ( .A1(n8632), .A2(n8631), .ZN(n8633) );
  XOR2_X1 U10030 ( .A(n8634), .B(n8633), .Z(n8641) );
  OAI22_X1 U10031 ( .A1(n9242), .A2(n8650), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8635), .ZN(n8636) );
  AOI21_X1 U10032 ( .B1(n9183), .B2(n8653), .A(n8636), .ZN(n8637) );
  OAI21_X1 U10033 ( .B1(n4275), .B2(n8638), .A(n8637), .ZN(n8639) );
  AOI21_X1 U10034 ( .B1(n9363), .B2(n8671), .A(n8639), .ZN(n8640) );
  OAI21_X1 U10035 ( .B1(n8641), .B2(n8645), .A(n8640), .ZN(P1_U3233) );
  INV_X1 U10036 ( .A(n8644), .ZN(n8649) );
  AOI21_X1 U10037 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(n8646) );
  NOR2_X1 U10038 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  OAI21_X1 U10039 ( .B1(n8649), .B2(n8648), .A(n8647), .ZN(n8655) );
  NAND2_X1 U10040 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9083) );
  OAI21_X1 U10041 ( .B1(n8650), .B2(n9276), .A(n9083), .ZN(n8652) );
  NOR2_X1 U10042 ( .A1(n4275), .A2(n9268), .ZN(n8651) );
  AOI211_X1 U10043 ( .C1(n8653), .C2(n8959), .A(n8652), .B(n8651), .ZN(n8654)
         );
  OAI211_X1 U10044 ( .C1(n9278), .C2(n8656), .A(n8655), .B(n8654), .ZN(
        P1_U3236) );
  INV_X1 U10045 ( .A(n8662), .ZN(n8659) );
  OAI21_X1 U10046 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n8675) );
  AOI21_X1 U10047 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8674) );
  OAI21_X1 U10048 ( .B1(n8664), .B2(n9290), .A(n8663), .ZN(n8665) );
  AOI21_X1 U10049 ( .B1(n8666), .B2(n8962), .A(n8665), .ZN(n8667) );
  OAI21_X1 U10050 ( .B1(n4275), .B2(n8668), .A(n8667), .ZN(n8670) );
  AOI21_X1 U10051 ( .B1(n8672), .B2(n8671), .A(n8670), .ZN(n8673) );
  OAI21_X1 U10052 ( .B1(n8675), .B2(n8674), .A(n8673), .ZN(P1_U3239) );
  INV_X1 U10053 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U10054 ( .A1(n8678), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8681) );
  INV_X1 U10055 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9101) );
  OR2_X1 U10056 ( .A1(n4280), .A2(n9101), .ZN(n8680) );
  OAI211_X1 U10057 ( .C1(n8683), .C2(n8682), .A(n8681), .B(n8680), .ZN(n9102)
         );
  INV_X1 U10058 ( .A(n9102), .ZN(n8684) );
  NAND2_X1 U10059 ( .A1(n8685), .A2(n6383), .ZN(n8689) );
  OR2_X1 U10060 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  INV_X1 U10061 ( .A(n8956), .ZN(n8690) );
  OR2_X1 U10062 ( .A1(n9108), .A2(n8690), .ZN(n8749) );
  NAND2_X1 U10063 ( .A1(n8939), .A2(n8749), .ZN(n8878) );
  NOR2_X1 U10064 ( .A1(n9322), .A2(n8956), .ZN(n8913) );
  INV_X1 U10065 ( .A(n8913), .ZN(n8747) );
  NAND2_X1 U10066 ( .A1(n8692), .A2(n8691), .ZN(n8826) );
  INV_X1 U10067 ( .A(n8817), .ZN(n8879) );
  AND2_X1 U10068 ( .A1(n8830), .A2(n8879), .ZN(n8693) );
  NOR2_X1 U10069 ( .A1(n8826), .A2(n8693), .ZN(n8831) );
  NAND2_X1 U10070 ( .A1(n8831), .A2(n8818), .ZN(n8721) );
  AND2_X1 U10071 ( .A1(n8809), .A2(n8810), .ZN(n8694) );
  NAND2_X1 U10072 ( .A1(n8751), .A2(n8694), .ZN(n8722) );
  NAND2_X1 U10073 ( .A1(n8696), .A2(n8695), .ZN(n8787) );
  NAND2_X1 U10074 ( .A1(n8787), .A2(n8788), .ZN(n8795) );
  INV_X1 U10075 ( .A(n8795), .ZN(n8727) );
  AND2_X1 U10076 ( .A1(n8773), .A2(n4476), .ZN(n8779) );
  INV_X1 U10077 ( .A(n8779), .ZN(n8697) );
  AND2_X1 U10078 ( .A1(n8697), .A2(n8782), .ZN(n8698) );
  NOR2_X1 U10079 ( .A1(n8699), .A2(n8698), .ZN(n8723) );
  NAND4_X1 U10080 ( .A1(n8727), .A2(n8723), .A3(n8776), .A4(n8766), .ZN(n8700)
         );
  NOR4_X1 U10081 ( .A1(n8721), .A2(n4474), .A3(n8722), .A4(n8700), .ZN(n8923)
         );
  AND2_X1 U10082 ( .A1(n8702), .A2(n8701), .ZN(n8885) );
  INV_X1 U10083 ( .A(n8885), .ZN(n8703) );
  OAI211_X1 U10084 ( .C1(n8704), .C2(n9634), .A(n8917), .B(n8703), .ZN(n8705)
         );
  NAND2_X1 U10085 ( .A1(n8705), .A2(n5886), .ZN(n8707) );
  OAI21_X1 U10086 ( .B1(n5925), .B2(n8707), .A(n8706), .ZN(n8709) );
  AOI22_X1 U10087 ( .A1(n8709), .A2(n8708), .B1(n9683), .B2(n8970), .ZN(n8720)
         );
  NAND2_X1 U10088 ( .A1(n8714), .A2(n8710), .ZN(n8759) );
  INV_X1 U10089 ( .A(n8759), .ZN(n8712) );
  AND2_X1 U10090 ( .A1(n8712), .A2(n8711), .ZN(n8761) );
  INV_X1 U10091 ( .A(n8761), .ZN(n8719) );
  NAND2_X1 U10092 ( .A1(n8714), .A2(n8713), .ZN(n8716) );
  AND2_X1 U10093 ( .A1(n8716), .A2(n8715), .ZN(n8763) );
  OR2_X1 U10094 ( .A1(n8759), .A2(n8754), .ZN(n8717) );
  AND2_X1 U10095 ( .A1(n8763), .A2(n8717), .ZN(n8758) );
  OAI211_X1 U10096 ( .C1(n8720), .C2(n8719), .A(n8758), .B(n8718), .ZN(n8738)
         );
  INV_X1 U10097 ( .A(n8721), .ZN(n8731) );
  INV_X1 U10098 ( .A(n8722), .ZN(n8730) );
  AND2_X1 U10099 ( .A1(n8782), .A2(n8777), .ZN(n8725) );
  INV_X1 U10100 ( .A(n8723), .ZN(n8724) );
  OAI211_X1 U10101 ( .C1(n8725), .C2(n8724), .A(n8786), .B(n8797), .ZN(n8726)
         );
  AOI21_X1 U10102 ( .B1(n8727), .B2(n8726), .A(n8801), .ZN(n8728) );
  OAI211_X1 U10103 ( .C1(n8728), .C2(n4474), .A(n8811), .B(n8806), .ZN(n8729)
         );
  NAND3_X1 U10104 ( .A1(n8731), .A2(n8730), .A3(n8729), .ZN(n8737) );
  NAND2_X1 U10105 ( .A1(n8844), .A2(n8836), .ZN(n8828) );
  INV_X1 U10106 ( .A(n8828), .ZN(n8736) );
  AND2_X1 U10107 ( .A1(n8818), .A2(n8751), .ZN(n8820) );
  INV_X1 U10108 ( .A(n8820), .ZN(n8733) );
  INV_X1 U10109 ( .A(n8815), .ZN(n8732) );
  NOR2_X1 U10110 ( .A1(n8880), .A2(n8732), .ZN(n8823) );
  OAI211_X1 U10111 ( .C1(n8753), .C2(n8733), .A(n8823), .B(n8830), .ZN(n8734)
         );
  NAND2_X1 U10112 ( .A1(n8831), .A2(n8734), .ZN(n8735) );
  NAND3_X1 U10113 ( .A1(n8737), .A2(n8736), .A3(n8735), .ZN(n8920) );
  AOI21_X1 U10114 ( .B1(n8923), .B2(n8738), .A(n8920), .ZN(n8739) );
  NAND2_X1 U10115 ( .A1(n8845), .A2(n8834), .ZN(n8840) );
  NAND2_X1 U10116 ( .A1(n9192), .A2(n9166), .ZN(n8919) );
  OAI21_X1 U10117 ( .B1(n8739), .B2(n8840), .A(n8919), .ZN(n8742) );
  NAND2_X1 U10118 ( .A1(n9153), .A2(n9142), .ZN(n8855) );
  INV_X1 U10119 ( .A(n8855), .ZN(n8740) );
  NOR3_X1 U10120 ( .A1(n8743), .A2(n8842), .A3(n8740), .ZN(n8929) );
  INV_X1 U10121 ( .A(n8929), .ZN(n8741) );
  AOI21_X1 U10122 ( .B1(n8848), .B2(n8742), .A(n8741), .ZN(n8745) );
  OAI211_X1 U10123 ( .C1(n8743), .C2(n8856), .A(n8859), .B(n8865), .ZN(n8927)
         );
  NAND2_X1 U10124 ( .A1(n8870), .A2(n8864), .ZN(n8932) );
  INV_X1 U10125 ( .A(n8932), .ZN(n8744) );
  OAI21_X1 U10126 ( .B1(n8745), .B2(n8927), .A(n8744), .ZN(n8746) );
  AND3_X1 U10127 ( .A1(n8747), .A2(n8930), .A3(n8746), .ZN(n8748) );
  OAI21_X1 U10128 ( .B1(n8878), .B2(n8748), .A(n8877), .ZN(n8947) );
  NAND2_X1 U10129 ( .A1(n8749), .A2(n9102), .ZN(n8750) );
  NAND2_X1 U10130 ( .A1(n8750), .A2(n9105), .ZN(n8936) );
  INV_X1 U10131 ( .A(n8869), .ZN(n8874) );
  AND2_X1 U10132 ( .A1(n8751), .A2(n8809), .ZN(n8752) );
  MUX2_X1 U10133 ( .A(n8753), .B(n8752), .S(n8874), .Z(n8814) );
  NAND2_X1 U10134 ( .A1(n8755), .A2(n8754), .ZN(n8756) );
  MUX2_X1 U10135 ( .A(n8757), .B(n8756), .S(n8869), .Z(n8762) );
  OAI21_X1 U10136 ( .B1(n8762), .B2(n8759), .A(n8758), .ZN(n8760) );
  AOI21_X1 U10137 ( .B1(n8760), .B2(n8766), .A(n8765), .ZN(n8770) );
  NAND2_X1 U10138 ( .A1(n8762), .A2(n8761), .ZN(n8768) );
  INV_X1 U10139 ( .A(n8763), .ZN(n8764) );
  NOR2_X1 U10140 ( .A1(n8765), .A2(n8764), .ZN(n8767) );
  AOI21_X1 U10141 ( .B1(n8768), .B2(n8767), .A(n4480), .ZN(n8769) );
  MUX2_X1 U10142 ( .A(n8770), .B(n8769), .S(n8869), .Z(n8778) );
  INV_X1 U10143 ( .A(n9594), .ZN(n8771) );
  OAI211_X1 U10144 ( .C1(n8778), .C2(n8771), .A(n4476), .B(n8776), .ZN(n8772)
         );
  NAND3_X1 U10145 ( .A1(n8772), .A2(n8782), .A3(n8882), .ZN(n8775) );
  NAND3_X1 U10146 ( .A1(n8775), .A2(n8774), .A3(n8773), .ZN(n8785) );
  OAI21_X1 U10147 ( .B1(n8778), .B2(n4481), .A(n8777), .ZN(n8780) );
  NAND2_X1 U10148 ( .A1(n8780), .A2(n8779), .ZN(n8783) );
  NAND3_X1 U10149 ( .A1(n8783), .A2(n8782), .A3(n8781), .ZN(n8784) );
  MUX2_X1 U10150 ( .A(n8785), .B(n8784), .S(n8874), .Z(n8793) );
  OR2_X1 U10151 ( .A1(n8801), .A2(n8874), .ZN(n8794) );
  NAND2_X1 U10152 ( .A1(n8786), .A2(n8797), .ZN(n8791) );
  NAND2_X1 U10153 ( .A1(n8787), .A2(n8874), .ZN(n8798) );
  NAND2_X1 U10154 ( .A1(n8789), .A2(n8788), .ZN(n8790) );
  OAI22_X1 U10155 ( .A1(n8794), .A2(n8791), .B1(n8798), .B2(n8790), .ZN(n8792)
         );
  OAI21_X1 U10156 ( .B1(n8793), .B2(n6587), .A(n8792), .ZN(n8804) );
  INV_X1 U10157 ( .A(n8794), .ZN(n8796) );
  NAND2_X1 U10158 ( .A1(n8796), .A2(n8795), .ZN(n8803) );
  INV_X1 U10159 ( .A(n8797), .ZN(n8800) );
  INV_X1 U10160 ( .A(n8798), .ZN(n8799) );
  OAI21_X1 U10161 ( .B1(n8801), .B2(n8800), .A(n8799), .ZN(n8802) );
  NAND4_X1 U10162 ( .A1(n8804), .A2(n8903), .A3(n8803), .A4(n8802), .ZN(n8808)
         );
  INV_X1 U10163 ( .A(n8906), .ZN(n9314) );
  MUX2_X1 U10164 ( .A(n8806), .B(n8805), .S(n8874), .Z(n8807) );
  NAND3_X1 U10165 ( .A1(n8808), .A2(n9314), .A3(n8807), .ZN(n8813) );
  NAND2_X1 U10166 ( .A1(n9271), .A2(n8809), .ZN(n8907) );
  MUX2_X1 U10167 ( .A(n8811), .B(n8810), .S(n8869), .Z(n8812) );
  NAND3_X1 U10168 ( .A1(n8821), .A2(n8816), .A3(n8815), .ZN(n8819) );
  NAND3_X1 U10169 ( .A1(n8819), .A2(n8818), .A3(n8817), .ZN(n8825) );
  NAND2_X1 U10170 ( .A1(n8821), .A2(n8820), .ZN(n8822) );
  NAND2_X1 U10171 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  AND2_X1 U10172 ( .A1(n8830), .A2(n4466), .ZN(n8827) );
  AOI21_X1 U10173 ( .B1(n8833), .B2(n8827), .A(n8826), .ZN(n8829) );
  NOR2_X1 U10174 ( .A1(n8829), .A2(n8828), .ZN(n8839) );
  INV_X1 U10175 ( .A(n8830), .ZN(n8832) );
  OAI21_X1 U10176 ( .B1(n8833), .B2(n8832), .A(n8831), .ZN(n8837) );
  INV_X1 U10177 ( .A(n8834), .ZN(n8835) );
  AOI21_X1 U10178 ( .B1(n8837), .B2(n8836), .A(n8835), .ZN(n8838) );
  NAND2_X1 U10179 ( .A1(n8847), .A2(n8919), .ZN(n8843) );
  NAND2_X1 U10180 ( .A1(n8840), .A2(n8919), .ZN(n8841) );
  AND2_X1 U10181 ( .A1(n8848), .A2(n8841), .ZN(n8924) );
  AOI21_X1 U10182 ( .B1(n8843), .B2(n8924), .A(n8842), .ZN(n8853) );
  NAND2_X1 U10183 ( .A1(n8919), .A2(n8844), .ZN(n8846) );
  OAI21_X1 U10184 ( .B1(n8847), .B2(n8846), .A(n8845), .ZN(n8851) );
  INV_X1 U10185 ( .A(n8848), .ZN(n8849) );
  AOI21_X1 U10186 ( .B1(n8851), .B2(n8850), .A(n8849), .ZN(n8852) );
  NAND2_X1 U10187 ( .A1(n8854), .A2(n9155), .ZN(n8858) );
  INV_X1 U10188 ( .A(n9139), .ZN(n9130) );
  MUX2_X1 U10189 ( .A(n8856), .B(n8855), .S(n8869), .Z(n8857) );
  INV_X1 U10190 ( .A(n9117), .ZN(n8862) );
  MUX2_X1 U10191 ( .A(n8860), .B(n8859), .S(n8869), .Z(n8861) );
  NAND3_X1 U10192 ( .A1(n8863), .A2(n8862), .A3(n8861), .ZN(n8867) );
  MUX2_X1 U10193 ( .A(n8865), .B(n8864), .S(n8869), .Z(n8866) );
  NAND2_X1 U10194 ( .A1(n8936), .A2(n8868), .ZN(n8872) );
  OR2_X1 U10195 ( .A1(n8870), .A2(n8869), .ZN(n8871) );
  NAND2_X1 U10196 ( .A1(n8872), .A2(n8871), .ZN(n8876) );
  NAND2_X1 U10197 ( .A1(n8956), .A2(n9102), .ZN(n8873) );
  AND2_X1 U10198 ( .A1(n9108), .A2(n8873), .ZN(n8940) );
  INV_X1 U10199 ( .A(n8940), .ZN(n8931) );
  INV_X1 U10200 ( .A(n8936), .ZN(n8875) );
  AOI22_X1 U10201 ( .A1(n8876), .A2(n8931), .B1(n8875), .B2(n8874), .ZN(n8945)
         );
  NAND3_X1 U10202 ( .A1(n8877), .A2(n8917), .A3(n5212), .ZN(n8944) );
  INV_X1 U10203 ( .A(n8878), .ZN(n8916) );
  INV_X1 U10204 ( .A(n9167), .ZN(n8911) );
  INV_X1 U10205 ( .A(n9213), .ZN(n9211) );
  INV_X1 U10206 ( .A(n9225), .ZN(n9227) );
  NOR2_X1 U10207 ( .A1(n8880), .A2(n8879), .ZN(n9239) );
  INV_X1 U10208 ( .A(n8881), .ZN(n8898) );
  INV_X1 U10209 ( .A(n8882), .ZN(n8884) );
  OR2_X1 U10210 ( .A1(n8884), .A2(n8883), .ZN(n9605) );
  NOR2_X1 U10211 ( .A1(n8886), .A2(n8885), .ZN(n9648) );
  NAND3_X1 U10212 ( .A1(n9648), .A2(n8888), .A3(n8887), .ZN(n8892) );
  NOR4_X1 U10213 ( .A1(n8892), .A2(n8891), .A3(n8890), .A4(n8889), .ZN(n8896)
         );
  INV_X1 U10214 ( .A(n9622), .ZN(n8895) );
  NAND4_X1 U10215 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8893), .ZN(n8897)
         );
  NOR4_X1 U10216 ( .A1(n8899), .A2(n8898), .A3(n9605), .A4(n8897), .ZN(n8901)
         );
  NAND4_X1 U10217 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), .ZN(n8905)
         );
  NOR4_X1 U10218 ( .A1(n8907), .A2(n8906), .A3(n8905), .A4(n8904), .ZN(n8908)
         );
  NAND4_X1 U10219 ( .A1(n9239), .A2(n4465), .A3(n9273), .A4(n8908), .ZN(n8909)
         );
  NOR4_X1 U10220 ( .A1(n9203), .A2(n9211), .A3(n9227), .A4(n8909), .ZN(n8910)
         );
  NAND3_X1 U10221 ( .A1(n8877), .A2(n8916), .A3(n8915), .ZN(n8918) );
  INV_X1 U10222 ( .A(n8919), .ZN(n8921) );
  AOI211_X1 U10223 ( .C1(n8923), .C2(n8922), .A(n8921), .B(n8920), .ZN(n8926)
         );
  INV_X1 U10224 ( .A(n8924), .ZN(n8925) );
  OR2_X1 U10225 ( .A1(n8926), .A2(n8925), .ZN(n8928) );
  AOI21_X1 U10226 ( .B1(n8929), .B2(n8928), .A(n8927), .ZN(n8933) );
  OAI211_X1 U10227 ( .C1(n8933), .C2(n8932), .A(n8931), .B(n8930), .ZN(n8935)
         );
  AOI211_X1 U10228 ( .C1(n8936), .C2(n8935), .A(n8934), .B(n8938), .ZN(n8937)
         );
  AOI211_X1 U10229 ( .C1(n8940), .C2(n8939), .A(n5219), .B(n8938), .ZN(n8942)
         );
  AOI21_X1 U10230 ( .B1(n8945), .B2(n8942), .A(n8941), .ZN(n8943) );
  NAND3_X1 U10231 ( .A1(n8950), .A2(n8949), .A3(n9557), .ZN(n8951) );
  OAI211_X1 U10232 ( .C1(n8952), .C2(n8954), .A(n8951), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8953) );
  OAI21_X1 U10233 ( .B1(n8955), .B2(n8954), .A(n8953), .ZN(P1_U3240) );
  MUX2_X1 U10234 ( .A(n9102), .B(P1_DATAO_REG_31__SCAN_IN), .S(n8972), .Z(
        P1_U3586) );
  MUX2_X1 U10235 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8956), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10236 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n7172), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10237 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n4490), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10238 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9142), .S(P1_U4006), .Z(
        P1_U3581) );
  INV_X1 U10239 ( .A(n8957), .ZN(n9184) );
  MUX2_X1 U10240 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9184), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10241 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9166), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10242 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9183), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10243 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9207), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10244 ( .A(n8958), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8972), .Z(
        P1_U3575) );
  MUX2_X1 U10245 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n8959), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10246 ( .A(n8960), .B(P1_DATAO_REG_18__SCAN_IN), .S(n8972), .Z(
        P1_U3573) );
  MUX2_X1 U10247 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9304), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10248 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8961), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10249 ( .A(n9303), .B(P1_DATAO_REG_15__SCAN_IN), .S(n8972), .Z(
        P1_U3570) );
  MUX2_X1 U10250 ( .A(n8962), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8972), .Z(
        P1_U3569) );
  MUX2_X1 U10251 ( .A(n8963), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8972), .Z(
        P1_U3568) );
  MUX2_X1 U10252 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8964), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10253 ( .A(n8965), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8972), .Z(
        P1_U3566) );
  MUX2_X1 U10254 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9597), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10255 ( .A(n8966), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8972), .Z(
        P1_U3564) );
  MUX2_X1 U10256 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9613), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10257 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8967), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10258 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9615), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10259 ( .A(n8968), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8972), .Z(
        P1_U3560) );
  MUX2_X1 U10260 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8969), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10261 ( .A(n8970), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8972), .Z(
        P1_U3558) );
  MUX2_X1 U10262 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8971), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10263 ( .A(n5380), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8972), .Z(
        P1_U3556) );
  NAND2_X1 U10264 ( .A1(n9579), .A2(n8973), .ZN(n8974) );
  OAI21_X1 U10265 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n8975), .A(n8974), .ZN(
        n8976) );
  AOI21_X1 U10266 ( .B1(n9564), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n8976), .ZN(
        n8988) );
  NAND2_X1 U10267 ( .A1(n9558), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8990) );
  INV_X1 U10268 ( .A(n8990), .ZN(n8980) );
  MUX2_X1 U10269 ( .A(n9645), .B(P1_REG2_REG_1__SCAN_IN), .S(n8977), .Z(n8979)
         );
  INV_X1 U10270 ( .A(n9005), .ZN(n8978) );
  OAI211_X1 U10271 ( .C1(n8980), .C2(n8979), .A(n9588), .B(n8978), .ZN(n8987)
         );
  INV_X1 U10272 ( .A(n8981), .ZN(n8985) );
  NOR2_X1 U10273 ( .A1(n8993), .A2(n9730), .ZN(n8984) );
  INV_X1 U10274 ( .A(n8982), .ZN(n8983) );
  OAI211_X1 U10275 ( .C1(n8985), .C2(n8984), .A(n9587), .B(n8983), .ZN(n8986)
         );
  NAND3_X1 U10276 ( .A1(n8988), .A2(n8987), .A3(n8986), .ZN(P1_U3242) );
  MUX2_X1 U10277 ( .A(n8990), .B(n8989), .S(n8991), .Z(n8996) );
  NOR2_X1 U10278 ( .A1(n8991), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8992) );
  OR2_X1 U10279 ( .A1(n4283), .A2(n8992), .ZN(n9555) );
  NAND2_X1 U10280 ( .A1(n9555), .A2(n8993), .ZN(n8994) );
  OAI211_X1 U10281 ( .C1(n8996), .C2(n4283), .A(P1_U4006), .B(n8994), .ZN(
        n9028) );
  OAI22_X1 U10282 ( .A1(n9422), .A2(n9006), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8997), .ZN(n8998) );
  AOI21_X1 U10283 ( .B1(n9564), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n8998), .ZN(
        n9013) );
  MUX2_X1 U10284 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n8999), .S(n9006), .Z(n9002)
         );
  INV_X1 U10285 ( .A(n9000), .ZN(n9001) );
  NAND2_X1 U10286 ( .A1(n9002), .A2(n9001), .ZN(n9004) );
  OAI211_X1 U10287 ( .C1(n9005), .C2(n9004), .A(n9588), .B(n9003), .ZN(n9012)
         );
  MUX2_X1 U10288 ( .A(n9732), .B(P1_REG1_REG_2__SCAN_IN), .S(n9006), .Z(n9010)
         );
  INV_X1 U10289 ( .A(n9007), .ZN(n9009) );
  OAI211_X1 U10290 ( .C1(n9010), .C2(n9009), .A(n9587), .B(n9008), .ZN(n9011)
         );
  NAND4_X1 U10291 ( .A1(n9028), .A2(n9013), .A3(n9012), .A4(n9011), .ZN(
        P1_U3243) );
  OAI21_X1 U10292 ( .B1(n9016), .B2(n9015), .A(n9014), .ZN(n9019) );
  INV_X1 U10293 ( .A(n9017), .ZN(n9018) );
  AOI22_X1 U10294 ( .A1(n9019), .A2(n9587), .B1(n9018), .B2(n9579), .ZN(n9027)
         );
  AOI21_X1 U10295 ( .B1(n9022), .B2(n9021), .A(n9020), .ZN(n9024) );
  OAI21_X1 U10296 ( .B1(n9571), .B2(n9024), .A(n9023), .ZN(n9025) );
  AOI21_X1 U10297 ( .B1(n9564), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9025), .ZN(
        n9026) );
  NAND3_X1 U10298 ( .A1(n9028), .A2(n9027), .A3(n9026), .ZN(P1_U3245) );
  OAI21_X1 U10299 ( .B1(n9031), .B2(n9030), .A(n9029), .ZN(n9036) );
  AOI211_X1 U10300 ( .C1(n9034), .C2(n9033), .A(n9032), .B(n9571), .ZN(n9035)
         );
  AOI21_X1 U10301 ( .B1(n9587), .B2(n9036), .A(n9035), .ZN(n9041) );
  NAND2_X1 U10302 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n9040) );
  NAND2_X1 U10303 ( .A1(n9579), .A2(n9037), .ZN(n9039) );
  NAND2_X1 U10304 ( .A1(n9564), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n9038) );
  NAND4_X1 U10305 ( .A1(n9041), .A2(n9040), .A3(n9039), .A4(n9038), .ZN(
        P1_U3251) );
  NOR2_X1 U10306 ( .A1(n9048), .A2(n9042), .ZN(n9044) );
  NAND2_X1 U10307 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9064), .ZN(n9045) );
  OAI21_X1 U10308 ( .B1(n9064), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9045), .ZN(
        n9046) );
  AOI211_X1 U10309 ( .C1(n4362), .C2(n9046), .A(n9060), .B(n9571), .ZN(n9059)
         );
  NOR2_X1 U10310 ( .A1(n9048), .A2(n9047), .ZN(n9050) );
  INV_X1 U10311 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9509) );
  NOR2_X1 U10312 ( .A1(n9064), .A2(n9509), .ZN(n9051) );
  AOI21_X1 U10313 ( .B1(n9064), .B2(n9509), .A(n9051), .ZN(n9052) );
  NOR2_X1 U10314 ( .A1(n9053), .A2(n9052), .ZN(n9063) );
  AOI211_X1 U10315 ( .C1(n9053), .C2(n9052), .A(n9063), .B(n9427), .ZN(n9058)
         );
  NAND2_X1 U10316 ( .A1(n9564), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9054) );
  OAI211_X1 U10317 ( .C1(n9422), .C2(n9056), .A(n9055), .B(n9054), .ZN(n9057)
         );
  OR3_X1 U10318 ( .A1(n9059), .A2(n9058), .A3(n9057), .ZN(P1_U3257) );
  AOI21_X1 U10319 ( .B1(n9064), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9060), .ZN(
        n9062) );
  XNOR2_X1 U10320 ( .A(n9077), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9061) );
  NOR2_X1 U10321 ( .A1(n9062), .A2(n9061), .ZN(n9076) );
  AOI211_X1 U10322 ( .C1(n9062), .C2(n9061), .A(n9076), .B(n9571), .ZN(n9072)
         );
  AOI21_X1 U10323 ( .B1(n9064), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9063), .ZN(
        n9066) );
  XNOR2_X1 U10324 ( .A(n9077), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9065) );
  NOR2_X1 U10325 ( .A1(n9066), .A2(n9065), .ZN(n9073) );
  AOI211_X1 U10326 ( .C1(n9066), .C2(n9065), .A(n9073), .B(n9427), .ZN(n9071)
         );
  INV_X1 U10327 ( .A(n9077), .ZN(n9069) );
  NAND2_X1 U10328 ( .A1(n9564), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9067) );
  OAI211_X1 U10329 ( .C1(n9422), .C2(n9069), .A(n9068), .B(n9067), .ZN(n9070)
         );
  OR3_X1 U10330 ( .A1(n9072), .A2(n9071), .A3(n9070), .ZN(P1_U3258) );
  INV_X1 U10331 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9087) );
  XOR2_X1 U10332 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9091), .Z(n9075) );
  NAND2_X1 U10333 ( .A1(n9075), .A2(n9074), .ZN(n9090) );
  OAI21_X1 U10334 ( .B1(n9075), .B2(n9074), .A(n9090), .ZN(n9082) );
  AOI21_X1 U10335 ( .B1(n9077), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9076), .ZN(
        n9080) );
  NAND2_X1 U10336 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9091), .ZN(n9078) );
  OAI21_X1 U10337 ( .B1(n9091), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9078), .ZN(
        n9079) );
  NOR2_X1 U10338 ( .A1(n9080), .A2(n9079), .ZN(n9088) );
  AOI211_X1 U10339 ( .C1(n9080), .C2(n9079), .A(n9088), .B(n9571), .ZN(n9081)
         );
  AOI21_X1 U10340 ( .B1(n9587), .B2(n9082), .A(n9081), .ZN(n9086) );
  INV_X1 U10341 ( .A(n9083), .ZN(n9084) );
  AOI21_X1 U10342 ( .B1(n9579), .B2(n9091), .A(n9084), .ZN(n9085) );
  OAI211_X1 U10343 ( .C1(n9593), .C2(n9087), .A(n9086), .B(n9085), .ZN(
        P1_U3259) );
  AOI21_X1 U10344 ( .B1(n9091), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9088), .ZN(
        n9089) );
  XNOR2_X1 U10345 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9089), .ZN(n9095) );
  OAI21_X1 U10346 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9091), .A(n9090), .ZN(
        n9092) );
  XNOR2_X1 U10347 ( .A(n9092), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9093) );
  AOI22_X1 U10348 ( .A1(n9095), .A2(n9588), .B1(n9587), .B2(n9093), .ZN(n9097)
         );
  INV_X1 U10349 ( .A(n9093), .ZN(n9096) );
  XNOR2_X1 U10350 ( .A(n9319), .B(n9099), .ZN(n9100) );
  NAND2_X1 U10351 ( .A1(n9100), .A2(n9625), .ZN(n9318) );
  NOR2_X1 U10352 ( .A1(n9644), .A2(n9101), .ZN(n9104) );
  NAND2_X1 U10353 ( .A1(n9103), .A2(n9102), .ZN(n9320) );
  NOR2_X1 U10354 ( .A1(n9660), .A2(n9320), .ZN(n9111) );
  AOI211_X1 U10355 ( .C1(n9105), .C2(n9620), .A(n9104), .B(n9111), .ZN(n9106)
         );
  OAI21_X1 U10356 ( .B1(n9318), .B2(n9310), .A(n9106), .ZN(P1_U3261) );
  XNOR2_X1 U10357 ( .A(n9108), .B(n9107), .ZN(n9109) );
  NAND2_X1 U10358 ( .A1(n9109), .A2(n9625), .ZN(n9321) );
  NOR2_X1 U10359 ( .A1(n9322), .A2(n9263), .ZN(n9110) );
  AOI211_X1 U10360 ( .C1(n9660), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9111), .B(
        n9110), .ZN(n9112) );
  OAI21_X1 U10361 ( .B1(n9321), .B2(n9310), .A(n9112), .ZN(P1_U3262) );
  OAI21_X1 U10362 ( .B1(n9114), .B2(n9117), .A(n9113), .ZN(n9335) );
  NOR2_X1 U10363 ( .A1(n9115), .A2(n9293), .ZN(n9120) );
  AOI211_X1 U10364 ( .C1(n9118), .C2(n9117), .A(n9289), .B(n9116), .ZN(n9119)
         );
  AOI211_X2 U10365 ( .C1(n9614), .C2(n4490), .A(n9120), .B(n9119), .ZN(n9334)
         );
  OR2_X1 U10366 ( .A1(n9334), .A2(n9660), .ZN(n9128) );
  AOI211_X1 U10367 ( .C1(n9332), .C2(n9131), .A(n9295), .B(n9121), .ZN(n9331)
         );
  NOR2_X1 U10368 ( .A1(n9122), .A2(n9263), .ZN(n9126) );
  OAI22_X1 U10369 ( .A1(n9641), .A2(n9124), .B1(n9123), .B2(n9306), .ZN(n9125)
         );
  AOI211_X1 U10370 ( .C1(n9331), .C2(n9628), .A(n9126), .B(n9125), .ZN(n9127)
         );
  OAI211_X1 U10371 ( .C1(n9335), .C2(n9301), .A(n9128), .B(n9127), .ZN(
        P1_U3263) );
  XNOR2_X1 U10372 ( .A(n9129), .B(n9130), .ZN(n9340) );
  INV_X1 U10373 ( .A(n9131), .ZN(n9132) );
  AOI211_X1 U10374 ( .C1(n9337), .C2(n9148), .A(n9295), .B(n9132), .ZN(n9336)
         );
  INV_X1 U10375 ( .A(n9133), .ZN(n9134) );
  AOI22_X1 U10376 ( .A1(n9660), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9134), .B2(
        n9661), .ZN(n9135) );
  OAI21_X1 U10377 ( .B1(n4491), .B2(n9263), .A(n9135), .ZN(n9144) );
  NOR2_X1 U10378 ( .A1(n9136), .A2(n9293), .ZN(n9141) );
  AOI211_X1 U10379 ( .C1(n9139), .C2(n9138), .A(n9289), .B(n9137), .ZN(n9140)
         );
  AOI211_X1 U10380 ( .C1(n9614), .C2(n9142), .A(n9141), .B(n9140), .ZN(n9339)
         );
  NOR2_X1 U10381 ( .A1(n9339), .A2(n9660), .ZN(n9143) );
  AOI211_X1 U10382 ( .C1(n9628), .C2(n9336), .A(n9144), .B(n9143), .ZN(n9145)
         );
  OAI21_X1 U10383 ( .B1(n9340), .B2(n9301), .A(n9145), .ZN(P1_U3264) );
  XOR2_X1 U10384 ( .A(n9155), .B(n9146), .Z(n9345) );
  OR2_X1 U10385 ( .A1(n9153), .A2(n9171), .ZN(n9147) );
  OAI22_X1 U10386 ( .A1(n9641), .A2(n9150), .B1(n9149), .B2(n9306), .ZN(n9151)
         );
  INV_X1 U10387 ( .A(n9151), .ZN(n9152) );
  OAI21_X1 U10388 ( .B1(n9153), .B2(n9263), .A(n9152), .ZN(n9159) );
  OAI21_X1 U10389 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9157) );
  AOI222_X1 U10390 ( .A1(n9617), .A2(n9157), .B1(n9184), .B2(n9614), .C1(n4490), .C2(n9649), .ZN(n9344) );
  NOR2_X1 U10391 ( .A1(n9344), .A2(n9660), .ZN(n9158) );
  AOI211_X1 U10392 ( .C1(n9341), .C2(n9628), .A(n9159), .B(n9158), .ZN(n9160)
         );
  OAI21_X1 U10393 ( .B1(n9345), .B2(n9301), .A(n9160), .ZN(P1_U3265) );
  NOR2_X1 U10394 ( .A1(n9161), .A2(n9293), .ZN(n9165) );
  AOI211_X1 U10395 ( .C1(n9167), .C2(n9163), .A(n9289), .B(n9162), .ZN(n9164)
         );
  AOI211_X1 U10396 ( .C1(n9614), .C2(n9166), .A(n9165), .B(n9164), .ZN(n9349)
         );
  XNOR2_X1 U10397 ( .A(n9168), .B(n9167), .ZN(n9346) );
  INV_X1 U10398 ( .A(n9301), .ZN(n9629) );
  NAND2_X1 U10399 ( .A1(n9346), .A2(n9629), .ZN(n9178) );
  OAI22_X1 U10400 ( .A1(n9644), .A2(n9170), .B1(n9169), .B2(n9306), .ZN(n9175)
         );
  INV_X1 U10401 ( .A(n9171), .ZN(n9172) );
  OAI211_X1 U10402 ( .C1(n9173), .C2(n9186), .A(n9172), .B(n9625), .ZN(n9347)
         );
  NOR2_X1 U10403 ( .A1(n9347), .A2(n9310), .ZN(n9174) );
  AOI211_X1 U10404 ( .C1(n9620), .C2(n9176), .A(n9175), .B(n9174), .ZN(n9177)
         );
  OAI211_X1 U10405 ( .C1(n9660), .C2(n9349), .A(n9178), .B(n9177), .ZN(
        P1_U3266) );
  XOR2_X1 U10406 ( .A(n9179), .B(n9181), .Z(n9355) );
  OAI21_X1 U10407 ( .B1(n9182), .B2(n9181), .A(n9180), .ZN(n9185) );
  AOI222_X1 U10408 ( .A1(n9617), .A2(n9185), .B1(n9184), .B2(n9649), .C1(n9183), .C2(n9614), .ZN(n9354) );
  INV_X1 U10409 ( .A(n9197), .ZN(n9187) );
  AOI211_X1 U10410 ( .C1(n9352), .C2(n9187), .A(n9295), .B(n9186), .ZN(n9351)
         );
  NAND2_X1 U10411 ( .A1(n9351), .A2(n9188), .ZN(n9189) );
  OAI211_X1 U10412 ( .C1(n9306), .C2(n9190), .A(n9354), .B(n9189), .ZN(n9194)
         );
  OAI22_X1 U10413 ( .A1(n9192), .A2(n9263), .B1(n9191), .B2(n9641), .ZN(n9193)
         );
  AOI21_X1 U10414 ( .B1(n9194), .B2(n9644), .A(n9193), .ZN(n9195) );
  OAI21_X1 U10415 ( .B1(n9355), .B2(n9301), .A(n9195), .ZN(P1_U3267) );
  XOR2_X1 U10416 ( .A(n9203), .B(n9196), .Z(n9360) );
  AOI211_X1 U10417 ( .C1(n9357), .C2(n9217), .A(n9295), .B(n9197), .ZN(n9356)
         );
  AOI22_X1 U10418 ( .A1(n9198), .A2(n9661), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9660), .ZN(n9199) );
  OAI21_X1 U10419 ( .B1(n9200), .B2(n9263), .A(n9199), .ZN(n9209) );
  NOR2_X1 U10420 ( .A1(n9201), .A2(n9293), .ZN(n9206) );
  AOI211_X1 U10421 ( .C1(n9204), .C2(n9203), .A(n9289), .B(n9202), .ZN(n9205)
         );
  AOI211_X1 U10422 ( .C1(n9614), .C2(n9207), .A(n9206), .B(n9205), .ZN(n9359)
         );
  NOR2_X1 U10423 ( .A1(n9359), .A2(n9660), .ZN(n9208) );
  AOI211_X1 U10424 ( .C1(n9356), .C2(n9628), .A(n9209), .B(n9208), .ZN(n9210)
         );
  OAI21_X1 U10425 ( .B1(n9360), .B2(n9301), .A(n9210), .ZN(P1_U3268) );
  XNOR2_X1 U10426 ( .A(n9212), .B(n9211), .ZN(n9365) );
  XNOR2_X1 U10427 ( .A(n9214), .B(n9213), .ZN(n9215) );
  OAI222_X1 U10428 ( .A1(n9291), .A2(n9242), .B1(n9293), .B2(n9216), .C1(n9215), .C2(n9289), .ZN(n9361) );
  INV_X1 U10429 ( .A(n9217), .ZN(n9218) );
  AOI211_X1 U10430 ( .C1(n9363), .C2(n4452), .A(n9295), .B(n9218), .ZN(n9362)
         );
  NAND2_X1 U10431 ( .A1(n9362), .A2(n9628), .ZN(n9221) );
  AOI22_X1 U10432 ( .A1(n9219), .A2(n9661), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9660), .ZN(n9220) );
  OAI211_X1 U10433 ( .C1(n9222), .C2(n9263), .A(n9221), .B(n9220), .ZN(n9223)
         );
  AOI21_X1 U10434 ( .B1(n9361), .B2(n9644), .A(n9223), .ZN(n9224) );
  OAI21_X1 U10435 ( .B1(n9365), .B2(n9301), .A(n9224), .ZN(P1_U3269) );
  XNOR2_X1 U10436 ( .A(n9226), .B(n9225), .ZN(n9370) );
  XNOR2_X1 U10437 ( .A(n9228), .B(n9227), .ZN(n9229) );
  OAI222_X1 U10438 ( .A1(n9291), .A2(n9256), .B1(n9293), .B2(n9230), .C1(n9289), .C2(n9229), .ZN(n9366) );
  AOI211_X1 U10439 ( .C1(n9368), .C2(n9243), .A(n9295), .B(n9231), .ZN(n9367)
         );
  NAND2_X1 U10440 ( .A1(n9367), .A2(n9628), .ZN(n9234) );
  AOI22_X1 U10441 ( .A1(n9232), .A2(n9661), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9660), .ZN(n9233) );
  OAI211_X1 U10442 ( .C1(n9235), .C2(n9263), .A(n9234), .B(n9233), .ZN(n9236)
         );
  AOI21_X1 U10443 ( .B1(n9366), .B2(n9644), .A(n9236), .ZN(n9237) );
  OAI21_X1 U10444 ( .B1(n9370), .B2(n9301), .A(n9237), .ZN(P1_U3270) );
  XNOR2_X1 U10445 ( .A(n9238), .B(n9239), .ZN(n9375) );
  XNOR2_X1 U10446 ( .A(n9240), .B(n9239), .ZN(n9241) );
  OAI222_X1 U10447 ( .A1(n9291), .A2(n9277), .B1(n9293), .B2(n9242), .C1(n9241), .C2(n9289), .ZN(n9371) );
  INV_X1 U10448 ( .A(n9243), .ZN(n9244) );
  AOI211_X1 U10449 ( .C1(n9373), .C2(n9257), .A(n9295), .B(n9244), .ZN(n9372)
         );
  NAND2_X1 U10450 ( .A1(n9372), .A2(n9628), .ZN(n9248) );
  INV_X1 U10451 ( .A(n9245), .ZN(n9246) );
  AOI22_X1 U10452 ( .A1(n9246), .A2(n9661), .B1(n9660), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9247) );
  OAI211_X1 U10453 ( .C1(n9249), .C2(n9263), .A(n9248), .B(n9247), .ZN(n9250)
         );
  AOI21_X1 U10454 ( .B1(n9371), .B2(n9641), .A(n9250), .ZN(n9251) );
  OAI21_X1 U10455 ( .B1(n9375), .B2(n9301), .A(n9251), .ZN(P1_U3271) );
  XNOR2_X1 U10456 ( .A(n4356), .B(n4465), .ZN(n9380) );
  AOI21_X1 U10457 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(n9255) );
  OAI222_X1 U10458 ( .A1(n9293), .A2(n9256), .B1(n9291), .B2(n9292), .C1(n9289), .C2(n9255), .ZN(n9376) );
  INV_X1 U10459 ( .A(n9279), .ZN(n9259) );
  INV_X1 U10460 ( .A(n9257), .ZN(n9258) );
  AOI211_X1 U10461 ( .C1(n9378), .C2(n9259), .A(n9295), .B(n9258), .ZN(n9377)
         );
  NAND2_X1 U10462 ( .A1(n9377), .A2(n9628), .ZN(n9262) );
  AOI22_X1 U10463 ( .A1(n9660), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9260), .B2(
        n9661), .ZN(n9261) );
  OAI211_X1 U10464 ( .C1(n9264), .C2(n9263), .A(n9262), .B(n9261), .ZN(n9265)
         );
  AOI21_X1 U10465 ( .B1(n9376), .B2(n9644), .A(n9265), .ZN(n9266) );
  OAI21_X1 U10466 ( .B1(n9380), .B2(n9301), .A(n9266), .ZN(P1_U3272) );
  NAND2_X1 U10467 ( .A1(n9267), .A2(n9273), .ZN(n9381) );
  NAND3_X1 U10468 ( .A1(n4751), .A2(n9629), .A3(n9381), .ZN(n9284) );
  OAI22_X1 U10469 ( .A1(n9644), .A2(n9269), .B1(n9268), .B2(n9306), .ZN(n9270)
         );
  AOI21_X1 U10470 ( .B1(n9384), .B2(n9620), .A(n9270), .ZN(n9283) );
  NAND2_X1 U10471 ( .A1(n9272), .A2(n9271), .ZN(n9274) );
  XNOR2_X1 U10472 ( .A(n9274), .B(n9273), .ZN(n9275) );
  OAI222_X1 U10473 ( .A1(n9293), .A2(n9277), .B1(n9291), .B2(n9276), .C1(n9289), .C2(n9275), .ZN(n9382) );
  NAND2_X1 U10474 ( .A1(n9382), .A2(n9641), .ZN(n9282) );
  OAI21_X1 U10475 ( .B1(n9294), .B2(n9278), .A(n9625), .ZN(n9280) );
  NOR2_X1 U10476 ( .A1(n9280), .A2(n9279), .ZN(n9383) );
  NAND2_X1 U10477 ( .A1(n9383), .A2(n9628), .ZN(n9281) );
  NAND4_X1 U10478 ( .A1(n9284), .A2(n9283), .A3(n9282), .A4(n9281), .ZN(
        P1_U3273) );
  XNOR2_X1 U10479 ( .A(n9285), .B(n9286), .ZN(n9392) );
  XNOR2_X1 U10480 ( .A(n9287), .B(n9286), .ZN(n9288) );
  OAI222_X1 U10481 ( .A1(n9293), .A2(n9292), .B1(n9291), .B2(n9290), .C1(n9289), .C2(n9288), .ZN(n9388) );
  AOI211_X1 U10482 ( .C1(n9390), .C2(n4292), .A(n9295), .B(n9294), .ZN(n9389)
         );
  INV_X1 U10483 ( .A(n9389), .ZN(n9297) );
  OAI22_X1 U10484 ( .A1(n9297), .A2(n9638), .B1(n9306), .B2(n9296), .ZN(n9298)
         );
  OAI21_X1 U10485 ( .B1(n9388), .B2(n9298), .A(n9644), .ZN(n9300) );
  AOI22_X1 U10486 ( .A1(n9390), .A2(n9620), .B1(n9660), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n9299) );
  OAI211_X1 U10487 ( .C1(n9392), .C2(n9301), .A(n9300), .B(n9299), .ZN(
        P1_U3274) );
  XNOR2_X1 U10488 ( .A(n9302), .B(n9314), .ZN(n9305) );
  AOI222_X1 U10489 ( .A1(n9617), .A2(n9305), .B1(n9304), .B2(n9649), .C1(n9303), .C2(n9614), .ZN(n9505) );
  OAI22_X1 U10490 ( .A1(n9641), .A2(n9308), .B1(n9307), .B2(n9306), .ZN(n9312)
         );
  INV_X1 U10491 ( .A(n9313), .ZN(n9506) );
  OAI211_X1 U10492 ( .C1(n4453), .C2(n9506), .A(n9625), .B(n4292), .ZN(n9504)
         );
  NOR2_X1 U10493 ( .A1(n9504), .A2(n9310), .ZN(n9311) );
  AOI211_X1 U10494 ( .C1(n9620), .C2(n9313), .A(n9312), .B(n9311), .ZN(n9317)
         );
  XNOR2_X1 U10495 ( .A(n9315), .B(n9314), .ZN(n9508) );
  NAND2_X1 U10496 ( .A1(n9508), .A2(n9629), .ZN(n9316) );
  OAI211_X1 U10497 ( .C1(n9505), .C2(n9660), .A(n9317), .B(n9316), .ZN(
        P1_U3275) );
  OAI211_X1 U10498 ( .C1(n9319), .C2(n9723), .A(n9318), .B(n9320), .ZN(n9397)
         );
  MUX2_X1 U10499 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9397), .S(n9748), .Z(
        P1_U3554) );
  OAI211_X1 U10500 ( .C1(n9322), .C2(n9723), .A(n9321), .B(n9320), .ZN(n9398)
         );
  MUX2_X1 U10501 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9398), .S(n9748), .Z(
        P1_U3553) );
  MUX2_X1 U10502 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9399), .S(n9748), .Z(
        P1_U3552) );
  AOI21_X1 U10503 ( .B1(n9332), .B2(n9689), .A(n9331), .ZN(n9333) );
  OAI211_X1 U10504 ( .C1(n9335), .C2(n9659), .A(n9334), .B(n9333), .ZN(n9400)
         );
  MUX2_X1 U10505 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9400), .S(n9748), .Z(
        P1_U3551) );
  AOI21_X1 U10506 ( .B1(n9337), .B2(n9689), .A(n9336), .ZN(n9338) );
  OAI211_X1 U10507 ( .C1(n9340), .C2(n9659), .A(n9339), .B(n9338), .ZN(n9401)
         );
  MUX2_X1 U10508 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9401), .S(n9748), .Z(
        P1_U3550) );
  AOI21_X1 U10509 ( .B1(n9342), .B2(n9689), .A(n9341), .ZN(n9343) );
  OAI211_X1 U10510 ( .C1(n9345), .C2(n9659), .A(n9344), .B(n9343), .ZN(n9402)
         );
  MUX2_X1 U10511 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9402), .S(n9748), .Z(
        P1_U3549) );
  INV_X1 U10512 ( .A(n9659), .ZN(n9725) );
  NAND2_X1 U10513 ( .A1(n9346), .A2(n9725), .ZN(n9350) );
  NAND4_X1 U10514 ( .A1(n9350), .A2(n9349), .A3(n9348), .A4(n9347), .ZN(n9403)
         );
  MUX2_X1 U10515 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9403), .S(n9748), .Z(
        P1_U3548) );
  AOI21_X1 U10516 ( .B1(n9352), .B2(n9689), .A(n9351), .ZN(n9353) );
  OAI211_X1 U10517 ( .C1(n9355), .C2(n9659), .A(n9354), .B(n9353), .ZN(n9404)
         );
  MUX2_X1 U10518 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9404), .S(n9748), .Z(
        P1_U3547) );
  AOI21_X1 U10519 ( .B1(n9357), .B2(n9689), .A(n9356), .ZN(n9358) );
  OAI211_X1 U10520 ( .C1(n9360), .C2(n9659), .A(n9359), .B(n9358), .ZN(n9405)
         );
  MUX2_X1 U10521 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9405), .S(n9748), .Z(
        P1_U3546) );
  AOI211_X1 U10522 ( .C1(n9363), .C2(n9689), .A(n9362), .B(n9361), .ZN(n9364)
         );
  OAI21_X1 U10523 ( .B1(n9365), .B2(n9659), .A(n9364), .ZN(n9406) );
  MUX2_X1 U10524 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9406), .S(n9748), .Z(
        P1_U3545) );
  AOI211_X1 U10525 ( .C1(n9368), .C2(n9689), .A(n9367), .B(n9366), .ZN(n9369)
         );
  OAI21_X1 U10526 ( .B1(n9370), .B2(n9659), .A(n9369), .ZN(n9407) );
  MUX2_X1 U10527 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9407), .S(n9748), .Z(
        P1_U3544) );
  AOI211_X1 U10528 ( .C1(n9373), .C2(n9689), .A(n9372), .B(n9371), .ZN(n9374)
         );
  OAI21_X1 U10529 ( .B1(n9375), .B2(n9659), .A(n9374), .ZN(n9408) );
  MUX2_X1 U10530 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9408), .S(n9748), .Z(
        P1_U3543) );
  AOI211_X1 U10531 ( .C1(n9378), .C2(n9689), .A(n9377), .B(n9376), .ZN(n9379)
         );
  OAI21_X1 U10532 ( .B1(n9659), .B2(n9380), .A(n9379), .ZN(n9409) );
  MUX2_X1 U10533 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9409), .S(n9748), .Z(
        P1_U3542) );
  NAND2_X1 U10534 ( .A1(n9381), .A2(n9725), .ZN(n9386) );
  AOI211_X1 U10535 ( .C1(n9384), .C2(n9689), .A(n9383), .B(n9382), .ZN(n9385)
         );
  OAI21_X1 U10536 ( .B1(n9387), .B2(n9386), .A(n9385), .ZN(n9410) );
  MUX2_X1 U10537 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9410), .S(n9748), .Z(
        P1_U3541) );
  AOI211_X1 U10538 ( .C1(n9390), .C2(n9689), .A(n9389), .B(n9388), .ZN(n9391)
         );
  OAI21_X1 U10539 ( .B1(n9659), .B2(n9392), .A(n9391), .ZN(n9411) );
  MUX2_X1 U10540 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9411), .S(n9748), .Z(
        P1_U3540) );
  NOR2_X1 U10541 ( .A1(n9394), .A2(n9393), .ZN(n9395) );
  AND2_X2 U10542 ( .A1(n9396), .A2(n9395), .ZN(n9729) );
  MUX2_X1 U10543 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9397), .S(n9729), .Z(
        P1_U3522) );
  MUX2_X1 U10544 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9398), .S(n9729), .Z(
        P1_U3521) );
  MUX2_X1 U10545 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9400), .S(n9729), .Z(
        P1_U3519) );
  MUX2_X1 U10546 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9401), .S(n9729), .Z(
        P1_U3518) );
  MUX2_X1 U10547 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9402), .S(n9729), .Z(
        P1_U3517) );
  MUX2_X1 U10548 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9403), .S(n9729), .Z(
        P1_U3516) );
  MUX2_X1 U10549 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9404), .S(n9729), .Z(
        P1_U3515) );
  MUX2_X1 U10550 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9405), .S(n9729), .Z(
        P1_U3514) );
  MUX2_X1 U10551 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9406), .S(n9729), .Z(
        P1_U3513) );
  MUX2_X1 U10552 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9407), .S(n9729), .Z(
        P1_U3512) );
  MUX2_X1 U10553 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9408), .S(n9729), .Z(
        P1_U3511) );
  MUX2_X1 U10554 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9409), .S(n9729), .Z(
        P1_U3510) );
  MUX2_X1 U10555 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9410), .S(n9729), .Z(
        P1_U3508) );
  MUX2_X1 U10556 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9411), .S(n9729), .Z(
        P1_U3505) );
  NAND4_X1 U10557 ( .A1(n5097), .A2(n9413), .A3(P1_IR_REG_31__SCAN_IN), .A4(
        P1_STATE_REG_SCAN_IN), .ZN(n9414) );
  OAI22_X1 U10558 ( .A1(n9412), .A2(n9414), .B1(n5125), .B2(n7361), .ZN(n9415)
         );
  INV_X1 U10559 ( .A(n9415), .ZN(n9416) );
  OAI21_X1 U10560 ( .B1(n9418), .B2(n9417), .A(n9416), .ZN(P1_U3322) );
  MUX2_X1 U10561 ( .A(n9419), .B(n9558), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  OAI22_X1 U10562 ( .A1(n9422), .A2(n9421), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9420), .ZN(n9423) );
  AOI21_X1 U10563 ( .B1(n9564), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9423), .ZN(
        n9434) );
  OAI211_X1 U10564 ( .C1(n9426), .C2(n9425), .A(n9588), .B(n9424), .ZN(n9433)
         );
  AOI211_X1 U10565 ( .C1(n9430), .C2(n9429), .A(n9428), .B(n9427), .ZN(n9431)
         );
  INV_X1 U10566 ( .A(n9431), .ZN(n9432) );
  NAND3_X1 U10567 ( .A1(n9434), .A2(n9433), .A3(n9432), .ZN(P1_U3244) );
  AOI22_X1 U10568 ( .A1(n9755), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9445) );
  NAND2_X1 U10569 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9437) );
  AOI211_X1 U10570 ( .C1(n9437), .C2(n9436), .A(n9435), .B(n9753), .ZN(n9442)
         );
  NAND2_X1 U10571 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9440) );
  AOI211_X1 U10572 ( .C1(n9440), .C2(n9439), .A(n9438), .B(n9449), .ZN(n9441)
         );
  AOI211_X1 U10573 ( .C1(n9456), .C2(n9443), .A(n9442), .B(n9441), .ZN(n9444)
         );
  NAND2_X1 U10574 ( .A1(n9445), .A2(n9444), .ZN(P2_U3246) );
  AOI22_X1 U10575 ( .A1(n9755), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9458) );
  AOI211_X1 U10576 ( .C1(n9448), .C2(n9447), .A(n9446), .B(n9753), .ZN(n9454)
         );
  AOI211_X1 U10577 ( .C1(n9452), .C2(n9451), .A(n9450), .B(n9449), .ZN(n9453)
         );
  AOI211_X1 U10578 ( .C1(n9456), .C2(n9455), .A(n9454), .B(n9453), .ZN(n9457)
         );
  NAND2_X1 U10579 ( .A1(n9458), .A2(n9457), .ZN(P2_U3247) );
  OAI21_X1 U10580 ( .B1(n9460), .B2(n9723), .A(n9459), .ZN(n9462) );
  AOI211_X1 U10581 ( .C1(n9463), .C2(n9725), .A(n9462), .B(n9461), .ZN(n9465)
         );
  AOI22_X1 U10582 ( .A1(n9729), .A2(n9465), .B1(n6404), .B2(n9727), .ZN(
        P1_U3484) );
  INV_X1 U10583 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9464) );
  AOI22_X1 U10584 ( .A1(n9748), .A2(n9465), .B1(n9464), .B2(n9745), .ZN(
        P1_U3533) );
  NOR2_X1 U10585 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9466) );
  AOI21_X1 U10586 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9466), .ZN(n9936) );
  NOR2_X1 U10587 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n9467) );
  AOI21_X1 U10588 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9467), .ZN(n9939) );
  NOR2_X1 U10589 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9468) );
  AOI21_X1 U10590 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9468), .ZN(n9942) );
  NOR2_X1 U10591 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9469) );
  AOI21_X1 U10592 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9469), .ZN(n9945) );
  NOR2_X1 U10593 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9470) );
  AOI21_X1 U10594 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9470), .ZN(n9948) );
  NOR2_X1 U10595 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9477) );
  XNOR2_X1 U10596 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9979) );
  NAND2_X1 U10597 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9475) );
  XOR2_X1 U10598 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n9977) );
  NAND2_X1 U10599 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9473) );
  XOR2_X1 U10600 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n9975) );
  AOI21_X1 U10601 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9928) );
  INV_X1 U10602 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9471) );
  NAND3_X1 U10603 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9930) );
  OAI21_X1 U10604 ( .B1(n9928), .B2(n9471), .A(n9930), .ZN(n9974) );
  NAND2_X1 U10605 ( .A1(n9975), .A2(n9974), .ZN(n9472) );
  NAND2_X1 U10606 ( .A1(n9473), .A2(n9472), .ZN(n9976) );
  NAND2_X1 U10607 ( .A1(n9977), .A2(n9976), .ZN(n9474) );
  NAND2_X1 U10608 ( .A1(n9475), .A2(n9474), .ZN(n9978) );
  NOR2_X1 U10609 ( .A1(n9979), .A2(n9978), .ZN(n9476) );
  NOR2_X1 U10610 ( .A1(n9477), .A2(n9476), .ZN(n9478) );
  NOR2_X1 U10611 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9478), .ZN(n9963) );
  AND2_X1 U10612 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9478), .ZN(n9962) );
  NOR2_X1 U10613 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9962), .ZN(n9479) );
  NOR2_X1 U10614 ( .A1(n9963), .A2(n9479), .ZN(n9480) );
  NAND2_X1 U10615 ( .A1(n9480), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9482) );
  XOR2_X1 U10616 ( .A(n9480), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9961) );
  NAND2_X1 U10617 ( .A1(n9961), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U10618 ( .A1(n9482), .A2(n9481), .ZN(n9483) );
  NAND2_X1 U10619 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9483), .ZN(n9485) );
  XOR2_X1 U10620 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9483), .Z(n9966) );
  NAND2_X1 U10621 ( .A1(n9966), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U10622 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  NAND2_X1 U10623 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9486), .ZN(n9488) );
  XOR2_X1 U10624 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9486), .Z(n9959) );
  NAND2_X1 U10625 ( .A1(n9959), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U10626 ( .A1(n9488), .A2(n9487), .ZN(n9489) );
  AND2_X1 U10627 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n9489), .ZN(n9490) );
  XNOR2_X1 U10628 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n9489), .ZN(n9972) );
  NOR2_X1 U10629 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  NAND2_X1 U10630 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9491) );
  OAI21_X1 U10631 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9491), .ZN(n9956) );
  AOI21_X1 U10632 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9955), .ZN(n9954) );
  NAND2_X1 U10633 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9492) );
  OAI21_X1 U10634 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9492), .ZN(n9953) );
  NOR2_X1 U10635 ( .A1(n9954), .A2(n9953), .ZN(n9952) );
  AOI21_X1 U10636 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9952), .ZN(n9951) );
  NOR2_X1 U10637 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9493) );
  AOI21_X1 U10638 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9493), .ZN(n9950) );
  NAND2_X1 U10639 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  OAI21_X1 U10640 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9949), .ZN(n9947) );
  NAND2_X1 U10641 ( .A1(n9948), .A2(n9947), .ZN(n9946) );
  OAI21_X1 U10642 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9946), .ZN(n9944) );
  NAND2_X1 U10643 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  OAI21_X1 U10644 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9943), .ZN(n9941) );
  NAND2_X1 U10645 ( .A1(n9942), .A2(n9941), .ZN(n9940) );
  OAI21_X1 U10646 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9940), .ZN(n9938) );
  NAND2_X1 U10647 ( .A1(n9939), .A2(n9938), .ZN(n9937) );
  OAI21_X1 U10648 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9937), .ZN(n9935) );
  NAND2_X1 U10649 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  OAI21_X1 U10650 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9934), .ZN(n9968) );
  NOR2_X1 U10651 ( .A1(n9969), .A2(n9968), .ZN(n9494) );
  NAND2_X1 U10652 ( .A1(n9969), .A2(n9968), .ZN(n9967) );
  OAI21_X1 U10653 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9494), .A(n9967), .ZN(
        n9496) );
  XOR2_X1 U10654 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n9495) );
  XNOR2_X1 U10655 ( .A(n9496), .B(n9495), .ZN(ADD_1071_U4) );
  OAI21_X1 U10656 ( .B1(n9498), .B2(n9900), .A(n9497), .ZN(n9499) );
  AOI21_X1 U10657 ( .B1(n9501), .B2(n9500), .A(n9499), .ZN(n9503) );
  AOI22_X1 U10658 ( .A1(n9927), .A2(n9503), .B1(n7521), .B2(n9925), .ZN(
        P2_U3550) );
  AOI22_X1 U10659 ( .A1(n9910), .A2(n9503), .B1(n9502), .B2(n9908), .ZN(
        P2_U3518) );
  OAI211_X1 U10660 ( .C1(n9506), .C2(n9723), .A(n9505), .B(n9504), .ZN(n9507)
         );
  AOI21_X1 U10661 ( .B1(n9508), .B2(n9725), .A(n9507), .ZN(n9544) );
  AOI22_X1 U10662 ( .A1(n9748), .A2(n9544), .B1(n9509), .B2(n9745), .ZN(
        P1_U3539) );
  OAI21_X1 U10663 ( .B1(n9511), .B2(n9723), .A(n9510), .ZN(n9512) );
  AOI21_X1 U10664 ( .B1(n9513), .B2(n9720), .A(n9512), .ZN(n9514) );
  AND2_X1 U10665 ( .A1(n9515), .A2(n9514), .ZN(n9546) );
  AOI22_X1 U10666 ( .A1(n9748), .A2(n9546), .B1(n9516), .B2(n9745), .ZN(
        P1_U3538) );
  OAI21_X1 U10667 ( .B1(n9518), .B2(n9723), .A(n9517), .ZN(n9520) );
  AOI211_X1 U10668 ( .C1(n9521), .C2(n9725), .A(n9520), .B(n9519), .ZN(n9548)
         );
  AOI22_X1 U10669 ( .A1(n9748), .A2(n9548), .B1(n9522), .B2(n9745), .ZN(
        P1_U3537) );
  INV_X1 U10670 ( .A(n9523), .ZN(n9525) );
  OAI21_X1 U10671 ( .B1(n9525), .B2(n9723), .A(n9524), .ZN(n9526) );
  AOI21_X1 U10672 ( .B1(n9527), .B2(n9720), .A(n9526), .ZN(n9528) );
  AND2_X1 U10673 ( .A1(n9529), .A2(n9528), .ZN(n9550) );
  AOI22_X1 U10674 ( .A1(n9748), .A2(n9550), .B1(n6602), .B2(n9745), .ZN(
        P1_U3536) );
  NAND2_X1 U10675 ( .A1(n9530), .A2(n9689), .ZN(n9531) );
  NAND2_X1 U10676 ( .A1(n9532), .A2(n9531), .ZN(n9533) );
  AOI21_X1 U10677 ( .B1(n9534), .B2(n9720), .A(n9533), .ZN(n9535) );
  AND2_X1 U10678 ( .A1(n9536), .A2(n9535), .ZN(n9552) );
  AOI22_X1 U10679 ( .A1(n9748), .A2(n9552), .B1(n6593), .B2(n9745), .ZN(
        P1_U3535) );
  INV_X1 U10680 ( .A(n9537), .ZN(n9542) );
  OAI21_X1 U10681 ( .B1(n9539), .B2(n9723), .A(n9538), .ZN(n9541) );
  AOI211_X1 U10682 ( .C1(n9720), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9554)
         );
  AOI22_X1 U10683 ( .A1(n9748), .A2(n9554), .B1(n9543), .B2(n9745), .ZN(
        P1_U3534) );
  AOI22_X1 U10684 ( .A1(n9729), .A2(n9544), .B1(n6879), .B2(n9727), .ZN(
        P1_U3502) );
  INV_X1 U10685 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9545) );
  AOI22_X1 U10686 ( .A1(n9729), .A2(n9546), .B1(n9545), .B2(n9727), .ZN(
        P1_U3499) );
  INV_X1 U10687 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9547) );
  AOI22_X1 U10688 ( .A1(n9729), .A2(n9548), .B1(n9547), .B2(n9727), .ZN(
        P1_U3496) );
  AOI22_X1 U10689 ( .A1(n9729), .A2(n9550), .B1(n9549), .B2(n9727), .ZN(
        P1_U3493) );
  INV_X1 U10690 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9551) );
  AOI22_X1 U10691 ( .A1(n9729), .A2(n9552), .B1(n9551), .B2(n9727), .ZN(
        P1_U3490) );
  INV_X1 U10692 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9553) );
  AOI22_X1 U10693 ( .A1(n9729), .A2(n9554), .B1(n9553), .B2(n9727), .ZN(
        P1_U3487) );
  XNOR2_X1 U10694 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10695 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10696 ( .A(n9555), .ZN(n9556) );
  OAI21_X1 U10697 ( .B1(n9557), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9556), .ZN(
        n9559) );
  XNOR2_X1 U10698 ( .A(n9559), .B(n9558), .ZN(n9561) );
  AOI22_X1 U10699 ( .A1(n9561), .A2(n9560), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3084), .ZN(n9562) );
  OAI21_X1 U10700 ( .B1(n9932), .B2(n9593), .A(n9562), .ZN(P1_U3241) );
  AOI22_X1 U10701 ( .A1(n9564), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9579), .B2(
        n9563), .ZN(n9576) );
  OAI211_X1 U10702 ( .C1(n9567), .C2(n9566), .A(n9565), .B(n9587), .ZN(n9574)
         );
  AOI21_X1 U10703 ( .B1(n9570), .B2(n9569), .A(n9568), .ZN(n9572) );
  OR2_X1 U10704 ( .A1(n9572), .A2(n9571), .ZN(n9573) );
  NAND4_X1 U10705 ( .A1(n9576), .A2(n9575), .A3(n9574), .A4(n9573), .ZN(
        P1_U3246) );
  INV_X1 U10706 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9592) );
  AOI21_X1 U10707 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9591) );
  OAI21_X1 U10708 ( .B1(n9582), .B2(n9581), .A(n9580), .ZN(n9589) );
  OAI21_X1 U10709 ( .B1(n9585), .B2(n9584), .A(n9583), .ZN(n9586) );
  AOI22_X1 U10710 ( .A1(n9589), .A2(n9588), .B1(n9587), .B2(n9586), .ZN(n9590)
         );
  OAI211_X1 U10711 ( .C1(n9593), .C2(n9592), .A(n9591), .B(n9590), .ZN(
        P1_U3252) );
  NAND2_X1 U10712 ( .A1(n9595), .A2(n9594), .ZN(n9596) );
  XNOR2_X1 U10713 ( .A(n9596), .B(n9605), .ZN(n9598) );
  AOI222_X1 U10714 ( .A1(n9617), .A2(n9598), .B1(n9597), .B2(n9649), .C1(n9613), .C2(n9614), .ZN(n9722) );
  INV_X1 U10715 ( .A(n9599), .ZN(n9600) );
  AOI222_X1 U10716 ( .A1(n9601), .A2(n9620), .B1(P1_REG2_REG_9__SCAN_IN), .B2(
        n9660), .C1(n9661), .C2(n9600), .ZN(n9611) );
  NAND2_X1 U10717 ( .A1(n9603), .A2(n9602), .ZN(n9604) );
  XOR2_X1 U10718 ( .A(n9605), .B(n9604), .Z(n9726) );
  INV_X1 U10719 ( .A(n9606), .ZN(n9608) );
  OAI211_X1 U10720 ( .C1(n9608), .C2(n4445), .A(n9625), .B(n9607), .ZN(n9721)
         );
  INV_X1 U10721 ( .A(n9721), .ZN(n9609) );
  AOI22_X1 U10722 ( .A1(n9726), .A2(n9629), .B1(n9628), .B2(n9609), .ZN(n9610)
         );
  OAI211_X1 U10723 ( .C1(n9660), .C2(n9722), .A(n9611), .B(n9610), .ZN(
        P1_U3282) );
  XNOR2_X1 U10724 ( .A(n9612), .B(n9622), .ZN(n9616) );
  AOI222_X1 U10725 ( .A1(n9617), .A2(n9616), .B1(n9615), .B2(n9614), .C1(n9613), .C2(n9649), .ZN(n9710) );
  INV_X1 U10726 ( .A(n9618), .ZN(n9619) );
  AOI222_X1 U10727 ( .A1(n9621), .A2(n9620), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9660), .C1(n9661), .C2(n9619), .ZN(n9631) );
  XNOR2_X1 U10728 ( .A(n9623), .B(n9622), .ZN(n9713) );
  OAI211_X1 U10729 ( .C1(n9626), .C2(n9711), .A(n9625), .B(n9624), .ZN(n9709)
         );
  INV_X1 U10730 ( .A(n9709), .ZN(n9627) );
  AOI22_X1 U10731 ( .A1(n9713), .A2(n9629), .B1(n9628), .B2(n9627), .ZN(n9630)
         );
  OAI211_X1 U10732 ( .C1(n9660), .C2(n9710), .A(n9631), .B(n9630), .ZN(
        P1_U3284) );
  INV_X1 U10733 ( .A(n9632), .ZN(n9636) );
  AOI22_X1 U10734 ( .A1(n9661), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9634), .B2(
        n9633), .ZN(n9635) );
  OAI211_X1 U10735 ( .C1(n9638), .C2(n9637), .A(n9636), .B(n9635), .ZN(n9642)
         );
  AOI22_X1 U10736 ( .A1(n9642), .A2(n9641), .B1(n9640), .B2(n9639), .ZN(n9643)
         );
  OAI21_X1 U10737 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(P1_U3290) );
  NAND2_X1 U10738 ( .A1(n9646), .A2(n9652), .ZN(n9647) );
  OR2_X1 U10739 ( .A1(n9648), .A2(n9647), .ZN(n9651) );
  NAND2_X1 U10740 ( .A1(n5380), .A2(n9649), .ZN(n9650) );
  AND2_X1 U10741 ( .A1(n9651), .A2(n9650), .ZN(n9656) );
  INV_X1 U10742 ( .A(n9656), .ZN(n9658) );
  INV_X1 U10743 ( .A(n9652), .ZN(n9653) );
  NAND2_X1 U10744 ( .A1(n9654), .A2(n9653), .ZN(n9655) );
  AND2_X1 U10745 ( .A1(n9656), .A2(n9655), .ZN(n9731) );
  INV_X1 U10746 ( .A(n9731), .ZN(n9657) );
  OAI21_X1 U10747 ( .B1(n9659), .B2(n9658), .A(n9657), .ZN(n9663) );
  AOI22_X1 U10748 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n9661), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n9660), .ZN(n9662) );
  OAI21_X1 U10749 ( .B1(n9660), .B2(n9663), .A(n9662), .ZN(P1_U3291) );
  AND2_X1 U10750 ( .A1(n9665), .A2(n9664), .ZN(n9671) );
  AND2_X1 U10751 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9672), .ZN(P1_U3292) );
  AND2_X1 U10752 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9672), .ZN(P1_U3293) );
  AND2_X1 U10753 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9672), .ZN(P1_U3294) );
  AND2_X1 U10754 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9672), .ZN(P1_U3295) );
  AND2_X1 U10755 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9672), .ZN(P1_U3296) );
  NOR2_X1 U10756 ( .A1(n9671), .A2(n9666), .ZN(P1_U3297) );
  AND2_X1 U10757 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9672), .ZN(P1_U3298) );
  AND2_X1 U10758 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9672), .ZN(P1_U3299) );
  AND2_X1 U10759 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9672), .ZN(P1_U3300) );
  AND2_X1 U10760 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9672), .ZN(P1_U3301) );
  AND2_X1 U10761 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9672), .ZN(P1_U3302) );
  AND2_X1 U10762 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9672), .ZN(P1_U3303) );
  AND2_X1 U10763 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9672), .ZN(P1_U3304) );
  AND2_X1 U10764 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9672), .ZN(P1_U3305) );
  AND2_X1 U10765 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9672), .ZN(P1_U3306) );
  AND2_X1 U10766 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9672), .ZN(P1_U3307) );
  NOR2_X1 U10767 ( .A1(n9671), .A2(n9667), .ZN(P1_U3308) );
  NOR2_X1 U10768 ( .A1(n9671), .A2(n9668), .ZN(P1_U3309) );
  AND2_X1 U10769 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9672), .ZN(P1_U3310) );
  AND2_X1 U10770 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9672), .ZN(P1_U3311) );
  NOR2_X1 U10771 ( .A1(n9671), .A2(n9669), .ZN(P1_U3312) );
  NOR2_X1 U10772 ( .A1(n9671), .A2(n9670), .ZN(P1_U3313) );
  AND2_X1 U10773 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9672), .ZN(P1_U3314) );
  AND2_X1 U10774 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9672), .ZN(P1_U3315) );
  AND2_X1 U10775 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9672), .ZN(P1_U3316) );
  AND2_X1 U10776 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9672), .ZN(P1_U3317) );
  AND2_X1 U10777 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9672), .ZN(P1_U3318) );
  AND2_X1 U10778 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9672), .ZN(P1_U3319) );
  AND2_X1 U10779 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9672), .ZN(P1_U3320) );
  AND2_X1 U10780 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9672), .ZN(P1_U3321) );
  AOI22_X1 U10781 ( .A1(n9729), .A2(n9731), .B1(n5106), .B2(n9727), .ZN(
        P1_U3454) );
  INV_X1 U10782 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9673) );
  AOI22_X1 U10783 ( .A1(n9729), .A2(n9674), .B1(n9673), .B2(n9727), .ZN(
        P1_U3457) );
  INV_X1 U10784 ( .A(n9675), .ZN(n9676) );
  OAI21_X1 U10785 ( .B1(n9677), .B2(n9723), .A(n9676), .ZN(n9679) );
  AOI211_X1 U10786 ( .C1(n9720), .C2(n9680), .A(n9679), .B(n9678), .ZN(n9733)
         );
  INV_X1 U10787 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9681) );
  AOI22_X1 U10788 ( .A1(n9729), .A2(n9733), .B1(n9681), .B2(n9727), .ZN(
        P1_U3460) );
  OAI21_X1 U10789 ( .B1(n9683), .B2(n9723), .A(n9682), .ZN(n9685) );
  AOI211_X1 U10790 ( .C1(n9720), .C2(n9686), .A(n9685), .B(n9684), .ZN(n9735)
         );
  INV_X1 U10791 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9687) );
  AOI22_X1 U10792 ( .A1(n9729), .A2(n9735), .B1(n9687), .B2(n9727), .ZN(
        P1_U3463) );
  AOI21_X1 U10793 ( .B1(n9690), .B2(n9689), .A(n9688), .ZN(n9691) );
  OAI211_X1 U10794 ( .C1(n9694), .C2(n9693), .A(n9692), .B(n9691), .ZN(n9695)
         );
  INV_X1 U10795 ( .A(n9695), .ZN(n9737) );
  AOI22_X1 U10796 ( .A1(n9729), .A2(n9737), .B1(n5529), .B2(n9727), .ZN(
        P1_U3466) );
  OAI21_X1 U10797 ( .B1(n9697), .B2(n9723), .A(n9696), .ZN(n9698) );
  AOI21_X1 U10798 ( .B1(n9699), .B2(n9725), .A(n9698), .ZN(n9701) );
  AND2_X1 U10799 ( .A1(n9701), .A2(n9700), .ZN(n9738) );
  INV_X1 U10800 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9702) );
  AOI22_X1 U10801 ( .A1(n9729), .A2(n9738), .B1(n9702), .B2(n9727), .ZN(
        P1_U3469) );
  OAI21_X1 U10802 ( .B1(n9704), .B2(n9723), .A(n9703), .ZN(n9706) );
  AOI211_X1 U10803 ( .C1(n9720), .C2(n9707), .A(n9706), .B(n9705), .ZN(n9740)
         );
  INV_X1 U10804 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9708) );
  AOI22_X1 U10805 ( .A1(n9729), .A2(n9740), .B1(n9708), .B2(n9727), .ZN(
        P1_U3472) );
  OAI211_X1 U10806 ( .C1(n9711), .C2(n9723), .A(n9710), .B(n9709), .ZN(n9712)
         );
  AOI21_X1 U10807 ( .B1(n9725), .B2(n9713), .A(n9712), .ZN(n9742) );
  INV_X1 U10808 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9714) );
  AOI22_X1 U10809 ( .A1(n9729), .A2(n9742), .B1(n9714), .B2(n9727), .ZN(
        P1_U3475) );
  INV_X1 U10810 ( .A(n9715), .ZN(n9719) );
  OAI21_X1 U10811 ( .B1(n4446), .B2(n9723), .A(n9716), .ZN(n9718) );
  AOI211_X1 U10812 ( .C1(n9720), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9744)
         );
  AOI22_X1 U10813 ( .A1(n9729), .A2(n9744), .B1(n6075), .B2(n9727), .ZN(
        P1_U3478) );
  OAI211_X1 U10814 ( .C1(n4445), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9724)
         );
  AOI21_X1 U10815 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(n9747) );
  AOI22_X1 U10816 ( .A1(n9729), .A2(n9747), .B1(n9728), .B2(n9727), .ZN(
        P1_U3481) );
  AOI22_X1 U10817 ( .A1(n9748), .A2(n9731), .B1(n9730), .B2(n9745), .ZN(
        P1_U3523) );
  AOI22_X1 U10818 ( .A1(n9748), .A2(n9733), .B1(n9732), .B2(n9745), .ZN(
        P1_U3525) );
  AOI22_X1 U10819 ( .A1(n9748), .A2(n9735), .B1(n9734), .B2(n9745), .ZN(
        P1_U3526) );
  AOI22_X1 U10820 ( .A1(n9748), .A2(n9737), .B1(n9736), .B2(n9745), .ZN(
        P1_U3527) );
  AOI22_X1 U10821 ( .A1(n9748), .A2(n9738), .B1(n5664), .B2(n9745), .ZN(
        P1_U3528) );
  AOI22_X1 U10822 ( .A1(n9748), .A2(n9740), .B1(n9739), .B2(n9745), .ZN(
        P1_U3529) );
  AOI22_X1 U10823 ( .A1(n9748), .A2(n9742), .B1(n9741), .B2(n9745), .ZN(
        P1_U3530) );
  INV_X1 U10824 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9743) );
  AOI22_X1 U10825 ( .A1(n9748), .A2(n9744), .B1(n9743), .B2(n9745), .ZN(
        P1_U3531) );
  INV_X1 U10826 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9746) );
  AOI22_X1 U10827 ( .A1(n9748), .A2(n9747), .B1(n9746), .B2(n9745), .ZN(
        P1_U3532) );
  AOI22_X1 U10828 ( .A1(n9750), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9749), .ZN(n9759) );
  NAND2_X1 U10829 ( .A1(n9750), .A2(n6151), .ZN(n9752) );
  OAI211_X1 U10830 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9753), .A(n9752), .B(
        n9751), .ZN(n9754) );
  INV_X1 U10831 ( .A(n9754), .ZN(n9757) );
  AOI22_X1 U10832 ( .A1(n9755), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9756) );
  OAI221_X1 U10833 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9759), .C1(n9758), .C2(
        n9757), .A(n9756), .ZN(P2_U3245) );
  NAND2_X1 U10834 ( .A1(n9761), .A2(n9777), .ZN(n9762) );
  NAND2_X1 U10835 ( .A1(n9760), .A2(n9762), .ZN(n9782) );
  INV_X1 U10836 ( .A(n9782), .ZN(n9891) );
  INV_X1 U10837 ( .A(n9798), .ZN(n9768) );
  INV_X1 U10838 ( .A(n9763), .ZN(n9764) );
  OAI21_X1 U10839 ( .B1(n9887), .B2(n9765), .A(n9764), .ZN(n9888) );
  INV_X1 U10840 ( .A(n9888), .ZN(n9766) );
  AOI22_X1 U10841 ( .A1(n9891), .A2(n9768), .B1(n9767), .B2(n9766), .ZN(n9790)
         );
  AOI22_X1 U10842 ( .A1(n9772), .A2(n9771), .B1(n9770), .B2(n9769), .ZN(n9780)
         );
  INV_X1 U10843 ( .A(n9774), .ZN(n9778) );
  OR2_X1 U10844 ( .A1(n9774), .A2(n9773), .ZN(n9775) );
  OAI211_X1 U10845 ( .C1(n9778), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9779)
         );
  OAI211_X1 U10846 ( .C1(n9782), .C2(n9781), .A(n9780), .B(n9779), .ZN(n9889)
         );
  NOR2_X1 U10847 ( .A1(n9795), .A2(n9887), .ZN(n9787) );
  OAI22_X1 U10848 ( .A1(n9785), .A2(n9784), .B1(n9783), .B2(n9792), .ZN(n9786)
         );
  AOI211_X1 U10849 ( .C1(n9889), .C2(n9788), .A(n9787), .B(n9786), .ZN(n9789)
         );
  NAND2_X1 U10850 ( .A1(n9790), .A2(n9789), .ZN(P2_U3286) );
  INV_X1 U10851 ( .A(n9791), .ZN(n9794) );
  OAI22_X1 U10852 ( .A1(n9794), .A2(n9793), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9792), .ZN(n9800) );
  OAI22_X1 U10853 ( .A1(n9798), .A2(n9797), .B1(n9796), .B2(n9795), .ZN(n9799)
         );
  AOI211_X1 U10854 ( .C1(P2_REG2_REG_3__SCAN_IN), .C2(n8399), .A(n9800), .B(
        n9799), .ZN(n9801) );
  OAI21_X1 U10855 ( .B1(n8399), .B2(n9802), .A(n9801), .ZN(P2_U3293) );
  INV_X1 U10856 ( .A(n9803), .ZN(n9805) );
  NOR2_X1 U10857 ( .A1(n9826), .A2(n9806), .ZN(P2_U3297) );
  INV_X1 U10858 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9807) );
  NOR2_X1 U10859 ( .A1(n9826), .A2(n9807), .ZN(P2_U3298) );
  INV_X1 U10860 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9808) );
  NOR2_X1 U10861 ( .A1(n9826), .A2(n9808), .ZN(P2_U3299) );
  INV_X1 U10862 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9809) );
  NOR2_X1 U10863 ( .A1(n9826), .A2(n9809), .ZN(P2_U3300) );
  INV_X1 U10864 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9810) );
  NOR2_X1 U10865 ( .A1(n9826), .A2(n9810), .ZN(P2_U3301) );
  INV_X1 U10866 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9811) );
  NOR2_X1 U10867 ( .A1(n9826), .A2(n9811), .ZN(P2_U3302) );
  INV_X1 U10868 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9812) );
  NOR2_X1 U10869 ( .A1(n9826), .A2(n9812), .ZN(P2_U3303) );
  INV_X1 U10870 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U10871 ( .A1(n9826), .A2(n9813), .ZN(P2_U3304) );
  INV_X1 U10872 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9814) );
  NOR2_X1 U10873 ( .A1(n9826), .A2(n9814), .ZN(P2_U3305) );
  INV_X1 U10874 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9815) );
  NOR2_X1 U10875 ( .A1(n9826), .A2(n9815), .ZN(P2_U3306) );
  INV_X1 U10876 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9816) );
  NOR2_X1 U10877 ( .A1(n9826), .A2(n9816), .ZN(P2_U3307) );
  INV_X1 U10878 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U10879 ( .A1(n9826), .A2(n9817), .ZN(P2_U3308) );
  INV_X1 U10880 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U10881 ( .A1(n9826), .A2(n9818), .ZN(P2_U3309) );
  INV_X1 U10882 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9819) );
  NOR2_X1 U10883 ( .A1(n9826), .A2(n9819), .ZN(P2_U3310) );
  INV_X1 U10884 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9820) );
  NOR2_X1 U10885 ( .A1(n9826), .A2(n9820), .ZN(P2_U3311) );
  INV_X1 U10886 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9821) );
  NOR2_X1 U10887 ( .A1(n9826), .A2(n9821), .ZN(P2_U3312) );
  NOR2_X1 U10888 ( .A1(n9826), .A2(n9822), .ZN(P2_U3313) );
  INV_X1 U10889 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U10890 ( .A1(n9826), .A2(n9823), .ZN(P2_U3314) );
  INV_X1 U10891 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U10892 ( .A1(n9826), .A2(n9824), .ZN(P2_U3315) );
  INV_X1 U10893 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9825) );
  NOR2_X1 U10894 ( .A1(n9826), .A2(n9825), .ZN(P2_U3316) );
  INV_X1 U10895 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9827) );
  NOR2_X1 U10896 ( .A1(n9826), .A2(n9827), .ZN(P2_U3317) );
  INV_X1 U10897 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U10898 ( .A1(n9826), .A2(n9828), .ZN(P2_U3318) );
  INV_X1 U10899 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9829) );
  NOR2_X1 U10900 ( .A1(n9826), .A2(n9829), .ZN(P2_U3319) );
  INV_X1 U10901 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U10902 ( .A1(n9826), .A2(n9830), .ZN(P2_U3320) );
  INV_X1 U10903 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9831) );
  NOR2_X1 U10904 ( .A1(n9826), .A2(n9831), .ZN(P2_U3321) );
  INV_X1 U10905 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9832) );
  NOR2_X1 U10906 ( .A1(n9826), .A2(n9832), .ZN(P2_U3322) );
  NOR2_X1 U10907 ( .A1(n9826), .A2(n9833), .ZN(P2_U3323) );
  INV_X1 U10908 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9834) );
  NOR2_X1 U10909 ( .A1(n9826), .A2(n9834), .ZN(P2_U3324) );
  INV_X1 U10910 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9835) );
  NOR2_X1 U10911 ( .A1(n9826), .A2(n9835), .ZN(P2_U3325) );
  NOR2_X1 U10912 ( .A1(n9826), .A2(n9836), .ZN(P2_U3326) );
  OAI22_X1 U10913 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9826), .B1(n9840), .B2(
        n9837), .ZN(n9838) );
  INV_X1 U10914 ( .A(n9838), .ZN(P2_U3437) );
  OAI22_X1 U10915 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9826), .B1(n9840), .B2(
        n9839), .ZN(n9841) );
  INV_X1 U10916 ( .A(n9841), .ZN(P2_U3438) );
  OAI21_X1 U10917 ( .B1(n9844), .B2(n9843), .A(n9842), .ZN(n9845) );
  AOI21_X1 U10918 ( .B1(n9907), .B2(n9846), .A(n9845), .ZN(n9912) );
  INV_X1 U10919 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9847) );
  AOI22_X1 U10920 ( .A1(n9910), .A2(n9912), .B1(n9847), .B2(n9908), .ZN(
        P2_U3451) );
  INV_X1 U10921 ( .A(n9848), .ZN(n9849) );
  OAI21_X1 U10922 ( .B1(n9850), .B2(n9900), .A(n9849), .ZN(n9851) );
  AOI211_X1 U10923 ( .C1(n9907), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9914)
         );
  INV_X1 U10924 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9854) );
  AOI22_X1 U10925 ( .A1(n9910), .A2(n9914), .B1(n9854), .B2(n9908), .ZN(
        P2_U3457) );
  OAI21_X1 U10926 ( .B1(n9856), .B2(n9900), .A(n9855), .ZN(n9858) );
  AOI211_X1 U10927 ( .C1(n9907), .C2(n9859), .A(n9858), .B(n9857), .ZN(n9915)
         );
  INV_X1 U10928 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9860) );
  AOI22_X1 U10929 ( .A1(n9910), .A2(n9915), .B1(n9860), .B2(n9908), .ZN(
        P2_U3466) );
  OAI22_X1 U10930 ( .A1(n9862), .A2(n9902), .B1(n9861), .B2(n9900), .ZN(n9864)
         );
  AOI211_X1 U10931 ( .C1(n9907), .C2(n9865), .A(n9864), .B(n9863), .ZN(n9916)
         );
  INV_X1 U10932 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9866) );
  AOI22_X1 U10933 ( .A1(n9910), .A2(n9916), .B1(n9866), .B2(n9908), .ZN(
        P2_U3469) );
  OAI211_X1 U10934 ( .C1(n9869), .C2(n9900), .A(n9868), .B(n9867), .ZN(n9870)
         );
  AOI21_X1 U10935 ( .B1(n9907), .B2(n9871), .A(n9870), .ZN(n9917) );
  AOI22_X1 U10936 ( .A1(n9910), .A2(n9917), .B1(n6019), .B2(n9908), .ZN(
        P2_U3472) );
  INV_X1 U10937 ( .A(n9872), .ZN(n9878) );
  INV_X1 U10938 ( .A(n9873), .ZN(n9874) );
  OAI22_X1 U10939 ( .A1(n9875), .A2(n9902), .B1(n9874), .B2(n9900), .ZN(n9877)
         );
  AOI211_X1 U10940 ( .C1(n9892), .C2(n9878), .A(n9877), .B(n9876), .ZN(n9919)
         );
  AOI22_X1 U10941 ( .A1(n9910), .A2(n9919), .B1(n9879), .B2(n9908), .ZN(
        P2_U3475) );
  INV_X1 U10942 ( .A(n9880), .ZN(n9885) );
  OAI22_X1 U10943 ( .A1(n9882), .A2(n9902), .B1(n9881), .B2(n9900), .ZN(n9884)
         );
  AOI211_X1 U10944 ( .C1(n9892), .C2(n9885), .A(n9884), .B(n9883), .ZN(n9921)
         );
  INV_X1 U10945 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9886) );
  AOI22_X1 U10946 ( .A1(n9910), .A2(n9921), .B1(n9886), .B2(n9908), .ZN(
        P2_U3478) );
  OAI22_X1 U10947 ( .A1(n9888), .A2(n9902), .B1(n9887), .B2(n9900), .ZN(n9890)
         );
  AOI211_X1 U10948 ( .C1(n9892), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9923)
         );
  INV_X1 U10949 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U10950 ( .A1(n9910), .A2(n9923), .B1(n9893), .B2(n9908), .ZN(
        P2_U3481) );
  OAI211_X1 U10951 ( .C1(n9896), .C2(n9900), .A(n9895), .B(n9894), .ZN(n9897)
         );
  AOI21_X1 U10952 ( .B1(n9898), .B2(n9907), .A(n9897), .ZN(n9924) );
  AOI22_X1 U10953 ( .A1(n9910), .A2(n9924), .B1(n9899), .B2(n9908), .ZN(
        P2_U3484) );
  OAI22_X1 U10954 ( .A1(n9903), .A2(n9902), .B1(n9901), .B2(n9900), .ZN(n9905)
         );
  AOI211_X1 U10955 ( .C1(n9907), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9926)
         );
  INV_X1 U10956 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U10957 ( .A1(n9910), .A2(n9926), .B1(n9909), .B2(n9908), .ZN(
        P2_U3487) );
  AOI22_X1 U10958 ( .A1(n9927), .A2(n9912), .B1(n9911), .B2(n9925), .ZN(
        P2_U3520) );
  AOI22_X1 U10959 ( .A1(n9927), .A2(n9914), .B1(n9913), .B2(n9925), .ZN(
        P2_U3522) );
  AOI22_X1 U10960 ( .A1(n9927), .A2(n9915), .B1(n5736), .B2(n9925), .ZN(
        P2_U3525) );
  AOI22_X1 U10961 ( .A1(n9927), .A2(n9916), .B1(n5824), .B2(n9925), .ZN(
        P2_U3526) );
  AOI22_X1 U10962 ( .A1(n9927), .A2(n9917), .B1(n5395), .B2(n9925), .ZN(
        P2_U3527) );
  AOI22_X1 U10963 ( .A1(n9927), .A2(n9919), .B1(n9918), .B2(n9925), .ZN(
        P2_U3528) );
  AOI22_X1 U10964 ( .A1(n9927), .A2(n9921), .B1(n9920), .B2(n9925), .ZN(
        P2_U3529) );
  AOI22_X1 U10965 ( .A1(n9927), .A2(n9923), .B1(n9922), .B2(n9925), .ZN(
        P2_U3530) );
  AOI22_X1 U10966 ( .A1(n9927), .A2(n9924), .B1(n6455), .B2(n9925), .ZN(
        P2_U3531) );
  AOI22_X1 U10967 ( .A1(n9927), .A2(n9926), .B1(n6497), .B2(n9925), .ZN(
        P2_U3532) );
  INV_X1 U10968 ( .A(n9928), .ZN(n9929) );
  NAND2_X1 U10969 ( .A1(n9930), .A2(n9929), .ZN(n9931) );
  XNOR2_X1 U10970 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9931), .ZN(ADD_1071_U5) );
  INV_X1 U10971 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9933) );
  AOI22_X1 U10972 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n9933), .B2(n9932), .ZN(ADD_1071_U46) );
  OAI21_X1 U10973 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(ADD_1071_U56) );
  OAI21_X1 U10974 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(ADD_1071_U57) );
  OAI21_X1 U10975 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(ADD_1071_U58) );
  OAI21_X1 U10976 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(ADD_1071_U59) );
  OAI21_X1 U10977 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(ADD_1071_U60) );
  OAI21_X1 U10978 ( .B1(n9951), .B2(n9950), .A(n9949), .ZN(ADD_1071_U61) );
  AOI21_X1 U10979 ( .B1(n9954), .B2(n9953), .A(n9952), .ZN(ADD_1071_U62) );
  AOI21_X1 U10980 ( .B1(n9957), .B2(n9956), .A(n9955), .ZN(ADD_1071_U63) );
  INV_X1 U10981 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9958) );
  XNOR2_X1 U10982 ( .A(n9959), .B(n9958), .ZN(ADD_1071_U48) );
  INV_X1 U10983 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9960) );
  XNOR2_X1 U10984 ( .A(n9961), .B(n9960), .ZN(ADD_1071_U50) );
  NOR2_X1 U10985 ( .A1(n9963), .A2(n9962), .ZN(n9964) );
  XOR2_X1 U10986 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9964), .Z(ADD_1071_U51) );
  INV_X1 U10987 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9965) );
  XNOR2_X1 U10988 ( .A(n9966), .B(n9965), .ZN(ADD_1071_U49) );
  OAI21_X1 U10989 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n9970) );
  XNOR2_X1 U10990 ( .A(n9970), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U10991 ( .B1(n9973), .B2(n9972), .A(n9971), .ZN(ADD_1071_U47) );
  XOR2_X1 U10992 ( .A(n9975), .B(n9974), .Z(ADD_1071_U54) );
  XOR2_X1 U10993 ( .A(n9977), .B(n9976), .Z(ADD_1071_U53) );
  XNOR2_X1 U10994 ( .A(n9979), .B(n9978), .ZN(ADD_1071_U52) );
  OR2_X2 U4821 ( .A1(n5219), .A2(n5218), .ZN(n9646) );
  INV_X1 U4816 ( .A(n7318), .ZN(n7290) );
  NAND2_X2 U4804 ( .A1(n8917), .A2(n6260), .ZN(n5281) );
  CLKBUF_X1 U4817 ( .A(n8550), .Z(n8551) );
  CLKBUF_X1 U4822 ( .A(n7318), .Z(n7283) );
  CLKBUF_X1 U4823 ( .A(n6027), .Z(n7517) );
  NAND2_X2 U4852 ( .A1(n8009), .A2(n5310), .ZN(n5466) );
  NAND3_X1 U4946 ( .A1(n8658), .A2(n8662), .A3(n4714), .ZN(n8591) );
  NAND2_X1 U9963 ( .A1(n8591), .A2(n7241), .ZN(n8600) );
endmodule

