

module b22_C_SARLock_k_64_7 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150;

  NAND2_X1 U7195 ( .A1(n7934), .A2(n7933), .ZN(n13320) );
  OAI22_X1 U7196 ( .A1(n11500), .A2(n6793), .B1(n11728), .B2(n6794), .ZN(
        n11735) );
  INV_X2 U7197 ( .A(n12834), .ZN(n6452) );
  INV_X2 U7198 ( .A(n11904), .ZN(n11834) );
  INV_X1 U7199 ( .A(n6451), .ZN(n13756) );
  INV_X1 U7200 ( .A(n10638), .ZN(n12381) );
  INV_X1 U7201 ( .A(n10466), .ZN(n12382) );
  NAND4_X2 U7203 ( .A1(n10241), .A2(n10240), .A3(n10239), .A4(n10238), .ZN(
        n14646) );
  CLKBUF_X1 U7204 ( .A(n7506), .Z(n8081) );
  INV_X1 U7205 ( .A(n12760), .ZN(n12383) );
  INV_X1 U7206 ( .A(n10532), .ZN(n13730) );
  INV_X2 U7207 ( .A(n9152), .ZN(n8080) );
  OAI211_X1 U7208 ( .C1(n10229), .C2(n9712), .A(n9711), .B(n9710), .ZN(n14734)
         );
  AND2_X2 U7209 ( .A1(n7472), .A2(n7471), .ZN(n7486) );
  INV_X1 U7210 ( .A(n10393), .ZN(n11810) );
  NAND2_X1 U7211 ( .A1(n12652), .A2(n8663), .ZN(n12638) );
  INV_X2 U7212 ( .A(n12915), .ZN(n12873) );
  OR2_X1 U7213 ( .A1(n13189), .A2(n13176), .ZN(n13174) );
  NOR2_X2 U7214 ( .A1(n7728), .A2(n7727), .ZN(n7749) );
  CLKBUF_X2 U7215 ( .A(n11842), .Z(n6459) );
  INV_X1 U7217 ( .A(n9970), .ZN(n9733) );
  INV_X1 U7219 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8361) );
  AND2_X2 U7220 ( .A1(n8158), .A2(n8104), .ZN(n8159) );
  INV_X2 U7221 ( .A(n7487), .ZN(n9148) );
  NAND2_X1 U7222 ( .A1(n7921), .A2(n7920), .ZN(n13176) );
  NAND2_X1 U7223 ( .A1(n9441), .A2(n11772), .ZN(n11895) );
  INV_X1 U7224 ( .A(n10532), .ZN(n12051) );
  INV_X1 U7225 ( .A(n14080), .ZN(n14212) );
  INV_X2 U7227 ( .A(n6452), .ZN(n13217) );
  BUF_X1 U7228 ( .A(n7964), .Z(n6463) );
  OR2_X1 U7230 ( .A1(n14280), .A2(n9400), .ZN(n9667) );
  NAND2_X1 U7231 ( .A1(n14273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9573) );
  XNOR2_X1 U7232 ( .A(n9432), .B(n9431), .ZN(n9561) );
  AOI21_X1 U7233 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n14375), .A(n14442), .ZN(
        n14391) );
  INV_X1 U7234 ( .A(n12564), .ZN(n7018) );
  INV_X1 U7235 ( .A(n10776), .ZN(n12380) );
  NAND4_X1 U7236 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n13844) );
  NOR2_X1 U7237 ( .A1(n13982), .A2(n13981), .ZN(n7436) );
  INV_X1 U7238 ( .A(n10743), .ZN(n6885) );
  AND2_X1 U7239 ( .A1(n9440), .A2(n9439), .ZN(n6446) );
  OR2_X2 U7240 ( .A1(n7169), .A2(n7172), .ZN(n7166) );
  OR2_X2 U7241 ( .A1(n12773), .A2(n12525), .ZN(n8766) );
  OAI21_X2 U7242 ( .B1(n7019), .B2(n8952), .A(n9730), .ZN(n8955) );
  OAI22_X2 U7243 ( .A1(n8761), .A2(n8760), .B1(P1_DATAO_REG_30__SCAN_IN), .B2(
        n12234), .ZN(n8749) );
  OR2_X2 U7244 ( .A1(n8109), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8110) );
  OAI21_X2 U7245 ( .B1(n12011), .B2(n14128), .A(n12010), .ZN(n14113) );
  NAND2_X2 U7246 ( .A1(n6832), .A2(n7077), .ZN(n11681) );
  NAND2_X1 U7247 ( .A1(n9265), .A2(n12769), .ZN(n9267) );
  NOR2_X2 U7248 ( .A1(n14366), .A2(n14365), .ZN(n14622) );
  XNOR2_X2 U7249 ( .A(n7842), .B(SI_20_), .ZN(n7840) );
  NAND2_X2 U7250 ( .A1(n7466), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7467) );
  NAND4_X2 U7251 ( .A1(n7492), .A2(n7491), .A3(n7490), .A4(n7489), .ZN(n8973)
         );
  OR2_X1 U7252 ( .A1(n6458), .A2(n9476), .ZN(n9710) );
  NOR2_X2 U7253 ( .A1(n12239), .A2(n12003), .ZN(n8198) );
  OAI21_X2 U7254 ( .B1(n14504), .B2(n7720), .A(n7719), .ZN(n11671) );
  INV_X4 U7255 ( .A(n13587), .ZN(n13768) );
  NAND2_X4 U7256 ( .A1(n7165), .A2(n13736), .ZN(n13587) );
  OAI22_X2 U7257 ( .A1(n14333), .A2(n14335), .B1(P1_ADDR_REG_1__SCAN_IN), .B2(
        n9782), .ZN(n7340) );
  NAND2_X1 U7258 ( .A1(n8795), .A2(n8794), .ZN(n10186) );
  NOR2_X1 U7259 ( .A1(n12239), .A2(n12003), .ZN(n6447) );
  NOR2_X1 U7260 ( .A1(n12239), .A2(n12003), .ZN(n6448) );
  NOR2_X2 U7261 ( .A1(n14337), .A2(n15148), .ZN(n14400) );
  INV_X4 U7262 ( .A(n8288), .ZN(n8762) );
  OAI21_X2 U7263 ( .B1(n8455), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n6771) );
  NOR2_X2 U7264 ( .A1(n10481), .A2(n10480), .ZN(n14771) );
  NOR2_X1 U7265 ( .A1(n8159), .A2(n8160), .ZN(n10014) );
  XNOR2_X2 U7266 ( .A(n8477), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n8476) );
  OAI21_X2 U7267 ( .B1(n8494), .B2(n8493), .A(n8495), .ZN(n8507) );
  NAND2_X2 U7268 ( .A1(n8479), .A2(n8478), .ZN(n8494) );
  AND4_X2 U7269 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), .ZN(n10466)
         );
  AOI21_X2 U7270 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14338), .A(n14399), .ZN(
        n15146) );
  NAND2_X1 U7271 ( .A1(n12937), .A2(n6999), .ZN(n13012) );
  NAND2_X1 U7272 ( .A1(n9147), .A2(n9146), .ZN(n13138) );
  AND2_X1 U7273 ( .A1(n12664), .A2(n8662), .ZN(n12653) );
  NAND2_X1 U7274 ( .A1(n13525), .A2(n13524), .ZN(n13523) );
  INV_X1 U7275 ( .A(n13193), .ZN(n8036) );
  OAI21_X1 U7276 ( .B1(n8076), .B2(n8075), .A(n8074), .ZN(n9136) );
  OR2_X1 U7277 ( .A1(n14212), .A2(n14086), .ZN(n14075) );
  NAND2_X1 U7278 ( .A1(n7200), .A2(n6534), .ZN(n12011) );
  NAND2_X1 U7279 ( .A1(n8655), .A2(n8654), .ZN(n11441) );
  XNOR2_X1 U7280 ( .A(n7897), .B(n12181), .ZN(n7896) );
  NAND2_X1 U7281 ( .A1(n7884), .A2(n7883), .ZN(n7897) );
  OAI21_X1 U7282 ( .B1(n11893), .B2(n7242), .A(n7866), .ZN(n7881) );
  NAND2_X1 U7283 ( .A1(n7845), .A2(n7844), .ZN(n13425) );
  XNOR2_X1 U7284 ( .A(n7865), .B(SI_22_), .ZN(n11893) );
  NAND2_X1 U7285 ( .A1(n7829), .A2(n7828), .ZN(n13367) );
  NAND2_X1 U7286 ( .A1(n7115), .A2(n7114), .ZN(n7113) );
  AND2_X1 U7287 ( .A1(n6849), .A2(n10722), .ZN(n10764) );
  NAND2_X1 U7288 ( .A1(n8805), .A2(n8806), .ZN(n10131) );
  INV_X1 U7289 ( .A(n13844), .ZN(n10623) );
  NAND2_X1 U7290 ( .A1(n10638), .A2(n10199), .ZN(n8806) );
  NAND2_X2 U7291 ( .A1(n8791), .A2(n9267), .ZN(n12765) );
  INV_X1 U7292 ( .A(n10831), .ZN(n10839) );
  INV_X1 U7293 ( .A(n13601), .ZN(n14768) );
  NOR2_X1 U7294 ( .A1(n15045), .A2(n10474), .ZN(n15044) );
  NAND4_X1 U7295 ( .A1(n7558), .A2(n7557), .A3(n7556), .A4(n7555), .ZN(n13044)
         );
  NAND4_X1 U7296 ( .A1(n7543), .A2(n7542), .A3(n7541), .A4(n7540), .ZN(n13045)
         );
  CLKBUF_X3 U7298 ( .A(n9713), .Z(n12222) );
  INV_X4 U7299 ( .A(n11904), .ZN(n11966) );
  INV_X1 U7300 ( .A(n14734), .ZN(n6664) );
  NAND2_X2 U7301 ( .A1(n8121), .A2(n12003), .ZN(n8163) );
  NAND2_X2 U7302 ( .A1(n12833), .A2(n12476), .ZN(n9734) );
  INV_X1 U7303 ( .A(n11895), .ZN(n11842) );
  AND2_X1 U7304 ( .A1(n9564), .A2(n13738), .ZN(n10547) );
  INV_X1 U7305 ( .A(n14155), .ZN(n13568) );
  XNOR2_X1 U7306 ( .A(n9435), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9564) );
  INV_X8 U7307 ( .A(n8134), .ZN(n9139) );
  INV_X2 U7308 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U7309 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8145) );
  OAI211_X1 U7310 ( .C1(n14177), .C2(n14769), .A(n6543), .B(n7436), .ZN(n14258) );
  NAND2_X1 U7311 ( .A1(n6611), .A2(n13985), .ZN(n14177) );
  AND2_X1 U7312 ( .A1(n12542), .A2(n6497), .ZN(n7169) );
  AOI21_X1 U7313 ( .B1(n6535), .B2(n6617), .A(n6616), .ZN(n13148) );
  AND2_X1 U7314 ( .A1(n6646), .A2(n13151), .ZN(n6645) );
  NAND2_X1 U7315 ( .A1(n8592), .A2(n8591), .ZN(n12544) );
  AND2_X1 U7316 ( .A1(n8026), .A2(n8025), .ZN(n8073) );
  OAI21_X1 U7317 ( .B1(n14166), .B2(n14126), .A(n12063), .ZN(n12064) );
  OR2_X1 U7318 ( .A1(n13157), .A2(n14530), .ZN(n6646) );
  AND2_X1 U7319 ( .A1(n13755), .A2(n7131), .ZN(n7130) );
  NAND2_X1 U7320 ( .A1(n9324), .A2(n9326), .ZN(n12320) );
  MUX2_X1 U7321 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n12216), .S(n15002), .Z(
        n11988) );
  AOI21_X1 U7322 ( .B1(n7356), .B2(n7358), .A(n6538), .ZN(n7355) );
  XNOR2_X1 U7323 ( .A(n12045), .B(n12044), .ZN(n14166) );
  AOI211_X1 U7324 ( .C1(n14182), .C2(n14784), .A(n14181), .B(n14180), .ZN(
        n14183) );
  AND2_X1 U7325 ( .A1(n6633), .A2(n6631), .ZN(n7134) );
  OAI21_X1 U7326 ( .B1(n8599), .B2(n8598), .A(n8601), .ZN(n8747) );
  AND2_X1 U7327 ( .A1(n12221), .A2(n7357), .ZN(n7356) );
  OR2_X1 U7328 ( .A1(n11986), .A2(n13217), .ZN(n13141) );
  NAND2_X1 U7329 ( .A1(n8021), .A2(n8020), .ZN(n13159) );
  NAND2_X1 U7330 ( .A1(n8559), .A2(n8558), .ZN(n9340) );
  NAND2_X1 U7331 ( .A1(n13012), .A2(n12888), .ZN(n12914) );
  XNOR2_X1 U7332 ( .A(n6684), .B(n10984), .ZN(n9248) );
  NAND2_X1 U7333 ( .A1(n8540), .A2(n8539), .ZN(n12709) );
  NAND2_X1 U7334 ( .A1(n6905), .A2(n6903), .ZN(n13317) );
  NAND2_X1 U7335 ( .A1(n8019), .A2(n8018), .ZN(n13182) );
  AND2_X1 U7336 ( .A1(n13747), .A2(n13746), .ZN(n13752) );
  NAND2_X1 U7337 ( .A1(n14012), .A2(n14011), .ZN(n14010) );
  NAND2_X1 U7338 ( .A1(n12297), .A2(n12607), .ZN(n12579) );
  OAI21_X1 U7339 ( .B1(n8570), .B2(n8569), .A(n8571), .ZN(n8588) );
  NAND2_X1 U7340 ( .A1(n12939), .A2(n12938), .ZN(n12937) );
  NAND2_X1 U7341 ( .A1(n12968), .A2(n12872), .ZN(n12939) );
  AOI21_X1 U7342 ( .B1(n7220), .B2(n14004), .A(n6525), .ZN(n7218) );
  NAND2_X1 U7343 ( .A1(n6943), .A2(n6946), .ZN(n14012) );
  XNOR2_X1 U7344 ( .A(n13138), .B(n13021), .ZN(n9247) );
  OAI21_X1 U7345 ( .B1(n13727), .B2(n6451), .A(n13729), .ZN(n13973) );
  OR2_X1 U7346 ( .A1(n12966), .A2(n12967), .ZN(n12968) );
  OAI21_X2 U7347 ( .B1(n13727), .B2(n7493), .A(n9190), .ZN(n13408) );
  AOI21_X1 U7348 ( .B1(n7364), .B2(n6783), .A(n6782), .ZN(n6781) );
  NAND2_X1 U7349 ( .A1(n14071), .A2(n12015), .ZN(n14051) );
  AND2_X1 U7350 ( .A1(n8100), .A2(n7958), .ZN(n9243) );
  NAND2_X1 U7351 ( .A1(n6670), .A2(n9189), .ZN(n13727) );
  AND2_X1 U7352 ( .A1(n9317), .A2(n12268), .ZN(n9318) );
  NOR2_X2 U7353 ( .A1(n13174), .A2(n13320), .ZN(n13163) );
  NAND2_X1 U7354 ( .A1(n13207), .A2(n7894), .ZN(n13185) );
  INV_X1 U7355 ( .A(n12924), .ZN(n13413) );
  NAND2_X1 U7356 ( .A1(n13523), .A2(n6528), .ZN(n13489) );
  INV_X1 U7357 ( .A(n14169), .ZN(n13742) );
  NAND2_X1 U7358 ( .A1(n8451), .A2(n8933), .ZN(n12670) );
  NAND2_X1 U7359 ( .A1(n7027), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7026) );
  NAND2_X1 U7360 ( .A1(n7205), .A2(n7204), .ZN(n14074) );
  AOI21_X1 U7361 ( .B1(n12034), .B2(n13756), .A(n6602), .ZN(n14169) );
  NAND2_X2 U7362 ( .A1(n12023), .A2(n12022), .ZN(n14174) );
  AND2_X1 U7363 ( .A1(n6948), .A2(n14035), .ZN(n12016) );
  XNOR2_X1 U7364 ( .A(n13998), .B(n12228), .ZN(n13995) );
  AND2_X1 U7365 ( .A1(n14025), .A2(n6950), .ZN(n6949) );
  XNOR2_X1 U7366 ( .A(n9144), .B(n9143), .ZN(n13757) );
  NAND2_X1 U7367 ( .A1(n7951), .A2(n7950), .ZN(n12924) );
  AND2_X1 U7368 ( .A1(n9316), .A2(n9315), .ZN(n12268) );
  OR2_X1 U7369 ( .A1(n9312), .A2(n12307), .ZN(n9316) );
  XNOR2_X1 U7370 ( .A(n14029), .B(n13824), .ZN(n14025) );
  NAND2_X2 U7371 ( .A1(n11958), .A2(n11957), .ZN(n13717) );
  NAND2_X1 U7372 ( .A1(n8510), .A2(n8509), .ZN(n12610) );
  NAND2_X1 U7373 ( .A1(n6705), .A2(n6703), .ZN(n13231) );
  NAND2_X1 U7374 ( .A1(n11777), .A2(n11776), .ZN(n13998) );
  OAI21_X1 U7375 ( .B1(n12928), .B2(n6970), .A(n6968), .ZN(n12867) );
  XNOR2_X1 U7376 ( .A(n9136), .B(n9135), .ZN(n12034) );
  OAI21_X1 U7377 ( .B1(n9136), .B2(n7274), .A(n7271), .ZN(n9144) );
  NAND2_X1 U7378 ( .A1(n12021), .A2(n13756), .ZN(n12023) );
  NAND2_X1 U7379 ( .A1(n6804), .A2(n6521), .ZN(n13481) );
  CLKBUF_X1 U7380 ( .A(n13339), .Z(n6644) );
  NOR2_X1 U7381 ( .A1(n13339), .A2(n6869), .ZN(n6868) );
  XNOR2_X1 U7382 ( .A(n8076), .B(n8075), .ZN(n12021) );
  NAND2_X1 U7383 ( .A1(n7887), .A2(n7886), .ZN(n13339) );
  XNOR2_X1 U7384 ( .A(n7946), .B(n7941), .ZN(n11775) );
  NAND2_X1 U7385 ( .A1(n13509), .A2(n7361), .ZN(n6804) );
  XNOR2_X1 U7386 ( .A(n7931), .B(n7930), .ZN(n13457) );
  XNOR2_X1 U7387 ( .A(n7885), .B(n7895), .ZN(n13465) );
  AOI21_X1 U7388 ( .B1(n14636), .B2(n7333), .A(n7332), .ZN(n7331) );
  NAND2_X1 U7389 ( .A1(n6712), .A2(n6894), .ZN(n13290) );
  NAND2_X1 U7390 ( .A1(n8469), .A2(n8468), .ZN(n12646) );
  AOI21_X1 U7391 ( .B1(n7094), .B2(n8009), .A(n6507), .ZN(n7093) );
  AND2_X1 U7392 ( .A1(n7898), .A2(n7270), .ZN(n7269) );
  NOR2_X1 U7393 ( .A1(n14571), .A2(n14570), .ZN(n11812) );
  NOR2_X1 U7394 ( .A1(n13261), .A2(n13425), .ZN(n13248) );
  NAND2_X1 U7395 ( .A1(n7896), .A2(n7895), .ZN(n7899) );
  NAND2_X1 U7396 ( .A1(n11913), .A2(n11912), .ZN(n14059) );
  AND2_X1 U7397 ( .A1(n11807), .A2(n11806), .ZN(n14571) );
  NAND2_X1 U7398 ( .A1(n11703), .A2(n11702), .ZN(n12007) );
  NAND2_X1 U7399 ( .A1(n7868), .A2(n7867), .ZN(n13345) );
  OR2_X1 U7400 ( .A1(n13277), .A2(n8008), .ZN(n8009) );
  NAND2_X1 U7401 ( .A1(n8435), .A2(n8434), .ZN(n8438) );
  NOR2_X1 U7402 ( .A1(n6480), .A2(n14369), .ZN(n14629) );
  OAI22_X1 U7403 ( .A1(n11758), .A2(n11757), .B1(n11756), .B2(n11755), .ZN(
        n14486) );
  AOI21_X1 U7404 ( .B1(n7215), .B2(n7214), .A(n6477), .ZN(n7213) );
  AOI21_X1 U7405 ( .B1(n7079), .B2(n7081), .A(n6530), .ZN(n7077) );
  XNOR2_X1 U7406 ( .A(n7804), .B(n7803), .ZN(n11841) );
  NAND2_X1 U7407 ( .A1(n11406), .A2(n8837), .ZN(n11331) );
  NAND2_X1 U7408 ( .A1(n11223), .A2(n11222), .ZN(n11381) );
  OR2_X2 U7409 ( .A1(n11338), .A2(n11337), .ZN(n11339) );
  NAND2_X1 U7410 ( .A1(n11828), .A2(n11827), .ZN(n14238) );
  NAND2_X1 U7411 ( .A1(n11221), .A2(n11220), .ZN(n11223) );
  NAND2_X1 U7412 ( .A1(n7014), .A2(n8410), .ZN(n8433) );
  NAND2_X1 U7413 ( .A1(n7790), .A2(n7789), .ZN(n13435) );
  NAND2_X1 U7414 ( .A1(n11474), .A2(n9232), .ZN(n7995) );
  NAND2_X2 U7415 ( .A1(n7772), .A2(n7771), .ZN(n13439) );
  NAND2_X1 U7416 ( .A1(n11496), .A2(n6790), .ZN(n11502) );
  XNOR2_X1 U7417 ( .A(n7820), .B(SI_18_), .ZN(n7799) );
  OR2_X1 U7418 ( .A1(n6788), .A2(n6787), .ZN(n11496) );
  NAND2_X1 U7419 ( .A1(n7236), .A2(n7783), .ZN(n7820) );
  OR2_X1 U7420 ( .A1(n14600), .A2(n11789), .ZN(n13664) );
  NAND2_X1 U7421 ( .A1(n7752), .A2(n7751), .ZN(n13399) );
  NAND2_X1 U7422 ( .A1(n10805), .A2(n7088), .ZN(n10804) );
  NAND2_X1 U7423 ( .A1(n7711), .A2(n7710), .ZN(n14503) );
  NAND2_X1 U7424 ( .A1(n7731), .A2(n7730), .ZN(n11767) );
  NAND2_X1 U7425 ( .A1(n10811), .A2(n8820), .ZN(n11040) );
  NAND2_X1 U7426 ( .A1(n7767), .A2(n7240), .ZN(n7236) );
  NAND2_X1 U7427 ( .A1(n11526), .A2(n11525), .ZN(n14600) );
  NAND2_X1 U7428 ( .A1(n7371), .A2(n7368), .ZN(n11348) );
  NAND2_X1 U7429 ( .A1(n7765), .A2(n7764), .ZN(n7767) );
  NAND2_X1 U7430 ( .A1(n7671), .A2(n7670), .ZN(n11565) );
  NAND2_X1 U7431 ( .A1(n11218), .A2(n11217), .ZN(n14564) );
  NAND2_X1 U7432 ( .A1(n7654), .A2(n7653), .ZN(n11467) );
  NAND2_X1 U7433 ( .A1(n7677), .A2(n7427), .ZN(n7679) );
  AND2_X1 U7434 ( .A1(n10966), .A2(n7087), .ZN(n7086) );
  NAND2_X1 U7435 ( .A1(n6848), .A2(n6847), .ZN(n11061) );
  INV_X2 U7436 ( .A(n15117), .ZN(n15119) );
  INV_X2 U7437 ( .A(n14991), .ZN(n10105) );
  BUF_X4 U7438 ( .A(n9203), .Z(n6462) );
  BUF_X4 U7439 ( .A(n9203), .Z(n6461) );
  NAND2_X1 U7440 ( .A1(n7597), .A2(n7596), .ZN(n11173) );
  AND2_X2 U7441 ( .A1(n8091), .A2(n13295), .ZN(n14951) );
  AND2_X1 U7442 ( .A1(n8802), .A2(n8801), .ZN(n10084) );
  INV_X1 U7443 ( .A(n10742), .ZN(n13046) );
  INV_X1 U7444 ( .A(n10475), .ZN(n10639) );
  AND2_X2 U7445 ( .A1(n7036), .A2(n10114), .ZN(n12764) );
  OAI211_X1 U7446 ( .C1(n9803), .C2(n13071), .A(n7104), .B(n7566), .ZN(n10855)
         );
  NOR2_X1 U7447 ( .A1(n15044), .A2(n7123), .ZN(n10022) );
  AND3_X1 U7448 ( .A1(n8197), .A2(n8196), .A3(n8195), .ZN(n10199) );
  OAI211_X1 U7449 ( .C1(n6449), .C2(n9500), .A(n8218), .B(n8217), .ZN(n10475)
         );
  AND2_X1 U7450 ( .A1(n6513), .A2(n7523), .ZN(n10742) );
  NAND2_X1 U7451 ( .A1(n7035), .A2(n8138), .ZN(n10114) );
  INV_X1 U7452 ( .A(n11311), .ZN(n8957) );
  OR2_X1 U7453 ( .A1(n10234), .A2(n10233), .ZN(n13601) );
  AND3_X1 U7454 ( .A1(n8180), .A2(n8179), .A3(n8178), .ZN(n10091) );
  NAND2_X1 U7455 ( .A1(n7504), .A2(n7503), .ZN(n10321) );
  INV_X2 U7456 ( .A(n11866), .ZN(n12027) );
  INV_X2 U7457 ( .A(n13542), .ZN(n13551) );
  AND2_X1 U7458 ( .A1(n13584), .A2(n9667), .ZN(n9713) );
  CLKBUF_X3 U7459 ( .A(n8182), .Z(n8756) );
  INV_X1 U7460 ( .A(n9910), .ZN(n11904) );
  INV_X1 U7461 ( .A(n10547), .ZN(n13584) );
  INV_X2 U7462 ( .A(n9734), .ZN(n8457) );
  NAND2_X1 U7463 ( .A1(n9803), .A2(n9139), .ZN(n7493) );
  INV_X1 U7464 ( .A(n7472), .ZN(n12215) );
  NAND2_X1 U7465 ( .A1(n7528), .A2(n7527), .ZN(n7069) );
  NAND2_X4 U7466 ( .A1(n13455), .A2(n8027), .ZN(n9803) );
  XNOR2_X1 U7467 ( .A(n7465), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7472) );
  INV_X1 U7468 ( .A(n11770), .ZN(n9574) );
  NAND2_X1 U7469 ( .A1(n7455), .A2(n7454), .ZN(n13455) );
  MUX2_X1 U7470 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7453), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n7455) );
  OAI21_X1 U7471 ( .B1(n14339), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6554), .ZN(
        n7339) );
  NAND2_X1 U7472 ( .A1(n9434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9435) );
  OR2_X1 U7473 ( .A1(n13443), .A2(n13444), .ZN(n7465) );
  NAND2_X1 U7474 ( .A1(n9430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9432) );
  MUX2_X1 U7475 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9570), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n9571) );
  XNOR2_X1 U7476 ( .A(n9397), .B(n9396), .ZN(n14281) );
  XNOR2_X1 U7477 ( .A(n14294), .B(n14293), .ZN(n14339) );
  AOI21_X1 U7478 ( .B1(n7547), .B2(n6843), .A(n6555), .ZN(n6842) );
  NAND2_X1 U7479 ( .A1(n8133), .A2(n8132), .ZN(n12476) );
  AND2_X1 U7480 ( .A1(n9540), .A2(n7342), .ZN(n9433) );
  AND2_X1 U7481 ( .A1(n8413), .A2(n8412), .ZN(n8417) );
  INV_X2 U7482 ( .A(n13451), .ZN(n13458) );
  OR2_X1 U7483 ( .A1(n7435), .A2(n9439), .ZN(n6655) );
  AND2_X1 U7484 ( .A1(n8396), .A2(n8395), .ZN(n8413) );
  INV_X2 U7485 ( .A(n14275), .ZN(n6454) );
  OAI21_X1 U7486 ( .B1(n9427), .B2(n9426), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9429) );
  NAND2_X2 U7487 ( .A1(n9139), .A2(P3_U3151), .ZN(n12829) );
  NOR2_X2 U7488 ( .A1(n8343), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8396) );
  AND3_X1 U7489 ( .A1(n9385), .A2(n7223), .A3(n10173), .ZN(n9440) );
  NAND2_X2 U7490 ( .A1(n8134), .A2(P1_U3086), .ZN(n14286) );
  XNOR2_X1 U7491 ( .A(n7549), .B(SI_4_), .ZN(n7547) );
  INV_X2 U7492 ( .A(n9582), .ZN(n8134) );
  NOR2_X1 U7493 ( .A1(n7559), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7668) );
  AND2_X1 U7494 ( .A1(n7417), .A2(n7450), .ZN(n7416) );
  NOR2_X1 U7495 ( .A1(n9392), .A2(n9391), .ZN(n9393) );
  AND2_X2 U7496 ( .A1(n7100), .A2(n7099), .ZN(n9582) );
  NAND4_X1 U7497 ( .A1(n13137), .A2(n13966), .A3(n7103), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7100) );
  AND2_X1 U7498 ( .A1(n7445), .A2(n7962), .ZN(n6902) );
  AND2_X1 U7499 ( .A1(n7449), .A2(n8048), .ZN(n7417) );
  NAND2_X1 U7500 ( .A1(n8135), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8154) );
  INV_X4 U7501 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7502 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9532) );
  INV_X1 U7503 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13966) );
  INV_X1 U7504 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9595) );
  INV_X1 U7505 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13137) );
  XNOR2_X1 U7506 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8155) );
  INV_X1 U7507 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9905) );
  INV_X1 U7508 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10096) );
  INV_X1 U7509 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7545) );
  INV_X1 U7510 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7445) );
  INV_X1 U7511 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9402) );
  NOR2_X1 U7512 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7444) );
  INV_X1 U7513 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8440) );
  NOR2_X1 U7514 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9378) );
  INV_X4 U7515 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U7516 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7517 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9431) );
  INV_X1 U7518 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8048) );
  INV_X1 U7519 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7449) );
  NAND2_X1 U7520 ( .A1(n13315), .A2(n6845), .ZN(n13410) );
  INV_X2 U7521 ( .A(n8120), .ZN(n12003) );
  NAND2_X2 U7522 ( .A1(n13489), .A2(n11892), .ZN(n13533) );
  INV_X1 U7523 ( .A(n10121), .ZN(n10374) );
  NOR2_X1 U7524 ( .A1(n11135), .A2(n11134), .ZN(n12386) );
  NAND2_X1 U7525 ( .A1(n11012), .A2(n13787), .ZN(n11118) );
  CLKBUF_X1 U7526 ( .A(n9441), .Z(n6455) );
  XNOR2_X1 U7527 ( .A(n9429), .B(n9428), .ZN(n9441) );
  AND2_X2 U7528 ( .A1(n9575), .A2(n11770), .ZN(n10235) );
  INV_X2 U7529 ( .A(n7471), .ZN(n7468) );
  INV_X1 U7530 ( .A(n11961), .ZN(n11866) );
  AND2_X4 U7531 ( .A1(n7472), .A2(n7468), .ZN(n7506) );
  CLKBUF_X2 U7532 ( .A(n14656), .Z(n6457) );
  OAI211_X1 U7533 ( .C1(n6451), .C2(n10228), .A(n10227), .B(n10226), .ZN(
        n14656) );
  NAND2_X2 U7534 ( .A1(n12517), .A2(n10371), .ZN(n9353) );
  INV_X4 U7535 ( .A(n8676), .ZN(n8606) );
  BUF_X8 U7536 ( .A(n13587), .Z(n13607) );
  INV_X4 U7537 ( .A(n8557), .ZN(n8243) );
  NAND2_X1 U7538 ( .A1(n9734), .A2(n8134), .ZN(n8557) );
  AND2_X2 U7539 ( .A1(n9575), .A2(n9574), .ZN(n11961) );
  XNOR2_X1 U7540 ( .A(n12484), .B(n14451), .ZN(n14447) );
  NAND2_X1 U7541 ( .A1(n9441), .A2(n11772), .ZN(n6458) );
  OAI21_X2 U7542 ( .B1(n8322), .B2(n8321), .A(n8323), .ZN(n8340) );
  OR2_X1 U7543 ( .A1(n14051), .A2(n14056), .ZN(n14034) );
  NOR2_X4 U7544 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7497) );
  AND3_X1 U7545 ( .A1(n9724), .A2(n9725), .A3(n9723), .ZN(n6512) );
  NAND2_X1 U7546 ( .A1(n7471), .A2(n12215), .ZN(n9152) );
  XNOR2_X2 U7547 ( .A(n7467), .B(P2_IR_REG_29__SCAN_IN), .ZN(n7471) );
  NAND2_X2 U7548 ( .A1(n12020), .A2(n12019), .ZN(n13996) );
  NAND2_X2 U7549 ( .A1(n6665), .A2(n6664), .ZN(n10258) );
  INV_X2 U7550 ( .A(n11109), .ZN(n12050) );
  OR2_X1 U7551 ( .A1(n9427), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n9395) );
  OAI211_X1 U7552 ( .C1(n10229), .C2(n9913), .A(n9912), .B(n9911), .ZN(n13581)
         );
  NAND2_X1 U7553 ( .A1(n11895), .A2(n8134), .ZN(n10229) );
  XNOR2_X2 U7554 ( .A(n10121), .B(n13048), .ZN(n10162) );
  OAI211_X2 U7555 ( .C1(n9803), .C2(n9815), .A(n7462), .B(n7461), .ZN(n10121)
         );
  AOI211_X1 U7556 ( .C1(n9250), .C2(n7968), .A(n9249), .B(n9248), .ZN(n9251)
         );
  OAI22_X2 U7557 ( .A1(n11701), .A2(n11700), .B1(n13834), .B2(n11799), .ZN(
        n11703) );
  AOI21_X2 U7558 ( .B1(n10589), .B2(n13780), .A(n6553), .ZN(n10713) );
  NOR2_X2 U7559 ( .A1(n14771), .A2(n10259), .ZN(n10589) );
  INV_X2 U7561 ( .A(n8981), .ZN(n9203) );
  INV_X2 U7562 ( .A(n9088), .ZN(n9126) );
  INV_X2 U7563 ( .A(n8981), .ZN(n9088) );
  NAND2_X1 U7564 ( .A1(n13048), .A2(n9203), .ZN(n8967) );
  AOI22_X1 U7565 ( .A1(n13048), .A2(n9126), .B1(n10121), .B2(n9088), .ZN(n8969) );
  OR2_X1 U7566 ( .A1(n12297), .A2(n12607), .ZN(n8780) );
  NAND2_X1 U7567 ( .A1(n7194), .A2(n7193), .ZN(n7192) );
  INV_X1 U7568 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U7569 ( .A1(n8078), .A2(n8077), .ZN(n13313) );
  NAND2_X1 U7570 ( .A1(n12034), .A2(n7612), .ZN(n8078) );
  NOR2_X1 U7571 ( .A1(n13717), .A2(n6861), .ZN(n6860) );
  OR2_X1 U7572 ( .A1(n14238), .A2(n12009), .ZN(n12038) );
  NOR2_X1 U7573 ( .A1(n9341), .A2(n12578), .ZN(n9342) );
  NAND2_X1 U7574 ( .A1(n8791), .A2(n12764), .ZN(n9262) );
  OR2_X1 U7575 ( .A1(n12739), .A2(n12681), .ZN(n8867) );
  INV_X1 U7576 ( .A(n8658), .ZN(n7183) );
  INV_X1 U7577 ( .A(n8144), .ZN(n8288) );
  NAND2_X1 U7578 ( .A1(n7912), .A2(n6906), .ZN(n6905) );
  NOR2_X1 U7579 ( .A1(n7929), .A2(n6907), .ZN(n6906) );
  INV_X1 U7580 ( .A(n7911), .ZN(n6907) );
  NAND2_X1 U7581 ( .A1(n11349), .A2(n11347), .ZN(n6789) );
  OR2_X1 U7582 ( .A1(n6537), .A2(n11347), .ZN(n6786) );
  OR2_X1 U7583 ( .A1(n14640), .A2(n7337), .ZN(n7336) );
  NAND2_X1 U7584 ( .A1(n8972), .A2(n8971), .ZN(n8979) );
  NAND2_X1 U7585 ( .A1(n6491), .A2(n6469), .ZN(n7409) );
  AOI21_X1 U7586 ( .B1(n7410), .B2(n7409), .A(n6569), .ZN(n7407) );
  NAND2_X1 U7587 ( .A1(n6608), .A2(n6607), .ZN(n13750) );
  NAND2_X1 U7588 ( .A1(n13740), .A2(n13768), .ZN(n6607) );
  NAND2_X1 U7589 ( .A1(n13973), .A2(n13607), .ZN(n6608) );
  AOI21_X1 U7590 ( .B1(n7237), .B2(n7239), .A(n7234), .ZN(n7233) );
  INV_X1 U7591 ( .A(n7827), .ZN(n7234) );
  NAND2_X1 U7592 ( .A1(n6842), .A2(n6844), .ZN(n6841) );
  INV_X1 U7593 ( .A(n15037), .ZN(n6729) );
  INV_X1 U7594 ( .A(n15038), .ZN(n6730) );
  OR2_X1 U7595 ( .A1(n10022), .A2(n10021), .ZN(n7122) );
  NAND2_X1 U7596 ( .A1(n7122), .A2(n7121), .ZN(n7120) );
  NAND2_X1 U7597 ( .A1(n10065), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7121) );
  INV_X1 U7598 ( .A(n12685), .ZN(n7178) );
  NOR2_X1 U7599 ( .A1(n12813), .A2(n12291), .ZN(n7175) );
  AND2_X1 U7600 ( .A1(n7196), .A2(n8106), .ZN(n7045) );
  NOR2_X1 U7601 ( .A1(n8115), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7196) );
  OR2_X1 U7602 ( .A1(n8265), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8268) );
  NOR2_X1 U7603 ( .A1(n12848), .A2(n7006), .ZN(n7004) );
  OR2_X1 U7604 ( .A1(n12946), .A2(n12846), .ZN(n12848) );
  AOI21_X1 U7605 ( .B1(n6839), .B2(n8012), .A(n13228), .ZN(n6837) );
  NAND2_X1 U7606 ( .A1(n11257), .A2(n7074), .ZN(n7070) );
  XNOR2_X1 U7607 ( .A(n8973), .B(n10321), .ZN(n9224) );
  INV_X1 U7608 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7415) );
  INV_X1 U7609 ( .A(n11825), .ZN(n7363) );
  AND2_X1 U7610 ( .A1(n13540), .A2(n7362), .ZN(n7361) );
  OR2_X1 U7611 ( .A1(n13510), .A2(n7363), .ZN(n7362) );
  AND2_X1 U7612 ( .A1(n6470), .A2(n6578), .ZN(n6802) );
  INV_X1 U7613 ( .A(n7153), .ZN(n7152) );
  AND2_X1 U7614 ( .A1(n14059), .A2(n12041), .ZN(n12042) );
  OAI21_X1 U7615 ( .B1(n6956), .B2(n6955), .A(n13789), .ZN(n6952) );
  AND2_X1 U7616 ( .A1(n7252), .A2(n7251), .ZN(n7250) );
  NAND2_X1 U7617 ( .A1(n7255), .A2(n7257), .ZN(n7252) );
  XNOR2_X1 U7618 ( .A(n7645), .B(SI_10_), .ZN(n7642) );
  INV_X1 U7619 ( .A(n7623), .ZN(n7624) );
  OAI22_X1 U7620 ( .A1(n14348), .A2(n14301), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14300), .ZN(n14302) );
  AOI21_X1 U7621 ( .B1(n12247), .B2(n7018), .A(n12242), .ZN(n9343) );
  AOI21_X1 U7622 ( .B1(n7308), .B2(n7306), .A(n6502), .ZN(n7305) );
  INV_X1 U7623 ( .A(n7311), .ZN(n7306) );
  AND2_X1 U7624 ( .A1(n12287), .A2(n12369), .ZN(n7299) );
  OR2_X1 U7625 ( .A1(n8400), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8424) );
  INV_X1 U7626 ( .A(n12376), .ZN(n11341) );
  BUF_X1 U7627 ( .A(n8163), .Z(n8753) );
  NAND2_X1 U7628 ( .A1(n15024), .A2(n15023), .ZN(n15022) );
  NAND2_X1 U7629 ( .A1(n6730), .A2(n6729), .ZN(n15035) );
  NAND2_X1 U7630 ( .A1(n8667), .A2(n7197), .ZN(n12588) );
  AND2_X1 U7631 ( .A1(n8938), .A2(n8666), .ZN(n7197) );
  AOI21_X1 U7632 ( .B1(n12620), .B2(n6516), .A(n7054), .ZN(n12591) );
  AND2_X1 U7633 ( .A1(n7055), .A2(n12592), .ZN(n7054) );
  INV_X1 U7634 ( .A(n7057), .ZN(n7055) );
  AND2_X1 U7635 ( .A1(n8780), .A2(n12579), .ZN(n12592) );
  AND3_X1 U7636 ( .A1(n8450), .A2(n8449), .A3(n8448), .ZN(n12681) );
  AOI21_X1 U7637 ( .B1(n7182), .B2(n7180), .A(n6539), .ZN(n7179) );
  INV_X1 U7638 ( .A(n6489), .ZN(n7180) );
  NAND2_X1 U7639 ( .A1(n8672), .A2(n9733), .ZN(n12683) );
  INV_X1 U7640 ( .A(n12666), .ZN(n12759) );
  INV_X1 U7641 ( .A(n12757), .ZN(n7036) );
  NAND2_X1 U7642 ( .A1(n8603), .A2(n8602), .ZN(n8767) );
  NAND2_X1 U7643 ( .A1(n8417), .A2(n8416), .ZN(n8455) );
  NAND2_X1 U7644 ( .A1(n8159), .A2(n8176), .ZN(n8212) );
  INV_X1 U7645 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8176) );
  XNOR2_X1 U7646 ( .A(n10317), .B(n10319), .ZN(n6972) );
  OR2_X1 U7647 ( .A1(n10161), .A2(n9891), .ZN(n10122) );
  INV_X1 U7648 ( .A(n13408), .ZN(n6872) );
  NAND2_X1 U7649 ( .A1(n13457), .A2(n7612), .ZN(n7921) );
  AOI21_X1 U7650 ( .B1(n6558), .B2(n6707), .A(n6704), .ZN(n6703) );
  NOR2_X1 U7651 ( .A1(n13425), .A2(n13031), .ZN(n6704) );
  OR2_X1 U7652 ( .A1(n10654), .A2(n10646), .ZN(n7984) );
  NAND2_X1 U7653 ( .A1(n10159), .A2(n7485), .ZN(n10205) );
  OR2_X1 U7654 ( .A1(n10162), .A2(n7484), .ZN(n10159) );
  INV_X1 U7655 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U7656 ( .A1(n10390), .A2(n7348), .ZN(n7347) );
  AOI21_X1 U7657 ( .B1(n7365), .B2(n7367), .A(n6531), .ZN(n7364) );
  INV_X1 U7658 ( .A(n7369), .ZN(n7368) );
  NAND2_X1 U7659 ( .A1(n10875), .A2(n7372), .ZN(n7371) );
  OAI21_X1 U7660 ( .B1(n7373), .B2(n7370), .A(n11288), .ZN(n7369) );
  AND2_X1 U7661 ( .A1(n13983), .A2(n7222), .ZN(n7220) );
  NAND2_X1 U7662 ( .A1(n13986), .A2(n12047), .ZN(n13987) );
  NAND2_X1 U7663 ( .A1(n11942), .A2(n11941), .ZN(n14029) );
  NAND2_X1 U7664 ( .A1(n14051), .A2(n12016), .ZN(n7201) );
  AOI21_X1 U7665 ( .B1(n12016), .B2(n14056), .A(n6495), .ZN(n7202) );
  AOI22_X1 U7666 ( .A1(n14095), .A2(n14098), .B1(n14225), .B2(n13829), .ZN(
        n14084) );
  AND2_X1 U7667 ( .A1(n12038), .A2(n12008), .ZN(n14128) );
  OR2_X1 U7668 ( .A1(n14564), .A2(n13837), .ZN(n11380) );
  NAND2_X1 U7669 ( .A1(n6932), .A2(n6931), .ZN(n10631) );
  AOI21_X1 U7670 ( .B1(n10627), .B2(n6930), .A(n6475), .ZN(n6931) );
  NAND2_X1 U7671 ( .A1(n10714), .A2(n6929), .ZN(n6932) );
  NAND2_X1 U7672 ( .A1(n10714), .A2(n6935), .ZN(n6934) );
  OAI21_X1 U7673 ( .B1(n14010), .B2(n6939), .A(n6936), .ZN(n12045) );
  AOI21_X1 U7674 ( .B1(n6938), .B2(n6942), .A(n6937), .ZN(n6936) );
  NAND2_X1 U7675 ( .A1(n9440), .A2(n9439), .ZN(n9569) );
  AOI21_X1 U7676 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14316), .A(n14315), .ZN(
        n14322) );
  OR2_X1 U7677 ( .A1(n14642), .A2(n6822), .ZN(n6817) );
  NAND2_X1 U7678 ( .A1(n14642), .A2(n6822), .ZN(n6818) );
  AOI21_X1 U7679 ( .B1(n6751), .B2(n9342), .A(n6559), .ZN(n6748) );
  AND2_X1 U7680 ( .A1(n6751), .A2(n6564), .ZN(n6749) );
  INV_X1 U7681 ( .A(n12683), .ZN(n12756) );
  NAND2_X1 U7682 ( .A1(n8459), .A2(n8458), .ZN(n12808) );
  XNOR2_X1 U7683 ( .A(n6720), .B(n8102), .ZN(n13311) );
  AOI21_X1 U7684 ( .B1(n7098), .B2(n14535), .A(n6589), .ZN(n13315) );
  INV_X1 U7685 ( .A(n9002), .ZN(n7398) );
  OR2_X1 U7686 ( .A1(n9010), .A2(n9011), .ZN(n9012) );
  OAI21_X1 U7687 ( .B1(n9003), .B2(n7397), .A(n7396), .ZN(n9010) );
  NAND2_X1 U7688 ( .A1(n9016), .A2(n9017), .ZN(n7413) );
  NAND2_X1 U7689 ( .A1(n13639), .A2(n13637), .ZN(n7140) );
  NAND2_X1 U7690 ( .A1(n7401), .A2(n6478), .ZN(n6662) );
  NAND2_X1 U7691 ( .A1(n13651), .A2(n7142), .ZN(n7141) );
  INV_X1 U7692 ( .A(n13650), .ZN(n7142) );
  NAND2_X1 U7693 ( .A1(n7145), .A2(n13663), .ZN(n7144) );
  AOI22_X1 U7694 ( .A1(n7404), .A2(n7406), .B1(n7408), .B2(n7410), .ZN(n7402)
         );
  INV_X1 U7695 ( .A(n7407), .ZN(n7406) );
  OR2_X1 U7696 ( .A1(n13685), .A2(n13684), .ZN(n7418) );
  NAND2_X1 U7697 ( .A1(n7124), .A2(n13691), .ZN(n6687) );
  INV_X1 U7698 ( .A(n13715), .ZN(n7157) );
  INV_X1 U7699 ( .A(n13714), .ZN(n7161) );
  INV_X1 U7700 ( .A(n7238), .ZN(n7237) );
  OAI21_X1 U7701 ( .B1(n7240), .B2(n7239), .A(n7819), .ZN(n7238) );
  MUX2_X1 U7702 ( .A(n8903), .B(n8902), .S(n9733), .Z(n8904) );
  AOI21_X1 U7703 ( .B1(n8437), .B2(n8452), .A(n6598), .ZN(n7025) );
  INV_X1 U7704 ( .A(n8452), .ZN(n7023) );
  OAI211_X1 U7705 ( .C1(n9174), .C2(n9173), .A(n6630), .B(n6629), .ZN(n9178)
         );
  NAND2_X1 U7706 ( .A1(n9170), .A2(n9169), .ZN(n6629) );
  NAND2_X1 U7707 ( .A1(n9172), .A2(n9171), .ZN(n6630) );
  NAND2_X1 U7708 ( .A1(n9155), .A2(n9154), .ZN(n9198) );
  NAND2_X1 U7709 ( .A1(n13711), .A2(n13710), .ZN(n6637) );
  AND2_X1 U7710 ( .A1(n6632), .A2(n7135), .ZN(n6631) );
  NAND2_X1 U7711 ( .A1(n13726), .A2(n7136), .ZN(n7135) );
  NAND2_X1 U7712 ( .A1(n7648), .A2(n12095), .ZN(n7661) );
  AND2_X1 U7713 ( .A1(n8700), .A2(n9257), .ZN(n7318) );
  INV_X1 U7714 ( .A(n9261), .ZN(n12240) );
  AND2_X1 U7715 ( .A1(n12773), .A2(n12525), .ZN(n8943) );
  NAND2_X1 U7716 ( .A1(n12388), .A2(n6594), .ZN(n12410) );
  AND2_X1 U7717 ( .A1(n6668), .A2(n12552), .ZN(n7172) );
  OR2_X1 U7718 ( .A1(n7063), .A2(n7067), .ZN(n7059) );
  INV_X1 U7719 ( .A(n8909), .ZN(n7063) );
  NAND2_X1 U7720 ( .A1(n12544), .A2(n9368), .ZN(n8909) );
  OR2_X1 U7721 ( .A1(n12544), .A2(n9368), .ZN(n8911) );
  NAND2_X1 U7722 ( .A1(n12588), .A2(n8668), .ZN(n12572) );
  OR2_X1 U7723 ( .A1(n8470), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8485) );
  OR2_X1 U7724 ( .A1(n12813), .A2(n12668), .ZN(n8870) );
  AND2_X1 U7725 ( .A1(n8848), .A2(n7042), .ZN(n7041) );
  NAND2_X1 U7726 ( .A1(n7043), .A2(n8843), .ZN(n7042) );
  INV_X1 U7727 ( .A(n8847), .ZN(n7039) );
  OR2_X1 U7728 ( .A1(n11630), .A2(n12371), .ZN(n8853) );
  INV_X1 U7729 ( .A(n8333), .ZN(n8332) );
  INV_X1 U7730 ( .A(n7051), .ZN(n7050) );
  OAI21_X1 U7731 ( .B1(n11039), .B2(n7052), .A(n8829), .ZN(n7051) );
  INV_X1 U7732 ( .A(n8825), .ZN(n7052) );
  INV_X1 U7733 ( .A(n10500), .ZN(n9258) );
  OR2_X1 U7734 ( .A1(n8325), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8343) );
  NOR2_X1 U7735 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n6741) );
  OR2_X1 U7736 ( .A1(n8212), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8214) );
  NOR2_X1 U7737 ( .A1(n8214), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8248) );
  NAND2_X1 U7738 ( .A1(n9197), .A2(n9196), .ZN(n9201) );
  INV_X1 U7739 ( .A(n7763), .ZN(n6898) );
  INV_X1 U7740 ( .A(n9220), .ZN(n6897) );
  INV_X1 U7741 ( .A(n7072), .ZN(n7071) );
  OAI21_X1 U7742 ( .B1(n6490), .B2(n7073), .A(n7991), .ZN(n7072) );
  NAND2_X1 U7743 ( .A1(n7088), .A2(n7986), .ZN(n7087) );
  INV_X1 U7744 ( .A(n7986), .ZN(n7089) );
  NAND2_X1 U7745 ( .A1(n13163), .A2(n13413), .ZN(n8092) );
  NAND2_X1 U7746 ( .A1(n13465), .A2(n7612), .ZN(n7887) );
  AND2_X1 U7747 ( .A1(n7748), .A2(n7768), .ZN(n7012) );
  INV_X1 U7748 ( .A(n7134), .ZN(n7133) );
  OR2_X1 U7749 ( .A1(n13573), .A2(n13738), .ZN(n7165) );
  NOR2_X1 U7750 ( .A1(n6693), .A2(n14200), .ZN(n6862) );
  INV_X1 U7751 ( .A(n6964), .ZN(n6963) );
  OAI21_X1 U7752 ( .B1(n12039), .B2(n6961), .A(n12038), .ZN(n6960) );
  NAND2_X1 U7753 ( .A1(n6965), .A2(n6964), .ZN(n6961) );
  NOR2_X1 U7754 ( .A1(n11710), .A2(n14575), .ZN(n6866) );
  OR2_X1 U7755 ( .A1(n11799), .A2(n11804), .ZN(n13672) );
  OR2_X1 U7756 ( .A1(n10626), .A2(n13616), .ZN(n6935) );
  NAND2_X1 U7757 ( .A1(n10764), .A2(n14776), .ZN(n10766) );
  AOI21_X1 U7758 ( .B1(n7930), .B2(n7268), .A(n7266), .ZN(n7265) );
  INV_X1 U7759 ( .A(n7932), .ZN(n7266) );
  AND2_X1 U7760 ( .A1(n7766), .A2(n7747), .ZN(n7764) );
  NAND2_X1 U7761 ( .A1(n7703), .A2(SI_13_), .ZN(n7704) );
  NOR2_X1 U7762 ( .A1(n7705), .A2(n7263), .ZN(n7262) );
  INV_X1 U7763 ( .A(n7678), .ZN(n7263) );
  INV_X1 U7764 ( .A(n7701), .ZN(n7705) );
  XNOR2_X1 U7765 ( .A(n7626), .B(SI_9_), .ZN(n7623) );
  INV_X1 U7766 ( .A(n7607), .ZN(n7608) );
  XNOR2_X1 U7767 ( .A(n7590), .B(SI_7_), .ZN(n7587) );
  AOI21_X1 U7768 ( .B1(n7579), .B2(n7246), .A(n6556), .ZN(n7245) );
  XNOR2_X1 U7769 ( .A(n7341), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n14333) );
  INV_X1 U7770 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n7341) );
  NOR2_X1 U7771 ( .A1(n14297), .A2(n14298), .ZN(n14299) );
  XNOR2_X1 U7772 ( .A(n14299), .B(n6812), .ZN(n14342) );
  AOI21_X1 U7773 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(n14351), .A(n14303), .ZN(
        n14354) );
  NAND2_X1 U7774 ( .A1(n14305), .A2(n6809), .ZN(n14307) );
  NAND2_X1 U7775 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(n6810), .ZN(n6809) );
  INV_X1 U7776 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U7777 ( .A1(n9343), .A2(n9342), .ZN(n7286) );
  INV_X1 U7778 ( .A(n9296), .ZN(n7309) );
  INV_X1 U7779 ( .A(n6754), .ZN(n6755) );
  OAI21_X1 U7780 ( .B1(n12298), .B2(n6760), .A(n12277), .ZN(n6754) );
  INV_X1 U7781 ( .A(n12370), .ZN(n11629) );
  NAND2_X1 U7782 ( .A1(n6639), .A2(n12299), .ZN(n6757) );
  NAND2_X1 U7783 ( .A1(n12298), .A2(n12364), .ZN(n6639) );
  NOR2_X1 U7784 ( .A1(n9297), .A2(n7312), .ZN(n7311) );
  INV_X1 U7785 ( .A(n9291), .ZN(n7312) );
  NAND2_X1 U7786 ( .A1(n6772), .A2(n6775), .ZN(n9323) );
  AND2_X1 U7787 ( .A1(n6776), .A2(n7278), .ZN(n6775) );
  AOI21_X1 U7788 ( .B1(n9318), .B2(n7280), .A(n7279), .ZN(n7278) );
  OAI211_X1 U7789 ( .C1(n6449), .C2(n9489), .A(n8162), .B(n8161), .ZN(n10183)
         );
  NAND2_X1 U7790 ( .A1(n8423), .A2(n8422), .ZN(n8444) );
  INV_X1 U7791 ( .A(n8424), .ZN(n8423) );
  NAND2_X1 U7792 ( .A1(n6768), .A2(n6767), .ZN(n7293) );
  NOR2_X1 U7793 ( .A1(n10382), .A2(n6769), .ZN(n6768) );
  AND2_X1 U7794 ( .A1(n10463), .A2(n7292), .ZN(n7291) );
  INV_X1 U7795 ( .A(n7422), .ZN(n7292) );
  NAND2_X1 U7796 ( .A1(n7290), .A2(n10635), .ZN(n7289) );
  INV_X1 U7797 ( .A(n9278), .ZN(n7290) );
  NAND2_X1 U7798 ( .A1(n6766), .A2(n7300), .ZN(n12349) );
  AOI21_X1 U7799 ( .B1(n7302), .B2(n7305), .A(n7301), .ZN(n7300) );
  NAND2_X1 U7800 ( .A1(n11339), .A2(n7303), .ZN(n6766) );
  NOR2_X1 U7801 ( .A1(n9299), .A2(n12371), .ZN(n7301) );
  OR2_X1 U7802 ( .A1(n15005), .A2(n9998), .ZN(n15003) );
  NAND2_X1 U7803 ( .A1(n15022), .A2(n6518), .ZN(n10020) );
  NOR2_X1 U7804 ( .A1(n6739), .A2(n15053), .ZN(n6735) );
  NAND2_X1 U7805 ( .A1(n6730), .A2(n6474), .ZN(n6732) );
  NAND2_X1 U7806 ( .A1(n10058), .A2(n6722), .ZN(n10297) );
  OR2_X1 U7807 ( .A1(n10060), .A2(n10059), .ZN(n6722) );
  INV_X1 U7808 ( .A(n7120), .ZN(n10304) );
  INV_X1 U7809 ( .A(n7113), .ZN(n10887) );
  OR2_X1 U7810 ( .A1(n15090), .A2(n15089), .ZN(n7119) );
  XNOR2_X1 U7811 ( .A(n11136), .B(n11143), .ZN(n10910) );
  NAND2_X1 U7812 ( .A1(n15082), .A2(n6721), .ZN(n11136) );
  OR2_X1 U7813 ( .A1(n15101), .A2(n10896), .ZN(n6721) );
  NAND2_X1 U7814 ( .A1(n7119), .A2(n7118), .ZN(n7117) );
  NAND2_X1 U7815 ( .A1(n10904), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7118) );
  NOR2_X1 U7816 ( .A1(n12386), .A2(n6591), .ZN(n12404) );
  XNOR2_X1 U7817 ( .A(n12410), .B(n12405), .ZN(n12389) );
  NAND2_X1 U7818 ( .A1(n12416), .A2(n12420), .ZN(n12435) );
  NAND2_X1 U7819 ( .A1(n12435), .A2(n12436), .ZN(n12456) );
  NAND2_X1 U7820 ( .A1(n7109), .A2(n12486), .ZN(n12506) );
  NAND2_X1 U7821 ( .A1(n7111), .A2(n7110), .ZN(n7109) );
  INV_X1 U7822 ( .A(n7432), .ZN(n7110) );
  OR2_X1 U7823 ( .A1(n8560), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U7824 ( .A1(n8529), .A2(n8528), .ZN(n8543) );
  NAND2_X1 U7825 ( .A1(n6562), .A2(n8779), .ZN(n7057) );
  NAND2_X1 U7826 ( .A1(n8783), .A2(n8888), .ZN(n7058) );
  AND2_X1 U7827 ( .A1(n8779), .A2(n8888), .ZN(n7056) );
  OAI21_X1 U7828 ( .B1(n12638), .B2(n7188), .A(n7186), .ZN(n12616) );
  INV_X1 U7829 ( .A(n7189), .ZN(n7188) );
  AOI21_X1 U7830 ( .B1(n7189), .B2(n7187), .A(n6541), .ZN(n7186) );
  AND2_X1 U7831 ( .A1(n8784), .A2(n8881), .ZN(n7046) );
  NOR2_X1 U7832 ( .A1(n12629), .A2(n7190), .ZN(n7189) );
  INV_X1 U7833 ( .A(n8664), .ZN(n7190) );
  OR2_X1 U7834 ( .A1(n12646), .A2(n12654), .ZN(n8881) );
  AND2_X1 U7835 ( .A1(n8784), .A2(n8785), .ZN(n12629) );
  NAND2_X1 U7836 ( .A1(n12638), .A2(n12645), .ZN(n12637) );
  OR2_X1 U7837 ( .A1(n8444), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8461) );
  AOI21_X1 U7838 ( .B1(n7176), .B2(n7179), .A(n7175), .ZN(n7174) );
  NAND2_X1 U7839 ( .A1(n7179), .A2(n7178), .ZN(n7177) );
  AND2_X1 U7840 ( .A1(n8870), .A2(n8868), .ZN(n12685) );
  INV_X1 U7841 ( .A(n11441), .ZN(n7185) );
  AND2_X1 U7842 ( .A1(n8853), .A2(n8852), .ZN(n11446) );
  NAND2_X1 U7843 ( .A1(n11331), .A2(n11330), .ZN(n11329) );
  INV_X1 U7844 ( .A(n11560), .ZN(n11409) );
  NAND2_X1 U7845 ( .A1(n10814), .A2(n6519), .ZN(n11041) );
  NAND2_X1 U7846 ( .A1(n11040), .A2(n11039), .ZN(n11038) );
  AND4_X1 U7847 ( .A1(n8260), .A2(n8259), .A3(n8258), .A4(n8257), .ZN(n11205)
         );
  NAND2_X1 U7848 ( .A1(n10816), .A2(n10815), .ZN(n10814) );
  NAND2_X1 U7849 ( .A1(n8820), .A2(n8821), .ZN(n10815) );
  NAND2_X1 U7850 ( .A1(n10427), .A2(n8634), .ZN(n10566) );
  OR2_X1 U7851 ( .A1(n8219), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U7852 ( .A1(n8806), .A2(n10131), .ZN(n6689) );
  INV_X1 U7853 ( .A(n10131), .ZN(n10138) );
  NAND2_X1 U7854 ( .A1(n10082), .A2(n8802), .ZN(n10139) );
  NAND2_X1 U7855 ( .A1(n10139), .A2(n10138), .ZN(n10137) );
  NAND2_X1 U7856 ( .A1(n10083), .A2(n10084), .ZN(n10082) );
  INV_X1 U7857 ( .A(n12680), .ZN(n12762) );
  AND2_X1 U7858 ( .A1(n9734), .A2(n9139), .ZN(n8144) );
  OR2_X1 U7859 ( .A1(n11324), .A2(n6449), .ZN(n8559) );
  INV_X1 U7860 ( .A(n14470), .ZN(n14467) );
  OAI22_X1 U7861 ( .A1(n8747), .A2(n8746), .B1(P2_DATAO_REG_29__SCAN_IN), .B2(
        n13448), .ZN(n8761) );
  AND2_X1 U7862 ( .A1(n8119), .A2(n12824), .ZN(n8120) );
  XNOR2_X1 U7863 ( .A(n8693), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U7864 ( .A1(n7316), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8693) );
  AND2_X1 U7865 ( .A1(n7314), .A2(n12094), .ZN(n7313) );
  NAND2_X1 U7866 ( .A1(n8555), .A2(n8554), .ZN(n8570) );
  OAI21_X1 U7867 ( .B1(n8537), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7026), .ZN(
        n8553) );
  NOR3_X1 U7868 ( .A1(n8325), .A2(n8110), .A3(P3_IR_REG_12__SCAN_IN), .ZN(
        n8617) );
  OR2_X1 U7869 ( .A1(n8438), .A2(n8437), .ZN(n8453) );
  AND2_X1 U7870 ( .A1(n8270), .A2(n8269), .ZN(n10906) );
  AND2_X1 U7871 ( .A1(n9501), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8244) );
  XNOR2_X1 U7872 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8261) );
  INV_X1 U7873 ( .A(n8207), .ZN(n8208) );
  INV_X1 U7874 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8104) );
  AOI21_X1 U7875 ( .B1(n6983), .B2(n6985), .A(n6560), .ZN(n6982) );
  INV_X1 U7876 ( .A(n10838), .ZN(n6983) );
  INV_X1 U7877 ( .A(n10946), .ZN(n6986) );
  NOR2_X1 U7878 ( .A1(n10947), .A2(n10847), .ZN(n6985) );
  AOI21_X1 U7879 ( .B1(n12862), .B2(n6969), .A(n6550), .ZN(n6968) );
  INV_X1 U7880 ( .A(n12862), .ZN(n6970) );
  INV_X1 U7881 ( .A(n12927), .ZN(n6969) );
  INV_X1 U7882 ( .A(n13002), .ZN(n6997) );
  NAND2_X1 U7883 ( .A1(n11275), .A2(n11276), .ZN(n11302) );
  NAND2_X1 U7884 ( .A1(n6988), .A2(n6511), .ZN(n11569) );
  INV_X1 U7885 ( .A(n11460), .ZN(n6987) );
  NAND2_X1 U7886 ( .A1(n6972), .A2(n6971), .ZN(n6975) );
  NAND2_X1 U7887 ( .A1(n12847), .A2(n7008), .ZN(n7001) );
  OR2_X1 U7888 ( .A1(n7004), .A2(n7000), .ZN(n6623) );
  NAND2_X1 U7889 ( .A1(n10837), .A2(n10838), .ZN(n10849) );
  OR2_X1 U7890 ( .A1(n7487), .A2(n10110), .ZN(n7479) );
  NAND2_X1 U7891 ( .A1(n13185), .A2(n7910), .ZN(n7912) );
  INV_X1 U7892 ( .A(n8012), .ZN(n6838) );
  NOR2_X1 U7893 ( .A1(n8007), .A2(n8010), .ZN(n7094) );
  NAND2_X1 U7894 ( .A1(n7096), .A2(n8009), .ZN(n7095) );
  INV_X1 U7895 ( .A(n8010), .ZN(n7096) );
  AOI21_X1 U7896 ( .B1(n6709), .B2(n6708), .A(n6506), .ZN(n6707) );
  INV_X1 U7897 ( .A(n7815), .ZN(n6708) );
  NOR2_X1 U7898 ( .A1(n6888), .A2(n13277), .ZN(n6887) );
  OR2_X1 U7899 ( .A1(n6889), .A2(n13367), .ZN(n6888) );
  NOR2_X1 U7900 ( .A1(n14505), .A2(n7083), .ZN(n7082) );
  INV_X1 U7901 ( .A(n9233), .ZN(n7083) );
  INV_X1 U7902 ( .A(n9237), .ZN(n11672) );
  AOI21_X1 U7903 ( .B1(n6716), .B2(n6718), .A(n6508), .ZN(n6715) );
  OAI22_X2 U7904 ( .A1(n11157), .A2(n7988), .B1(n11319), .B2(n13041), .ZN(
        n11257) );
  NAND2_X1 U7905 ( .A1(n10804), .A2(n6492), .ZN(n10969) );
  NOR2_X1 U7906 ( .A1(n11162), .A2(n11316), .ZN(n11263) );
  AND2_X1 U7907 ( .A1(n10502), .A2(n7982), .ZN(n10645) );
  NOR2_X1 U7908 ( .A1(n8960), .A2(n8956), .ZN(n10161) );
  INV_X1 U7909 ( .A(n12921), .ZN(n6616) );
  NOR2_X1 U7910 ( .A1(n8073), .A2(n13371), .ZN(n6617) );
  INV_X1 U7911 ( .A(n7919), .ZN(n7808) );
  INV_X1 U7912 ( .A(n9803), .ZN(n7807) );
  OR3_X2 U7913 ( .A1(n7452), .A2(P2_IR_REG_28__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n7466) );
  INV_X1 U7914 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7448) );
  NAND2_X1 U7915 ( .A1(n7447), .A2(n7667), .ZN(n6901) );
  INV_X1 U7916 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7748) );
  INV_X1 U7917 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U7918 ( .A1(n11004), .A2(n11003), .ZN(n13640) );
  AOI21_X1 U7919 ( .B1(n7361), .B2(n7363), .A(n6533), .ZN(n7360) );
  OR2_X1 U7920 ( .A1(n13550), .A2(n7358), .ZN(n7357) );
  MUX2_X1 U7921 ( .A(n10393), .B(n9718), .S(n9717), .Z(n9719) );
  AND2_X1 U7922 ( .A1(n13471), .A2(n7366), .ZN(n7365) );
  OR2_X1 U7923 ( .A1(n13534), .A2(n7367), .ZN(n7366) );
  INV_X1 U7924 ( .A(n14650), .ZN(n7345) );
  AOI21_X1 U7925 ( .B1(n12223), .B2(n13846), .A(n9715), .ZN(n9716) );
  AOI21_X1 U7926 ( .B1(n6464), .B2(n6802), .A(n6540), .ZN(n6801) );
  AND4_X1 U7927 ( .A1(n10616), .A2(n10615), .A3(n10614), .A4(n10613), .ZN(
        n11290) );
  NAND2_X1 U7928 ( .A1(n9385), .A2(n10173), .ZN(n10880) );
  NOR2_X1 U7929 ( .A1(n13987), .A2(n13742), .ZN(n13974) );
  NAND2_X1 U7930 ( .A1(n14179), .A2(n12228), .ZN(n7222) );
  OR2_X1 U7931 ( .A1(n14174), .A2(n12024), .ZN(n12025) );
  INV_X1 U7932 ( .A(n13995), .ZN(n14004) );
  AND2_X1 U7933 ( .A1(n6860), .A2(n6572), .ZN(n13986) );
  AND2_X1 U7934 ( .A1(n6949), .A2(n12042), .ZN(n6944) );
  XNOR2_X1 U7935 ( .A(n13717), .B(n12018), .ZN(n14008) );
  INV_X1 U7936 ( .A(n14025), .ZN(n7203) );
  NAND2_X1 U7937 ( .A1(n12046), .A2(n13825), .ZN(n6950) );
  NOR2_X1 U7938 ( .A1(n14054), .A2(n12042), .ZN(n14039) );
  NAND2_X1 U7939 ( .A1(n14038), .A2(n14039), .ZN(n14037) );
  OAI21_X1 U7940 ( .B1(n14067), .B2(n13696), .A(n13699), .ZN(n14057) );
  AND2_X1 U7941 ( .A1(n14057), .A2(n14056), .ZN(n14054) );
  XNOR2_X1 U7942 ( .A(n14059), .B(n13826), .ZN(n14056) );
  OR2_X1 U7943 ( .A1(n7207), .A2(n12013), .ZN(n7204) );
  NOR2_X1 U7944 ( .A1(n7209), .A2(n7208), .ZN(n7207) );
  NOR2_X1 U7945 ( .A1(n14115), .A2(n14105), .ZN(n14099) );
  AND2_X1 U7946 ( .A1(n14233), .A2(n13577), .ZN(n12040) );
  NAND2_X1 U7947 ( .A1(n6866), .A2(n6865), .ZN(n14151) );
  NAND2_X1 U7948 ( .A1(n13682), .A2(n6966), .ZN(n6964) );
  NAND2_X1 U7949 ( .A1(n13683), .A2(n6967), .ZN(n6966) );
  INV_X1 U7950 ( .A(n12036), .ZN(n6967) );
  NAND2_X1 U7951 ( .A1(n13682), .A2(n13796), .ZN(n6965) );
  AND2_X1 U7952 ( .A1(n14575), .A2(n13677), .ZN(n12036) );
  NOR2_X1 U7953 ( .A1(n11699), .A2(n11702), .ZN(n12037) );
  NAND2_X1 U7954 ( .A1(n11584), .A2(n11700), .ZN(n11698) );
  NAND2_X1 U7955 ( .A1(n11382), .A2(n13793), .ZN(n11529) );
  NOR2_X1 U7956 ( .A1(n13793), .A2(n6920), .ZN(n6919) );
  NOR2_X1 U7957 ( .A1(n13791), .A2(n6921), .ZN(n6920) );
  INV_X1 U7958 ( .A(n11373), .ZN(n6921) );
  NAND2_X1 U7959 ( .A1(n11219), .A2(n13791), .ZN(n11374) );
  OR2_X1 U7960 ( .A1(n13649), .A2(n13838), .ZN(n11220) );
  NAND2_X1 U7961 ( .A1(n6953), .A2(n6951), .ZN(n11214) );
  INV_X1 U7962 ( .A(n6952), .ZN(n6951) );
  NOR2_X1 U7963 ( .A1(n6955), .A2(n11053), .ZN(n6954) );
  AND2_X1 U7964 ( .A1(n11060), .A2(n14800), .ZN(n11121) );
  NOR2_X1 U7965 ( .A1(n11061), .A2(n14698), .ZN(n11060) );
  NAND2_X1 U7966 ( .A1(n11016), .A2(n13788), .ZN(n11055) );
  AND2_X1 U7967 ( .A1(n13616), .A2(n13843), .ZN(n6657) );
  NAND2_X1 U7968 ( .A1(n10626), .A2(n13616), .ZN(n6933) );
  INV_X1 U7969 ( .A(n13783), .ZN(n10757) );
  NAND2_X1 U7970 ( .A1(n10625), .A2(n10624), .ZN(n10714) );
  NAND2_X1 U7971 ( .A1(n11895), .A2(n6916), .ZN(n9711) );
  AND2_X1 U7972 ( .A1(n9139), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U7973 ( .A1(n6805), .A2(n13569), .ZN(n14789) );
  NOR2_X1 U7974 ( .A1(n9187), .A2(n7276), .ZN(n7275) );
  INV_X1 U7975 ( .A(n9138), .ZN(n7276) );
  AND2_X1 U7976 ( .A1(n9393), .A2(n6571), .ZN(n7223) );
  NAND2_X1 U7977 ( .A1(n7267), .A2(n7913), .ZN(n7931) );
  NAND2_X1 U7978 ( .A1(n7899), .A2(n7269), .ZN(n7267) );
  INV_X1 U7979 ( .A(n7864), .ZN(n7242) );
  NAND2_X1 U7980 ( .A1(n7865), .A2(SI_22_), .ZN(n7866) );
  XNOR2_X1 U7981 ( .A(n7853), .B(n7852), .ZN(n11880) );
  OAI21_X1 U7982 ( .B1(n7840), .B2(n7232), .A(n7843), .ZN(n7853) );
  NOR2_X2 U7983 ( .A1(n10880), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n9540) );
  XNOR2_X1 U7984 ( .A(n14342), .B(n7330), .ZN(n14344) );
  INV_X1 U7985 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7330) );
  NOR2_X1 U7986 ( .A1(n14309), .A2(n6826), .ZN(n14325) );
  AND2_X1 U7987 ( .A1(n14310), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n6826) );
  NOR2_X1 U7988 ( .A1(n14364), .A2(n14363), .ZN(n14309) );
  AOI21_X1 U7989 ( .B1(n14623), .B2(n7323), .A(n7322), .ZN(n7321) );
  NOR2_X1 U7990 ( .A1(n7324), .A2(n7325), .ZN(n7322) );
  OAI21_X1 U7991 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n14318), .A(n14317), .ZN(
        n14373) );
  AND3_X1 U7992 ( .A1(n6747), .A2(n12251), .A3(n6746), .ZN(n6743) );
  NAND2_X1 U7993 ( .A1(n6748), .A2(n6752), .ZN(n6746) );
  NAND2_X1 U7994 ( .A1(n6749), .A2(n9342), .ZN(n6747) );
  NOR2_X1 U7995 ( .A1(n9271), .A2(n10033), .ZN(n10031) );
  NAND2_X1 U7996 ( .A1(n9264), .A2(n9263), .ZN(n9271) );
  INV_X1 U7997 ( .A(n12365), .ZN(n12628) );
  NAND2_X1 U7998 ( .A1(n12350), .A2(n6763), .ZN(n12289) );
  OR2_X1 U7999 ( .A1(n9301), .A2(n11629), .ZN(n6763) );
  INV_X1 U8000 ( .A(n12654), .ZN(n12367) );
  NAND4_X1 U8001 ( .A1(n8279), .A2(n8278), .A3(n8277), .A4(n8276), .ZN(n12376)
         );
  XNOR2_X1 U8002 ( .A(n10297), .B(n10305), .ZN(n10061) );
  NAND2_X1 U8003 ( .A1(n10061), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n10299) );
  NAND2_X1 U8004 ( .A1(n15083), .A2(n15084), .ZN(n15082) );
  XNOR2_X1 U8005 ( .A(n7117), .B(n11137), .ZN(n10889) );
  NOR2_X1 U8006 ( .A1(n10889), .A2(n11411), .ZN(n11132) );
  NAND2_X1 U8007 ( .A1(n11140), .A2(n11141), .ZN(n12388) );
  XNOR2_X1 U8008 ( .A(n12456), .B(n12462), .ZN(n12437) );
  NAND2_X1 U8009 ( .A1(n12459), .A2(n12460), .ZN(n12492) );
  OR2_X1 U8010 ( .A1(n12515), .A2(n6728), .ZN(n6727) );
  AND2_X1 U8011 ( .A1(n14425), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n6728) );
  OAI21_X1 U8012 ( .B1(n8684), .B2(n12680), .A(n8683), .ZN(n12529) );
  NOR2_X1 U8013 ( .A1(n8682), .A2(n8681), .ZN(n8683) );
  NAND2_X1 U8014 ( .A1(n12541), .A2(n12540), .ZN(n12699) );
  OR3_X1 U8015 ( .A1(n12538), .A2(n12537), .A3(n12680), .ZN(n12541) );
  AND2_X1 U8016 ( .A1(n7170), .A2(n7169), .ZN(n12538) );
  NAND2_X1 U8017 ( .A1(n8667), .A2(n8666), .ZN(n12590) );
  NAND2_X1 U8018 ( .A1(n12670), .A2(n8867), .ZN(n12659) );
  NAND2_X1 U8019 ( .A1(n8399), .A2(n8398), .ZN(n12747) );
  INV_X1 U8020 ( .A(n12778), .ZN(n6668) );
  AOI21_X1 U8021 ( .B1(n12534), .B2(n14475), .A(n12529), .ZN(n8741) );
  NAND2_X1 U8022 ( .A1(n9803), .A2(n7375), .ZN(n7461) );
  OR2_X1 U8023 ( .A1(n7919), .A2(n9478), .ZN(n7462) );
  NOR2_X1 U8024 ( .A1(n9712), .A2(n8134), .ZN(n7375) );
  AND2_X1 U8025 ( .A1(n6973), .A2(n6976), .ZN(n10738) );
  INV_X1 U8026 ( .A(n10324), .ZN(n6973) );
  OR2_X1 U8027 ( .A1(n10521), .A2(n7493), .ZN(n7104) );
  NAND2_X1 U8028 ( .A1(n14930), .A2(n6658), .ZN(n13100) );
  OR2_X1 U8029 ( .A1(n14936), .A2(n13099), .ZN(n6658) );
  XNOR2_X1 U8030 ( .A(n13144), .B(n13138), .ZN(n11986) );
  AOI21_X1 U8031 ( .B1(n13312), .B2(n14509), .A(n8097), .ZN(n8098) );
  AND2_X1 U8032 ( .A1(n7502), .A2(n7433), .ZN(n7503) );
  AND2_X1 U8033 ( .A1(n6672), .A2(n6671), .ZN(n13314) );
  NAND2_X1 U8034 ( .A1(n6799), .A2(n11973), .ZN(n6798) );
  NAND2_X1 U8035 ( .A1(n13549), .A2(n13550), .ZN(n6799) );
  INV_X1 U8036 ( .A(n12221), .ZN(n6797) );
  INV_X1 U8037 ( .A(n11354), .ZN(n6787) );
  NAND2_X1 U8038 ( .A1(n11500), .A2(n11499), .ZN(n11721) );
  AOI21_X1 U8039 ( .B1(n6781), .B2(n6784), .A(n6532), .ZN(n6778) );
  NAND2_X1 U8040 ( .A1(n6796), .A2(n11720), .ZN(n6793) );
  AND2_X1 U8041 ( .A1(n14562), .A2(n6795), .ZN(n6794) );
  AND2_X1 U8042 ( .A1(n9672), .A2(n9671), .ZN(n14657) );
  INV_X1 U8043 ( .A(n11799), .ZN(n14594) );
  INV_X1 U8044 ( .A(n12011), .ZN(n14129) );
  NAND2_X1 U8045 ( .A1(n6458), .A2(n6915), .ZN(n9912) );
  AND2_X1 U8046 ( .A1(n9139), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U8047 ( .A1(n14173), .A2(n6697), .ZN(n14257) );
  NAND2_X1 U8048 ( .A1(n14623), .A2(n14896), .ZN(n14621) );
  XNOR2_X1 U8049 ( .A(n14325), .B(n6825), .ZN(n14625) );
  INV_X1 U8050 ( .A(n14326), .ZN(n6825) );
  NOR2_X1 U8051 ( .A1(n14372), .A2(n14371), .ZN(n14634) );
  INV_X1 U8052 ( .A(n14640), .ZN(n7335) );
  AND2_X1 U8053 ( .A1(n7336), .A2(n6510), .ZN(n7332) );
  AND2_X1 U8054 ( .A1(n7336), .A2(n14637), .ZN(n7333) );
  OR2_X1 U8055 ( .A1(n13776), .A2(n13584), .ZN(n13586) );
  INV_X1 U8056 ( .A(n10258), .ZN(n13589) );
  OR2_X1 U8057 ( .A1(n13617), .A2(n13619), .ZN(n7162) );
  NAND2_X1 U8058 ( .A1(n7398), .A2(n6488), .ZN(n7396) );
  AOI21_X1 U8059 ( .B1(n7397), .B2(n7396), .A(n7394), .ZN(n7393) );
  INV_X1 U8060 ( .A(n9011), .ZN(n7394) );
  NAND2_X1 U8061 ( .A1(n7414), .A2(n7412), .ZN(n7411) );
  INV_X1 U8062 ( .A(n9017), .ZN(n7412) );
  NAND2_X1 U8063 ( .A1(n13638), .A2(n7139), .ZN(n7138) );
  INV_X1 U8064 ( .A(n13637), .ZN(n7139) );
  NAND2_X1 U8065 ( .A1(n13652), .A2(n13650), .ZN(n7143) );
  INV_X1 U8066 ( .A(n9046), .ZN(n7400) );
  AND2_X1 U8067 ( .A1(n7409), .A2(n6569), .ZN(n7408) );
  AOI21_X1 U8068 ( .B1(n7407), .B2(n7405), .A(n9061), .ZN(n7404) );
  INV_X1 U8069 ( .A(n7409), .ZN(n7405) );
  NOR2_X1 U8070 ( .A1(n6491), .A2(n6469), .ZN(n7410) );
  NAND2_X1 U8071 ( .A1(n13662), .A2(n7147), .ZN(n7146) );
  AND2_X1 U8072 ( .A1(n7391), .A2(n9087), .ZN(n7390) );
  NAND2_X1 U8073 ( .A1(n9085), .A2(n7392), .ZN(n7391) );
  INV_X1 U8074 ( .A(n7390), .ZN(n7389) );
  NAND2_X1 U8075 ( .A1(n9084), .A2(n9080), .ZN(n7388) );
  OAI22_X1 U8076 ( .A1(n9069), .A2(n9068), .B1(n9073), .B2(n9072), .ZN(n9077)
         );
  AOI21_X1 U8077 ( .B1(n13798), .B2(n13689), .A(n13688), .ZN(n7125) );
  MUX2_X1 U8078 ( .A(n12579), .B(n8782), .S(n9970), .Z(n8896) );
  NAND2_X1 U8079 ( .A1(n9162), .A2(n9161), .ZN(n9167) );
  AOI21_X1 U8080 ( .B1(n7382), .B2(n9103), .A(n9102), .ZN(n7377) );
  NAND2_X1 U8081 ( .A1(n6641), .A2(n6640), .ZN(n13744) );
  NAND2_X1 U8082 ( .A1(n13820), .A2(n13768), .ZN(n6640) );
  NAND2_X1 U8083 ( .A1(n13742), .A2(n13607), .ZN(n6641) );
  NAND2_X1 U8084 ( .A1(n13744), .A2(n13745), .ZN(n6632) );
  INV_X1 U8085 ( .A(n7783), .ZN(n7239) );
  NAND2_X1 U8086 ( .A1(n7704), .A2(n7261), .ZN(n7260) );
  INV_X1 U8087 ( .A(n7259), .ZN(n7258) );
  OAI21_X1 U8088 ( .B1(n7262), .B2(n7260), .A(n7721), .ZN(n7259) );
  INV_X1 U8089 ( .A(n9318), .ZN(n7281) );
  NOR2_X1 U8090 ( .A1(n7159), .A2(n6546), .ZN(n7155) );
  NOR2_X1 U8091 ( .A1(n7160), .A2(n13718), .ZN(n7159) );
  INV_X1 U8092 ( .A(n13719), .ZN(n7160) );
  AOI21_X1 U8093 ( .B1(n7155), .B2(n7156), .A(n7154), .ZN(n7153) );
  NOR2_X1 U8094 ( .A1(n7161), .A2(n7157), .ZN(n7156) );
  NOR2_X1 U8095 ( .A1(n7158), .A2(n13719), .ZN(n7154) );
  INV_X1 U8096 ( .A(n13718), .ZN(n7158) );
  AOI21_X1 U8097 ( .B1(n7153), .B2(n7151), .A(n7150), .ZN(n7149) );
  INV_X1 U8098 ( .A(n13723), .ZN(n7150) );
  INV_X1 U8099 ( .A(n7155), .ZN(n7151) );
  NOR2_X1 U8100 ( .A1(n13726), .A2(n7136), .ZN(n7132) );
  INV_X1 U8101 ( .A(n14112), .ZN(n13798) );
  INV_X1 U8102 ( .A(n7913), .ZN(n7268) );
  NOR2_X1 U8103 ( .A1(n7784), .A2(n7241), .ZN(n7240) );
  INV_X1 U8104 ( .A(n7766), .ZN(n7241) );
  INV_X1 U8105 ( .A(n7256), .ZN(n7255) );
  OAI21_X1 U8106 ( .B1(n7262), .B2(n7257), .A(SI_14_), .ZN(n7256) );
  INV_X1 U8107 ( .A(n7704), .ZN(n7257) );
  OR2_X1 U8108 ( .A1(n7255), .A2(n7258), .ZN(n7253) );
  NAND2_X1 U8109 ( .A1(n7258), .A2(n7260), .ZN(n7251) );
  NAND2_X1 U8110 ( .A1(n7724), .A2(n7723), .ZN(n7741) );
  NOR2_X1 U8111 ( .A1(n7247), .A2(n7244), .ZN(n7243) );
  INV_X1 U8112 ( .A(n7561), .ZN(n7244) );
  INV_X1 U8113 ( .A(n7579), .ZN(n7247) );
  INV_X1 U8114 ( .A(n7565), .ZN(n7246) );
  INV_X1 U8115 ( .A(n7339), .ZN(n14296) );
  INV_X1 U8116 ( .A(n9309), .ZN(n7280) );
  INV_X1 U8117 ( .A(n9319), .ZN(n7279) );
  NOR2_X1 U8118 ( .A1(n7281), .A2(n6774), .ZN(n6773) );
  INV_X1 U8119 ( .A(n9308), .ZN(n6774) );
  OR2_X1 U8120 ( .A1(n7281), .A2(n6504), .ZN(n6776) );
  NOR2_X1 U8121 ( .A1(n9300), .A2(n7304), .ZN(n7303) );
  INV_X1 U8122 ( .A(n7305), .ZN(n7304) );
  NOR2_X1 U8123 ( .A1(n7308), .A2(n9300), .ZN(n7302) );
  AND2_X1 U8124 ( .A1(n8911), .A2(n8910), .ZN(n6614) );
  NAND2_X1 U8125 ( .A1(n12492), .A2(n6601), .ZN(n12495) );
  NAND2_X1 U8126 ( .A1(n8484), .A2(n8483), .ZN(n8498) );
  AND2_X1 U8127 ( .A1(n7178), .A2(n7181), .ZN(n7176) );
  NAND2_X1 U8128 ( .A1(n12382), .A2(n10385), .ZN(n8801) );
  INV_X1 U8129 ( .A(SI_12_), .ZN(n8327) );
  INV_X1 U8130 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n12101) );
  AND2_X1 U8131 ( .A1(n8685), .A2(n8687), .ZN(n7315) );
  AND2_X1 U8132 ( .A1(n7315), .A2(n8112), .ZN(n7314) );
  AOI21_X1 U8133 ( .B1(n7025), .B2(n7023), .A(n6595), .ZN(n7022) );
  INV_X1 U8134 ( .A(n7025), .ZN(n7024) );
  AND2_X1 U8135 ( .A1(n12861), .A2(n12988), .ZN(n12862) );
  OR2_X1 U8136 ( .A1(n12991), .A2(n12863), .ZN(n12861) );
  INV_X1 U8137 ( .A(n11171), .ZN(n6980) );
  INV_X1 U8138 ( .A(n12847), .ZN(n7000) );
  AND2_X1 U8139 ( .A1(n9184), .A2(n9180), .ZN(n7437) );
  NAND2_X1 U8140 ( .A1(n7227), .A2(n7229), .ZN(n6621) );
  NAND2_X1 U8141 ( .A1(n7228), .A2(n9186), .ZN(n7227) );
  NAND2_X1 U8142 ( .A1(n7224), .A2(n9247), .ZN(n6620) );
  INV_X1 U8143 ( .A(n9184), .ZN(n7226) );
  NAND2_X1 U8144 ( .A1(n9185), .A2(n9183), .ZN(n7225) );
  INV_X1 U8145 ( .A(n6870), .ZN(n6869) );
  NOR2_X1 U8146 ( .A1(n13345), .A2(n13421), .ZN(n6870) );
  AND2_X1 U8147 ( .A1(n6707), .A2(n13255), .ZN(n6706) );
  OR2_X1 U8148 ( .A1(n13435), .A2(n13439), .ZN(n6889) );
  INV_X1 U8149 ( .A(n7080), .ZN(n7079) );
  INV_X1 U8150 ( .A(n6486), .ZN(n7081) );
  NOR2_X1 U8151 ( .A1(n11565), .A2(n11467), .ZN(n6878) );
  NAND2_X1 U8152 ( .A1(n7076), .A2(n6490), .ZN(n7075) );
  AND2_X1 U8153 ( .A1(n6717), .A2(n11156), .ZN(n6716) );
  OR2_X1 U8154 ( .A1(n6492), .A2(n6718), .ZN(n6717) );
  INV_X1 U8155 ( .A(n7606), .ZN(n6718) );
  AND2_X1 U8156 ( .A1(n6885), .A2(n14965), .ZN(n6884) );
  INV_X1 U8157 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7450) );
  INV_X1 U8158 ( .A(n10876), .ZN(n7370) );
  INV_X1 U8159 ( .A(n7373), .ZN(n7372) );
  INV_X1 U8160 ( .A(n10236), .ZN(n10532) );
  INV_X1 U8161 ( .A(n12235), .ZN(n9575) );
  INV_X1 U8162 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9379) );
  INV_X1 U8163 ( .A(n14085), .ZN(n7208) );
  INV_X1 U8164 ( .A(n6499), .ZN(n7209) );
  AND2_X1 U8165 ( .A1(n6472), .A2(n7211), .ZN(n7206) );
  OR2_X1 U8166 ( .A1(n14212), .A2(n12014), .ZN(n13700) );
  NAND2_X1 U8167 ( .A1(n11121), .A2(n6473), .ZN(n6859) );
  NOR2_X1 U8168 ( .A1(n14564), .A2(n13649), .ZN(n6858) );
  INV_X1 U8169 ( .A(n11102), .ZN(n6955) );
  AND2_X1 U8170 ( .A1(n6935), .A2(n10627), .ZN(n6929) );
  INV_X1 U8171 ( .A(n6933), .ZN(n6930) );
  INV_X1 U8172 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10533) );
  NOR2_X1 U8173 ( .A1(n10245), .A2(n10244), .ZN(n10260) );
  NAND2_X1 U8174 ( .A1(n10220), .A2(n14734), .ZN(n13590) );
  INV_X1 U8175 ( .A(n12043), .ZN(n6937) );
  XOR2_X1 U8176 ( .A(n13741), .B(n13742), .Z(n13804) );
  INV_X1 U8177 ( .A(n6866), .ZN(n14153) );
  NOR2_X1 U8178 ( .A1(n9564), .A2(n6806), .ZN(n6805) );
  INV_X1 U8179 ( .A(n7275), .ZN(n7274) );
  AOI21_X1 U8180 ( .B1(n7275), .B2(n7273), .A(n7272), .ZN(n7271) );
  INV_X1 U8181 ( .A(n9141), .ZN(n7272) );
  INV_X1 U8182 ( .A(n9135), .ZN(n7273) );
  INV_X1 U8183 ( .A(n7914), .ZN(n7270) );
  AND2_X1 U8184 ( .A1(n7932), .A2(n7918), .ZN(n7930) );
  AOI21_X1 U8185 ( .B1(n7843), .B2(n7232), .A(n7852), .ZN(n7230) );
  AND2_X1 U8186 ( .A1(n9386), .A2(n9538), .ZN(n7342) );
  INV_X1 U8187 ( .A(n7841), .ZN(n7232) );
  XNOR2_X1 U8188 ( .A(n7702), .B(SI_13_), .ZN(n7701) );
  NAND2_X1 U8189 ( .A1(n7664), .A2(n8327), .ZN(n7678) );
  OR3_X1 U8190 ( .A1(n9613), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        P1_IR_REG_10__SCAN_IN), .ZN(n9677) );
  INV_X1 U8191 ( .A(n7642), .ZN(n7643) );
  NAND2_X1 U8192 ( .A1(n7661), .A2(n7650), .ZN(n7662) );
  NOR2_X1 U8193 ( .A1(n9526), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9533) );
  XNOR2_X1 U8194 ( .A(n7610), .B(SI_8_), .ZN(n7607) );
  INV_X1 U8195 ( .A(n7531), .ZN(n6843) );
  INV_X1 U8196 ( .A(n7547), .ZN(n6844) );
  OAI21_X1 U8197 ( .B1(n9582), .B2(n6699), .A(n6698), .ZN(n7515) );
  NAND2_X1 U8198 ( .A1(n9582), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6698) );
  OAI21_X1 U8199 ( .B1(P2_DATAO_REG_1__SCAN_IN), .B2(n9582), .A(n7458), .ZN(
        n7494) );
  NAND2_X1 U8200 ( .A1(n9582), .A2(n9478), .ZN(n7458) );
  AND2_X1 U8201 ( .A1(n6815), .A2(n6813), .ZN(n14294) );
  NAND2_X1 U8202 ( .A1(n7340), .A2(n6814), .ZN(n6813) );
  INV_X1 U8203 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6814) );
  XNOR2_X1 U8204 ( .A(n7339), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14329) );
  INV_X1 U8205 ( .A(n6823), .ZN(n14327) );
  OAI21_X1 U8206 ( .B1(n14354), .B2(n14355), .A(n6824), .ZN(n6823) );
  NAND2_X1 U8207 ( .A1(n14304), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6824) );
  NOR2_X1 U8208 ( .A1(n6807), .A2(n14308), .ZN(n14364) );
  NOR2_X1 U8209 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14362), .ZN(n6807) );
  NOR2_X1 U8210 ( .A1(n14625), .A2(n7327), .ZN(n7324) );
  NAND2_X1 U8211 ( .A1(n14625), .A2(n7327), .ZN(n7325) );
  INV_X1 U8212 ( .A(n7324), .ZN(n7320) );
  NOR2_X1 U8213 ( .A1(n7324), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7323) );
  OAI21_X1 U8214 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14312), .A(n14311), .ZN(
        n14368) );
  AOI21_X1 U8215 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n14314), .A(n14313), .ZN(
        n14324) );
  NOR2_X1 U8216 ( .A1(n14368), .A2(n14367), .ZN(n14313) );
  OAI21_X1 U8217 ( .B1(n14320), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n14319), .ZN(
        n14376) );
  OR2_X1 U8218 ( .A1(n14374), .A2(n14373), .ZN(n14319) );
  INV_X1 U8219 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10384) );
  NAND2_X1 U8220 ( .A1(n12306), .A2(n9309), .ZN(n12269) );
  INV_X1 U8221 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10637) );
  NAND2_X1 U8222 ( .A1(n7298), .A2(n12682), .ZN(n7297) );
  INV_X1 U8223 ( .A(n12287), .ZN(n7298) );
  OR2_X1 U8224 ( .A1(n8511), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8530) );
  INV_X1 U8225 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U8226 ( .A1(n7293), .A2(n7291), .ZN(n10461) );
  OR2_X1 U8227 ( .A1(n11203), .A2(n11204), .ZN(n11201) );
  NAND2_X1 U8228 ( .A1(n8273), .A2(n12142), .ZN(n8289) );
  INV_X1 U8229 ( .A(n8274), .ZN(n8273) );
  NAND2_X1 U8230 ( .A1(n9323), .A2(n9322), .ZN(n9326) );
  NAND2_X1 U8231 ( .A1(n11339), .A2(n9291), .ZN(n11636) );
  NAND2_X1 U8232 ( .A1(n7296), .A2(n7294), .ZN(n12328) );
  NOR2_X1 U8233 ( .A1(n11989), .A2(n7295), .ZN(n7294) );
  INV_X1 U8234 ( .A(n7297), .ZN(n7295) );
  INV_X1 U8235 ( .A(n8383), .ZN(n8382) );
  INV_X1 U8236 ( .A(n8943), .ZN(n8771) );
  AND4_X2 U8237 ( .A1(n8153), .A2(n8152), .A3(n8151), .A4(n8150), .ZN(n12760)
         );
  NAND2_X1 U8238 ( .A1(n9779), .A2(n9986), .ZN(n9778) );
  AOI21_X1 U8239 ( .B1(n10019), .B2(n10005), .A(n15029), .ZN(n15050) );
  AND2_X1 U8240 ( .A1(n10020), .A2(n15053), .ZN(n7123) );
  INV_X1 U8241 ( .A(n7122), .ZN(n10064) );
  XNOR2_X1 U8242 ( .A(n7120), .B(n10298), .ZN(n10066) );
  INV_X1 U8243 ( .A(n7115), .ZN(n10885) );
  NAND2_X1 U8244 ( .A1(n10886), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7114) );
  OAI21_X1 U8245 ( .B1(n15095), .B2(n15094), .A(n15093), .ZN(n15098) );
  OR2_X1 U8246 ( .A1(n6481), .A2(n12422), .ZN(n7106) );
  OR2_X1 U8247 ( .A1(n12387), .A2(n7107), .ZN(n7105) );
  OR2_X1 U8248 ( .A1(n12422), .A2(n8352), .ZN(n7107) );
  OR2_X1 U8249 ( .A1(n12387), .A2(n8352), .ZN(n7108) );
  NAND2_X1 U8250 ( .A1(n12411), .A2(n12412), .ZN(n12416) );
  NOR3_X1 U8251 ( .A1(n12424), .A2(n12423), .A3(n12425), .ZN(n12438) );
  NOR2_X1 U8252 ( .A1(n12441), .A2(n12442), .ZN(n12461) );
  AND3_X2 U8253 ( .A1(n7105), .A2(n6596), .A3(n7106), .ZN(n12451) );
  NOR2_X1 U8254 ( .A1(n12483), .A2(n7112), .ZN(n12484) );
  NOR2_X1 U8255 ( .A1(n12494), .A2(n12464), .ZN(n7112) );
  OR2_X2 U8256 ( .A1(n14447), .A2(n14448), .ZN(n7111) );
  XNOR2_X1 U8257 ( .A(n12495), .B(n14451), .ZN(n14450) );
  AOI21_X1 U8258 ( .B1(n12480), .B2(n14398), .A(n14455), .ZN(n12510) );
  NOR2_X1 U8259 ( .A1(n7172), .A2(n12555), .ZN(n7168) );
  NOR2_X1 U8260 ( .A1(n9368), .A2(n12683), .ZN(n8682) );
  NOR2_X1 U8261 ( .A1(n7064), .A2(n7063), .ZN(n7062) );
  INV_X1 U8262 ( .A(n7065), .ZN(n7064) );
  XNOR2_X1 U8263 ( .A(n8767), .B(n12539), .ZN(n8944) );
  NOR2_X1 U8264 ( .A1(n7067), .A2(n7066), .ZN(n7065) );
  INV_X1 U8265 ( .A(n8903), .ZN(n7066) );
  INV_X1 U8266 ( .A(n8908), .ZN(n7067) );
  NAND2_X1 U8267 ( .A1(n12551), .A2(n12550), .ZN(n7170) );
  AOI21_X1 U8268 ( .B1(n7170), .B2(n6497), .A(n12542), .ZN(n12537) );
  AND2_X1 U8269 ( .A1(n8550), .A2(n8549), .ZN(n12594) );
  NAND2_X1 U8270 ( .A1(n8542), .A2(n8541), .ZN(n8560) );
  INV_X1 U8271 ( .A(n8543), .ZN(n8542) );
  NAND2_X1 U8272 ( .A1(n8779), .A2(n8519), .ZN(n12608) );
  AND2_X1 U8273 ( .A1(n8887), .A2(n8888), .ZN(n12619) );
  NAND2_X1 U8274 ( .A1(n12653), .A2(n12658), .ZN(n12652) );
  NAND2_X1 U8275 ( .A1(n8460), .A2(n12262), .ZN(n8470) );
  AND2_X1 U8276 ( .A1(n8857), .A2(n8856), .ZN(n11665) );
  AOI21_X1 U8277 ( .B1(n7041), .B2(n7044), .A(n7039), .ZN(n7038) );
  INV_X1 U8278 ( .A(n8843), .ZN(n7044) );
  NAND2_X1 U8279 ( .A1(n8349), .A2(n11515), .ZN(n8365) );
  OR2_X1 U8280 ( .A1(n8365), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8383) );
  AOI21_X1 U8281 ( .B1(n7050), .B2(n7052), .A(n7048), .ZN(n7047) );
  INV_X1 U8282 ( .A(n8828), .ZN(n7048) );
  NAND2_X1 U8283 ( .A1(n8234), .A2(n10062), .ZN(n8254) );
  NAND2_X1 U8284 ( .A1(n7033), .A2(n7034), .ZN(n7031) );
  AND2_X1 U8285 ( .A1(n8817), .A2(n8816), .ZN(n10565) );
  NAND2_X1 U8286 ( .A1(n10130), .A2(n8632), .ZN(n10425) );
  AND2_X1 U8287 ( .A1(n8633), .A2(n8632), .ZN(n7198) );
  NAND2_X1 U8288 ( .A1(n10384), .A2(n10465), .ZN(n8200) );
  NAND2_X1 U8289 ( .A1(n8527), .A2(n8526), .ZN(n12297) );
  NAND2_X1 U8290 ( .A1(n8380), .A2(n8379), .ZN(n11666) );
  NAND2_X1 U8291 ( .A1(n8699), .A2(n8698), .ZN(n8701) );
  AND2_X1 U8292 ( .A1(n9732), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9490) );
  MUX2_X1 U8293 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8131), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n8133) );
  NAND2_X1 U8294 ( .A1(n7026), .A2(n8525), .ZN(n8537) );
  NAND2_X1 U8295 ( .A1(n8375), .A2(n8374), .ZN(n8392) );
  AND2_X1 U8296 ( .A1(n9695), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8321) );
  NOR2_X1 U8297 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8105) );
  NOR2_X1 U8298 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n6742) );
  NOR2_X1 U8299 ( .A1(n8268), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8284) );
  XNOR2_X1 U8300 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8280) );
  INV_X1 U8301 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8247) );
  XNOR2_X1 U8302 ( .A(n8231), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10060) );
  INV_X1 U8303 ( .A(n8226), .ZN(n8227) );
  XNOR2_X1 U8304 ( .A(n9503), .B(P2_DATAO_REG_5__SCAN_IN), .ZN(n8226) );
  XNOR2_X1 U8305 ( .A(n9504), .B(P2_DATAO_REG_4__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U8306 ( .A1(n9502), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8191) );
  INV_X1 U8307 ( .A(n8188), .ZN(n8189) );
  XNOR2_X1 U8308 ( .A(n9502), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n8188) );
  XNOR2_X1 U8309 ( .A(n9505), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n8169) );
  OAI22_X1 U8310 ( .A1(n8158), .A2(n7116), .B1(P3_IR_REG_31__SCAN_IN), .B2(
        P3_IR_REG_2__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U8311 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7116) );
  OAI22_X1 U8312 ( .A1(n7007), .A2(n12841), .B1(n12839), .B2(n12840), .ZN(
        n7006) );
  INV_X1 U8313 ( .A(n14487), .ZN(n7007) );
  INV_X1 U8314 ( .A(n12841), .ZN(n7008) );
  OR2_X1 U8315 ( .A1(n7634), .A2(n7633), .ZN(n7655) );
  AOI21_X1 U8316 ( .B1(n6991), .B2(n6990), .A(n6561), .ZN(n6989) );
  INV_X1 U8317 ( .A(n11276), .ZN(n6990) );
  INV_X1 U8318 ( .A(n11454), .ZN(n6992) );
  NAND2_X1 U8319 ( .A1(n6624), .A2(n6991), .ZN(n6988) );
  INV_X1 U8320 ( .A(n11275), .ZN(n6624) );
  AOI21_X1 U8321 ( .B1(n9820), .B2(P2_REG2_REG_3__SCAN_IN), .A(n13057), .ZN(
        n14849) );
  AOI21_X1 U8322 ( .B1(n9848), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9855), .ZN(
        n9863) );
  AOI21_X1 U8323 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n9955), .A(n9954), .ZN(
        n14891) );
  NAND2_X1 U8324 ( .A1(n14906), .A2(n10279), .ZN(n13092) );
  NOR2_X1 U8325 ( .A1(n12924), .A2(n12891), .ZN(n6669) );
  XNOR2_X1 U8326 ( .A(n13313), .B(n13023), .ZN(n9244) );
  NAND2_X1 U8327 ( .A1(n8016), .A2(n8015), .ZN(n13187) );
  NAND2_X1 U8328 ( .A1(n6487), .A2(n6910), .ZN(n6909) );
  NAND2_X1 U8329 ( .A1(n13228), .A2(n6487), .ZN(n6911) );
  NAND2_X1 U8330 ( .A1(n7878), .A2(n7863), .ZN(n6910) );
  NAND2_X1 U8331 ( .A1(n13248), .A2(n6870), .ZN(n13218) );
  AOI21_X1 U8332 ( .B1(n6837), .B2(n6838), .A(n6527), .ZN(n6834) );
  NAND2_X1 U8333 ( .A1(n6912), .A2(n13228), .ZN(n13230) );
  NAND2_X1 U8334 ( .A1(n13248), .A2(n13235), .ZN(n13234) );
  NOR2_X1 U8335 ( .A1(n11743), .A2(n6889), .ZN(n13293) );
  AOI21_X1 U8336 ( .B1(n6896), .B2(n11691), .A(n6895), .ZN(n6894) );
  NAND2_X1 U8337 ( .A1(n11690), .A2(n6896), .ZN(n6712) );
  INV_X1 U8338 ( .A(n9221), .ZN(n6895) );
  OR2_X1 U8339 ( .A1(n11686), .A2(n13399), .ZN(n11743) );
  NOR2_X1 U8340 ( .A1(n11743), .A2(n13439), .ZN(n13292) );
  AND2_X1 U8341 ( .A1(n11265), .A2(n6874), .ZN(n14506) );
  NOR2_X1 U8342 ( .A1(n14503), .A2(n6876), .ZN(n6874) );
  AOI21_X1 U8343 ( .B1(n7700), .B2(n6465), .A(n6515), .ZN(n6892) );
  NAND2_X1 U8344 ( .A1(n11265), .A2(n6878), .ZN(n11475) );
  NAND2_X1 U8345 ( .A1(n7071), .A2(n7070), .ZN(n11427) );
  NAND2_X1 U8346 ( .A1(n11265), .A2(n14987), .ZN(n11434) );
  AND2_X1 U8347 ( .A1(n7075), .A2(n6503), .ZN(n11242) );
  NAND2_X1 U8348 ( .A1(n7075), .A2(n7074), .ZN(n11240) );
  AND2_X1 U8349 ( .A1(n11263), .A2(n14977), .ZN(n11265) );
  AOI21_X1 U8350 ( .B1(n7086), .B2(n7089), .A(n6522), .ZN(n7085) );
  OR2_X1 U8351 ( .A1(n10978), .A2(n11173), .ZN(n11162) );
  NAND2_X1 U8352 ( .A1(n10802), .A2(n7986), .ZN(n10971) );
  NAND2_X1 U8353 ( .A1(n10804), .A2(n7586), .ZN(n10967) );
  NAND2_X1 U8354 ( .A1(n6676), .A2(n9229), .ZN(n10802) );
  NAND2_X1 U8355 ( .A1(n6882), .A2(n6880), .ZN(n10978) );
  AND2_X1 U8356 ( .A1(n6881), .A2(n6884), .ZN(n6880) );
  AND2_X1 U8357 ( .A1(n10927), .A2(n10839), .ZN(n6881) );
  OR2_X1 U8358 ( .A1(n10667), .A2(n6883), .ZN(n10656) );
  NAND2_X1 U8359 ( .A1(n10839), .A2(n6885), .ZN(n6883) );
  NOR2_X1 U8360 ( .A1(n10667), .A2(n6879), .ZN(n10806) );
  NAND2_X1 U8361 ( .A1(n6884), .A2(n10839), .ZN(n6879) );
  INV_X1 U8362 ( .A(n10502), .ZN(n10668) );
  OR2_X1 U8363 ( .A1(n10667), .A2(n10743), .ZN(n10665) );
  AND2_X1 U8364 ( .A1(n7012), .A2(n7786), .ZN(n7011) );
  INV_X1 U8365 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7010) );
  AND2_X1 U8366 ( .A1(n8035), .A2(n10450), .ZN(n10405) );
  NAND2_X1 U8367 ( .A1(n13313), .A2(n13398), .ZN(n6671) );
  OR2_X1 U8368 ( .A1(n6873), .A2(n6673), .ZN(n6672) );
  INV_X1 U8369 ( .A(n6674), .ZN(n6673) );
  NAND2_X1 U8370 ( .A1(n11775), .A2(n7612), .ZN(n7934) );
  INV_X1 U8371 ( .A(n14535), .ZN(n13371) );
  NOR2_X1 U8372 ( .A1(n8051), .A2(n13460), .ZN(n14952) );
  INV_X1 U8373 ( .A(n8037), .ZN(n8042) );
  AND2_X1 U8374 ( .A1(n7749), .A2(n7012), .ZN(n7787) );
  OR2_X1 U8375 ( .A1(n7592), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7594) );
  OR2_X1 U8376 ( .A1(n7594), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7615) );
  NAND3_X1 U8377 ( .A1(n7511), .A2(n7497), .A3(n7013), .ZN(n7559) );
  AND2_X1 U8378 ( .A1(n7525), .A2(n7445), .ZN(n7013) );
  NOR2_X1 U8379 ( .A1(n11845), .A2(n13485), .ZN(n11864) );
  NAND2_X1 U8380 ( .A1(n10937), .A2(n7374), .ZN(n7373) );
  INV_X1 U8381 ( .A(n10935), .ZN(n7374) );
  OR2_X1 U8382 ( .A1(n10534), .A2(n10533), .ZN(n10600) );
  NAND2_X1 U8383 ( .A1(n11864), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11883) );
  INV_X1 U8384 ( .A(n7365), .ZN(n6783) );
  INV_X1 U8385 ( .A(n13517), .ZN(n6782) );
  INV_X1 U8386 ( .A(n7364), .ZN(n6784) );
  NAND2_X1 U8387 ( .A1(n11914), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11944) );
  AND2_X1 U8388 ( .A1(n11586), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11704) );
  NAND2_X1 U8389 ( .A1(n11897), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11929) );
  INV_X1 U8390 ( .A(n11944), .ZN(n11928) );
  NAND2_X1 U8391 ( .A1(n11503), .A2(n11720), .ZN(n6795) );
  NOR2_X1 U8392 ( .A1(n11105), .A2(n11104), .ZN(n11226) );
  NAND2_X1 U8393 ( .A1(n13533), .A2(n13534), .ZN(n13532) );
  OR2_X1 U8394 ( .A1(n11020), .A2(n11504), .ZN(n11105) );
  NAND2_X1 U8395 ( .A1(n11704), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11830) );
  OR2_X1 U8396 ( .A1(n11830), .A2(n11829), .ZN(n11845) );
  NAND2_X1 U8397 ( .A1(n13509), .A2(n13510), .ZN(n13508) );
  NAND2_X1 U8398 ( .A1(n11928), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11960) );
  INV_X1 U8399 ( .A(n12223), .ZN(n11803) );
  OR2_X1 U8400 ( .A1(n11385), .A2(n11384), .ZN(n11533) );
  INV_X1 U8401 ( .A(n13806), .ZN(n7129) );
  NAND2_X1 U8402 ( .A1(n11961), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9724) );
  OR2_X1 U8403 ( .A1(n9520), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U8404 ( .A1(n14010), .A2(n6941), .ZN(n6940) );
  OR2_X1 U8405 ( .A1(n14187), .A2(n13823), .ZN(n7424) );
  NAND2_X1 U8406 ( .A1(n14043), .A2(n6860), .ZN(n14013) );
  NAND2_X1 U8407 ( .A1(n14043), .A2(n12046), .ZN(n14044) );
  NAND2_X1 U8408 ( .A1(n6864), .A2(n6863), .ZN(n14115) );
  NAND2_X1 U8409 ( .A1(n6863), .A2(n13577), .ZN(n7212) );
  XNOR2_X1 U8411 ( .A(n14233), .B(n13577), .ZN(n14112) );
  INV_X1 U8412 ( .A(n6960), .ZN(n6959) );
  NOR2_X1 U8413 ( .A1(n12039), .A2(n6963), .ZN(n6962) );
  NOR2_X1 U8414 ( .A1(n14110), .A2(n14112), .ZN(n14109) );
  INV_X1 U8415 ( .A(n13794), .ZN(n11700) );
  NOR2_X2 U8416 ( .A1(n6859), .A2(n14600), .ZN(n11597) );
  AOI21_X1 U8417 ( .B1(n6919), .B2(n6921), .A(n6549), .ZN(n6917) );
  NAND2_X1 U8418 ( .A1(n11121), .A2(n6858), .ZN(n11383) );
  NAND2_X1 U8419 ( .A1(n11121), .A2(n14607), .ZN(n11224) );
  OR2_X1 U8420 ( .A1(n13640), .A2(n13839), .ZN(n11117) );
  INV_X1 U8421 ( .A(n11017), .ZN(n6957) );
  OR2_X1 U8422 ( .A1(n14787), .A2(n13841), .ZN(n10994) );
  OR2_X1 U8423 ( .A1(n10600), .A2(n10599), .ZN(n10609) );
  NOR2_X1 U8424 ( .A1(n10243), .A2(n6924), .ZN(n6923) );
  INV_X1 U8425 ( .A(n10230), .ZN(n6924) );
  OAI22_X1 U8426 ( .A1(n14704), .A2(n14706), .B1(n6457), .B2(n13845), .ZN(
        n10481) );
  NAND2_X1 U8427 ( .A1(n9585), .A2(n10257), .ZN(n14722) );
  XNOR2_X1 U8429 ( .A(n7915), .B(n7914), .ZN(n13462) );
  XNOR2_X1 U8430 ( .A(n7785), .B(n7780), .ZN(n11816) );
  NAND2_X1 U8431 ( .A1(n7767), .A2(n7766), .ZN(n7785) );
  NAND2_X1 U8432 ( .A1(n7254), .A2(n7704), .ZN(n7722) );
  NAND2_X1 U8433 ( .A1(n7679), .A2(n7262), .ZN(n7254) );
  XNOR2_X1 U8434 ( .A(n7706), .B(n7701), .ZN(n11375) );
  NAND2_X1 U8435 ( .A1(n7679), .A2(n7678), .ZN(n7706) );
  XNOR2_X1 U8436 ( .A(n7563), .B(SI_5_), .ZN(n7561) );
  INV_X1 U8437 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9383) );
  INV_X1 U8438 ( .A(n9412), .ZN(n9384) );
  XNOR2_X1 U8439 ( .A(n7494), .B(SI_1_), .ZN(n7496) );
  NAND2_X1 U8440 ( .A1(n8134), .A2(n7459), .ZN(n9584) );
  NAND2_X1 U8441 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n9511), .ZN(n14335) );
  INV_X1 U8442 ( .A(n7340), .ZN(n14331) );
  XNOR2_X1 U8443 ( .A(n14329), .B(n7338), .ZN(n14330) );
  INV_X1 U8444 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U8445 ( .A1(n15137), .A2(n14345), .ZN(n14346) );
  AND2_X1 U8446 ( .A1(n6811), .A2(n6573), .ZN(n14348) );
  OR2_X1 U8447 ( .A1(n14342), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6811) );
  NOR2_X1 U8448 ( .A1(n15141), .A2(n14353), .ZN(n14356) );
  XNOR2_X1 U8449 ( .A(n14307), .B(n6808), .ZN(n14362) );
  AND2_X1 U8450 ( .A1(n7328), .A2(n14429), .ZN(n14366) );
  OAI21_X1 U8451 ( .B1(n14430), .B2(n14431), .A(n7329), .ZN(n7328) );
  INV_X1 U8452 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7329) );
  NOR2_X1 U8453 ( .A1(n14629), .A2(n14370), .ZN(n14371) );
  INV_X1 U8454 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7337) );
  AND4_X1 U8455 ( .A1(n8225), .A2(n8224), .A3(n8223), .A4(n8222), .ZN(n10862)
         );
  NOR2_X1 U8456 ( .A1(n6520), .A2(n7284), .ZN(n7283) );
  INV_X1 U8457 ( .A(n7286), .ZN(n7284) );
  NAND2_X1 U8458 ( .A1(n7286), .A2(n7287), .ZN(n7285) );
  INV_X1 U8459 ( .A(n9343), .ZN(n7287) );
  OAI21_X1 U8460 ( .B1(n11339), .B2(n7307), .A(n7305), .ZN(n11627) );
  AND2_X1 U8461 ( .A1(n8536), .A2(n8535), .ZN(n12607) );
  NAND2_X1 U8462 ( .A1(n6767), .A2(n6770), .ZN(n10381) );
  AND2_X1 U8463 ( .A1(n6777), .A2(n6504), .ZN(n12306) );
  NAND2_X1 U8464 ( .A1(n12328), .A2(n9308), .ZN(n6777) );
  NAND2_X1 U8465 ( .A1(n9266), .A2(n12384), .ZN(n9270) );
  INV_X1 U8466 ( .A(n9268), .ZN(n9266) );
  NAND2_X1 U8467 ( .A1(n8482), .A2(n8481), .ZN(n12631) );
  NAND2_X1 U8468 ( .A1(n10461), .A2(n9278), .ZN(n10636) );
  NAND2_X1 U8469 ( .A1(n7296), .A2(n7297), .ZN(n11990) );
  INV_X1 U8470 ( .A(n6757), .ZN(n6759) );
  NAND2_X1 U8471 ( .A1(n7310), .A2(n9296), .ZN(n11513) );
  NAND2_X1 U8472 ( .A1(n11339), .A2(n7311), .ZN(n7310) );
  NAND2_X1 U8473 ( .A1(n8497), .A2(n8496), .ZN(n12324) );
  AND4_X1 U8474 ( .A1(n8310), .A2(n8309), .A3(n8308), .A4(n8307), .ZN(n11646)
         );
  INV_X1 U8475 ( .A(n10183), .ZN(n10078) );
  INV_X1 U8476 ( .A(n12354), .ZN(n12311) );
  NAND2_X1 U8477 ( .A1(n7289), .A2(n6526), .ZN(n7288) );
  AND2_X1 U8478 ( .A1(n9348), .A2(n15111), .ZN(n12360) );
  NAND2_X1 U8479 ( .A1(n9360), .A2(n9359), .ZN(n12356) );
  NAND2_X1 U8480 ( .A1(n6765), .A2(n6764), .ZN(n12350) );
  INV_X1 U8481 ( .A(n12348), .ZN(n6764) );
  NAND2_X1 U8482 ( .A1(n8922), .A2(n8923), .ZN(n7020) );
  OR2_X1 U8483 ( .A1(n8922), .A2(n15109), .ZN(n7021) );
  NAND2_X1 U8484 ( .A1(n8567), .A2(n8566), .ZN(n12578) );
  INV_X1 U8485 ( .A(n12594), .ZN(n12362) );
  INV_X1 U8486 ( .A(n11646), .ZN(n12374) );
  NAND4_X2 U8487 ( .A1(n8126), .A2(n8125), .A3(n8124), .A4(n8123), .ZN(n12757)
         );
  OAI21_X1 U8488 ( .B1(n6493), .B2(n10010), .A(n6731), .ZN(n10012) );
  NOR2_X1 U8489 ( .A1(n6737), .A2(n15057), .ZN(n6733) );
  NAND2_X1 U8490 ( .A1(n10299), .A2(n10300), .ZN(n10303) );
  NAND2_X1 U8491 ( .A1(n15076), .A2(n10909), .ZN(n15083) );
  INV_X1 U8492 ( .A(n7119), .ZN(n15088) );
  NAND2_X1 U8493 ( .A1(n11138), .A2(n11139), .ZN(n11140) );
  NOR2_X1 U8494 ( .A1(n11132), .A2(n11133), .ZN(n11135) );
  INV_X1 U8495 ( .A(n7117), .ZN(n11131) );
  XNOR2_X1 U8496 ( .A(n12404), .B(n12405), .ZN(n12387) );
  NAND2_X1 U8497 ( .A1(n7105), .A2(n7106), .ZN(n12432) );
  AND2_X1 U8498 ( .A1(n7108), .A2(n6481), .ZN(n12409) );
  NAND2_X1 U8499 ( .A1(n12457), .A2(n12458), .ZN(n12459) );
  INV_X1 U8500 ( .A(n7111), .ZN(n14446) );
  INV_X1 U8501 ( .A(n12516), .ZN(n6726) );
  NAND2_X1 U8502 ( .A1(n12556), .A2(n12555), .ZN(n12554) );
  NAND2_X1 U8503 ( .A1(n7053), .A2(n7057), .ZN(n12593) );
  NAND2_X1 U8504 ( .A1(n12620), .A2(n7056), .ZN(n7053) );
  NAND2_X1 U8505 ( .A1(n12637), .A2(n8664), .ZN(n12626) );
  NAND2_X1 U8506 ( .A1(n12642), .A2(n8881), .ZN(n12630) );
  NAND2_X1 U8507 ( .A1(n8443), .A2(n8442), .ZN(n12739) );
  NAND2_X1 U8508 ( .A1(n7173), .A2(n7179), .ZN(n12678) );
  NAND2_X1 U8509 ( .A1(n11441), .A2(n7182), .ZN(n7173) );
  NAND2_X1 U8510 ( .A1(n7184), .A2(n8658), .ZN(n11602) );
  NAND2_X1 U8511 ( .A1(n7185), .A2(n6489), .ZN(n7184) );
  NAND2_X1 U8512 ( .A1(n11329), .A2(n8843), .ZN(n11490) );
  AND2_X1 U8513 ( .A1(n11041), .A2(n8639), .ZN(n11072) );
  NAND2_X1 U8514 ( .A1(n11038), .A2(n8825), .ZN(n11069) );
  AND2_X1 U8515 ( .A1(n10814), .A2(n8638), .ZN(n11043) );
  NAND2_X1 U8516 ( .A1(n10137), .A2(n8806), .ZN(n10422) );
  OR2_X1 U8517 ( .A1(n9983), .A2(n9978), .ZN(n12689) );
  INV_X1 U8518 ( .A(n12689), .ZN(n14463) );
  AND3_X1 U8519 ( .A1(n8253), .A2(n8252), .A3(n8251), .ZN(n10820) );
  NOR2_X1 U8520 ( .A1(n12525), .A2(n12524), .ZN(n14466) );
  INV_X1 U8521 ( .A(n12324), .ZN(n12796) );
  AND2_X1 U8522 ( .A1(n12736), .A2(n12735), .ZN(n12806) );
  NAND2_X1 U8523 ( .A1(n8421), .A2(n8420), .ZN(n12813) );
  NAND2_X1 U8524 ( .A1(n8364), .A2(n8363), .ZN(n11630) );
  AND2_X1 U8525 ( .A1(n8320), .A2(n8319), .ZN(n11560) );
  OAI211_X1 U8526 ( .C1(n8288), .C2(SI_9_), .A(n8287), .B(n8286), .ZN(n11206)
         );
  INV_X1 U8527 ( .A(n11092), .ZN(n11094) );
  INV_X1 U8528 ( .A(n10114), .ZN(n12001) );
  AND2_X1 U8529 ( .A1(n8701), .A2(n8700), .ZN(n12822) );
  CLKBUF_X1 U8530 ( .A(n12476), .Z(n6622) );
  INV_X1 U8531 ( .A(n8717), .ZN(n11325) );
  NAND2_X1 U8532 ( .A1(n8616), .A2(n8615), .ZN(n10500) );
  NAND2_X1 U8533 ( .A1(n8453), .A2(n8452), .ZN(n8467) );
  NAND2_X1 U8534 ( .A1(n7029), .A2(n8358), .ZN(n8357) );
  NOR2_X1 U8535 ( .A1(n8159), .A2(n8361), .ZN(n8174) );
  OAI21_X1 U8536 ( .B1(n10837), .B2(n6984), .A(n6982), .ZN(n11172) );
  NOR2_X1 U8537 ( .A1(n14486), .A2(n14487), .ZN(n14485) );
  XNOR2_X1 U8538 ( .A(n12867), .B(n12865), .ZN(n12896) );
  NAND2_X1 U8539 ( .A1(n11302), .A2(n11301), .ZN(n11456) );
  NAND2_X1 U8540 ( .A1(n6996), .A2(n6995), .ZN(n12906) );
  AND2_X1 U8541 ( .A1(n6996), .A2(n6509), .ZN(n12908) );
  NAND2_X1 U8542 ( .A1(n6997), .A2(n6998), .ZN(n6996) );
  INV_X1 U8543 ( .A(n6972), .ZN(n10124) );
  NAND2_X1 U8544 ( .A1(n12928), .A2(n12927), .ZN(n12989) );
  NAND2_X1 U8545 ( .A1(n7005), .A2(n7003), .ZN(n12945) );
  INV_X1 U8546 ( .A(n7006), .ZN(n7003) );
  NAND2_X1 U8547 ( .A1(n14486), .A2(n7008), .ZN(n7005) );
  INV_X1 U8548 ( .A(n14490), .ZN(n12957) );
  NAND2_X1 U8549 ( .A1(n6993), .A2(n6994), .ZN(n12980) );
  AOI21_X1 U8550 ( .B1(n6995), .B2(n13001), .A(n12855), .ZN(n6994) );
  NAND2_X1 U8551 ( .A1(n6988), .A2(n6989), .ZN(n11461) );
  NAND2_X1 U8552 ( .A1(n10849), .A2(n10848), .ZN(n10948) );
  NOR2_X1 U8553 ( .A1(n13009), .A2(n12876), .ZN(n6999) );
  NAND2_X1 U8554 ( .A1(n12937), .A2(n12877), .ZN(n13010) );
  INV_X1 U8555 ( .A(n11418), .ZN(n6643) );
  NAND2_X1 U8556 ( .A1(n9148), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7540) );
  OR2_X1 U8557 ( .A1(n7487), .A2(n7488), .ZN(n7490) );
  OR2_X1 U8558 ( .A1(n9152), .A2(n7470), .ZN(n7475) );
  OR2_X1 U8559 ( .A1(n9152), .A2(n10119), .ZN(n7480) );
  NAND2_X1 U8560 ( .A1(n7506), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7477) );
  OAI21_X1 U8561 ( .B1(n14863), .B2(n13073), .A(n9795), .ZN(n13076) );
  XNOR2_X1 U8562 ( .A(n13092), .B(n6659), .ZN(n10280) );
  NAND2_X1 U8563 ( .A1(n13100), .A2(n13101), .ZN(n13105) );
  NOR2_X1 U8564 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13107), .ZN(n13126) );
  NOR2_X1 U8565 ( .A1(n6908), .A2(n6904), .ZN(n6903) );
  INV_X1 U8566 ( .A(n7928), .ZN(n6904) );
  NAND2_X1 U8567 ( .A1(n6905), .A2(n7928), .ZN(n13160) );
  NAND2_X1 U8568 ( .A1(n7912), .A2(n7911), .ZN(n13172) );
  INV_X1 U8569 ( .A(n6836), .ZN(n13229) );
  AOI21_X1 U8570 ( .B1(n7090), .B2(n7091), .A(n6838), .ZN(n6836) );
  OAI21_X1 U8571 ( .B1(n13279), .B2(n7095), .A(n7093), .ZN(n13256) );
  NAND2_X1 U8572 ( .A1(n6702), .A2(n6707), .ZN(n13244) );
  OR2_X1 U8573 ( .A1(n13273), .A2(n6710), .ZN(n6702) );
  NAND2_X1 U8574 ( .A1(n6711), .A2(n7816), .ZN(n13269) );
  NAND2_X1 U8575 ( .A1(n13273), .A2(n7815), .ZN(n6711) );
  NAND2_X1 U8576 ( .A1(n7092), .A2(n8009), .ZN(n13260) );
  NAND2_X1 U8577 ( .A1(n13279), .A2(n8007), .ZN(n7092) );
  NAND2_X1 U8578 ( .A1(n11841), .A2(n7612), .ZN(n7810) );
  NAND2_X1 U8579 ( .A1(n7762), .A2(n7761), .ZN(n13401) );
  NAND2_X1 U8580 ( .A1(n7078), .A2(n6486), .ZN(n11673) );
  NAND2_X1 U8581 ( .A1(n7995), .A2(n7082), .ZN(n7078) );
  NAND2_X1 U8582 ( .A1(n7995), .A2(n9233), .ZN(n14496) );
  OR2_X1 U8583 ( .A1(n11239), .A2(n6465), .ZN(n11471) );
  NAND2_X1 U8584 ( .A1(n6846), .A2(n7630), .ZN(n11308) );
  NAND2_X1 U8585 ( .A1(n11001), .A2(n7612), .ZN(n6846) );
  NAND2_X1 U8586 ( .A1(n10969), .A2(n7606), .ZN(n11155) );
  INV_X1 U8587 ( .A(n13205), .ZN(n14502) );
  INV_X1 U8588 ( .A(n14509), .ZN(n13302) );
  OR2_X1 U8589 ( .A1(n9884), .A2(n14961), .ZN(n13295) );
  NAND2_X1 U8590 ( .A1(n7618), .A2(n7617), .ZN(n11316) );
  NAND2_X1 U8591 ( .A1(n13148), .A2(n6645), .ZN(n13411) );
  INV_X1 U8592 ( .A(n10954), .ZN(n10927) );
  NOR2_X1 U8593 ( .A1(n9886), .A2(P2_U3088), .ZN(n14959) );
  INV_X1 U8594 ( .A(n14959), .ZN(n14961) );
  NAND2_X1 U8595 ( .A1(n7463), .A2(n6914), .ZN(n6913) );
  NOR2_X1 U8596 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6914) );
  NAND2_X1 U8597 ( .A1(n7452), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7453) );
  OAI21_X1 U8598 ( .B1(n6901), .B2(n6900), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7969) );
  INV_X1 U8599 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10472) );
  INV_X1 U8600 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10459) );
  AND2_X1 U8601 ( .A1(n7749), .A2(n7748), .ZN(n7769) );
  INV_X1 U8602 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10178) );
  INV_X1 U8603 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9840) );
  INV_X1 U8604 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9692) );
  INV_X1 U8605 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9501) );
  INV_X1 U8606 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9503) );
  INV_X1 U8607 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U8608 ( .A1(n7524), .A2(n7511), .ZN(n7544) );
  INV_X1 U8609 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9502) );
  INV_X2 U8610 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9505) );
  XNOR2_X1 U8611 ( .A(n7457), .B(n7456), .ZN(n9815) );
  NAND2_X1 U8612 ( .A1(n6803), .A2(n10873), .ZN(n10875) );
  NOR2_X1 U8613 ( .A1(n10875), .A2(n10876), .ZN(n10936) );
  NAND2_X1 U8614 ( .A1(n13532), .A2(n11910), .ZN(n13470) );
  NAND2_X1 U8615 ( .A1(n6804), .A2(n7360), .ZN(n13480) );
  NAND2_X1 U8616 ( .A1(n7355), .A2(n7351), .ZN(n7350) );
  NAND2_X1 U8617 ( .A1(n12227), .A2(n7352), .ZN(n7351) );
  INV_X1 U8618 ( .A(n7356), .ZN(n7352) );
  NAND2_X1 U8619 ( .A1(n7355), .A2(n12227), .ZN(n7354) );
  OR2_X1 U8620 ( .A1(n10936), .A2(n7373), .ZN(n11289) );
  NAND2_X1 U8621 ( .A1(n13523), .A2(n11879), .ZN(n13491) );
  OAI21_X1 U8622 ( .B1(n14650), .B2(n6464), .A(n6470), .ZN(n10520) );
  NAND2_X1 U8623 ( .A1(n13533), .A2(n7365), .ZN(n6780) );
  NAND2_X2 U8624 ( .A1(n11927), .A2(n11926), .ZN(n14200) );
  NAND2_X1 U8625 ( .A1(n13465), .A2(n13756), .ZN(n11927) );
  NAND2_X1 U8626 ( .A1(n7345), .A2(n7344), .ZN(n10389) );
  NOR2_X1 U8627 ( .A1(n10340), .A2(n7348), .ZN(n7344) );
  INV_X1 U8628 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11504) );
  NAND2_X1 U8629 ( .A1(n6792), .A2(n6791), .ZN(n6790) );
  INV_X1 U8630 ( .A(n11497), .ZN(n6792) );
  OR2_X1 U8631 ( .A1(n9919), .A2(n9918), .ZN(n9920) );
  NAND2_X1 U8632 ( .A1(n13508), .A2(n11825), .ZN(n13541) );
  NAND2_X1 U8633 ( .A1(n6801), .A2(n6800), .ZN(n10874) );
  NAND2_X1 U8634 ( .A1(n13457), .A2(n13756), .ZN(n11958) );
  INV_X1 U8635 ( .A(n14578), .ZN(n14649) );
  AND2_X1 U8636 ( .A1(n13810), .A2(n13811), .ZN(n6688) );
  NAND2_X1 U8637 ( .A1(n6855), .A2(n14730), .ZN(n14161) );
  XNOR2_X1 U8638 ( .A(n13967), .B(n6856), .ZN(n6855) );
  INV_X1 U8639 ( .A(n13973), .ZN(n14164) );
  INV_X1 U8640 ( .A(n12064), .ZN(n12065) );
  NAND2_X1 U8641 ( .A1(n7221), .A2(n7220), .ZN(n13985) );
  INV_X1 U8642 ( .A(n7222), .ZN(n6690) );
  NAND2_X1 U8643 ( .A1(n7201), .A2(n7202), .ZN(n14024) );
  NAND2_X1 U8644 ( .A1(n14037), .A2(n6950), .ZN(n14021) );
  NAND2_X1 U8645 ( .A1(n14288), .A2(n6458), .ZN(n14080) );
  NAND2_X1 U8646 ( .A1(n11882), .A2(n11881), .ZN(n14090) );
  NAND2_X1 U8647 ( .A1(n11863), .A2(n11862), .ZN(n14105) );
  OAI21_X1 U8648 ( .B1(n11699), .B2(n6965), .A(n6964), .ZN(n14127) );
  NOR2_X1 U8649 ( .A1(n12037), .A2(n12036), .ZN(n14147) );
  INV_X1 U8650 ( .A(n7200), .ZN(n14143) );
  NAND2_X1 U8651 ( .A1(n11697), .A2(n11696), .ZN(n14575) );
  NAND2_X1 U8652 ( .A1(n11583), .A2(n11582), .ZN(n11799) );
  NAND2_X1 U8653 ( .A1(n11529), .A2(n7215), .ZN(n7431) );
  OAI21_X1 U8654 ( .B1(n11219), .B2(n6921), .A(n6919), .ZN(n11522) );
  NAND2_X1 U8655 ( .A1(n11374), .A2(n11373), .ZN(n11379) );
  NAND2_X1 U8656 ( .A1(n11055), .A2(n11017), .ZN(n11018) );
  NAND2_X1 U8657 ( .A1(n10999), .A2(n10998), .ZN(n14698) );
  NAND2_X1 U8658 ( .A1(n10593), .A2(n10592), .ZN(n13620) );
  NAND2_X1 U8659 ( .A1(n6934), .A2(n6933), .ZN(n10758) );
  NAND2_X1 U8660 ( .A1(n14116), .A2(n12057), .ZN(n14120) );
  INV_X1 U8661 ( .A(n14728), .ZN(n14116) );
  INV_X1 U8662 ( .A(n14160), .ZN(n14124) );
  NAND2_X1 U8663 ( .A1(n14161), .A2(n6853), .ZN(n14255) );
  INV_X1 U8664 ( .A(n6854), .ZN(n6853) );
  OAI21_X1 U8665 ( .B1(n6856), .B2(n14799), .A(n14162), .ZN(n6854) );
  INV_X1 U8666 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U8667 ( .A1(n7277), .A2(n7275), .ZN(n9189) );
  NOR2_X1 U8668 ( .A1(n9568), .A2(n6548), .ZN(n6654) );
  NAND2_X1 U8669 ( .A1(n9540), .A2(n9386), .ZN(n7343) );
  INV_X1 U8670 ( .A(n9540), .ZN(n9541) );
  INV_X1 U8671 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10436) );
  INV_X1 U8672 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10176) );
  INV_X1 U8673 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9695) );
  INV_X1 U8674 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9599) );
  INV_X1 U8675 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9529) );
  INV_X1 U8676 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9522) );
  INV_X1 U8677 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9496) );
  INV_X1 U8678 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9493) );
  INV_X1 U8679 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10232) );
  INV_X1 U8680 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9492) );
  XNOR2_X1 U8681 ( .A(n14330), .B(n14853), .ZN(n15136) );
  XNOR2_X1 U8682 ( .A(n6681), .B(n14344), .ZN(n15139) );
  INV_X1 U8683 ( .A(n14343), .ZN(n6681) );
  NAND2_X1 U8684 ( .A1(n15139), .A2(n15138), .ZN(n15137) );
  XNOR2_X1 U8685 ( .A(n14346), .B(n6682), .ZN(n14412) );
  XNOR2_X1 U8686 ( .A(n14352), .B(n14881), .ZN(n15142) );
  NOR2_X1 U8687 ( .A1(n15142), .A2(n15143), .ZN(n15141) );
  XNOR2_X1 U8688 ( .A(n14356), .B(n6685), .ZN(n14420) );
  INV_X1 U8689 ( .A(n14357), .ZN(n6685) );
  NAND2_X1 U8690 ( .A1(n14420), .A2(n9846), .ZN(n14419) );
  INV_X1 U8691 ( .A(n6821), .ZN(n14443) );
  AND2_X1 U8692 ( .A1(n6821), .A2(n6820), .ZN(n14442) );
  OAI211_X1 U8693 ( .C1(n6750), .C2(n6745), .A(n6744), .B(n6743), .ZN(P3_U3160) );
  INV_X1 U8694 ( .A(n6749), .ZN(n6745) );
  NAND2_X1 U8695 ( .A1(n6750), .A2(n6748), .ZN(n6744) );
  AOI21_X1 U8696 ( .B1(n6725), .B2(n15086), .A(n6723), .ZN(n12522) );
  XNOR2_X1 U8697 ( .A(n6727), .B(n6726), .ZN(n6725) );
  NOR2_X1 U8698 ( .A1(n6514), .A2(n6649), .ZN(n6648) );
  NOR2_X1 U8699 ( .A1(n15133), .A2(n8742), .ZN(n6649) );
  AOI21_X1 U8700 ( .B1(n6668), .B2(n8743), .A(n6667), .ZN(n6666) );
  NOR2_X1 U8701 ( .A1(n15133), .A2(n12700), .ZN(n6667) );
  NOR2_X1 U8702 ( .A1(n6517), .A2(n6652), .ZN(n6651) );
  NOR2_X1 U8703 ( .A1(n15129), .A2(n8726), .ZN(n6652) );
  OAI21_X1 U8704 ( .B1(n12777), .B2(n15127), .A(n6552), .ZN(P3_U3455) );
  NAND2_X1 U8705 ( .A1(n15127), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n6625) );
  INV_X1 U8706 ( .A(n6976), .ZN(n10325) );
  INV_X1 U8707 ( .A(n8099), .ZN(n8103) );
  OAI21_X1 U8708 ( .B1(n13315), .B2(n14951), .A(n8098), .ZN(n8099) );
  NAND2_X1 U8709 ( .A1(n6604), .A2(n6603), .ZN(P2_U3530) );
  NAND2_X1 U8710 ( .A1(n13138), .A2(n8070), .ZN(n6603) );
  INV_X1 U8711 ( .A(n11988), .ZN(n6604) );
  NAND2_X1 U8712 ( .A1(n13410), .A2(n15002), .ZN(n6619) );
  INV_X1 U8713 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U8714 ( .A1(n6606), .A2(n6605), .ZN(P2_U3498) );
  NAND2_X1 U8715 ( .A1(n13138), .A2(n13440), .ZN(n6605) );
  INV_X1 U8716 ( .A(n12217), .ZN(n6606) );
  MUX2_X1 U8717 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n12216), .S(n10105), .Z(
        n12217) );
  NAND2_X1 U8718 ( .A1(n14991), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U8719 ( .A1(n13410), .A2(n10105), .ZN(n6891) );
  XNOR2_X1 U8720 ( .A(n6798), .B(n6797), .ZN(n11985) );
  NAND2_X1 U8721 ( .A1(n11721), .A2(n11720), .ZN(n14563) );
  OR2_X1 U8722 ( .A1(n14819), .A2(n6927), .ZN(n6926) );
  INV_X1 U8723 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6927) );
  INV_X1 U8724 ( .A(n6850), .ZN(P1_U3527) );
  AOI21_X1 U8725 ( .B1(n14255), .B2(n14807), .A(n6851), .ZN(n6850) );
  NOR2_X1 U8726 ( .A1(n14807), .A2(n6852), .ZN(n6851) );
  INV_X1 U8727 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U8728 ( .A1(n14626), .A2(n14625), .ZN(n14624) );
  NAND2_X1 U8729 ( .A1(n7326), .A2(n14621), .ZN(n14626) );
  NAND2_X1 U8730 ( .A1(n14633), .A2(n14635), .ZN(n14639) );
  AND3_X1 U8731 ( .A1(n14633), .A2(n14635), .A3(n7335), .ZN(n14638) );
  NAND2_X1 U8732 ( .A1(n7331), .A2(n7334), .ZN(n14643) );
  INV_X2 U8733 ( .A(n9088), .ZN(n9204) );
  NAND2_X1 U8734 ( .A1(n10339), .A2(n7347), .ZN(n6464) );
  INV_X1 U8735 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13444) );
  OAI211_X1 U8736 ( .C1(n9803), .C2(n14858), .A(n7552), .B(n7551), .ZN(n10831)
         );
  OR2_X1 U8737 ( .A1(n11421), .A2(n7698), .ZN(n6465) );
  INV_X1 U8738 ( .A(n10341), .ZN(n7348) );
  INV_X1 U8739 ( .A(n10010), .ZN(n15053) );
  AND2_X1 U8740 ( .A1(n6762), .A2(n12618), .ZN(n6466) );
  AND2_X1 U8741 ( .A1(n6675), .A2(n7984), .ZN(n6467) );
  NAND2_X1 U8742 ( .A1(n13995), .A2(n6498), .ZN(n6468) );
  AND2_X1 U8743 ( .A1(n9055), .A2(n9054), .ZN(n6469) );
  INV_X1 U8744 ( .A(n14038), .ZN(n6948) );
  OR2_X1 U8745 ( .A1(n14243), .A2(n13543), .ZN(n13682) );
  OR2_X1 U8746 ( .A1(n10390), .A2(n7348), .ZN(n6470) );
  OR2_X1 U8747 ( .A1(n12610), .A2(n12618), .ZN(n8779) );
  AND2_X1 U8748 ( .A1(n6499), .A2(n7210), .ZN(n6471) );
  AND2_X1 U8749 ( .A1(n13800), .A2(n7212), .ZN(n6472) );
  NAND2_X2 U8750 ( .A1(n8957), .A2(n9249), .ZN(n8981) );
  INV_X1 U8751 ( .A(n13001), .ZN(n6998) );
  NAND2_X1 U8752 ( .A1(n8881), .A2(n8882), .ZN(n12645) );
  INV_X1 U8753 ( .A(n12645), .ZN(n7187) );
  AND2_X1 U8754 ( .A1(n6858), .A2(n6857), .ZN(n6473) );
  AND2_X1 U8755 ( .A1(n6729), .A2(n15053), .ZN(n6474) );
  AND2_X1 U8756 ( .A1(n13620), .A2(n10628), .ZN(n6475) );
  INV_X1 U8757 ( .A(n13663), .ZN(n7147) );
  INV_X1 U8758 ( .A(n9925), .ZN(n11109) );
  NAND2_X1 U8759 ( .A1(n7416), .A2(n7415), .ZN(n6476) );
  NOR2_X1 U8760 ( .A1(n11585), .A2(n11789), .ZN(n6477) );
  INV_X1 U8761 ( .A(n13669), .ZN(n7217) );
  AND2_X1 U8762 ( .A1(n9031), .A2(n9030), .ZN(n6478) );
  INV_X1 U8763 ( .A(n14145), .ZN(n6680) );
  AND2_X1 U8764 ( .A1(n11055), .A2(n6956), .ZN(n6479) );
  CLKBUF_X1 U8765 ( .A(n14734), .Z(n6656) );
  AND2_X1 U8766 ( .A1(n7321), .A2(n7319), .ZN(n6480) );
  INV_X1 U8767 ( .A(n13822), .ZN(n12228) );
  NAND2_X1 U8768 ( .A1(n7317), .A2(n9260), .ZN(n9283) );
  INV_X1 U8769 ( .A(n9229), .ZN(n7088) );
  OR2_X1 U8770 ( .A1(n12405), .A2(n12404), .ZN(n6481) );
  INV_X1 U8771 ( .A(n13717), .ZN(n14187) );
  NAND2_X1 U8772 ( .A1(n8617), .A2(n8111), .ZN(n8613) );
  AND2_X1 U8773 ( .A1(n6758), .A2(n6759), .ZN(n6482) );
  AND2_X1 U8774 ( .A1(n6687), .A2(n6686), .ZN(n6483) );
  AND2_X1 U8775 ( .A1(n14043), .A2(n6862), .ZN(n6484) );
  NAND2_X1 U8776 ( .A1(n7965), .A2(n7449), .ZN(n6485) );
  INV_X1 U8777 ( .A(n12555), .ZN(n12550) );
  OR2_X1 U8778 ( .A1(n14523), .A2(n13037), .ZN(n6486) );
  OR2_X1 U8779 ( .A1(n13345), .A2(n13029), .ZN(n6487) );
  AND2_X1 U8780 ( .A1(n9001), .A2(n9000), .ZN(n6488) );
  NOR2_X1 U8781 ( .A1(n11446), .A2(n7434), .ZN(n6489) );
  OR2_X1 U8782 ( .A1(n13640), .A2(n11351), .ZN(n11102) );
  AND2_X1 U8783 ( .A1(n8216), .A2(n8215), .ZN(n10010) );
  NAND2_X1 U8784 ( .A1(n11308), .A2(n7989), .ZN(n6490) );
  INV_X1 U8785 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7511) );
  INV_X1 U8786 ( .A(n12227), .ZN(n7359) );
  NAND2_X1 U8787 ( .A1(n9057), .A2(n9056), .ZN(n6491) );
  AND2_X1 U8788 ( .A1(n7497), .A2(n7445), .ZN(n7524) );
  AND2_X1 U8789 ( .A1(n10970), .A2(n7586), .ZN(n6492) );
  AND2_X1 U8790 ( .A1(n15035), .A2(n6738), .ZN(n6493) );
  AND2_X1 U8791 ( .A1(n12016), .A2(n14034), .ZN(n6494) );
  AND2_X1 U8792 ( .A1(n12046), .A2(n13574), .ZN(n6495) );
  OR2_X1 U8793 ( .A1(n12778), .A2(n12818), .ZN(n6496) );
  NAND2_X1 U8794 ( .A1(n6780), .A2(n7364), .ZN(n13516) );
  OR2_X1 U8795 ( .A1(n12701), .A2(n7018), .ZN(n6497) );
  NAND2_X1 U8796 ( .A1(n13998), .A2(n12228), .ZN(n6498) );
  OR2_X1 U8797 ( .A1(n14225), .A2(n12012), .ZN(n6499) );
  INV_X1 U8798 ( .A(n6710), .ZN(n6709) );
  NAND2_X1 U8799 ( .A1(n7816), .A2(n6505), .ZN(n6710) );
  XNOR2_X1 U8800 ( .A(n13320), .B(n8022), .ZN(n13158) );
  INV_X1 U8801 ( .A(n13158), .ZN(n6908) );
  NAND2_X1 U8802 ( .A1(n13760), .A2(n13759), .ZN(n13970) );
  INV_X1 U8803 ( .A(n13970), .ZN(n6856) );
  AND2_X1 U8804 ( .A1(n8585), .A2(n8584), .ZN(n12564) );
  MUX2_X1 U8805 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13469), .S(n9803), .Z(n10165)
         );
  NAND2_X1 U8806 ( .A1(n11101), .A2(n11100), .ZN(n13649) );
  AND4_X1 U8807 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n7030), .ZN(n6500)
         );
  OR2_X1 U8808 ( .A1(n10623), .A2(n13608), .ZN(n6501) );
  AND2_X1 U8809 ( .A1(n11511), .A2(n12372), .ZN(n6502) );
  OR2_X1 U8810 ( .A1(n11308), .A2(n7989), .ZN(n6503) );
  OR2_X1 U8811 ( .A1(n9307), .A2(n12329), .ZN(n6504) );
  OR2_X1 U8812 ( .A1(n13367), .A2(n13032), .ZN(n6505) );
  INV_X1 U8813 ( .A(n13743), .ZN(n7136) );
  AND2_X1 U8814 ( .A1(n13367), .A2(n13032), .ZN(n6506) );
  AND2_X1 U8815 ( .A1(n13367), .A2(n9219), .ZN(n6507) );
  INV_X1 U8816 ( .A(n13796), .ZN(n11702) );
  NOR2_X1 U8817 ( .A1(n8092), .A2(n13313), .ZN(n6873) );
  AND2_X1 U8818 ( .A1(n11316), .A2(n13041), .ZN(n6508) );
  NAND2_X1 U8819 ( .A1(n12852), .A2(n12851), .ZN(n6509) );
  AND2_X1 U8820 ( .A1(n14640), .A2(n7337), .ZN(n6510) );
  XNOR2_X1 U8821 ( .A(n13044), .B(n10855), .ZN(n10648) );
  AND2_X1 U8822 ( .A1(n6989), .A2(n6987), .ZN(n6511) );
  AND3_X1 U8823 ( .A1(n7522), .A2(n7521), .A3(n7520), .ZN(n6513) );
  AND2_X1 U8824 ( .A1(n8767), .A2(n8743), .ZN(n6514) );
  AOI21_X1 U8825 ( .B1(n7093), .B2(n7095), .A(n13255), .ZN(n7091) );
  AND2_X1 U8826 ( .A1(n14527), .A2(n14483), .ZN(n6515) );
  NAND2_X1 U8827 ( .A1(n9384), .A2(n9383), .ZN(n9417) );
  AND2_X1 U8828 ( .A1(n12592), .A2(n7056), .ZN(n6516) );
  AND2_X1 U8829 ( .A1(n8767), .A2(n8727), .ZN(n6517) );
  OR2_X1 U8830 ( .A1(n10019), .A2(n10018), .ZN(n6518) );
  AND2_X1 U8831 ( .A1(n11042), .A2(n8638), .ZN(n6519) );
  NOR2_X1 U8832 ( .A1(n9343), .A2(n9342), .ZN(n6520) );
  AND2_X1 U8833 ( .A1(n11856), .A2(n7360), .ZN(n6521) );
  AND2_X1 U8834 ( .A1(n14970), .A2(n13042), .ZN(n6522) );
  CLKBUF_X1 U8835 ( .A(n10220), .Z(n13846) );
  INV_X1 U8836 ( .A(n10220), .ZN(n6665) );
  INV_X1 U8837 ( .A(n7308), .ZN(n7307) );
  NOR2_X1 U8838 ( .A1(n9298), .A2(n7309), .ZN(n7308) );
  AND2_X1 U8839 ( .A1(n13610), .A2(n13609), .ZN(n6523) );
  INV_X1 U8840 ( .A(n6752), .ZN(n6751) );
  OAI21_X1 U8841 ( .B1(n12340), .B2(n9342), .A(n9343), .ZN(n6752) );
  NOR2_X1 U8842 ( .A1(n11455), .A2(n11300), .ZN(n6991) );
  NOR2_X1 U8843 ( .A1(n6898), .A2(n6897), .ZN(n6896) );
  AND2_X1 U8844 ( .A1(n12637), .A2(n7189), .ZN(n6524) );
  AND2_X1 U8845 ( .A1(n14174), .A2(n13821), .ZN(n6525) );
  NAND2_X1 U8846 ( .A1(n9280), .A2(n10776), .ZN(n6526) );
  AND2_X1 U8847 ( .A1(n13421), .A2(n12901), .ZN(n6527) );
  INV_X1 U8848 ( .A(n6942), .ZN(n6941) );
  NAND2_X1 U8849 ( .A1(n7424), .A2(n6498), .ZN(n6942) );
  AND2_X1 U8850 ( .A1(n11889), .A2(n11879), .ZN(n6528) );
  OR2_X1 U8851 ( .A1(n8987), .A2(n8986), .ZN(n6529) );
  INV_X1 U8852 ( .A(n6739), .ZN(n6738) );
  NOR2_X1 U8853 ( .A1(n10019), .A2(n10009), .ZN(n6739) );
  INV_X1 U8854 ( .A(n8933), .ZN(n8661) );
  AND2_X1 U8855 ( .A1(n8867), .A2(n8872), .ZN(n8933) );
  AND2_X1 U8856 ( .A1(n11767), .A2(n7997), .ZN(n6530) );
  AND2_X1 U8857 ( .A1(n11925), .A2(n11924), .ZN(n6531) );
  AND2_X1 U8858 ( .A1(n11940), .A2(n11939), .ZN(n6532) );
  AND2_X1 U8859 ( .A1(n11840), .A2(n11839), .ZN(n6533) );
  NAND2_X1 U8860 ( .A1(n14243), .A2(n13832), .ZN(n6534) );
  OR2_X1 U8861 ( .A1(n8026), .A2(n8025), .ZN(n6535) );
  NAND2_X1 U8862 ( .A1(n7378), .A2(n7377), .ZN(n6536) );
  INV_X1 U8863 ( .A(n7074), .ZN(n7073) );
  AND2_X1 U8864 ( .A1(n11241), .A2(n6503), .ZN(n7074) );
  INV_X1 U8865 ( .A(n6737), .ZN(n6736) );
  NOR2_X1 U8866 ( .A1(n6738), .A2(n10010), .ZN(n6737) );
  AND2_X1 U8867 ( .A1(n11349), .A2(n11292), .ZN(n6537) );
  AND2_X1 U8868 ( .A1(n12220), .A2(n12219), .ZN(n6538) );
  NOR2_X1 U8869 ( .A1(n12747), .A2(n12369), .ZN(n6539) );
  INV_X1 U8870 ( .A(n12299), .ZN(n6760) );
  AND2_X1 U8871 ( .A1(n12277), .A2(n9334), .ZN(n12299) );
  NOR2_X1 U8872 ( .A1(n10519), .A2(n10518), .ZN(n6540) );
  NOR2_X1 U8873 ( .A1(n12631), .A2(n12366), .ZN(n6541) );
  INV_X1 U8874 ( .A(n11728), .ZN(n6796) );
  AND2_X1 U8875 ( .A1(n12269), .A2(n9318), .ZN(n6542) );
  AND2_X1 U8876 ( .A1(n14175), .A2(n14176), .ZN(n6543) );
  NAND2_X1 U8877 ( .A1(n10320), .A2(n10319), .ZN(n6544) );
  AND3_X1 U8878 ( .A1(n7476), .A2(n7473), .A3(n7474), .ZN(n6545) );
  INV_X1 U8879 ( .A(n8806), .ZN(n7034) );
  AND2_X1 U8880 ( .A1(n7161), .A2(n7157), .ZN(n6546) );
  AND4_X1 U8881 ( .A1(n7446), .A2(n6902), .A3(n7448), .A4(n7497), .ZN(n6547)
         );
  AND2_X1 U8882 ( .A1(n9439), .A2(n14272), .ZN(n6548) );
  NOR2_X1 U8883 ( .A1(n13661), .A2(n11732), .ZN(n6549) );
  NOR2_X1 U8884 ( .A1(n12864), .A2(n12990), .ZN(n6550) );
  INV_X1 U8885 ( .A(n6876), .ZN(n6875) );
  NAND2_X1 U8886 ( .A1(n6878), .A2(n6877), .ZN(n6876) );
  AND2_X1 U8887 ( .A1(n13580), .A2(n14753), .ZN(n6551) );
  AND2_X1 U8888 ( .A1(n6496), .A2(n6625), .ZN(n6552) );
  INV_X1 U8889 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8111) );
  XNOR2_X1 U8890 ( .A(n14090), .B(n13693), .ZN(n14085) );
  AND2_X1 U8891 ( .A1(n10588), .A2(n10623), .ZN(n6553) );
  OR2_X1 U8892 ( .A1(n14294), .A2(n14293), .ZN(n6554) );
  INV_X1 U8893 ( .A(n7216), .ZN(n7215) );
  NAND2_X1 U8894 ( .A1(n7217), .A2(n11528), .ZN(n7216) );
  INV_X1 U8895 ( .A(n6985), .ZN(n6984) );
  AND2_X1 U8896 ( .A1(n7550), .A2(SI_4_), .ZN(n6555) );
  AND2_X1 U8897 ( .A1(n7582), .A2(SI_6_), .ZN(n6556) );
  INV_X1 U8898 ( .A(n7382), .ZN(n7381) );
  NOR2_X1 U8899 ( .A1(n9098), .A2(n9099), .ZN(n7382) );
  NAND2_X1 U8900 ( .A1(n11170), .A2(n11169), .ZN(n6557) );
  AND2_X1 U8901 ( .A1(n6710), .A2(n13255), .ZN(n6558) );
  NAND2_X1 U8902 ( .A1(n12248), .A2(n6753), .ZN(n6559) );
  AND2_X1 U8903 ( .A1(n10945), .A2(n6986), .ZN(n6560) );
  AND2_X1 U8904 ( .A1(n11453), .A2(n6992), .ZN(n6561) );
  INV_X1 U8905 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U8906 ( .A1(n8891), .A2(n7058), .ZN(n6562) );
  INV_X1 U8907 ( .A(n9032), .ZN(n7401) );
  INV_X1 U8908 ( .A(n13662), .ZN(n7145) );
  AND2_X1 U8909 ( .A1(n11071), .A2(n8639), .ZN(n6563) );
  AND2_X1 U8910 ( .A1(n12241), .A2(n12341), .ZN(n6564) );
  AND3_X1 U8911 ( .A1(n7334), .A2(n7331), .A3(n6819), .ZN(n6565) );
  AND2_X1 U8912 ( .A1(n7291), .A2(n10635), .ZN(n6566) );
  OR2_X1 U8913 ( .A1(n12555), .A2(n7067), .ZN(n6567) );
  AND2_X1 U8914 ( .A1(n13401), .A2(n7763), .ZN(n6568) );
  AND2_X1 U8915 ( .A1(n9060), .A2(n9059), .ZN(n6569) );
  AND2_X1 U8916 ( .A1(n13230), .A2(n7863), .ZN(n6570) );
  AND2_X1 U8917 ( .A1(n9438), .A2(n9437), .ZN(n6571) );
  AND2_X1 U8918 ( .A1(n14179), .A2(n14043), .ZN(n6572) );
  OR2_X1 U8919 ( .A1(n14299), .A2(n6812), .ZN(n6573) );
  OR2_X1 U8920 ( .A1(n7494), .A2(n9469), .ZN(n6574) );
  AND2_X1 U8921 ( .A1(n8877), .A2(n8867), .ZN(n6575) );
  OR2_X1 U8922 ( .A1(n7404), .A2(n7408), .ZN(n6576) );
  AND2_X1 U8923 ( .A1(n9179), .A2(n9134), .ZN(n6577) );
  NAND2_X1 U8924 ( .A1(n6868), .A2(n13248), .ZN(n6871) );
  NAND2_X1 U8925 ( .A1(n12025), .A2(n12043), .ZN(n13983) );
  NAND2_X1 U8926 ( .A1(n10519), .A2(n10518), .ZN(n6578) );
  AND2_X1 U8927 ( .A1(n7356), .A2(n7359), .ZN(n6579) );
  AND2_X1 U8928 ( .A1(n9383), .A2(n9418), .ZN(n6580) );
  AND2_X1 U8929 ( .A1(n13700), .A2(n13699), .ZN(n14073) );
  OR2_X1 U8930 ( .A1(n9046), .A2(n9042), .ZN(n6581) );
  OR2_X1 U8931 ( .A1(n7400), .A2(n9043), .ZN(n6582) );
  NOR2_X1 U8932 ( .A1(n14193), .A2(n13824), .ZN(n6583) );
  AND2_X1 U8933 ( .A1(n7011), .A2(n7010), .ZN(n6584) );
  AND2_X1 U8934 ( .A1(n12907), .A2(n6509), .ZN(n6995) );
  NOR2_X1 U8935 ( .A1(n7384), .A2(n7383), .ZN(n6585) );
  INV_X1 U8936 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9538) );
  OR2_X1 U8937 ( .A1(n7401), .A2(n6478), .ZN(n6586) );
  INV_X1 U8938 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7525) );
  INV_X1 U8939 ( .A(n8110), .ZN(n7194) );
  INV_X1 U8940 ( .A(n9234), .ZN(n11426) );
  INV_X1 U8941 ( .A(n12298), .ZN(n6761) );
  INV_X1 U8942 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8266) );
  AND2_X1 U8943 ( .A1(n8843), .A2(n8842), .ZN(n11330) );
  INV_X1 U8944 ( .A(n11330), .ZN(n7043) );
  INV_X1 U8945 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7030) );
  NAND2_X1 U8946 ( .A1(n11844), .A2(n11843), .ZN(n14233) );
  INV_X1 U8947 ( .A(n14233), .ZN(n6863) );
  AND2_X1 U8948 ( .A1(n8518), .A2(n8517), .ZN(n12618) );
  NAND2_X1 U8949 ( .A1(n6893), .A2(n6892), .ZN(n14504) );
  INV_X1 U8950 ( .A(n12277), .ZN(n6756) );
  NAND2_X1 U8951 ( .A1(n6713), .A2(n7740), .ZN(n11690) );
  OR3_X1 U8952 ( .A1(n11743), .A2(n13277), .A3(n6889), .ZN(n6587) );
  AND4_X1 U8953 ( .A1(n8242), .A2(n8241), .A3(n8240), .A4(n8239), .ZN(n10960)
         );
  INV_X1 U8954 ( .A(n10960), .ZN(n12378) );
  AND4_X1 U8955 ( .A1(n8295), .A2(n8294), .A3(n8293), .A4(n8292), .ZN(n11405)
         );
  INV_X1 U8956 ( .A(n11405), .ZN(n12375) );
  INV_X1 U8957 ( .A(n6864), .ZN(n14134) );
  NOR2_X1 U8958 ( .A1(n14151), .A2(n14238), .ZN(n6864) );
  AND2_X1 U8959 ( .A1(n11529), .A2(n11528), .ZN(n6588) );
  INV_X1 U8960 ( .A(n7182), .ZN(n7181) );
  NOR2_X1 U8961 ( .A1(n8659), .A2(n7183), .ZN(n7182) );
  INV_X1 U8962 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6812) );
  NAND2_X1 U8963 ( .A1(n8087), .A2(n8086), .ZN(n6589) );
  INV_X1 U8964 ( .A(n14622), .ZN(n7326) );
  INV_X1 U8965 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n12094) );
  INV_X1 U8966 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9909) );
  NAND2_X2 U8967 ( .A1(n13571), .A2(n13584), .ZN(n10393) );
  INV_X1 U8968 ( .A(n11109), .ZN(n11930) );
  INV_X1 U8969 ( .A(n13793), .ZN(n7214) );
  NAND2_X1 U8970 ( .A1(n11378), .A2(n11377), .ZN(n13661) );
  INV_X1 U8971 ( .A(n13661), .ZN(n6857) );
  AND2_X1 U8972 ( .A1(n8725), .A2(n8724), .ZN(n15127) );
  NAND2_X1 U8973 ( .A1(n7965), .A2(n7416), .ZN(n8040) );
  INV_X1 U8974 ( .A(SI_14_), .ZN(n7261) );
  NOR2_X1 U8975 ( .A1(n13787), .A2(n6957), .ZN(n6956) );
  AND2_X1 U8976 ( .A1(n11265), .A2(n6875), .ZN(n6590) );
  INV_X1 U8977 ( .A(n10667), .ZN(n6882) );
  AND2_X1 U8978 ( .A1(n14406), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U8979 ( .A1(n6922), .A2(n10242), .ZN(n10622) );
  NAND2_X1 U8980 ( .A1(n7686), .A2(n7685), .ZN(n14527) );
  INV_X1 U8981 ( .A(n14527), .ZN(n6877) );
  OR2_X1 U8982 ( .A1(n10529), .A2(n10528), .ZN(n6592) );
  NAND2_X1 U8983 ( .A1(n11818), .A2(n11817), .ZN(n14243) );
  INV_X1 U8984 ( .A(n14243), .ZN(n6865) );
  OR2_X1 U8985 ( .A1(n15002), .A2(n6618), .ZN(n6593) );
  NAND2_X1 U8986 ( .A1(n7749), .A2(n7011), .ZN(n7805) );
  OR2_X1 U8987 ( .A1(n12393), .A2(n14476), .ZN(n6594) );
  INV_X1 U8988 ( .A(n6849), .ZN(n10720) );
  NOR2_X1 U8989 ( .A1(n10482), .A2(n13608), .ZN(n6849) );
  INV_X1 U8990 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6682) );
  AND2_X1 U8991 ( .A1(n12129), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8992 ( .A1(n12440), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n6596) );
  OAI21_X1 U8993 ( .B1(n14650), .B2(n10340), .A(n7348), .ZN(n7346) );
  NAND2_X1 U8994 ( .A1(n7965), .A2(n7417), .ZN(n6597) );
  AND2_X1 U8995 ( .A1(n10986), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U8996 ( .A1(n8686), .A2(n8685), .ZN(n6599) );
  NOR2_X1 U8997 ( .A1(n10936), .A2(n10935), .ZN(n6600) );
  NAND2_X1 U8998 ( .A1(n6975), .A2(n6544), .ZN(n6976) );
  XNOR2_X1 U8999 ( .A(n9539), .B(n9538), .ZN(n13738) );
  INV_X1 U9000 ( .A(n13738), .ZN(n6806) );
  INV_X1 U9001 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6808) );
  OR2_X1 U9002 ( .A1(n12494), .A2(n12493), .ZN(n6601) );
  NAND2_X1 U9003 ( .A1(n6925), .A2(n10230), .ZN(n10479) );
  NAND2_X1 U9004 ( .A1(n10598), .A2(n10597), .ZN(n14787) );
  INV_X1 U9005 ( .A(n14787), .ZN(n6847) );
  AND2_X1 U9006 ( .A1(n13728), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U9007 ( .A1(n7968), .A2(n11369), .ZN(n11311) );
  INV_X1 U9008 ( .A(n13093), .ZN(n6659) );
  INV_X1 U9009 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U9010 ( .A1(n6829), .A2(n7516), .ZN(n7528) );
  NAND2_X1 U9011 ( .A1(n6831), .A2(n6574), .ZN(n7097) );
  OAI21_X2 U9012 ( .B1(n6835), .B2(n6833), .A(n6834), .ZN(n13214) );
  NAND2_X1 U9013 ( .A1(n6660), .A2(n7245), .ZN(n7589) );
  NAND2_X1 U9014 ( .A1(n6619), .A2(n6593), .ZN(P2_U3528) );
  NAND4_X1 U9015 ( .A1(n9247), .A2(n9246), .A3(n9245), .A4(n9244), .ZN(n6684)
         );
  NAND2_X1 U9016 ( .A1(n14022), .A2(n12017), .ZN(n14009) );
  NAND3_X1 U9017 ( .A1(n7202), .A2(n7201), .A3(n7203), .ZN(n14022) );
  NAND2_X1 U9018 ( .A1(n7219), .A2(n7218), .ZN(n12035) );
  OAI21_X1 U9019 ( .B1(n7743), .B2(n7742), .A(n7741), .ZN(n7765) );
  NAND2_X1 U9020 ( .A1(n6918), .A2(n6917), .ZN(n11527) );
  OAI21_X1 U9021 ( .B1(n7663), .B2(n7662), .A(n7661), .ZN(n7677) );
  NAND2_X1 U9022 ( .A1(n7235), .A2(n7233), .ZN(n7842) );
  NAND2_X1 U9023 ( .A1(n6683), .A2(n7591), .ZN(n7609) );
  NAND2_X1 U9024 ( .A1(n13749), .A2(n13750), .ZN(n6633) );
  NAND2_X1 U9025 ( .A1(n6610), .A2(n6609), .ZN(P1_U3525) );
  OR2_X1 U9026 ( .A1(n14807), .A2(n12029), .ZN(n6609) );
  NAND2_X1 U9027 ( .A1(n14257), .A2(n14807), .ZN(n6610) );
  NAND2_X1 U9028 ( .A1(n7609), .A2(n7608), .ZN(n6828) );
  AOI21_X1 U9029 ( .B1(n7130), .B2(n7133), .A(n7129), .ZN(n7128) );
  OAI21_X1 U9030 ( .B1(n7002), .B2(n7001), .A(n6623), .ZN(n12954) );
  NAND2_X1 U9031 ( .A1(n13002), .A2(n6995), .ZN(n6993) );
  OAI21_X2 U9032 ( .B1(n12980), .B2(n12976), .A(n12977), .ZN(n12928) );
  INV_X1 U9033 ( .A(n11910), .ZN(n7367) );
  NAND2_X1 U9034 ( .A1(n6779), .A2(n6778), .ZN(n13499) );
  OAI21_X2 U9035 ( .B1(n6691), .B2(n6690), .A(n13984), .ZN(n6611) );
  INV_X1 U9036 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7101) );
  INV_X1 U9037 ( .A(n6939), .ZN(n6938) );
  INV_X1 U9038 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7103) );
  NAND2_X1 U9039 ( .A1(n11775), .A2(n13756), .ZN(n11777) );
  INV_X1 U9040 ( .A(n6612), .ZN(n6697) );
  OAI21_X1 U9041 ( .B1(n14166), .B2(n14795), .A(n14172), .ZN(n6612) );
  NAND3_X1 U9042 ( .A1(n7437), .A2(n6613), .A3(n9247), .ZN(n9200) );
  NAND2_X1 U9043 ( .A1(n9115), .A2(n6577), .ZN(n6613) );
  NOR2_X1 U9044 ( .A1(n9094), .A2(n6585), .ZN(n7380) );
  NAND3_X1 U9045 ( .A1(n9012), .A2(n7413), .A3(n9013), .ZN(n6627) );
  NAND2_X2 U9046 ( .A1(n6545), .A2(n7475), .ZN(n13048) );
  NAND2_X1 U9047 ( .A1(n8901), .A2(n12565), .ZN(n8905) );
  NAND2_X1 U9048 ( .A1(n8157), .A2(n8156), .ZN(n8171) );
  NAND2_X1 U9049 ( .A1(n8192), .A2(n8191), .ZN(n8209) );
  NAND2_X1 U9050 ( .A1(n8906), .A2(n12555), .ZN(n8912) );
  OAI21_X2 U9051 ( .B1(n8340), .B2(n8339), .A(n8341), .ZN(n8342) );
  OAI21_X2 U9052 ( .B1(n8245), .B2(n8244), .A(n8246), .ZN(n8262) );
  NAND2_X1 U9053 ( .A1(n8907), .A2(n8914), .ZN(n6615) );
  NAND2_X1 U9054 ( .A1(n6615), .A2(n6614), .ZN(n8917) );
  AOI21_X1 U9055 ( .B1(n13159), .B2(n6908), .A(n8023), .ZN(n8026) );
  OAI21_X1 U9056 ( .B1(n13411), .B2(n14991), .A(n7421), .ZN(n13412) );
  NAND3_X1 U9057 ( .A1(n7130), .A2(n13725), .A3(n13724), .ZN(n7127) );
  INV_X1 U9058 ( .A(n11973), .ZN(n7358) );
  NAND2_X1 U9059 ( .A1(n7249), .A2(n7250), .ZN(n7743) );
  OAI21_X1 U9060 ( .B1(n7355), .B2(n7359), .A(n7350), .ZN(n7349) );
  NAND2_X1 U9061 ( .A1(n6828), .A2(n7611), .ZN(n7625) );
  NAND3_X1 U9062 ( .A1(n9200), .A2(n6621), .A3(n6620), .ZN(n9210) );
  NAND2_X1 U9063 ( .A1(n6873), .A2(n6872), .ZN(n13144) );
  NAND2_X1 U9064 ( .A1(n12521), .A2(n15055), .ZN(n6724) );
  NAND2_X1 U9065 ( .A1(n6724), .A2(n12520), .ZN(n6723) );
  NAND2_X1 U9066 ( .A1(n11612), .A2(n11611), .ZN(n11758) );
  NAND2_X4 U9067 ( .A1(n11255), .A2(n10120), .ZN(n12915) );
  OR2_X2 U9068 ( .A1(n7971), .A2(n6463), .ZN(n11255) );
  NAND2_X2 U9069 ( .A1(n12582), .A2(n8897), .ZN(n12566) );
  NAND2_X1 U9070 ( .A1(n10813), .A2(n10812), .ZN(n10811) );
  BUF_X2 U9071 ( .A(n8121), .Z(n12239) );
  BUF_X4 U9072 ( .A(n8198), .Z(n8604) );
  AND2_X2 U9073 ( .A1(n6689), .A2(n10424), .ZN(n7033) );
  NAND2_X2 U9074 ( .A1(n8491), .A2(n8785), .ZN(n12620) );
  OR2_X1 U9075 ( .A1(n9038), .A2(n9037), .ZN(n7438) );
  NAND2_X1 U9076 ( .A1(n7395), .A2(n7393), .ZN(n9009) );
  NAND2_X1 U9077 ( .A1(n6661), .A2(n6529), .ZN(n8994) );
  NAND2_X1 U9078 ( .A1(n6627), .A2(n7411), .ZN(n9024) );
  NAND2_X1 U9079 ( .A1(n6626), .A2(n6536), .ZN(n9109) );
  OR2_X1 U9080 ( .A1(n9104), .A2(n9103), .ZN(n6626) );
  INV_X1 U9081 ( .A(n8985), .ZN(n6661) );
  AOI21_X1 U9082 ( .B1(n9109), .B2(n9108), .A(n9107), .ZN(n9114) );
  NAND2_X1 U9083 ( .A1(n8994), .A2(n8995), .ZN(n8993) );
  NAND2_X1 U9084 ( .A1(n7376), .A2(n7381), .ZN(n9104) );
  AOI21_X1 U9085 ( .B1(n6628), .B2(n13980), .A(n14795), .ZN(n13982) );
  NAND2_X1 U9086 ( .A1(n13979), .A2(n13983), .ZN(n6628) );
  NAND2_X1 U9087 ( .A1(n9124), .A2(n9123), .ZN(n9164) );
  AOI21_X1 U9088 ( .B1(n6949), .B2(n6948), .A(n6583), .ZN(n6947) );
  NAND2_X1 U9089 ( .A1(n6634), .A2(n7146), .ZN(n13670) );
  NAND3_X1 U9090 ( .A1(n13660), .A2(n7144), .A3(n13659), .ZN(n6634) );
  NAND2_X1 U9091 ( .A1(n6635), .A2(n13818), .ZN(P1_U3242) );
  NAND3_X1 U9092 ( .A1(n13813), .A2(n6688), .A3(n13812), .ZN(n6635) );
  NAND3_X1 U9093 ( .A1(n13594), .A2(n14706), .A3(n13595), .ZN(n13599) );
  OR2_X1 U9094 ( .A1(n13722), .A2(n13723), .ZN(n13724) );
  NAND2_X1 U9095 ( .A1(n13585), .A2(n13586), .ZN(n13591) );
  OAI21_X1 U9096 ( .B1(n7124), .B2(n13691), .A(n13692), .ZN(n6686) );
  AOI21_X1 U9097 ( .B1(n13680), .B2(n13679), .A(n6680), .ZN(n6679) );
  INV_X1 U9098 ( .A(n13773), .ZN(n13767) );
  NAND2_X1 U9099 ( .A1(n7127), .A2(n7128), .ZN(n13773) );
  NAND2_X1 U9100 ( .A1(n6636), .A2(n7143), .ZN(n13655) );
  NAND3_X1 U9101 ( .A1(n13648), .A2(n13647), .A3(n7141), .ZN(n6636) );
  NAND2_X1 U9102 ( .A1(n9136), .A2(n9135), .ZN(n7277) );
  NOR2_X1 U9103 ( .A1(n13591), .A2(n13590), .ZN(n13592) );
  NAND2_X1 U9104 ( .A1(n13716), .A2(n7155), .ZN(n7148) );
  NAND2_X1 U9105 ( .A1(n13712), .A2(n6637), .ZN(n13716) );
  NAND2_X1 U9106 ( .A1(n9433), .A2(n9389), .ZN(n9430) );
  NAND2_X1 U9107 ( .A1(n7126), .A2(n7125), .ZN(n7124) );
  NAND2_X1 U9108 ( .A1(n13570), .A2(n13571), .ZN(n13573) );
  AOI22_X1 U9109 ( .A1(n13708), .A2(n13707), .B1(n13706), .B2(n13705), .ZN(
        n13711) );
  NOR2_X1 U9110 ( .A1(n13676), .A2(n13675), .ZN(n13680) );
  NAND2_X1 U9111 ( .A1(n13681), .A2(n6679), .ZN(n13687) );
  NAND2_X2 U9112 ( .A1(n12566), .A2(n8902), .ZN(n8568) );
  NAND2_X1 U9113 ( .A1(n6638), .A2(n12338), .ZN(n12342) );
  NAND2_X1 U9114 ( .A1(n12339), .A2(n12340), .ZN(n12338) );
  OR2_X1 U9115 ( .A1(n12339), .A2(n12340), .ZN(n6638) );
  AOI21_X1 U9116 ( .B1(n6566), .B2(n7293), .A(n7288), .ZN(n10775) );
  OAI21_X1 U9117 ( .B1(n7195), .B2(n8110), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8131) );
  INV_X1 U9118 ( .A(n12349), .ZN(n6765) );
  NAND2_X1 U9119 ( .A1(n6642), .A2(n9256), .ZN(P2_U3328) );
  OAI21_X1 U9120 ( .B1(n9252), .B2(n9251), .A(n6643), .ZN(n6642) );
  NAND2_X1 U9121 ( .A1(n6647), .A2(n8155), .ZN(n8157) );
  INV_X1 U9122 ( .A(n8154), .ZN(n6647) );
  NAND2_X1 U9123 ( .A1(n6650), .A2(n6648), .ZN(P3_U3488) );
  OR2_X1 U9124 ( .A1(n8741), .A2(n15131), .ZN(n6650) );
  NAND2_X1 U9125 ( .A1(n6653), .A2(n6651), .ZN(P3_U3456) );
  OR2_X1 U9126 ( .A1(n8741), .A2(n15127), .ZN(n6653) );
  NOR2_X1 U9127 ( .A1(n8073), .A2(n6669), .ZN(n8079) );
  NAND2_X2 U9128 ( .A1(n6655), .A2(n6654), .ZN(n11772) );
  AOI21_X2 U9129 ( .B1(n10577), .B2(n10578), .A(n6551), .ZN(n14704) );
  AOI21_X2 U9130 ( .B1(n10713), .B2(n10590), .A(n6657), .ZN(n10756) );
  OAI22_X1 U9131 ( .A1(n9202), .A2(n9201), .B1(n9199), .B2(n9198), .ZN(n7229)
         );
  NAND2_X1 U9132 ( .A1(n6468), .A2(n13984), .ZN(n6939) );
  NAND2_X1 U9133 ( .A1(n9198), .A2(n9199), .ZN(n9184) );
  NOR2_X1 U9134 ( .A1(n15063), .A2(n10888), .ZN(n15090) );
  MUX2_X1 U9135 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14255), .S(n14819), .Z(
        P1_U3559) );
  INV_X1 U9136 ( .A(n6862), .ZN(n6861) );
  NAND3_X1 U9137 ( .A1(n6840), .A2(n6841), .A3(n7243), .ZN(n6660) );
  NOR2_X1 U9138 ( .A1(n7226), .A2(n7225), .ZN(n7224) );
  NAND2_X2 U9139 ( .A1(n8037), .A2(n7451), .ZN(n7452) );
  OR2_X2 U9140 ( .A1(n8979), .A2(n8978), .ZN(n7430) );
  OR2_X1 U9141 ( .A1(n9052), .A2(n9051), .ZN(n7419) );
  NOR2_X2 U9142 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7442) );
  NAND2_X1 U9143 ( .A1(n6694), .A2(n6547), .ZN(n6899) );
  NAND2_X1 U9144 ( .A1(n6663), .A2(n6662), .ZN(n9038) );
  NAND3_X1 U9145 ( .A1(n9039), .A2(n7438), .A3(n6581), .ZN(n7399) );
  NAND3_X1 U9146 ( .A1(n9029), .A2(n9028), .A3(n6586), .ZN(n6663) );
  INV_X1 U9147 ( .A(n6901), .ZN(n6694) );
  NAND2_X1 U9148 ( .A1(n7403), .A2(n7402), .ZN(n9069) );
  NAND2_X1 U9149 ( .A1(n7380), .A2(n7379), .ZN(n7376) );
  NAND2_X2 U9150 ( .A1(n13590), .A2(n10258), .ZN(n10256) );
  NAND2_X1 U9151 ( .A1(n11070), .A2(n8640), .ZN(n11191) );
  NAND2_X1 U9152 ( .A1(n8127), .A2(n12101), .ZN(n8129) );
  NAND2_X1 U9153 ( .A1(n7028), .A2(n8229), .ZN(n8245) );
  NAND2_X1 U9154 ( .A1(n8645), .A2(n8644), .ZN(n11326) );
  OAI21_X1 U9155 ( .B1(n11441), .B2(n7177), .A(n7174), .ZN(n8660) );
  OAI21_X1 U9156 ( .B1(n12777), .B2(n15131), .A(n6666), .ZN(P3_U3487) );
  OAI22_X1 U9157 ( .A1(n12616), .A2(n8665), .B1(n12796), .B2(n12628), .ZN(
        n12605) );
  NAND2_X1 U9158 ( .A1(n6940), .A2(n6938), .ZN(n13980) );
  INV_X1 U9159 ( .A(n6947), .ZN(n6945) );
  NAND2_X1 U9160 ( .A1(n9188), .A2(n9187), .ZN(n6670) );
  NAND2_X1 U9161 ( .A1(n7134), .A2(n7132), .ZN(n7131) );
  NAND2_X1 U9162 ( .A1(n6891), .A2(n6890), .ZN(P2_U3496) );
  INV_X1 U9163 ( .A(n6719), .ZN(n6845) );
  INV_X1 U9164 ( .A(n6672), .ZN(n13312) );
  AOI21_X1 U9165 ( .B1(n8092), .B2(n13313), .A(n13217), .ZN(n6674) );
  NAND2_X1 U9166 ( .A1(n6677), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7029) );
  OAI21_X2 U9167 ( .B1(n8438), .B2(n7024), .A(n7022), .ZN(n8477) );
  NAND2_X2 U9168 ( .A1(n8911), .A2(n8909), .ZN(n12542) );
  NAND3_X1 U9169 ( .A1(n10501), .A2(n10645), .A3(n10648), .ZN(n6675) );
  INV_X1 U9170 ( .A(n7487), .ZN(n7469) );
  NAND2_X2 U9171 ( .A1(n7468), .A2(n12215), .ZN(n7487) );
  NAND2_X1 U9172 ( .A1(n11430), .A2(n7993), .ZN(n11474) );
  OAI21_X1 U9173 ( .B1(n11681), .B2(n7761), .A(n7999), .ZN(n11742) );
  NAND2_X1 U9174 ( .A1(n8006), .A2(n8005), .ZN(n13279) );
  INV_X1 U9175 ( .A(n10799), .ZN(n6676) );
  NAND2_X1 U9176 ( .A1(n6676), .A2(n7086), .ZN(n7084) );
  OR2_X1 U9177 ( .A1(n9225), .A2(n7977), .ZN(n7978) );
  XNOR2_X1 U9178 ( .A(n8588), .B(n8573), .ZN(n11450) );
  INV_X1 U9179 ( .A(n8342), .ZN(n6677) );
  NAND3_X1 U9180 ( .A1(n7029), .A2(P1_DATAO_REG_13__SCAN_IN), .A3(n8358), .ZN(
        n8359) );
  NAND2_X1 U9181 ( .A1(n8950), .A2(n9257), .ZN(n8951) );
  NAND2_X1 U9182 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  NAND2_X1 U9183 ( .A1(n8315), .A2(n8314), .ZN(n8322) );
  XNOR2_X1 U9184 ( .A(n7171), .B(n8944), .ZN(n8684) );
  NAND2_X1 U9185 ( .A1(n8521), .A2(n8520), .ZN(n8523) );
  NAND2_X1 U9186 ( .A1(n8264), .A2(n8263), .ZN(n8281) );
  OR2_X1 U9187 ( .A1(n7981), .A2(n7980), .ZN(n7983) );
  OAI21_X1 U9188 ( .B1(n6523), .B2(n6678), .A(n7163), .ZN(n13623) );
  NAND2_X1 U9189 ( .A1(n13615), .A2(n7162), .ZN(n6678) );
  NAND3_X1 U9190 ( .A1(n7070), .A2(n7071), .A3(n9234), .ZN(n11430) );
  NAND2_X1 U9191 ( .A1(n11742), .A2(n8000), .ZN(n8003) );
  NAND2_X1 U9192 ( .A1(n13606), .A2(n13605), .ZN(n13611) );
  NAND2_X1 U9193 ( .A1(n14292), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6815) );
  NOR2_X1 U9194 ( .A1(n14426), .A2(n14361), .ZN(n14430) );
  NAND2_X1 U9195 ( .A1(n7068), .A2(n8014), .ZN(n13198) );
  NAND2_X1 U9196 ( .A1(n7589), .A2(n7588), .ZN(n6683) );
  NAND2_X1 U9197 ( .A1(n7767), .A2(n7237), .ZN(n7235) );
  NAND2_X1 U9198 ( .A1(n7277), .A2(n9138), .ZN(n9188) );
  NAND2_X1 U9199 ( .A1(n14430), .A2(n14431), .ZN(n14429) );
  NAND2_X1 U9200 ( .A1(n10607), .A2(n10630), .ZN(n10995) );
  XNOR2_X2 U9201 ( .A(n14647), .B(n6453), .ZN(n13777) );
  NAND2_X2 U9202 ( .A1(n9722), .A2(n6512), .ZN(n14647) );
  NAND2_X1 U9203 ( .A1(n7137), .A2(n7140), .ZN(n13643) );
  NAND2_X1 U9204 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  NAND2_X1 U9205 ( .A1(n13628), .A2(n13627), .ZN(n13631) );
  OAI21_X1 U9206 ( .B1(n13604), .B2(n13603), .A(n13602), .ZN(n13606) );
  NAND2_X1 U9207 ( .A1(n7148), .A2(n7153), .ZN(n13722) );
  OAI21_X2 U9208 ( .B1(n10256), .B2(n14721), .A(n10258), .ZN(n10577) );
  OR2_X2 U9209 ( .A1(n14144), .A2(n14145), .ZN(n7200) );
  NAND2_X1 U9210 ( .A1(n6696), .A2(n13696), .ZN(n14071) );
  NAND2_X1 U9211 ( .A1(n12007), .A2(n12006), .ZN(n14144) );
  OAI21_X2 U9212 ( .B1(n11382), .B2(n7216), .A(n7213), .ZN(n11701) );
  NAND2_X1 U9213 ( .A1(n11118), .A2(n11117), .ZN(n11120) );
  NAND2_X1 U9214 ( .A1(n10995), .A2(n10994), .ZN(n11051) );
  NAND2_X1 U9215 ( .A1(n10755), .A2(n10594), .ZN(n10607) );
  NAND2_X1 U9216 ( .A1(n10756), .A2(n10757), .ZN(n10755) );
  OR2_X1 U9217 ( .A1(n11866), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9928) );
  NAND2_X1 U9218 ( .A1(n13462), .A2(n7612), .ZN(n7904) );
  XNOR2_X2 U9219 ( .A(n13193), .B(n13027), .ZN(n13186) );
  INV_X1 U9220 ( .A(n8169), .ZN(n8170) );
  NAND2_X1 U9221 ( .A1(n8173), .A2(n8172), .ZN(n8190) );
  NAND2_X1 U9222 ( .A1(n8211), .A2(n8210), .ZN(n8228) );
  NAND2_X1 U9223 ( .A1(n8373), .A2(n8372), .ZN(n8375) );
  NAND2_X1 U9224 ( .A1(n8313), .A2(n8312), .ZN(n8315) );
  NAND2_X1 U9225 ( .A1(n8433), .A2(n8432), .ZN(n8435) );
  NAND2_X1 U9226 ( .A1(n8262), .A2(n8261), .ZN(n8264) );
  OAI21_X2 U9227 ( .B1(n8507), .B2(n8506), .A(n8508), .ZN(n8521) );
  NOR2_X2 U9228 ( .A1(n7195), .A2(n7192), .ZN(n8127) );
  NAND2_X1 U9229 ( .A1(n7060), .A2(n6567), .ZN(n12543) );
  NAND3_X2 U9230 ( .A1(n8159), .A2(n6500), .A3(n8105), .ZN(n8325) );
  NAND2_X1 U9231 ( .A1(n7049), .A2(n7047), .ZN(n11195) );
  NAND2_X1 U9232 ( .A1(n7040), .A2(n7038), .ZN(n11445) );
  INV_X1 U9233 ( .A(n7221), .ZN(n6691) );
  AND2_X1 U9234 ( .A1(n13848), .A2(n10257), .ZN(n14721) );
  NAND2_X1 U9235 ( .A1(n14113), .A2(n14112), .ZN(n14111) );
  INV_X1 U9236 ( .A(n6692), .ZN(n9783) );
  NAND2_X1 U9237 ( .A1(n6692), .A2(n9740), .ZN(n9741) );
  OR2_X1 U9238 ( .A1(n9784), .A2(n9744), .ZN(n6692) );
  XNOR2_X1 U9239 ( .A(n7113), .B(n15071), .ZN(n15064) );
  NOR2_X1 U9240 ( .A1(n10306), .A2(n10307), .ZN(n10309) );
  XNOR2_X2 U9241 ( .A(n8145), .B(P3_IR_REG_1__SCAN_IN), .ZN(n9762) );
  INV_X1 U9242 ( .A(n6837), .ZN(n6835) );
  NAND2_X1 U9243 ( .A1(n6467), .A2(n7985), .ZN(n10799) );
  XNOR2_X1 U9244 ( .A(n13046), .B(n10743), .ZN(n10502) );
  NAND2_X1 U9245 ( .A1(n11041), .A2(n6563), .ZN(n11070) );
  NAND2_X1 U9246 ( .A1(n10130), .A2(n7198), .ZN(n10427) );
  NAND2_X1 U9247 ( .A1(n7191), .A2(n7045), .ZN(n7195) );
  NAND2_X1 U9248 ( .A1(n8626), .A2(n8625), .ZN(n10185) );
  NOR2_X4 U9249 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8158) );
  INV_X1 U9250 ( .A(n6873), .ZN(n13142) );
  NAND2_X1 U9251 ( .A1(n6940), .A2(n6468), .ZN(n13979) );
  NAND2_X1 U9252 ( .A1(n7647), .A2(n7646), .ZN(n7663) );
  NAND2_X1 U9253 ( .A1(n6827), .A2(n7627), .ZN(n7644) );
  NOR2_X1 U9254 ( .A1(n6945), .A2(n6944), .ZN(n6943) );
  NAND2_X1 U9255 ( .A1(n8359), .A2(n8358), .ZN(n8373) );
  NAND2_X1 U9256 ( .A1(n7016), .A2(n8300), .ZN(n8313) );
  NAND2_X1 U9257 ( .A1(n8228), .A2(n8227), .ZN(n7028) );
  INV_X1 U9258 ( .A(n8524), .ZN(n7027) );
  NAND2_X1 U9259 ( .A1(n7015), .A2(n8393), .ZN(n8409) );
  NAND2_X1 U9260 ( .A1(n7017), .A2(n8282), .ZN(n8298) );
  AOI21_X2 U9261 ( .B1(n8921), .B2(n8945), .A(n8943), .ZN(n8922) );
  NAND2_X1 U9262 ( .A1(n7995), .A2(n7079), .ZN(n6832) );
  NOR2_X1 U9263 ( .A1(n7464), .A2(n13444), .ZN(n6867) );
  NAND2_X1 U9264 ( .A1(n14257), .A2(n14819), .ZN(n6928) );
  INV_X1 U9265 ( .A(n14074), .ZN(n6696) );
  XNOR2_X2 U9266 ( .A(n9573), .B(n9572), .ZN(n12235) );
  NAND2_X1 U9267 ( .A1(n6928), .A2(n6926), .ZN(P1_U3557) );
  XNOR2_X1 U9268 ( .A(n7515), .B(SI_2_), .ZN(n7514) );
  NAND2_X2 U9269 ( .A1(n11381), .A2(n11380), .ZN(n11382) );
  XNOR2_X1 U9270 ( .A(n7548), .B(n7547), .ZN(n10231) );
  AND2_X2 U9271 ( .A1(n6701), .A2(n6700), .ZN(n7446) );
  NOR2_X2 U9272 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6700) );
  NOR2_X2 U9273 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6701) );
  NAND2_X1 U9274 ( .A1(n13273), .A2(n6706), .ZN(n6705) );
  INV_X1 U9275 ( .A(n11690), .ZN(n7762) );
  NAND2_X1 U9276 ( .A1(n11671), .A2(n9237), .ZN(n6713) );
  NAND2_X1 U9277 ( .A1(n10804), .A2(n6716), .ZN(n6714) );
  NAND2_X1 U9278 ( .A1(n6714), .A2(n6715), .ZN(n11253) );
  OAI21_X1 U9279 ( .B1(n13311), .B2(n14530), .A(n13314), .ZN(n6719) );
  NAND2_X1 U9280 ( .A1(n8101), .A2(n8100), .ZN(n6720) );
  NAND2_X1 U9281 ( .A1(n8039), .A2(n7452), .ZN(n13460) );
  NAND2_X1 U9282 ( .A1(n15035), .A2(n6735), .ZN(n6734) );
  NAND3_X1 U9283 ( .A1(n6734), .A2(n6736), .A3(n6732), .ZN(n15058) );
  NAND3_X1 U9284 ( .A1(n6734), .A2(n6733), .A3(n6732), .ZN(n6731) );
  NOR2_X2 U9285 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n6740) );
  INV_X1 U9286 ( .A(n12339), .ZN(n6750) );
  AND2_X1 U9287 ( .A1(n12243), .A2(n12341), .ZN(n6753) );
  INV_X1 U9288 ( .A(n12256), .ZN(n6762) );
  OAI21_X1 U9289 ( .B1(n12256), .B2(n6757), .A(n6755), .ZN(n9338) );
  NAND2_X1 U9290 ( .A1(n12256), .A2(n12298), .ZN(n6758) );
  INV_X1 U9291 ( .A(n6770), .ZN(n6769) );
  OR2_X1 U9292 ( .A1(n9274), .A2(n12383), .ZN(n6770) );
  OR2_X1 U9293 ( .A1(n10075), .A2(n10076), .ZN(n6767) );
  INV_X1 U9294 ( .A(n7293), .ZN(n10380) );
  XNOR2_X2 U9295 ( .A(n6771), .B(n8456), .ZN(n12517) );
  NAND2_X1 U9296 ( .A1(n12328), .A2(n6773), .ZN(n6772) );
  INV_X1 U9297 ( .A(n9323), .ZN(n9320) );
  NAND2_X1 U9298 ( .A1(n13533), .A2(n6781), .ZN(n6779) );
  NAND2_X1 U9299 ( .A1(n11348), .A2(n6786), .ZN(n6785) );
  OAI21_X1 U9300 ( .B1(n11348), .B2(n6789), .A(n6785), .ZN(n6788) );
  INV_X1 U9301 ( .A(n6788), .ZN(n11355) );
  XNOR2_X1 U9302 ( .A(n11348), .B(n11292), .ZN(n11350) );
  INV_X1 U9303 ( .A(n11498), .ZN(n6791) );
  NAND2_X1 U9304 ( .A1(n11735), .A2(n11734), .ZN(n14552) );
  NAND2_X2 U9305 ( .A1(n11956), .A2(n11955), .ZN(n13549) );
  NAND2_X1 U9306 ( .A1(n14650), .A2(n6802), .ZN(n6800) );
  NAND3_X1 U9307 ( .A1(n6801), .A2(n6800), .A3(n6592), .ZN(n6803) );
  NAND3_X1 U9308 ( .A1(n6805), .A2(n9561), .A3(n14155), .ZN(n11394) );
  NAND2_X1 U9309 ( .A1(n13569), .A2(n13738), .ZN(n13761) );
  AND2_X2 U9310 ( .A1(n11394), .A2(n9713), .ZN(n12223) );
  NAND3_X1 U9311 ( .A1(n7334), .A2(n7331), .A3(n6818), .ZN(n6816) );
  NAND2_X1 U9312 ( .A1(n6816), .A2(n6817), .ZN(n6821) );
  INV_X1 U9313 ( .A(n14642), .ZN(n6819) );
  INV_X1 U9314 ( .A(n14444), .ZN(n6820) );
  INV_X1 U9315 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U9316 ( .A1(n7625), .A2(n7624), .ZN(n6827) );
  NAND2_X1 U9317 ( .A1(n7097), .A2(n6830), .ZN(n6829) );
  INV_X1 U9318 ( .A(n7514), .ZN(n6830) );
  NAND2_X1 U9319 ( .A1(n7496), .A2(n7495), .ZN(n6831) );
  INV_X1 U9320 ( .A(n7090), .ZN(n6833) );
  INV_X1 U9321 ( .A(n7091), .ZN(n6839) );
  NAND2_X1 U9322 ( .A1(n7069), .A2(n6842), .ZN(n6840) );
  OAI21_X1 U9323 ( .B1(n7069), .B2(n6844), .A(n6842), .ZN(n7562) );
  NAND2_X1 U9324 ( .A1(n7069), .A2(n7531), .ZN(n7548) );
  INV_X1 U9325 ( .A(n10766), .ZN(n6848) );
  INV_X1 U9326 ( .A(n6859), .ZN(n11530) );
  XNOR2_X2 U9327 ( .A(n6867), .B(P2_IR_REG_28__SCAN_IN), .ZN(n8027) );
  NOR2_X2 U9328 ( .A1(n7452), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7464) );
  NAND3_X1 U9329 ( .A1(n8036), .A2(n6868), .A3(n13248), .ZN(n13189) );
  INV_X1 U9330 ( .A(n6871), .ZN(n13188) );
  INV_X1 U9331 ( .A(n11743), .ZN(n6886) );
  NAND2_X1 U9332 ( .A1(n6886), .A2(n6887), .ZN(n13261) );
  NAND2_X1 U9333 ( .A1(n11239), .A2(n7700), .ZN(n6893) );
  NOR2_X2 U9334 ( .A1(n6899), .A2(n6476), .ZN(n8037) );
  INV_X1 U9335 ( .A(n6899), .ZN(n7965) );
  NAND3_X1 U9336 ( .A1(n7446), .A2(n6902), .A3(n7497), .ZN(n6900) );
  OAI21_X1 U9337 ( .B1(n13231), .B2(n6911), .A(n6909), .ZN(n13209) );
  INV_X1 U9338 ( .A(n13231), .ZN(n6912) );
  NOR2_X1 U9339 ( .A1(n7452), .A2(n6913), .ZN(n13443) );
  NAND2_X2 U9340 ( .A1(n11895), .A2(n9139), .ZN(n13758) );
  NAND2_X1 U9341 ( .A1(n13728), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n10227) );
  NAND3_X1 U9342 ( .A1(n9385), .A2(n9393), .A3(n10173), .ZN(n9427) );
  AND2_X2 U9343 ( .A1(n9384), .A2(n6580), .ZN(n10173) );
  AND2_X2 U9344 ( .A1(n10174), .A2(n9382), .ZN(n9385) );
  NOR2_X2 U9345 ( .A1(n9381), .A2(n9380), .ZN(n10174) );
  NAND2_X1 U9346 ( .A1(n11219), .A2(n6919), .ZN(n6918) );
  NAND2_X1 U9347 ( .A1(n14705), .A2(n14706), .ZN(n6925) );
  NAND3_X1 U9348 ( .A1(n6922), .A2(n10242), .A3(n6501), .ZN(n10625) );
  NAND2_X1 U9349 ( .A1(n6923), .A2(n6925), .ZN(n6922) );
  NAND2_X1 U9350 ( .A1(n14010), .A2(n7424), .ZN(n14005) );
  NAND2_X1 U9351 ( .A1(n14054), .A2(n6949), .ZN(n6946) );
  NAND2_X1 U9352 ( .A1(n11016), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U9353 ( .A1(n11699), .A2(n6962), .ZN(n6958) );
  NAND2_X1 U9354 ( .A1(n6958), .A2(n6959), .ZN(n14110) );
  NAND2_X1 U9355 ( .A1(n10736), .A2(n10324), .ZN(n6974) );
  INV_X1 U9356 ( .A(n6975), .ZN(n10318) );
  INV_X1 U9357 ( .A(n10123), .ZN(n6971) );
  OAI21_X1 U9358 ( .B1(n10737), .B2(n6976), .A(n6974), .ZN(n10794) );
  INV_X1 U9359 ( .A(n6977), .ZN(n11177) );
  OAI21_X1 U9360 ( .B1(n10837), .B2(n6981), .A(n6978), .ZN(n6977) );
  INV_X1 U9361 ( .A(n6979), .ZN(n6978) );
  OAI21_X1 U9362 ( .B1(n6982), .B2(n6980), .A(n6557), .ZN(n6979) );
  NAND2_X1 U9363 ( .A1(n6985), .A2(n11171), .ZN(n6981) );
  INV_X1 U9364 ( .A(n14486), .ZN(n7002) );
  NAND2_X1 U9365 ( .A1(n7749), .A2(n6584), .ZN(n7009) );
  NAND2_X1 U9366 ( .A1(n7009), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7806) );
  INV_X1 U9367 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U9368 ( .A1(n8409), .A2(n8408), .ZN(n7014) );
  NAND2_X1 U9369 ( .A1(n8392), .A2(n8391), .ZN(n7015) );
  NAND2_X1 U9370 ( .A1(n8298), .A2(n8297), .ZN(n7016) );
  NAND2_X1 U9371 ( .A1(n8281), .A2(n8280), .ZN(n7017) );
  XNOR2_X2 U9372 ( .A(n12701), .B(n7018), .ZN(n12555) );
  NAND2_X2 U9373 ( .A1(n8575), .A2(n8574), .ZN(n12701) );
  NAND3_X1 U9374 ( .A1(n8951), .A2(n7021), .A3(n7020), .ZN(n7019) );
  NAND2_X1 U9375 ( .A1(n8342), .A2(n9909), .ZN(n8358) );
  OAI21_X1 U9376 ( .B1(n10139), .B2(n7034), .A(n7033), .ZN(n10421) );
  NAND3_X1 U9377 ( .A1(n7032), .A2(n7031), .A3(n8809), .ZN(n10564) );
  NAND2_X1 U9378 ( .A1(n7033), .A2(n10139), .ZN(n7032) );
  OAI21_X1 U9379 ( .B1(n8288), .B2(n9581), .A(n8137), .ZN(n7037) );
  INV_X1 U9380 ( .A(n7037), .ZN(n7035) );
  NAND2_X1 U9381 ( .A1(n11331), .A2(n7041), .ZN(n7040) );
  NAND2_X1 U9382 ( .A1(n12670), .A2(n6575), .ZN(n8466) );
  NAND2_X1 U9383 ( .A1(n12642), .A2(n7046), .ZN(n8491) );
  NAND2_X2 U9384 ( .A1(n8475), .A2(n7187), .ZN(n12642) );
  NAND2_X1 U9385 ( .A1(n11040), .A2(n7050), .ZN(n7049) );
  OAI21_X1 U9386 ( .B1(n12620), .B2(n8783), .A(n8888), .ZN(n12609) );
  OAI21_X1 U9387 ( .B1(n7059), .B2(n12555), .A(n8911), .ZN(n7061) );
  NAND2_X1 U9388 ( .A1(n8568), .A2(n7065), .ZN(n7060) );
  NAND2_X1 U9389 ( .A1(n8568), .A2(n8903), .ZN(n12556) );
  AOI21_X2 U9390 ( .B1(n8568), .B2(n7062), .A(n7061), .ZN(n8744) );
  NAND2_X1 U9391 ( .A1(n8553), .A2(n8552), .ZN(n8555) );
  NAND2_X1 U9392 ( .A1(n8190), .A2(n8189), .ZN(n8192) );
  NAND2_X1 U9393 ( .A1(n8171), .A2(n8170), .ZN(n8173) );
  NAND2_X1 U9394 ( .A1(n9405), .A2(n7199), .ZN(n9412) );
  XNOR2_X1 U9395 ( .A(n7514), .B(n7513), .ZN(n9913) );
  NAND2_X1 U9396 ( .A1(n13198), .A2(n13197), .ZN(n8016) );
  NAND2_X1 U9397 ( .A1(n13214), .A2(n13223), .ZN(n7068) );
  INV_X1 U9398 ( .A(n11257), .ZN(n7076) );
  OAI21_X1 U9399 ( .B1(n7082), .B2(n7081), .A(n11672), .ZN(n7080) );
  NAND2_X1 U9400 ( .A1(n7084), .A2(n7085), .ZN(n11157) );
  NAND2_X1 U9401 ( .A1(n13279), .A2(n7093), .ZN(n7090) );
  INV_X1 U9402 ( .A(n7097), .ZN(n7513) );
  NAND2_X1 U9403 ( .A1(n9584), .A2(n7482), .ZN(n7495) );
  XNOR2_X1 U9404 ( .A(n8079), .B(n9244), .ZN(n7098) );
  NAND4_X1 U9405 ( .A1(n7102), .A2(n7101), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7099) );
  INV_X1 U9406 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7102) );
  XNOR2_X1 U9407 ( .A(n7580), .B(n7579), .ZN(n10521) );
  INV_X1 U9408 ( .A(n7108), .ZN(n12406) );
  OR2_X2 U9409 ( .A1(n10309), .A2(n10308), .ZN(n7115) );
  NAND2_X1 U9410 ( .A1(n13687), .A2(n7426), .ZN(n7126) );
  NAND3_X1 U9411 ( .A1(n13636), .A2(n7138), .A3(n13635), .ZN(n7137) );
  OAI21_X1 U9412 ( .B1(n13716), .B2(n7152), .A(n7149), .ZN(n13721) );
  OR2_X1 U9413 ( .A1(n13618), .A2(n7164), .ZN(n7163) );
  INV_X1 U9414 ( .A(n13617), .ZN(n7164) );
  NOR2_X2 U9415 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8107) );
  NAND2_X1 U9416 ( .A1(n7167), .A2(n7166), .ZN(n7171) );
  NAND2_X1 U9417 ( .A1(n12551), .A2(n7168), .ZN(n7167) );
  INV_X1 U9418 ( .A(n8325), .ZN(n7191) );
  NAND2_X1 U9419 ( .A1(n10132), .A2(n10131), .ZN(n10130) );
  INV_X1 U9420 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7199) );
  NOR2_X2 U9421 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9405) );
  NAND2_X1 U9422 ( .A1(n6695), .A2(n6472), .ZN(n7210) );
  NAND2_X1 U9423 ( .A1(n14111), .A2(n7206), .ZN(n7205) );
  NAND2_X1 U9424 ( .A1(n6695), .A2(n7212), .ZN(n14097) );
  INV_X1 U9425 ( .A(n7210), .ZN(n14096) );
  INV_X1 U9426 ( .A(n12013), .ZN(n7211) );
  NAND2_X1 U9427 ( .A1(n13996), .A2(n7220), .ZN(n7219) );
  OR2_X2 U9428 ( .A1(n13996), .A2(n14004), .ZN(n7221) );
  MUX2_X1 U9429 ( .A(n13021), .B(n6462), .S(n13138), .Z(n7228) );
  NAND2_X1 U9430 ( .A1(n7231), .A2(n7230), .ZN(n7856) );
  NAND2_X1 U9431 ( .A1(n7840), .A2(n7843), .ZN(n7231) );
  NAND2_X1 U9432 ( .A1(n7562), .A2(n7561), .ZN(n7248) );
  NAND2_X1 U9433 ( .A1(n7248), .A2(n7565), .ZN(n7580) );
  NAND2_X1 U9434 ( .A1(n7679), .A2(n7253), .ZN(n7249) );
  NAND3_X1 U9435 ( .A1(n7899), .A2(n7930), .A3(n7269), .ZN(n7264) );
  NAND2_X1 U9436 ( .A1(n7264), .A2(n7265), .ZN(n7946) );
  NAND2_X1 U9437 ( .A1(n7899), .A2(n7898), .ZN(n7915) );
  NAND2_X1 U9438 ( .A1(n12338), .A2(n7283), .ZN(n7282) );
  OAI211_X1 U9439 ( .C1(n12338), .C2(n7285), .A(n12341), .B(n7282), .ZN(n9373)
         );
  NOR2_X1 U9440 ( .A1(n10380), .A2(n7422), .ZN(n10462) );
  OR2_X2 U9441 ( .A1(n12289), .A2(n7299), .ZN(n7296) );
  NAND2_X1 U9442 ( .A1(n8686), .A2(n7314), .ZN(n8692) );
  NAND2_X1 U9443 ( .A1(n8686), .A2(n7313), .ZN(n7316) );
  NAND2_X1 U9444 ( .A1(n8686), .A2(n7315), .ZN(n8720) );
  INV_X2 U9445 ( .A(n9283), .ZN(n9261) );
  NAND2_X1 U9446 ( .A1(n7318), .A2(n8701), .ZN(n7317) );
  NAND2_X1 U9447 ( .A1(n14622), .A2(n7320), .ZN(n7319) );
  INV_X1 U9448 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7327) );
  NOR2_X2 U9449 ( .A1(n15134), .A2(n14341), .ZN(n14343) );
  INV_X1 U9450 ( .A(n14634), .ZN(n14635) );
  NAND2_X1 U9451 ( .A1(n14636), .A2(n14637), .ZN(n14633) );
  NAND2_X1 U9452 ( .A1(n14634), .A2(n7336), .ZN(n7334) );
  NOR2_X2 U9453 ( .A1(n14410), .A2(n14350), .ZN(n14352) );
  NAND2_X1 U9454 ( .A1(n7343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9539) );
  NOR2_X2 U9455 ( .A1(n14653), .A2(n14652), .ZN(n14650) );
  NAND2_X1 U9456 ( .A1(n13549), .A2(n6579), .ZN(n7353) );
  OAI211_X1 U9457 ( .C1(n13549), .C2(n7354), .A(n7353), .B(n7349), .ZN(n12233)
         );
  NAND4_X1 U9458 ( .A1(n7447), .A2(n7524), .A3(n7667), .A4(n7446), .ZN(n7961)
         );
  NAND3_X1 U9459 ( .A1(n7380), .A2(n7379), .A3(n9103), .ZN(n7378) );
  INV_X1 U9460 ( .A(n9095), .ZN(n7379) );
  INV_X1 U9461 ( .A(n9099), .ZN(n7383) );
  INV_X1 U9462 ( .A(n9098), .ZN(n7384) );
  NAND2_X1 U9463 ( .A1(n7385), .A2(n7386), .ZN(n9093) );
  NAND2_X1 U9464 ( .A1(n9081), .A2(n7387), .ZN(n7385) );
  NAND2_X1 U9465 ( .A1(n7390), .A2(n9084), .ZN(n7386) );
  NAND2_X1 U9466 ( .A1(n7389), .A2(n7388), .ZN(n7387) );
  INV_X1 U9467 ( .A(n9080), .ZN(n7392) );
  NAND2_X1 U9468 ( .A1(n9003), .A2(n7396), .ZN(n7395) );
  NOR2_X1 U9469 ( .A1(n7398), .A2(n6488), .ZN(n7397) );
  NAND2_X1 U9470 ( .A1(n7399), .A2(n6582), .ZN(n9052) );
  AOI21_X1 U9471 ( .B1(n9038), .B2(n9037), .A(n9035), .ZN(n9036) );
  NAND2_X1 U9472 ( .A1(n9058), .A2(n6576), .ZN(n7403) );
  INV_X1 U9473 ( .A(n9016), .ZN(n7414) );
  NAND2_X1 U9474 ( .A1(n13411), .A2(n15002), .ZN(n8072) );
  NOR2_X1 U9475 ( .A1(n12699), .A2(n12698), .ZN(n12777) );
  AND2_X1 U9476 ( .A1(n12697), .A2(n14475), .ZN(n12698) );
  INV_X1 U9477 ( .A(n8127), .ZN(n8132) );
  NAND2_X1 U9478 ( .A1(n11191), .A2(n11190), .ZN(n11402) );
  XNOR2_X1 U9479 ( .A(n7528), .B(n7527), .ZN(n10228) );
  INV_X1 U9480 ( .A(n9265), .ZN(n8148) );
  NAND2_X1 U9481 ( .A1(n13767), .A2(n7429), .ZN(n13813) );
  AND2_X2 U9482 ( .A1(n8617), .A2(n7428), .ZN(n8686) );
  NAND2_X1 U9483 ( .A1(n8744), .A2(n8919), .ZN(n8774) );
  NAND2_X1 U9484 ( .A1(n9325), .A2(n7425), .ZN(n9329) );
  OR2_X1 U9485 ( .A1(n9327), .A2(n9326), .ZN(n9328) );
  NAND2_X1 U9486 ( .A1(n12279), .A2(n9339), .ZN(n12339) );
  NOR2_X1 U9487 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n14329), .ZN(n14297) );
  NAND2_X1 U9488 ( .A1(n10859), .A2(n9285), .ZN(n10959) );
  NAND4_X1 U9489 ( .A1(n9590), .A2(n9589), .A3(n9588), .A4(n9587), .ZN(n10220)
         );
  INV_X2 U9490 ( .A(n7486), .ZN(n8029) );
  OR2_X1 U9491 ( .A1(n9283), .A2(n10036), .ZN(n9268) );
  OR2_X1 U9492 ( .A1(n14789), .A2(n14155), .ZN(n10354) );
  NAND2_X1 U9493 ( .A1(n8960), .A2(n8956), .ZN(n8959) );
  INV_X1 U9494 ( .A(n9024), .ZN(n9027) );
  OAI21_X2 U9495 ( .B1(n12562), .B2(n8671), .A(n8670), .ZN(n12551) );
  INV_X1 U9496 ( .A(n14128), .ZN(n12039) );
  NAND2_X1 U9497 ( .A1(n15133), .A2(n14467), .ZN(n12755) );
  INV_X1 U9498 ( .A(n12755), .ZN(n8743) );
  OR2_X1 U9499 ( .A1(n15127), .A2(n14470), .ZN(n12818) );
  INV_X1 U9500 ( .A(n12818), .ZN(n8727) );
  INV_X1 U9501 ( .A(n14043), .ZN(n14058) );
  AND2_X1 U9502 ( .A1(n8956), .A2(n12915), .ZN(n7420) );
  OR2_X1 U9503 ( .A1(n10105), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7421) );
  AND2_X1 U9504 ( .A1(n9276), .A2(n12382), .ZN(n7422) );
  OR2_X1 U9505 ( .A1(n13311), .A2(n13224), .ZN(n7423) );
  NOR2_X1 U9506 ( .A1(n12365), .A2(n9327), .ZN(n7425) );
  AND3_X1 U9507 ( .A1(n13798), .A2(n13686), .A3(n7418), .ZN(n7426) );
  INV_X1 U9508 ( .A(n14200), .ZN(n12046) );
  AND2_X1 U9509 ( .A1(n7678), .A2(n7666), .ZN(n7427) );
  INV_X1 U9510 ( .A(n13378), .ZN(n8070) );
  NOR2_X1 U9511 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), .ZN(
        n7428) );
  AND2_X1 U9512 ( .A1(n13766), .A2(n13765), .ZN(n7429) );
  INV_X1 U9513 ( .A(n13749), .ZN(n13748) );
  INV_X1 U9514 ( .A(n14951), .ZN(n13298) );
  NOR2_X1 U9515 ( .A1(n12484), .A2(n14451), .ZN(n7432) );
  OR2_X1 U9516 ( .A1(n10104), .A2(n10103), .ZN(n14991) );
  OR2_X1 U9517 ( .A1(n9803), .A2(n9818), .ZN(n7433) );
  NOR2_X1 U9518 ( .A1(n11666), .A2(n12370), .ZN(n7434) );
  INV_X1 U9519 ( .A(n11691), .ZN(n7761) );
  OR2_X1 U9520 ( .A1(n9440), .A2(n14272), .ZN(n7435) );
  INV_X1 U9521 ( .A(n8767), .ZN(n12532) );
  INV_X1 U9522 ( .A(n13788), .ZN(n11053) );
  INV_X1 U9523 ( .A(n13986), .ZN(n13997) );
  INV_X1 U9524 ( .A(n10165), .ZN(n8956) );
  NAND2_X1 U9525 ( .A1(n8981), .A2(n10165), .ZN(n8958) );
  OAI21_X1 U9526 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n8972) );
  AOI21_X1 U9527 ( .B1(n8979), .B2(n8978), .A(n8976), .ZN(n8977) );
  NAND2_X1 U9528 ( .A1(n8999), .A2(n8998), .ZN(n9003) );
  INV_X1 U9529 ( .A(n9025), .ZN(n9026) );
  AOI21_X1 U9530 ( .B1(n9052), .B2(n9051), .A(n9049), .ZN(n9050) );
  OAI21_X1 U9531 ( .B1(n9077), .B2(n9076), .A(n9075), .ZN(n9081) );
  INV_X1 U9532 ( .A(n14073), .ZN(n13696) );
  INV_X1 U9533 ( .A(n9086), .ZN(n9087) );
  OAI21_X1 U9534 ( .B1(n13711), .B2(n13710), .A(n13709), .ZN(n13712) );
  INV_X1 U9535 ( .A(n9088), .ZN(n9192) );
  INV_X1 U9536 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9390) );
  AND2_X1 U9537 ( .A1(n8651), .A2(n8650), .ZN(n8652) );
  INV_X1 U9538 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8106) );
  INV_X1 U9539 ( .A(n9243), .ZN(n8025) );
  OR2_X1 U9540 ( .A1(n13661), .A2(n13836), .ZN(n11528) );
  INV_X1 U9541 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9389) );
  INV_X1 U9542 ( .A(n8350), .ZN(n8349) );
  AND2_X1 U9543 ( .A1(n9353), .A2(n9259), .ZN(n9260) );
  NAND2_X1 U9544 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  INV_X1 U9545 ( .A(n8485), .ZN(n8484) );
  INV_X1 U9546 ( .A(n8578), .ZN(n8577) );
  INV_X1 U9547 ( .A(n10424), .ZN(n8633) );
  INV_X1 U9548 ( .A(n10084), .ZN(n8629) );
  AND2_X1 U9549 ( .A1(n7732), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7753) );
  INV_X1 U9550 ( .A(n10970), .ZN(n10966) );
  NAND2_X1 U9551 ( .A1(n13022), .A2(n11987), .ZN(n8086) );
  NAND2_X1 U9552 ( .A1(n11286), .A2(n11287), .ZN(n11288) );
  AND2_X1 U9553 ( .A1(n13753), .A2(n13754), .ZN(n13755) );
  INV_X1 U9554 ( .A(n14174), .ZN(n12047) );
  INV_X1 U9555 ( .A(n7587), .ZN(n7588) );
  INV_X1 U9556 ( .A(n8235), .ZN(n8234) );
  INV_X1 U9557 ( .A(n8461), .ZN(n8460) );
  INV_X1 U9558 ( .A(n8530), .ZN(n8529) );
  OR2_X1 U9559 ( .A1(n8498), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U9560 ( .A1(n8332), .A2(n8331), .ZN(n8350) );
  NAND2_X1 U9561 ( .A1(n8577), .A2(n8576), .ZN(n8593) );
  INV_X1 U9562 ( .A(n8200), .ZN(n8199) );
  NAND2_X1 U9563 ( .A1(n10560), .A2(n9258), .ZN(n9970) );
  NAND2_X1 U9564 ( .A1(n8476), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8479) );
  OR2_X1 U9565 ( .A1(n7655), .A2(n11462), .ZN(n7690) );
  INV_X1 U9566 ( .A(n9244), .ZN(n8102) );
  NAND2_X1 U9567 ( .A1(n11718), .A2(n11719), .ZN(n11720) );
  OR2_X1 U9568 ( .A1(n14575), .A2(n13833), .ZN(n12006) );
  INV_X1 U9569 ( .A(n13835), .ZN(n11789) );
  AND2_X1 U9570 ( .A1(n14646), .A2(n13601), .ZN(n10259) );
  OR2_X1 U9571 ( .A1(n13620), .A2(n13842), .ZN(n10594) );
  NAND2_X1 U9572 ( .A1(n7897), .A2(SI_24_), .ZN(n7898) );
  NOR2_X1 U9573 ( .A1(n14324), .A2(n14323), .ZN(n14315) );
  INV_X1 U9574 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10062) );
  OR2_X1 U9575 ( .A1(n8289), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8304) );
  AND2_X1 U9576 ( .A1(n9339), .A2(n9337), .ZN(n12278) );
  NAND2_X1 U9577 ( .A1(n9277), .A2(n10638), .ZN(n9278) );
  OR2_X1 U9578 ( .A1(n8304), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U9579 ( .A1(n8382), .A2(n8381), .ZN(n8400) );
  INV_X1 U9580 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n12142) );
  OR2_X1 U9581 ( .A1(n8593), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12526) );
  AND2_X1 U9582 ( .A1(n8837), .A2(n8838), .ZN(n11407) );
  OR2_X1 U9583 ( .A1(n8254), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U9584 ( .A1(n8199), .A2(n10637), .ZN(n8219) );
  INV_X1 U9585 ( .A(n12517), .ZN(n8947) );
  AND2_X1 U9586 ( .A1(n8734), .A2(n8776), .ZN(n12680) );
  INV_X1 U9587 ( .A(n10820), .ZN(n10988) );
  AND2_X1 U9588 ( .A1(n9376), .A2(n9490), .ZN(n9731) );
  NAND2_X1 U9589 ( .A1(n8694), .A2(n8717), .ZN(n8697) );
  NAND2_X1 U9590 ( .A1(n8209), .A2(n8208), .ZN(n8211) );
  OR2_X1 U9591 ( .A1(n7792), .A2(n7791), .ZN(n7834) );
  INV_X1 U9592 ( .A(n11173), .ZN(n14970) );
  OR2_X1 U9593 ( .A1(n7888), .A2(n12972), .ZN(n7924) );
  NOR2_X1 U9594 ( .A1(n8956), .A2(n12834), .ZN(n9891) );
  OR2_X1 U9595 ( .A1(n7846), .A2(n12931), .ZN(n7870) );
  INV_X1 U9596 ( .A(n9213), .ZN(n9218) );
  OR2_X1 U9597 ( .A1(n9952), .A2(n9953), .ZN(n10283) );
  INV_X1 U9598 ( .A(n13255), .ZN(n13245) );
  INV_X1 U9599 ( .A(n9238), .ZN(n13289) );
  NAND2_X1 U9600 ( .A1(n10742), .A2(n10743), .ZN(n10503) );
  INV_X1 U9601 ( .A(n8055), .ZN(n10108) );
  INV_X1 U9602 ( .A(n14503), .ZN(n14523) );
  INV_X1 U9603 ( .A(n10648), .ZN(n10654) );
  OR2_X1 U9604 ( .A1(n8054), .A2(n8055), .ZN(n9884) );
  INV_X1 U9605 ( .A(n11929), .ZN(n11914) );
  INV_X1 U9606 ( .A(n13479), .ZN(n11856) );
  NOR2_X1 U9607 ( .A1(n11883), .A2(n13494), .ZN(n11896) );
  INV_X1 U9608 ( .A(n11960), .ZN(n11943) );
  INV_X1 U9609 ( .A(n11915), .ZN(n11897) );
  NOR2_X1 U9610 ( .A1(n11533), .A2(n11532), .ZN(n11586) );
  OR2_X1 U9611 ( .A1(n14281), .A2(n14284), .ZN(n9400) );
  INV_X1 U9612 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10599) );
  INV_X1 U9613 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11294) );
  AND2_X1 U9614 ( .A1(n13682), .A2(n13683), .ZN(n14145) );
  OR2_X1 U9615 ( .A1(n14564), .A2(n11372), .ZN(n11373) );
  NOR2_X1 U9616 ( .A1(n10609), .A2(n11294), .ZN(n11005) );
  AND2_X1 U9617 ( .A1(n9566), .A2(n10393), .ZN(n10364) );
  OR2_X1 U9618 ( .A1(n14739), .A2(n10361), .ZN(n14712) );
  INV_X1 U9619 ( .A(n13785), .ZN(n10630) );
  INV_X1 U9620 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U9621 ( .A1(n7741), .A2(n7726), .ZN(n7742) );
  NAND2_X1 U9622 ( .A1(n10861), .A2(n10860), .ZN(n10859) );
  NAND2_X1 U9623 ( .A1(n9270), .A2(n9272), .ZN(n10033) );
  INV_X1 U9624 ( .A(n12360), .ZN(n12334) );
  AND2_X1 U9625 ( .A1(n9344), .A2(n9731), .ZN(n12341) );
  AND2_X1 U9626 ( .A1(n8759), .A2(n8758), .ZN(n12525) );
  AND3_X1 U9627 ( .A1(n8474), .A2(n8473), .A3(n8472), .ZN(n12654) );
  AND4_X1 U9628 ( .A1(n8356), .A2(n8355), .A3(n8354), .A4(n8353), .ZN(n11328)
         );
  INV_X1 U9629 ( .A(n10015), .ZN(n15016) );
  INV_X1 U9630 ( .A(n15040), .ZN(n15086) );
  XNOR2_X1 U9631 ( .A(n8744), .B(n8944), .ZN(n12534) );
  AND2_X1 U9632 ( .A1(n8679), .A2(n9733), .ZN(n12666) );
  NAND2_X1 U9633 ( .A1(n15114), .A2(n10136), .ZN(n12691) );
  INV_X1 U9634 ( .A(n15111), .ZN(n12687) );
  XNOR2_X1 U9635 ( .A(n8612), .B(P3_IR_REG_22__SCAN_IN), .ZN(n10560) );
  XNOR2_X1 U9636 ( .A(n12924), .B(n12917), .ZN(n12918) );
  NOR2_X1 U9637 ( .A1(n10122), .A2(n7420), .ZN(n10123) );
  OR2_X1 U9638 ( .A1(n9899), .A2(n9897), .ZN(n14491) );
  OR2_X1 U9639 ( .A1(n9152), .A2(n7539), .ZN(n7541) );
  OR2_X1 U9640 ( .A1(n9805), .A2(n9804), .ZN(n9809) );
  INV_X1 U9641 ( .A(n13224), .ZN(n14510) );
  AND2_X1 U9642 ( .A1(n14948), .A2(n10984), .ZN(n14509) );
  NAND2_X1 U9643 ( .A1(n8960), .A2(n10165), .ZN(n10158) );
  AND2_X1 U9644 ( .A1(n11311), .A2(n11255), .ZN(n14530) );
  AND2_X1 U9645 ( .A1(n9897), .A2(n10108), .ZN(n13398) );
  INV_X1 U9646 ( .A(n14530), .ZN(n14983) );
  INV_X1 U9647 ( .A(n14651), .ZN(n14576) );
  AND4_X1 U9648 ( .A1(n12033), .A2(n12032), .A3(n12031), .A4(n12030), .ZN(
        n13741) );
  INV_X1 U9649 ( .A(n13956), .ZN(n14690) );
  INV_X1 U9650 ( .A(n13800), .ZN(n14098) );
  AND2_X1 U9651 ( .A1(n13664), .A2(n13665), .ZN(n13669) );
  INV_X1 U9652 ( .A(n14712), .ZN(n14735) );
  AND2_X1 U9653 ( .A1(n9559), .A2(n9558), .ZN(n10355) );
  OR2_X1 U9654 ( .A1(n9565), .A2(n9657), .ZN(n14799) );
  INV_X1 U9655 ( .A(n14803), .ZN(n14769) );
  AND2_X1 U9656 ( .A1(n9563), .A2(n9562), .ZN(n14795) );
  INV_X1 U9657 ( .A(n14795), .ZN(n14784) );
  AND2_X1 U9658 ( .A1(n10358), .A2(n9556), .ZN(n10219) );
  OR2_X1 U9659 ( .A1(n9518), .A2(n9661), .ZN(n10353) );
  INV_X1 U9660 ( .A(n9561), .ZN(n9565) );
  XNOR2_X1 U9661 ( .A(n7581), .B(SI_6_), .ZN(n7579) );
  INV_X1 U9662 ( .A(n9371), .ZN(n9372) );
  INV_X1 U9663 ( .A(n12341), .ZN(n12347) );
  INV_X1 U9664 ( .A(n12618), .ZN(n12364) );
  INV_X1 U9665 ( .A(n11328), .ZN(n12372) );
  INV_X1 U9666 ( .A(n15055), .ZN(n15096) );
  AND2_X1 U9667 ( .A1(n12657), .A2(n12656), .ZN(n12736) );
  NAND2_X1 U9668 ( .A1(n9983), .A2(n15111), .ZN(n15117) );
  INV_X1 U9669 ( .A(n15133), .ZN(n15131) );
  INV_X1 U9670 ( .A(n9512), .ZN(n9513) );
  AND2_X1 U9671 ( .A1(n8696), .A2(n8695), .ZN(n12820) );
  INV_X1 U9672 ( .A(SI_11_), .ZN(n12095) );
  INV_X1 U9673 ( .A(n15101), .ZN(n10904) );
  INV_X1 U9674 ( .A(n10060), .ZN(n10065) );
  INV_X1 U9675 ( .A(n13014), .ZN(n14488) );
  OR2_X1 U9676 ( .A1(n9899), .A2(n9895), .ZN(n14490) );
  OR2_X1 U9677 ( .A1(n9255), .A2(n9254), .ZN(n9256) );
  AND2_X1 U9678 ( .A1(n11433), .A2(n11432), .ZN(n14542) );
  AOI21_X1 U9679 ( .B1(n12924), .B2(n8070), .A(n8069), .ZN(n8071) );
  OR2_X1 U9680 ( .A1(n10104), .A2(n14958), .ZN(n14999) );
  INV_X1 U9681 ( .A(n13277), .ZN(n13432) );
  AND2_X1 U9682 ( .A1(n14542), .A2(n14541), .ZN(n14551) );
  AND2_X1 U9683 ( .A1(n14974), .A2(n14973), .ZN(n14996) );
  INV_X1 U9684 ( .A(n14955), .ZN(n14956) );
  INV_X1 U9685 ( .A(n6463), .ZN(n10984) );
  INV_X1 U9686 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9856) );
  INV_X1 U9687 ( .A(n14105), .ZN(n14225) );
  INV_X1 U9688 ( .A(n14657), .ZN(n13567) );
  NAND4_X1 U9689 ( .A1(n11965), .A2(n11964), .A3(n11963), .A4(n11962), .ZN(
        n13823) );
  INV_X1 U9690 ( .A(n11290), .ZN(n13840) );
  OR2_X1 U9691 ( .A1(n14739), .A2(n10365), .ZN(n14160) );
  OR2_X1 U9692 ( .A1(n14739), .A2(n14795), .ZN(n14126) );
  INV_X1 U9693 ( .A(n14819), .ZN(n14816) );
  INV_X1 U9694 ( .A(n14807), .ZN(n14805) );
  OR2_X1 U9695 ( .A1(n10353), .A2(n9516), .ZN(n14744) );
  INV_X1 U9696 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10496) );
  INV_X1 U9697 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9842) );
  INV_X1 U9698 ( .A(n12385), .ZN(P3_U3897) );
  NAND2_X1 U9699 ( .A1(n8103), .A2(n7423), .ZN(P2_U3236) );
  NAND2_X1 U9700 ( .A1(n8072), .A2(n8071), .ZN(P2_U3527) );
  NOR2_X1 U9701 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n7441) );
  NOR2_X2 U9702 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7440) );
  NOR2_X2 U9703 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7439) );
  AND4_X2 U9704 ( .A1(n7441), .A2(n7440), .A3(n7439), .A4(n7545), .ZN(n7447)
         );
  NOR2_X2 U9705 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7443) );
  AND3_X2 U9706 ( .A1(n7444), .A2(n7443), .A3(n7442), .ZN(n7667) );
  INV_X1 U9707 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7451) );
  INV_X1 U9708 ( .A(n7464), .ZN(n7454) );
  INV_X1 U9709 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7457) );
  NAND2_X1 U9710 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7456) );
  NAND2_X2 U9711 ( .A1(n9803), .A2(n8134), .ZN(n7919) );
  INV_X1 U9712 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9478) );
  INV_X1 U9713 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9477) );
  AND2_X1 U9714 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7459) );
  AND2_X1 U9715 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7460) );
  NAND2_X1 U9716 ( .A1(n9582), .A2(n7460), .ZN(n7482) );
  XNOR2_X1 U9717 ( .A(n7496), .B(n7495), .ZN(n9712) );
  NAND2_X1 U9718 ( .A1(n7469), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7476) );
  INV_X1 U9719 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7470) );
  NAND2_X1 U9720 ( .A1(n7506), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U9721 ( .A1(n7486), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7473) );
  INV_X1 U9722 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10119) );
  INV_X1 U9723 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10110) );
  NAND2_X1 U9724 ( .A1(n7486), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7478) );
  NAND4_X2 U9725 ( .A1(n7480), .A2(n7479), .A3(n7478), .A4(n7477), .ZN(n8960)
         );
  NAND2_X1 U9726 ( .A1(n9139), .A2(SI_0_), .ZN(n7481) );
  NAND2_X1 U9727 ( .A1(n7481), .A2(n8135), .ZN(n7483) );
  AND2_X1 U9728 ( .A1(n7483), .A2(n7482), .ZN(n13469) );
  INV_X1 U9729 ( .A(n10158), .ZN(n7484) );
  OR2_X1 U9730 ( .A1(n13048), .A2(n10121), .ZN(n7485) );
  NAND2_X1 U9731 ( .A1(n8080), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U9732 ( .A1(n7486), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7491) );
  INV_X1 U9733 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7488) );
  NAND2_X1 U9734 ( .A1(n7506), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7489) );
  OR2_X1 U9735 ( .A1(n7919), .A2(n9505), .ZN(n7504) );
  INV_X1 U9736 ( .A(SI_1_), .ZN(n9469) );
  OR2_X1 U9737 ( .A1(n7493), .A2(n9913), .ZN(n7502) );
  NOR2_X1 U9738 ( .A1(n7497), .A2(n13444), .ZN(n7498) );
  MUX2_X1 U9739 ( .A(n13444), .B(n7498), .S(P2_IR_REG_2__SCAN_IN), .Z(n7499)
         );
  INV_X1 U9740 ( .A(n7499), .ZN(n7501) );
  INV_X1 U9741 ( .A(n7524), .ZN(n7500) );
  NAND2_X1 U9742 ( .A1(n7501), .A2(n7500), .ZN(n9818) );
  INV_X1 U9743 ( .A(n9224), .ZN(n10207) );
  NAND2_X1 U9744 ( .A1(n10205), .A2(n10207), .ZN(n10204) );
  OR2_X1 U9745 ( .A1(n8973), .A2(n10321), .ZN(n7505) );
  NAND2_X1 U9746 ( .A1(n10204), .A2(n7505), .ZN(n10404) );
  OR2_X1 U9747 ( .A1(n8029), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U9748 ( .A1(n8080), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U9749 ( .A1(n9148), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7508) );
  NAND2_X1 U9750 ( .A1(n8081), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7507) );
  NAND4_X2 U9751 ( .A1(n7507), .A2(n7509), .A3(n7508), .A4(n7510), .ZN(n13047)
         );
  OR2_X1 U9752 ( .A1(n7524), .A2(n13444), .ZN(n7512) );
  XNOR2_X1 U9753 ( .A(n7512), .B(n7511), .ZN(n13051) );
  NAND2_X1 U9754 ( .A1(n7515), .A2(SI_2_), .ZN(n7516) );
  MUX2_X1 U9755 ( .A(n9492), .B(n9502), .S(n9582), .Z(n7529) );
  XNOR2_X1 U9756 ( .A(n7529), .B(SI_3_), .ZN(n7527) );
  OR2_X1 U9757 ( .A1(n7493), .A2(n10228), .ZN(n7518) );
  OR2_X1 U9758 ( .A1(n7919), .A2(n9502), .ZN(n7517) );
  OAI211_X1 U9759 ( .C1(n9803), .C2(n13051), .A(n7518), .B(n7517), .ZN(n14939)
         );
  XNOR2_X1 U9760 ( .A(n13047), .B(n14939), .ZN(n9225) );
  INV_X1 U9761 ( .A(n9225), .ZN(n10409) );
  NAND2_X1 U9762 ( .A1(n10404), .A2(n10409), .ZN(n10403) );
  INV_X1 U9763 ( .A(n13047), .ZN(n7974) );
  INV_X1 U9764 ( .A(n14939), .ZN(n10417) );
  NAND2_X1 U9765 ( .A1(n7974), .A2(n10417), .ZN(n7519) );
  NAND2_X1 U9766 ( .A1(n10403), .A2(n7519), .ZN(n10664) );
  NAND2_X1 U9767 ( .A1(n8080), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7522) );
  AND2_X1 U9768 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7535) );
  INV_X1 U9769 ( .A(n7535), .ZN(n7537) );
  OAI21_X1 U9770 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7537), .ZN(n10749) );
  OR2_X1 U9771 ( .A1(n8029), .A2(n10749), .ZN(n7521) );
  NAND2_X1 U9772 ( .A1(n8081), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U9773 ( .A1(n9148), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U9774 ( .A1(n7544), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7526) );
  XNOR2_X1 U9775 ( .A(n7526), .B(n7525), .ZN(n9823) );
  INV_X1 U9776 ( .A(n7529), .ZN(n7530) );
  NAND2_X1 U9777 ( .A1(n7530), .A2(SI_3_), .ZN(n7531) );
  MUX2_X1 U9778 ( .A(n10232), .B(n9504), .S(n9582), .Z(n7549) );
  OR2_X1 U9779 ( .A1(n7493), .A2(n10231), .ZN(n7533) );
  OR2_X1 U9780 ( .A1(n7919), .A2(n9504), .ZN(n7532) );
  OAI211_X1 U9781 ( .C1(n9803), .C2(n9823), .A(n7533), .B(n7532), .ZN(n10743)
         );
  NAND2_X1 U9782 ( .A1(n10664), .A2(n10668), .ZN(n10663) );
  NAND2_X1 U9783 ( .A1(n10742), .A2(n6885), .ZN(n7534) );
  NAND2_X1 U9784 ( .A1(n10663), .A2(n7534), .ZN(n10508) );
  NAND2_X1 U9785 ( .A1(n7535), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7571) );
  INV_X1 U9786 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7536) );
  NAND2_X1 U9787 ( .A1(n7537), .A2(n7536), .ZN(n7538) );
  NAND2_X1 U9788 ( .A1(n7571), .A2(n7538), .ZN(n10842) );
  OR2_X1 U9789 ( .A1(n8029), .A2(n10842), .ZN(n7543) );
  NAND2_X1 U9790 ( .A1(n7506), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7542) );
  INV_X1 U9791 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7539) );
  NAND2_X1 U9792 ( .A1(n7559), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7546) );
  XNOR2_X1 U9793 ( .A(n7546), .B(n7545), .ZN(n14858) );
  INV_X1 U9794 ( .A(n7549), .ZN(n7550) );
  MUX2_X1 U9795 ( .A(n9493), .B(n9503), .S(n9582), .Z(n7563) );
  XNOR2_X1 U9796 ( .A(n7562), .B(n7561), .ZN(n10251) );
  OR2_X1 U9797 ( .A1(n7493), .A2(n10251), .ZN(n7552) );
  OR2_X1 U9798 ( .A1(n7919), .A2(n9503), .ZN(n7551) );
  XNOR2_X1 U9799 ( .A(n13045), .B(n10831), .ZN(n9228) );
  INV_X1 U9800 ( .A(n9228), .ZN(n10507) );
  NAND2_X1 U9801 ( .A1(n10508), .A2(n10507), .ZN(n10506) );
  INV_X1 U9802 ( .A(n13045), .ZN(n7553) );
  NAND2_X1 U9803 ( .A1(n7553), .A2(n10839), .ZN(n7554) );
  NAND2_X1 U9804 ( .A1(n10506), .A2(n7554), .ZN(n10655) );
  NAND2_X1 U9805 ( .A1(n8081), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9806 ( .A1(n8080), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7557) );
  XNOR2_X1 U9807 ( .A(n7571), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n10850) );
  NAND2_X1 U9808 ( .A1(n7486), .A2(n10850), .ZN(n7556) );
  NAND2_X1 U9809 ( .A1(n9148), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7555) );
  OR2_X1 U9810 ( .A1(n7668), .A2(n13444), .ZN(n7560) );
  INV_X1 U9811 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7577) );
  XNOR2_X1 U9812 ( .A(n7560), .B(n7577), .ZN(n13071) );
  INV_X1 U9813 ( .A(n7563), .ZN(n7564) );
  NAND2_X1 U9814 ( .A1(n7564), .A2(SI_5_), .ZN(n7565) );
  MUX2_X1 U9815 ( .A(n9496), .B(n9501), .S(n9582), .Z(n7581) );
  OR2_X1 U9816 ( .A1(n7919), .A2(n9501), .ZN(n7566) );
  NAND2_X1 U9817 ( .A1(n10655), .A2(n10654), .ZN(n10653) );
  OR2_X1 U9818 ( .A1(n13044), .A2(n10855), .ZN(n7567) );
  NAND2_X1 U9819 ( .A1(n10653), .A2(n7567), .ZN(n10805) );
  INV_X1 U9820 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7569) );
  INV_X1 U9821 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7568) );
  OAI21_X1 U9822 ( .B1(n7571), .B2(n7569), .A(n7568), .ZN(n7572) );
  NAND2_X1 U9823 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n7570) );
  NOR2_X1 U9824 ( .A1(n7571), .A2(n7570), .ZN(n7598) );
  INV_X1 U9825 ( .A(n7598), .ZN(n7600) );
  NAND2_X1 U9826 ( .A1(n7572), .A2(n7600), .ZN(n10952) );
  OR2_X1 U9827 ( .A1(n8029), .A2(n10952), .ZN(n7576) );
  NAND2_X1 U9828 ( .A1(n8080), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U9829 ( .A1(n8081), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7574) );
  NAND2_X1 U9830 ( .A1(n9148), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7573) );
  NAND4_X1 U9831 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(n13043)
         );
  NAND2_X1 U9832 ( .A1(n7668), .A2(n7577), .ZN(n7592) );
  NAND2_X1 U9833 ( .A1(n7592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7578) );
  XNOR2_X1 U9834 ( .A(n7578), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14873) );
  AOI22_X1 U9835 ( .A1(n7808), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7807), .B2(
        n14873), .ZN(n7584) );
  INV_X1 U9836 ( .A(n7581), .ZN(n7582) );
  MUX2_X1 U9837 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9139), .Z(n7590) );
  XNOR2_X1 U9838 ( .A(n7589), .B(n7587), .ZN(n10591) );
  INV_X2 U9839 ( .A(n7493), .ZN(n7612) );
  NAND2_X1 U9840 ( .A1(n10591), .A2(n7612), .ZN(n7583) );
  NAND2_X1 U9841 ( .A1(n7584), .A2(n7583), .ZN(n10954) );
  XNOR2_X1 U9842 ( .A(n13043), .B(n10954), .ZN(n9229) );
  INV_X1 U9843 ( .A(n13043), .ZN(n7585) );
  NAND2_X1 U9844 ( .A1(n7585), .A2(n10927), .ZN(n7586) );
  NAND2_X1 U9845 ( .A1(n7590), .A2(SI_7_), .ZN(n7591) );
  MUX2_X1 U9846 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9139), .Z(n7610) );
  XNOR2_X1 U9847 ( .A(n7609), .B(n7607), .ZN(n10595) );
  NAND2_X1 U9848 ( .A1(n10595), .A2(n7612), .ZN(n7597) );
  NAND2_X1 U9849 ( .A1(n7594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7593) );
  INV_X1 U9850 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n12106) );
  MUX2_X1 U9851 ( .A(n7593), .B(P2_IR_REG_31__SCAN_IN), .S(n12106), .Z(n7595)
         );
  NAND2_X1 U9852 ( .A1(n7595), .A2(n7615), .ZN(n9829) );
  INV_X1 U9853 ( .A(n9829), .ZN(n9848) );
  AOI22_X1 U9854 ( .A1(n7808), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7807), .B2(
        n9848), .ZN(n7596) );
  NAND2_X1 U9855 ( .A1(n7598), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7634) );
  INV_X1 U9856 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7599) );
  NAND2_X1 U9857 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  NAND2_X1 U9858 ( .A1(n7634), .A2(n7601), .ZN(n11181) );
  OR2_X1 U9859 ( .A1(n8029), .A2(n11181), .ZN(n7605) );
  NAND2_X1 U9860 ( .A1(n7506), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U9861 ( .A1(n8080), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9862 ( .A1(n9148), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7602) );
  NAND4_X1 U9863 ( .A1(n7605), .A2(n7604), .A3(n7603), .A4(n7602), .ZN(n13042)
         );
  XNOR2_X1 U9864 ( .A(n14970), .B(n13042), .ZN(n10970) );
  NAND2_X1 U9865 ( .A1(n13042), .A2(n11173), .ZN(n7606) );
  NAND2_X1 U9866 ( .A1(n7610), .A2(SI_8_), .ZN(n7611) );
  MUX2_X1 U9867 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9139), .Z(n7626) );
  XNOR2_X1 U9868 ( .A(n7625), .B(n7623), .ZN(n10996) );
  NAND2_X1 U9869 ( .A1(n10996), .A2(n7612), .ZN(n7618) );
  NAND2_X1 U9870 ( .A1(n7615), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7613) );
  MUX2_X1 U9871 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7613), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7614) );
  INV_X1 U9872 ( .A(n7614), .ZN(n7616) );
  NOR2_X1 U9873 ( .A1(n7615), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7628) );
  NOR2_X1 U9874 ( .A1(n7616), .A2(n7628), .ZN(n9864) );
  AOI22_X1 U9875 ( .A1(n7808), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7807), .B2(
        n9864), .ZN(n7617) );
  NAND2_X1 U9876 ( .A1(n8080), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7622) );
  NAND2_X1 U9877 ( .A1(n9148), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7621) );
  XNOR2_X1 U9878 ( .A(n7634), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n11277) );
  NAND2_X1 U9879 ( .A1(n7486), .A2(n11277), .ZN(n7620) );
  NAND2_X1 U9880 ( .A1(n7506), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7619) );
  NAND4_X1 U9881 ( .A1(n7622), .A2(n7621), .A3(n7620), .A4(n7619), .ZN(n13041)
         );
  INV_X1 U9882 ( .A(n13041), .ZN(n7987) );
  XNOR2_X1 U9883 ( .A(n11316), .B(n7987), .ZN(n11156) );
  NAND2_X1 U9884 ( .A1(n7626), .A2(SI_9_), .ZN(n7627) );
  MUX2_X1 U9885 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9139), .Z(n7645) );
  XNOR2_X1 U9886 ( .A(n7644), .B(n7642), .ZN(n11001) );
  INV_X1 U9887 ( .A(n7628), .ZN(n7651) );
  NAND2_X1 U9888 ( .A1(n7651), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7629) );
  XNOR2_X1 U9889 ( .A(n7629), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U9890 ( .A1(n7808), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7807), .B2(
        n9955), .ZN(n7630) );
  INV_X1 U9891 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7632) );
  INV_X1 U9892 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7631) );
  OAI21_X1 U9893 ( .B1(n7634), .B2(n7632), .A(n7631), .ZN(n7635) );
  NAND2_X1 U9894 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n7633) );
  NAND2_X1 U9895 ( .A1(n7635), .A2(n7655), .ZN(n11306) );
  OR2_X1 U9896 ( .A1(n8029), .A2(n11306), .ZN(n7639) );
  NAND2_X1 U9897 ( .A1(n7506), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9898 ( .A1(n8080), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7637) );
  NAND2_X1 U9899 ( .A1(n9148), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7636) );
  NAND4_X1 U9900 ( .A1(n7639), .A2(n7638), .A3(n7637), .A4(n7636), .ZN(n13040)
         );
  INV_X1 U9901 ( .A(n13040), .ZN(n7989) );
  XNOR2_X1 U9902 ( .A(n11308), .B(n7989), .ZN(n11254) );
  NAND2_X1 U9903 ( .A1(n11253), .A2(n11254), .ZN(n7641) );
  NAND2_X1 U9904 ( .A1(n11308), .A2(n13040), .ZN(n7640) );
  NAND2_X1 U9905 ( .A1(n7641), .A2(n7640), .ZN(n11239) );
  NAND2_X1 U9906 ( .A1(n7644), .A2(n7643), .ZN(n7647) );
  NAND2_X1 U9907 ( .A1(n7645), .A2(SI_10_), .ZN(n7646) );
  MUX2_X1 U9908 ( .A(n9695), .B(n9692), .S(n9139), .Z(n7648) );
  INV_X1 U9909 ( .A(n7648), .ZN(n7649) );
  NAND2_X1 U9910 ( .A1(n7649), .A2(SI_11_), .ZN(n7650) );
  XNOR2_X1 U9911 ( .A(n7663), .B(n7662), .ZN(n11098) );
  NAND2_X1 U9912 ( .A1(n11098), .A2(n7612), .ZN(n7654) );
  OAI21_X1 U9913 ( .B1(n7651), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7652) );
  XNOR2_X1 U9914 ( .A(n7652), .B(P2_IR_REG_11__SCAN_IN), .ZN(n14888) );
  AOI22_X1 U9915 ( .A1(n7808), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7807), .B2(
        n14888), .ZN(n7653) );
  INV_X1 U9916 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11462) );
  NAND2_X1 U9917 ( .A1(n7655), .A2(n11462), .ZN(n7656) );
  NAND2_X1 U9918 ( .A1(n7690), .A2(n7656), .ZN(n11465) );
  OR2_X1 U9919 ( .A1(n8029), .A2(n11465), .ZN(n7660) );
  NAND2_X1 U9920 ( .A1(n7506), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U9921 ( .A1(n8080), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U9922 ( .A1(n9148), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7657) );
  NAND4_X1 U9923 ( .A1(n7660), .A2(n7659), .A3(n7658), .A4(n7657), .ZN(n13039)
         );
  AND2_X1 U9924 ( .A1(n11467), .A2(n13039), .ZN(n11421) );
  MUX2_X1 U9925 ( .A(n9842), .B(n9840), .S(n9139), .Z(n7664) );
  INV_X1 U9926 ( .A(n7664), .ZN(n7665) );
  NAND2_X1 U9927 ( .A1(n7665), .A2(SI_12_), .ZN(n7666) );
  XNOR2_X1 U9928 ( .A(n7677), .B(n7427), .ZN(n11215) );
  NAND2_X1 U9929 ( .A1(n11215), .A2(n7612), .ZN(n7671) );
  NAND2_X1 U9930 ( .A1(n7668), .A2(n7667), .ZN(n7680) );
  NAND2_X1 U9931 ( .A1(n7680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7669) );
  XNOR2_X1 U9932 ( .A(n7669), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U9933 ( .A1(n7808), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7807), .B2(
        n9959), .ZN(n7670) );
  NAND2_X1 U9934 ( .A1(n7506), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9935 ( .A1(n8080), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7674) );
  XNOR2_X1 U9936 ( .A(n7690), .B(P2_REG3_REG_12__SCAN_IN), .ZN(n11573) );
  NAND2_X1 U9937 ( .A1(n7486), .A2(n11573), .ZN(n7673) );
  NAND2_X1 U9938 ( .A1(n9148), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7672) );
  NAND4_X1 U9939 ( .A1(n7675), .A2(n7674), .A3(n7673), .A4(n7672), .ZN(n13038)
         );
  OR2_X1 U9940 ( .A1(n11565), .A2(n13038), .ZN(n7696) );
  INV_X1 U9941 ( .A(n7696), .ZN(n7676) );
  XNOR2_X1 U9942 ( .A(n11565), .B(n13038), .ZN(n9234) );
  NOR2_X1 U9943 ( .A1(n7676), .A2(n11426), .ZN(n7698) );
  MUX2_X1 U9944 ( .A(n9909), .B(n9856), .S(n9139), .Z(n7702) );
  NAND2_X1 U9945 ( .A1(n11375), .A2(n7612), .ZN(n7686) );
  INV_X1 U9946 ( .A(n7680), .ZN(n7682) );
  NAND2_X1 U9947 ( .A1(n7682), .A2(n7681), .ZN(n7728) );
  NAND2_X1 U9948 ( .A1(n7728), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7683) );
  MUX2_X1 U9949 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7683), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n7684) );
  OR2_X1 U9950 ( .A1(n7728), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U9951 ( .A1(n7684), .A2(n7708), .ZN(n14911) );
  INV_X1 U9952 ( .A(n14911), .ZN(n10286) );
  AOI22_X1 U9953 ( .A1(n7808), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7807), .B2(
        n10286), .ZN(n7685) );
  NAND2_X1 U9954 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n7687) );
  NOR2_X1 U9955 ( .A1(n7690), .A2(n7687), .ZN(n7712) );
  INV_X1 U9956 ( .A(n7712), .ZN(n7713) );
  INV_X1 U9957 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7689) );
  INV_X1 U9958 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7688) );
  OAI21_X1 U9959 ( .B1(n7690), .B2(n7689), .A(n7688), .ZN(n7691) );
  NAND2_X1 U9960 ( .A1(n7713), .A2(n7691), .ZN(n11613) );
  OR2_X1 U9961 ( .A1(n8029), .A2(n11613), .ZN(n7695) );
  NAND2_X1 U9962 ( .A1(n8080), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7694) );
  NAND2_X1 U9963 ( .A1(n9148), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U9964 ( .A1(n7506), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7692) );
  NAND4_X1 U9965 ( .A1(n7695), .A2(n7694), .A3(n7693), .A4(n7692), .ZN(n14483)
         );
  OR2_X1 U9966 ( .A1(n14527), .A2(n14483), .ZN(n7699) );
  OR2_X1 U9967 ( .A1(n11467), .A2(n13039), .ZN(n11422) );
  AND2_X1 U9968 ( .A1(n11422), .A2(n7696), .ZN(n7697) );
  OR2_X1 U9969 ( .A1(n7698), .A2(n7697), .ZN(n11470) );
  AND2_X1 U9970 ( .A1(n7699), .A2(n11470), .ZN(n7700) );
  INV_X1 U9971 ( .A(n7702), .ZN(n7703) );
  MUX2_X1 U9972 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9139), .Z(n7721) );
  XNOR2_X1 U9973 ( .A(n7721), .B(SI_14_), .ZN(n7707) );
  XNOR2_X1 U9974 ( .A(n7722), .B(n7707), .ZN(n11523) );
  NAND2_X1 U9975 ( .A1(n11523), .A2(n7612), .ZN(n7711) );
  NAND2_X1 U9976 ( .A1(n7708), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7709) );
  XNOR2_X1 U9977 ( .A(n7709), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U9978 ( .A1(n7808), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7807), .B2(
        n13093), .ZN(n7710) );
  NAND2_X1 U9979 ( .A1(n7712), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7734) );
  INV_X1 U9980 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10281) );
  NAND2_X1 U9981 ( .A1(n7713), .A2(n10281), .ZN(n7714) );
  NAND2_X1 U9982 ( .A1(n7734), .A2(n7714), .ZN(n14500) );
  OR2_X1 U9983 ( .A1(n8029), .A2(n14500), .ZN(n7718) );
  NAND2_X1 U9984 ( .A1(n8080), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U9985 ( .A1(n7506), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U9986 ( .A1(n9148), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7715) );
  NAND4_X1 U9987 ( .A1(n7718), .A2(n7717), .A3(n7716), .A4(n7715), .ZN(n13037)
         );
  AND2_X1 U9988 ( .A1(n14503), .A2(n13037), .ZN(n7720) );
  OR2_X1 U9989 ( .A1(n14503), .A2(n13037), .ZN(n7719) );
  MUX2_X1 U9990 ( .A(n10176), .B(n10178), .S(n9139), .Z(n7724) );
  INV_X1 U9991 ( .A(SI_15_), .ZN(n7723) );
  INV_X1 U9992 ( .A(n7724), .ZN(n7725) );
  NAND2_X1 U9993 ( .A1(n7725), .A2(SI_15_), .ZN(n7726) );
  XNOR2_X1 U9994 ( .A(n7743), .B(n7742), .ZN(n11581) );
  NAND2_X1 U9995 ( .A1(n11581), .A2(n7612), .ZN(n7731) );
  OR2_X1 U9996 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7727) );
  OR2_X1 U9997 ( .A1(n7749), .A2(n13444), .ZN(n7729) );
  XNOR2_X1 U9998 ( .A(n7729), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U9999 ( .A1(n7808), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7807), .B2(
        n13096), .ZN(n7730) );
  INV_X1 U10000 ( .A(n7734), .ZN(n7732) );
  INV_X1 U10001 ( .A(n7753), .ZN(n7755) );
  INV_X1 U10002 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U10003 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  NAND2_X1 U10004 ( .A1(n7755), .A2(n7735), .ZN(n11764) );
  OR2_X1 U10005 ( .A1(n8029), .A2(n11764), .ZN(n7739) );
  NAND2_X1 U10006 ( .A1(n7506), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10007 ( .A1(n8080), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10008 ( .A1(n9148), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7736) );
  NAND4_X1 U10009 ( .A1(n7739), .A2(n7738), .A3(n7737), .A4(n7736), .ZN(n14482) );
  INV_X1 U10010 ( .A(n14482), .ZN(n7997) );
  XNOR2_X1 U10011 ( .A(n11767), .B(n7997), .ZN(n9237) );
  OR2_X1 U10012 ( .A1(n11767), .A2(n14482), .ZN(n7740) );
  MUX2_X1 U10013 ( .A(n10436), .B(n10459), .S(n9139), .Z(n7745) );
  INV_X1 U10014 ( .A(SI_16_), .ZN(n7744) );
  NAND2_X1 U10015 ( .A1(n7745), .A2(n7744), .ZN(n7766) );
  INV_X1 U10016 ( .A(n7745), .ZN(n7746) );
  NAND2_X1 U10017 ( .A1(n7746), .A2(SI_16_), .ZN(n7747) );
  XNOR2_X1 U10018 ( .A(n7765), .B(n7764), .ZN(n11695) );
  NAND2_X1 U10019 ( .A1(n11695), .A2(n7612), .ZN(n7752) );
  OR2_X1 U10020 ( .A1(n7769), .A2(n13444), .ZN(n7750) );
  XNOR2_X1 U10021 ( .A(n7750), .B(n7768), .ZN(n14936) );
  INV_X1 U10022 ( .A(n14936), .ZN(n13084) );
  AOI22_X1 U10023 ( .A1(n7808), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7807), 
        .B2(n13084), .ZN(n7751) );
  NAND2_X1 U10024 ( .A1(n7753), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7774) );
  INV_X1 U10025 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7754) );
  NAND2_X1 U10026 ( .A1(n7755), .A2(n7754), .ZN(n7756) );
  NAND2_X1 U10027 ( .A1(n7774), .A2(n7756), .ZN(n12948) );
  OR2_X1 U10028 ( .A1(n8029), .A2(n12948), .ZN(n7760) );
  NAND2_X1 U10029 ( .A1(n7506), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U10030 ( .A1(n8080), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U10031 ( .A1(n9148), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7757) );
  NAND4_X1 U10032 ( .A1(n7760), .A2(n7759), .A3(n7758), .A4(n7757), .ZN(n13036) );
  XNOR2_X1 U10033 ( .A(n13399), .B(n13036), .ZN(n11691) );
  NAND2_X1 U10034 ( .A1(n13399), .A2(n13036), .ZN(n7763) );
  MUX2_X1 U10035 ( .A(n10496), .B(n10472), .S(n9139), .Z(n7781) );
  XNOR2_X1 U10036 ( .A(n7781), .B(SI_17_), .ZN(n7780) );
  NAND2_X1 U10037 ( .A1(n11816), .A2(n7612), .ZN(n7772) );
  OR2_X1 U10038 ( .A1(n7787), .A2(n13444), .ZN(n7770) );
  XNOR2_X1 U10039 ( .A(n7770), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13110) );
  AOI22_X1 U10040 ( .A1(n7808), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7807), 
        .B2(n13110), .ZN(n7771) );
  INV_X1 U10041 ( .A(n7774), .ZN(n7773) );
  NAND2_X1 U10042 ( .A1(n7773), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7792) );
  INV_X1 U10043 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12960) );
  NAND2_X1 U10044 ( .A1(n7774), .A2(n12960), .ZN(n7775) );
  NAND2_X1 U10045 ( .A1(n7792), .A2(n7775), .ZN(n12959) );
  OR2_X1 U10046 ( .A1(n8029), .A2(n12959), .ZN(n7779) );
  NAND2_X1 U10047 ( .A1(n7506), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U10048 ( .A1(n8080), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7777) );
  NAND2_X1 U10049 ( .A1(n9148), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7776) );
  NAND4_X1 U10050 ( .A1(n7779), .A2(n7778), .A3(n7777), .A4(n7776), .ZN(n13035) );
  NAND2_X1 U10051 ( .A1(n13439), .A2(n13035), .ZN(n9220) );
  OR2_X1 U10052 ( .A1(n13439), .A2(n13035), .ZN(n9221) );
  INV_X1 U10053 ( .A(n7780), .ZN(n7784) );
  INV_X1 U10054 ( .A(n7781), .ZN(n7782) );
  NAND2_X1 U10055 ( .A1(n7782), .A2(SI_17_), .ZN(n7783) );
  MUX2_X1 U10056 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9139), .Z(n7821) );
  XNOR2_X1 U10057 ( .A(n7799), .B(n7821), .ZN(n11826) );
  NAND2_X1 U10058 ( .A1(n11826), .A2(n7612), .ZN(n7790) );
  INV_X1 U10059 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U10060 ( .A1(n7805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7788) );
  XNOR2_X1 U10061 ( .A(n7788), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U10062 ( .A1(n7808), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7807), 
        .B2(n13124), .ZN(n7789) );
  INV_X1 U10063 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U10064 ( .A1(n7792), .A2(n7791), .ZN(n7793) );
  NAND2_X1 U10065 ( .A1(n7834), .A2(n7793), .ZN(n13296) );
  OR2_X1 U10066 ( .A1(n8029), .A2(n13296), .ZN(n7797) );
  NAND2_X1 U10067 ( .A1(n7506), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U10068 ( .A1(n8080), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U10069 ( .A1(n9148), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7794) );
  NAND4_X1 U10070 ( .A1(n7797), .A2(n7796), .A3(n7795), .A4(n7794), .ZN(n13034) );
  XNOR2_X1 U10071 ( .A(n13435), .B(n13034), .ZN(n9238) );
  NAND2_X1 U10072 ( .A1(n13290), .A2(n13289), .ZN(n13288) );
  OR2_X1 U10073 ( .A1(n13435), .A2(n13034), .ZN(n7798) );
  NAND2_X1 U10074 ( .A1(n13288), .A2(n7798), .ZN(n13273) );
  INV_X1 U10075 ( .A(n7799), .ZN(n7800) );
  NAND2_X1 U10076 ( .A1(n7800), .A2(n7821), .ZN(n7802) );
  NAND2_X1 U10077 ( .A1(n7820), .A2(SI_18_), .ZN(n7801) );
  NAND2_X1 U10078 ( .A1(n7802), .A2(n7801), .ZN(n7804) );
  MUX2_X1 U10079 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9139), .Z(n7824) );
  XNOR2_X1 U10080 ( .A(n7824), .B(SI_19_), .ZN(n7803) );
  XNOR2_X1 U10081 ( .A(n7806), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7964) );
  AOI22_X1 U10082 ( .A1(n7808), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6463), 
        .B2(n7807), .ZN(n7809) );
  NAND2_X2 U10083 ( .A1(n7810), .A2(n7809), .ZN(n13277) );
  NAND2_X1 U10084 ( .A1(n7506), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U10085 ( .A1(n8080), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7813) );
  XNOR2_X1 U10086 ( .A(n7834), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U10087 ( .A1(n7486), .A2(n13274), .ZN(n7812) );
  NAND2_X1 U10088 ( .A1(n9148), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7811) );
  NAND4_X1 U10089 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n13033) );
  NAND2_X1 U10090 ( .A1(n13277), .A2(n13033), .ZN(n7815) );
  OR2_X1 U10091 ( .A1(n13277), .A2(n13033), .ZN(n7816) );
  INV_X1 U10092 ( .A(n7824), .ZN(n7817) );
  INV_X1 U10093 ( .A(SI_19_), .ZN(n10073) );
  NAND2_X1 U10094 ( .A1(n7817), .A2(n10073), .ZN(n7825) );
  OAI21_X1 U10095 ( .B1(SI_18_), .B2(n7821), .A(n7825), .ZN(n7818) );
  INV_X1 U10096 ( .A(n7818), .ZN(n7819) );
  INV_X1 U10097 ( .A(n7821), .ZN(n7823) );
  INV_X1 U10098 ( .A(SI_18_), .ZN(n7822) );
  NOR2_X1 U10099 ( .A1(n7823), .A2(n7822), .ZN(n7826) );
  AOI22_X1 U10100 ( .A1(n7826), .A2(n7825), .B1(n7824), .B2(SI_19_), .ZN(n7827) );
  MUX2_X1 U10101 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9139), .Z(n7841) );
  XNOR2_X1 U10102 ( .A(n7840), .B(n7841), .ZN(n11861) );
  NAND2_X1 U10103 ( .A1(n11861), .A2(n7612), .ZN(n7829) );
  INV_X1 U10104 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11037) );
  OR2_X1 U10105 ( .A1(n7919), .A2(n11037), .ZN(n7828) );
  INV_X1 U10106 ( .A(n7834), .ZN(n7831) );
  AND2_X1 U10107 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n7830) );
  NAND2_X1 U10108 ( .A1(n7831), .A2(n7830), .ZN(n7846) );
  INV_X1 U10109 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7833) );
  INV_X1 U10110 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7832) );
  OAI21_X1 U10111 ( .B1(n7834), .B2(n7833), .A(n7832), .ZN(n7835) );
  NAND2_X1 U10112 ( .A1(n7846), .A2(n7835), .ZN(n13263) );
  OR2_X1 U10113 ( .A1(n8029), .A2(n13263), .ZN(n7839) );
  NAND2_X1 U10114 ( .A1(n8080), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10115 ( .A1(n7506), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10116 ( .A1(n9148), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7836) );
  NAND4_X1 U10117 ( .A1(n7839), .A2(n7838), .A3(n7837), .A4(n7836), .ZN(n13032) );
  NAND2_X1 U10118 ( .A1(n7842), .A2(SI_20_), .ZN(n7843) );
  MUX2_X1 U10119 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9139), .Z(n7854) );
  XNOR2_X1 U10120 ( .A(n7854), .B(SI_21_), .ZN(n7852) );
  NAND2_X1 U10121 ( .A1(n11880), .A2(n7612), .ZN(n7845) );
  INV_X1 U10122 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11189) );
  OR2_X1 U10123 ( .A1(n7919), .A2(n11189), .ZN(n7844) );
  INV_X1 U10124 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12931) );
  NAND2_X1 U10125 ( .A1(n7846), .A2(n12931), .ZN(n7847) );
  NAND2_X1 U10126 ( .A1(n7870), .A2(n7847), .ZN(n13249) );
  OR2_X1 U10127 ( .A1(n8029), .A2(n13249), .ZN(n7851) );
  NAND2_X1 U10128 ( .A1(n8080), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U10129 ( .A1(n9148), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U10130 ( .A1(n8081), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7848) );
  NAND4_X1 U10131 ( .A1(n7851), .A2(n7850), .A3(n7849), .A4(n7848), .ZN(n13031) );
  INV_X1 U10132 ( .A(n13031), .ZN(n8011) );
  XNOR2_X1 U10133 ( .A(n13425), .B(n8011), .ZN(n13255) );
  NAND2_X1 U10134 ( .A1(n7854), .A2(SI_21_), .ZN(n7855) );
  NAND2_X1 U10135 ( .A1(n7856), .A2(n7855), .ZN(n7865) );
  MUX2_X1 U10136 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9139), .Z(n7864) );
  XNOR2_X1 U10137 ( .A(n11893), .B(n7864), .ZN(n11368) );
  NAND2_X1 U10138 ( .A1(n11368), .A2(n7612), .ZN(n7858) );
  INV_X1 U10139 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11371) );
  OR2_X1 U10140 ( .A1(n7919), .A2(n11371), .ZN(n7857) );
  NAND2_X2 U10141 ( .A1(n7858), .A2(n7857), .ZN(n13421) );
  NAND2_X1 U10142 ( .A1(n7506), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U10143 ( .A1(n8080), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7861) );
  XNOR2_X1 U10144 ( .A(n7870), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U10145 ( .A1(n7486), .A2(n13236), .ZN(n7860) );
  NAND2_X1 U10146 ( .A1(n9148), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7859) );
  NAND4_X1 U10147 ( .A1(n7862), .A2(n7861), .A3(n7860), .A4(n7859), .ZN(n13030) );
  INV_X1 U10148 ( .A(n13030), .ZN(n12901) );
  XNOR2_X1 U10149 ( .A(n13421), .B(n12901), .ZN(n13228) );
  INV_X1 U10150 ( .A(n13228), .ZN(n13232) );
  NAND2_X1 U10151 ( .A1(n13421), .A2(n13030), .ZN(n7863) );
  MUX2_X1 U10152 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9139), .Z(n7882) );
  XNOR2_X1 U10153 ( .A(n7882), .B(SI_23_), .ZN(n7879) );
  XNOR2_X1 U10154 ( .A(n7881), .B(n7879), .ZN(n11911) );
  NAND2_X1 U10155 ( .A1(n11911), .A2(n7612), .ZN(n7868) );
  INV_X1 U10156 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11420) );
  OR2_X1 U10157 ( .A1(n7919), .A2(n11420), .ZN(n7867) );
  INV_X1 U10158 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12996) );
  INV_X1 U10159 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7869) );
  OAI21_X1 U10160 ( .B1(n7870), .B2(n12996), .A(n7869), .ZN(n7873) );
  INV_X1 U10161 ( .A(n7870), .ZN(n7872) );
  AND2_X1 U10162 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n7871) );
  NAND2_X1 U10163 ( .A1(n7872), .A2(n7871), .ZN(n7888) );
  NAND2_X1 U10164 ( .A1(n7873), .A2(n7888), .ZN(n13222) );
  OR2_X1 U10165 ( .A1(n8029), .A2(n13222), .ZN(n7877) );
  NAND2_X1 U10166 ( .A1(n7506), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10167 ( .A1(n8080), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10168 ( .A1(n9148), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7874) );
  NAND4_X1 U10169 ( .A1(n7877), .A2(n7876), .A3(n7875), .A4(n7874), .ZN(n13029) );
  NAND2_X1 U10170 ( .A1(n13345), .A2(n13029), .ZN(n7878) );
  INV_X1 U10171 ( .A(n7879), .ZN(n7880) );
  NAND2_X1 U10172 ( .A1(n7881), .A2(n7880), .ZN(n7884) );
  NAND2_X1 U10173 ( .A1(n7882), .A2(SI_23_), .ZN(n7883) );
  INV_X1 U10174 ( .A(SI_24_), .ZN(n12181) );
  INV_X1 U10175 ( .A(n7896), .ZN(n7885) );
  MUX2_X1 U10176 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9139), .Z(n7895) );
  INV_X1 U10177 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13468) );
  OR2_X1 U10178 ( .A1(n7919), .A2(n13468), .ZN(n7886) );
  INV_X1 U10179 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12972) );
  NAND2_X1 U10180 ( .A1(n7888), .A2(n12972), .ZN(n7889) );
  NAND2_X1 U10181 ( .A1(n7924), .A2(n7889), .ZN(n13200) );
  OR2_X1 U10182 ( .A1(n13200), .A2(n8029), .ZN(n7893) );
  NAND2_X1 U10183 ( .A1(n8080), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U10184 ( .A1(n9148), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U10185 ( .A1(n7506), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7890) );
  NAND4_X1 U10186 ( .A1(n7893), .A2(n7892), .A3(n7891), .A4(n7890), .ZN(n13028) );
  XNOR2_X1 U10187 ( .A(n13339), .B(n13028), .ZN(n13197) );
  INV_X1 U10188 ( .A(n13197), .ZN(n13208) );
  NAND2_X1 U10189 ( .A1(n13209), .A2(n13208), .ZN(n13207) );
  NAND2_X1 U10190 ( .A1(n6644), .A2(n13028), .ZN(n7894) );
  INV_X1 U10191 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14283) );
  INV_X1 U10192 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13464) );
  MUX2_X1 U10193 ( .A(n14283), .B(n13464), .S(n9139), .Z(n7900) );
  INV_X1 U10194 ( .A(SI_25_), .ZN(n12254) );
  NAND2_X1 U10195 ( .A1(n7900), .A2(n12254), .ZN(n7913) );
  INV_X1 U10196 ( .A(n7900), .ZN(n7901) );
  NAND2_X1 U10197 ( .A1(n7901), .A2(SI_25_), .ZN(n7902) );
  NAND2_X1 U10198 ( .A1(n7913), .A2(n7902), .ZN(n7914) );
  OR2_X1 U10199 ( .A1(n7919), .A2(n13464), .ZN(n7903) );
  NAND2_X2 U10200 ( .A1(n7904), .A2(n7903), .ZN(n13193) );
  INV_X1 U10201 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U10202 ( .A1(n7506), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U10203 ( .A1(n8080), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n7905) );
  AND2_X1 U10204 ( .A1(n7906), .A2(n7905), .ZN(n7908) );
  XNOR2_X1 U10205 ( .A(n7924), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n13190) );
  NAND2_X1 U10206 ( .A1(n13190), .A2(n7486), .ZN(n7907) );
  OAI211_X1 U10207 ( .C1(n7487), .C2(n7909), .A(n7908), .B(n7907), .ZN(n13027)
         );
  OR2_X1 U10208 ( .A1(n13193), .A2(n13027), .ZN(n7910) );
  NAND2_X1 U10209 ( .A1(n13193), .A2(n13027), .ZN(n7911) );
  INV_X1 U10210 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14278) );
  INV_X1 U10211 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13459) );
  MUX2_X1 U10212 ( .A(n14278), .B(n13459), .S(n9139), .Z(n7916) );
  INV_X1 U10213 ( .A(SI_26_), .ZN(n11323) );
  NAND2_X1 U10214 ( .A1(n7916), .A2(n11323), .ZN(n7932) );
  INV_X1 U10215 ( .A(n7916), .ZN(n7917) );
  NAND2_X1 U10216 ( .A1(n7917), .A2(SI_26_), .ZN(n7918) );
  OR2_X1 U10217 ( .A1(n7919), .A2(n13459), .ZN(n7920) );
  INV_X1 U10218 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12940) );
  INV_X1 U10219 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7922) );
  OAI21_X1 U10220 ( .B1(n7924), .B2(n12940), .A(n7922), .ZN(n7925) );
  NAND2_X1 U10221 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n7923) );
  NOR2_X1 U10222 ( .A1(n7924), .A2(n7923), .ZN(n7935) );
  INV_X1 U10223 ( .A(n7935), .ZN(n7936) );
  NAND2_X1 U10224 ( .A1(n7925), .A2(n7936), .ZN(n13015) );
  AOI22_X1 U10225 ( .A1(n8080), .A2(P2_REG1_REG_26__SCAN_IN), .B1(n9148), .B2(
        P2_REG0_REG_26__SCAN_IN), .ZN(n7927) );
  NAND2_X1 U10226 ( .A1(n7506), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7926) );
  OAI211_X1 U10227 ( .C1(n13015), .C2(n8029), .A(n7927), .B(n7926), .ZN(n13026) );
  AND2_X1 U10228 ( .A1(n13176), .A2(n13026), .ZN(n7929) );
  OR2_X1 U10229 ( .A1(n13176), .A2(n13026), .ZN(n7928) );
  INV_X1 U10230 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11774) );
  INV_X1 U10231 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13454) );
  MUX2_X1 U10232 ( .A(n11774), .B(n13454), .S(n9139), .Z(n7942) );
  XNOR2_X1 U10233 ( .A(n7942), .B(SI_27_), .ZN(n7941) );
  OR2_X1 U10234 ( .A1(n7919), .A2(n13454), .ZN(n7933) );
  NAND2_X1 U10235 ( .A1(n7935), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7953) );
  INV_X1 U10236 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U10237 ( .A1(n7936), .A2(n12892), .ZN(n7937) );
  NAND2_X1 U10238 ( .A1(n7953), .A2(n7937), .ZN(n13164) );
  AOI22_X1 U10239 ( .A1(n8080), .A2(P2_REG1_REG_27__SCAN_IN), .B1(n7506), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10240 ( .A1(n9148), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7938) );
  OAI211_X1 U10241 ( .C1(n13164), .C2(n8029), .A(n7939), .B(n7938), .ZN(n13025) );
  INV_X1 U10242 ( .A(n13025), .ZN(n8022) );
  NAND2_X1 U10243 ( .A1(n13320), .A2(n13025), .ZN(n7940) );
  NAND2_X1 U10244 ( .A1(n13317), .A2(n7940), .ZN(n7959) );
  INV_X1 U10245 ( .A(n7941), .ZN(n7945) );
  INV_X1 U10246 ( .A(n7942), .ZN(n7943) );
  NAND2_X1 U10247 ( .A1(n7943), .A2(SI_27_), .ZN(n7944) );
  OAI21_X2 U10248 ( .B1(n7946), .B2(n7945), .A(n7944), .ZN(n8076) );
  INV_X1 U10249 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11773) );
  INV_X1 U10250 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8600) );
  MUX2_X1 U10251 ( .A(n11773), .B(n8600), .S(n9139), .Z(n7947) );
  INV_X1 U10252 ( .A(SI_28_), .ZN(n12830) );
  NAND2_X1 U10253 ( .A1(n7947), .A2(n12830), .ZN(n8074) );
  INV_X1 U10254 ( .A(n7947), .ZN(n7948) );
  NAND2_X1 U10255 ( .A1(n7948), .A2(SI_28_), .ZN(n7949) );
  NAND2_X1 U10256 ( .A1(n8074), .A2(n7949), .ZN(n8075) );
  NAND2_X1 U10257 ( .A1(n12021), .A2(n7612), .ZN(n7951) );
  OR2_X1 U10258 ( .A1(n7919), .A2(n8600), .ZN(n7950) );
  INV_X1 U10259 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7957) );
  INV_X1 U10260 ( .A(n7953), .ZN(n7952) );
  NAND2_X1 U10261 ( .A1(n7952), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8093) );
  INV_X1 U10262 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U10263 ( .A1(n7953), .A2(n12920), .ZN(n7954) );
  NAND2_X1 U10264 ( .A1(n8093), .A2(n7954), .ZN(n13149) );
  OR2_X1 U10265 ( .A1(n13149), .A2(n8029), .ZN(n7956) );
  AOI22_X1 U10266 ( .A1(n8080), .A2(P2_REG1_REG_28__SCAN_IN), .B1(n7506), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n7955) );
  OAI211_X1 U10267 ( .C1(n7487), .C2(n7957), .A(n7956), .B(n7955), .ZN(n13024)
         );
  NAND2_X1 U10268 ( .A1(n12924), .A2(n13024), .ZN(n8100) );
  OR2_X1 U10269 ( .A1(n12924), .A2(n13024), .ZN(n7958) );
  NAND2_X1 U10270 ( .A1(n7959), .A2(n9243), .ZN(n8101) );
  OR2_X1 U10271 ( .A1(n7959), .A2(n9243), .ZN(n7960) );
  NAND2_X1 U10272 ( .A1(n8101), .A2(n7960), .ZN(n13157) );
  NAND2_X1 U10273 ( .A1(n7961), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7963) );
  INV_X1 U10274 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7962) );
  XNOR2_X1 U10275 ( .A(n7963), .B(n7962), .ZN(n11035) );
  NAND2_X1 U10276 ( .A1(n7964), .A2(n11035), .ZN(n8054) );
  INV_X1 U10277 ( .A(n8054), .ZN(n7968) );
  NAND2_X1 U10278 ( .A1(n6899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7966) );
  MUX2_X1 U10279 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7966), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n7967) );
  NAND2_X1 U10280 ( .A1(n7967), .A2(n6485), .ZN(n11369) );
  INV_X1 U10281 ( .A(n11369), .ZN(n9253) );
  MUX2_X1 U10282 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7969), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n7970) );
  NAND2_X1 U10283 ( .A1(n7970), .A2(n6899), .ZN(n11187) );
  INV_X1 U10284 ( .A(n11187), .ZN(n9249) );
  NAND2_X1 U10285 ( .A1(n9249), .A2(n11035), .ZN(n10120) );
  XNOR2_X1 U10286 ( .A(n10120), .B(n11369), .ZN(n7971) );
  NAND2_X1 U10287 ( .A1(n13045), .A2(n10839), .ZN(n7982) );
  NAND2_X1 U10288 ( .A1(n10162), .A2(n10161), .ZN(n7973) );
  OR2_X1 U10289 ( .A1(n13048), .A2(n10374), .ZN(n7972) );
  NAND2_X1 U10290 ( .A1(n7973), .A2(n7972), .ZN(n10208) );
  NAND2_X1 U10291 ( .A1(n10208), .A2(n9224), .ZN(n10408) );
  INV_X1 U10292 ( .A(n10321), .ZN(n10450) );
  OR2_X1 U10293 ( .A1(n8973), .A2(n10450), .ZN(n10407) );
  NAND2_X1 U10294 ( .A1(n7974), .A2(n14939), .ZN(n7976) );
  AND2_X1 U10295 ( .A1(n7976), .A2(n10407), .ZN(n7975) );
  NAND2_X1 U10296 ( .A1(n10408), .A2(n7975), .ZN(n7979) );
  INV_X1 U10297 ( .A(n7976), .ZN(n7977) );
  AND2_X1 U10298 ( .A1(n7979), .A2(n7978), .ZN(n10501) );
  INV_X1 U10299 ( .A(n10503), .ZN(n7981) );
  NOR2_X1 U10300 ( .A1(n13045), .A2(n10839), .ZN(n7980) );
  NAND2_X1 U10301 ( .A1(n7983), .A2(n7982), .ZN(n10646) );
  INV_X1 U10302 ( .A(n10855), .ZN(n14965) );
  OR2_X1 U10303 ( .A1(n13044), .A2(n14965), .ZN(n7985) );
  NAND2_X1 U10304 ( .A1(n13043), .A2(n10927), .ZN(n7986) );
  NOR2_X1 U10305 ( .A1(n11316), .A2(n7987), .ZN(n7988) );
  INV_X1 U10306 ( .A(n11316), .ZN(n11319) );
  XNOR2_X1 U10307 ( .A(n11467), .B(n13039), .ZN(n11241) );
  INV_X1 U10308 ( .A(n13039), .ZN(n7990) );
  NAND2_X1 U10309 ( .A1(n11467), .A2(n7990), .ZN(n7991) );
  INV_X1 U10310 ( .A(n13038), .ZN(n7992) );
  OR2_X1 U10311 ( .A1(n11565), .A2(n7992), .ZN(n7993) );
  INV_X1 U10312 ( .A(n14483), .ZN(n7994) );
  NAND2_X1 U10313 ( .A1(n14527), .A2(n7994), .ZN(n9232) );
  OR2_X1 U10314 ( .A1(n14527), .A2(n7994), .ZN(n9233) );
  INV_X1 U10315 ( .A(n13037), .ZN(n7996) );
  XNOR2_X1 U10316 ( .A(n14503), .B(n7996), .ZN(n14505) );
  INV_X1 U10317 ( .A(n13036), .ZN(n7998) );
  OR2_X1 U10318 ( .A1(n13399), .A2(n7998), .ZN(n7999) );
  INV_X1 U10319 ( .A(n13035), .ZN(n8001) );
  NAND2_X1 U10320 ( .A1(n13439), .A2(n8001), .ZN(n8000) );
  OR2_X1 U10321 ( .A1(n13439), .A2(n8001), .ZN(n8002) );
  NAND2_X1 U10322 ( .A1(n8003), .A2(n8002), .ZN(n13287) );
  INV_X1 U10323 ( .A(n13034), .ZN(n12835) );
  NAND2_X1 U10324 ( .A1(n13435), .A2(n12835), .ZN(n8004) );
  NAND2_X1 U10325 ( .A1(n13287), .A2(n8004), .ZN(n8006) );
  OR2_X1 U10326 ( .A1(n13435), .A2(n12835), .ZN(n8005) );
  INV_X1 U10327 ( .A(n13033), .ZN(n8008) );
  NAND2_X1 U10328 ( .A1(n13277), .A2(n8008), .ZN(n8007) );
  INV_X1 U10329 ( .A(n13032), .ZN(n9219) );
  NOR2_X1 U10330 ( .A1(n13367), .A2(n9219), .ZN(n8010) );
  NAND2_X1 U10331 ( .A1(n13425), .A2(n8011), .ZN(n8012) );
  XNOR2_X1 U10332 ( .A(n13345), .B(n13029), .ZN(n13223) );
  INV_X1 U10333 ( .A(n13029), .ZN(n8013) );
  NAND2_X1 U10334 ( .A1(n13345), .A2(n8013), .ZN(n8014) );
  INV_X1 U10335 ( .A(n13028), .ZN(n12899) );
  NAND2_X1 U10336 ( .A1(n13339), .A2(n12899), .ZN(n8015) );
  NAND2_X1 U10337 ( .A1(n13187), .A2(n13186), .ZN(n8019) );
  INV_X1 U10338 ( .A(n13027), .ZN(n8017) );
  NAND2_X1 U10339 ( .A1(n13193), .A2(n8017), .ZN(n8018) );
  INV_X1 U10340 ( .A(n13026), .ZN(n12890) );
  XNOR2_X1 U10341 ( .A(n13176), .B(n12890), .ZN(n13173) );
  INV_X1 U10342 ( .A(n13173), .ZN(n13181) );
  NAND2_X1 U10343 ( .A1(n13182), .A2(n13181), .ZN(n8021) );
  NAND2_X1 U10344 ( .A1(n13176), .A2(n12890), .ZN(n8020) );
  AND2_X1 U10345 ( .A1(n13320), .A2(n8022), .ZN(n8023) );
  NAND2_X1 U10346 ( .A1(n6463), .A2(n9253), .ZN(n8024) );
  INV_X1 U10347 ( .A(n11035), .ZN(n9223) );
  NAND2_X1 U10348 ( .A1(n9249), .A2(n9223), .ZN(n9212) );
  NAND2_X1 U10349 ( .A1(n8024), .A2(n9212), .ZN(n14535) );
  INV_X1 U10350 ( .A(n8027), .ZN(n8028) );
  NOR2_X1 U10351 ( .A1(n11369), .A2(n11187), .ZN(n9894) );
  NAND2_X1 U10352 ( .A1(n8028), .A2(n9894), .ZN(n12900) );
  INV_X2 U10353 ( .A(n12900), .ZN(n14484) );
  NAND2_X1 U10354 ( .A1(n13025), .A2(n14484), .ZN(n8034) );
  INV_X1 U10355 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8032) );
  OR2_X1 U10356 ( .A1(n8093), .A2(n8029), .ZN(n8031) );
  AOI22_X1 U10357 ( .A1(n8080), .A2(P2_REG1_REG_29__SCAN_IN), .B1(n7506), .B2(
        P2_REG2_REG_29__SCAN_IN), .ZN(n8030) );
  OAI211_X1 U10358 ( .C1(n7487), .C2(n8032), .A(n8031), .B(n8030), .ZN(n13023)
         );
  AND2_X1 U10359 ( .A1(n8027), .A2(n9894), .ZN(n14481) );
  INV_X1 U10360 ( .A(n14481), .ZN(n12898) );
  INV_X1 U10361 ( .A(n12898), .ZN(n13013) );
  NAND2_X1 U10362 ( .A1(n13023), .A2(n13013), .ZN(n8033) );
  AND2_X1 U10363 ( .A1(n8034), .A2(n8033), .ZN(n12921) );
  INV_X1 U10364 ( .A(n13421), .ZN(n13235) );
  NOR2_X1 U10365 ( .A1(n10121), .A2(n10165), .ZN(n8035) );
  NAND2_X1 U10366 ( .A1(n10405), .A2(n10417), .ZN(n10667) );
  INV_X1 U10367 ( .A(n11308), .ZN(n14977) );
  INV_X1 U10368 ( .A(n11467), .ZN(n14987) );
  INV_X1 U10369 ( .A(n11767), .ZN(n14516) );
  NAND2_X1 U10370 ( .A1(n14506), .A2(n14516), .ZN(n11686) );
  INV_X1 U10371 ( .A(n13435), .ZN(n13291) );
  NAND2_X1 U10372 ( .A1(n11369), .A2(n11187), .ZN(n8055) );
  NAND2_X1 U10373 ( .A1(n10108), .A2(n11035), .ZN(n12834) );
  OAI211_X1 U10374 ( .C1(n13413), .C2(n13163), .A(n6452), .B(n8092), .ZN(
        n13151) );
  NAND2_X1 U10375 ( .A1(n8042), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8038) );
  MUX2_X1 U10376 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8038), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8039) );
  INV_X1 U10377 ( .A(n13460), .ZN(n8047) );
  NAND2_X1 U10378 ( .A1(n8040), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8041) );
  MUX2_X1 U10379 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8041), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8043) );
  NAND2_X1 U10380 ( .A1(n8043), .A2(n8042), .ZN(n13463) );
  NAND2_X1 U10381 ( .A1(n6597), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8044) );
  MUX2_X1 U10382 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8044), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8045) );
  NAND2_X1 U10383 ( .A1(n8045), .A2(n8040), .ZN(n13466) );
  NOR2_X1 U10384 ( .A1(n13463), .A2(n13466), .ZN(n8046) );
  NAND2_X1 U10385 ( .A1(n8047), .A2(n8046), .ZN(n9375) );
  NAND2_X1 U10386 ( .A1(n6485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8049) );
  XNOR2_X1 U10387 ( .A(n8049), .B(n8048), .ZN(n9801) );
  NAND2_X1 U10388 ( .A1(n9375), .A2(n9801), .ZN(n9886) );
  XNOR2_X1 U10389 ( .A(n13466), .B(P2_B_REG_SCAN_IN), .ZN(n8050) );
  AND2_X1 U10390 ( .A1(n8050), .A2(n13463), .ZN(n8051) );
  INV_X1 U10391 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14962) );
  NAND2_X1 U10392 ( .A1(n14952), .A2(n14962), .ZN(n8053) );
  NAND2_X1 U10393 ( .A1(n13460), .A2(n13463), .ZN(n8052) );
  NAND2_X1 U10394 ( .A1(n8053), .A2(n8052), .ZN(n8089) );
  AND2_X1 U10395 ( .A1(n14959), .A2(n8089), .ZN(n14960) );
  NAND2_X1 U10396 ( .A1(n10984), .A2(n11035), .ZN(n9897) );
  NAND2_X1 U10397 ( .A1(n9897), .A2(n9894), .ZN(n9888) );
  NOR4_X1 U10398 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8059) );
  NOR4_X1 U10399 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8058) );
  NOR4_X1 U10400 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8057) );
  NOR4_X1 U10401 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8056) );
  NAND4_X1 U10402 ( .A1(n8059), .A2(n8058), .A3(n8057), .A4(n8056), .ZN(n8065)
         );
  NOR2_X1 U10403 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .ZN(
        n8063) );
  NOR4_X1 U10404 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8062) );
  NOR4_X1 U10405 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n8061) );
  NOR4_X1 U10406 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8060) );
  NAND4_X1 U10407 ( .A1(n8063), .A2(n8062), .A3(n8061), .A4(n8060), .ZN(n8064)
         );
  OAI21_X1 U10408 ( .B1(n8065), .B2(n8064), .A(n14952), .ZN(n8088) );
  NAND4_X1 U10409 ( .A1(n14960), .A2(n9884), .A3(n9888), .A4(n8088), .ZN(
        n10104) );
  INV_X1 U10410 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14957) );
  NAND2_X1 U10411 ( .A1(n14952), .A2(n14957), .ZN(n8067) );
  NAND2_X1 U10412 ( .A1(n13460), .A2(n13466), .ZN(n8066) );
  NAND2_X1 U10413 ( .A1(n8067), .A2(n8066), .ZN(n14958) );
  INV_X2 U10414 ( .A(n14999), .ZN(n15002) );
  NAND2_X1 U10415 ( .A1(n15002), .A2(n13398), .ZN(n13378) );
  INV_X1 U10416 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8068) );
  NOR2_X1 U10417 ( .A1(n15002), .A2(n8068), .ZN(n8069) );
  INV_X1 U10418 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11771) );
  INV_X1 U10419 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13448) );
  MUX2_X1 U10420 ( .A(n11771), .B(n13448), .S(n9139), .Z(n9137) );
  XNOR2_X1 U10421 ( .A(n9137), .B(SI_29_), .ZN(n9135) );
  OR2_X1 U10422 ( .A1(n7919), .A2(n13448), .ZN(n8077) );
  NAND2_X1 U10423 ( .A1(n13024), .A2(n14484), .ZN(n8087) );
  NAND2_X1 U10424 ( .A1(n8080), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8084) );
  NAND2_X1 U10425 ( .A1(n7506), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8083) );
  NAND2_X1 U10426 ( .A1(n9148), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8082) );
  AND3_X1 U10427 ( .A1(n8084), .A2(n8083), .A3(n8082), .ZN(n9193) );
  INV_X1 U10428 ( .A(n9193), .ZN(n13022) );
  INV_X1 U10429 ( .A(n13455), .ZN(n9834) );
  NAND2_X1 U10430 ( .A1(n9834), .A2(P2_B_REG_SCAN_IN), .ZN(n8085) );
  AND2_X1 U10431 ( .A1(n14481), .A2(n8085), .ZN(n11987) );
  INV_X1 U10432 ( .A(n8088), .ZN(n8090) );
  OR2_X1 U10433 ( .A1(n8090), .A2(n8089), .ZN(n9885) );
  INV_X1 U10434 ( .A(n9885), .ZN(n9892) );
  NAND4_X1 U10435 ( .A1(n9892), .A2(n14959), .A3(n9888), .A4(n14958), .ZN(
        n8091) );
  INV_X1 U10436 ( .A(n14951), .ZN(n14948) );
  INV_X1 U10437 ( .A(n13313), .ZN(n8096) );
  NAND2_X1 U10438 ( .A1(n10108), .A2(n9223), .ZN(n9898) );
  INV_X1 U10439 ( .A(n9898), .ZN(n14940) );
  NAND2_X1 U10440 ( .A1(n13298), .A2(n14940), .ZN(n13205) );
  INV_X1 U10441 ( .A(n8093), .ZN(n8094) );
  INV_X1 U10442 ( .A(n13295), .ZN(n14941) );
  AOI22_X1 U10443 ( .A1(n8094), .A2(n14941), .B1(n14951), .B2(
        P2_REG2_REG_29__SCAN_IN), .ZN(n8095) );
  OAI21_X1 U10444 ( .B1(n8096), .B2(n13205), .A(n8095), .ZN(n8097) );
  OR2_X1 U10445 ( .A1(n8054), .A2(n11187), .ZN(n10437) );
  NAND2_X1 U10446 ( .A1(n10437), .A2(n11255), .ZN(n14947) );
  NAND2_X1 U10447 ( .A1(n13298), .A2(n14947), .ZN(n13224) );
  INV_X1 U10448 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8726) );
  NOR2_X1 U10449 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n8108) );
  INV_X2 U10450 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n12100) );
  NAND4_X1 U10451 ( .A1(n8108), .A2(n8107), .A3(n12100), .A4(n8440), .ZN(n8109) );
  NOR2_X1 U10452 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), 
        .ZN(n8114) );
  NOR2_X1 U10453 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), 
        .ZN(n8113) );
  INV_X1 U10454 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8112) );
  NAND4_X1 U10455 ( .A1(n8114), .A2(n8113), .A3(n12094), .A4(n8112), .ZN(n8115) );
  OR2_X2 U10456 ( .A1(n8129), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n12824) );
  NAND2_X2 U10457 ( .A1(n12824), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8117) );
  INV_X1 U10458 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8116) );
  XNOR2_X2 U10459 ( .A(n8117), .B(n8116), .ZN(n8121) );
  NAND2_X1 U10460 ( .A1(n8129), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8118) );
  MUX2_X1 U10461 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8118), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8119) );
  AND2_X2 U10462 ( .A1(n8121), .A2(n8120), .ZN(n8513) );
  NAND2_X1 U10463 ( .A1(n8513), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U10464 ( .A1(n8198), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8125) );
  INV_X1 U10465 ( .A(n8121), .ZN(n8122) );
  NAND2_X2 U10466 ( .A1(n8122), .A2(n12003), .ZN(n8182) );
  INV_X1 U10467 ( .A(n8182), .ZN(n8426) );
  NAND2_X1 U10468 ( .A1(n8426), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8124) );
  INV_X4 U10469 ( .A(n8163), .ZN(n8673) );
  NAND2_X1 U10470 ( .A1(n8673), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10471 ( .A1(n8132), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8128) );
  MUX2_X1 U10472 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8128), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8130) );
  NAND2_X1 U10473 ( .A1(n8130), .A2(n8129), .ZN(n12833) );
  INV_X1 U10474 ( .A(SI_0_), .ZN(n9581) );
  INV_X1 U10475 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9580) );
  NAND2_X1 U10476 ( .A1(n9580), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U10477 ( .A1(n8154), .A2(n8136), .ZN(n9494) );
  NAND2_X1 U10478 ( .A1(n8243), .A2(n9494), .ZN(n8138) );
  NAND2_X1 U10479 ( .A1(n8457), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10480 ( .A1(n8513), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U10481 ( .A1(n6447), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8142) );
  INV_X1 U10482 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8139) );
  OR2_X1 U10483 ( .A1(n8163), .A2(n8139), .ZN(n8141) );
  INV_X1 U10484 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9744) );
  OR2_X1 U10485 ( .A1(n8182), .A2(n9744), .ZN(n8140) );
  AND4_X2 U10486 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n9265)
         );
  XNOR2_X1 U10487 ( .A(n8155), .B(n8154), .ZN(n9468) );
  NAND2_X1 U10488 ( .A1(n8144), .A2(SI_1_), .ZN(n8147) );
  NAND2_X1 U10489 ( .A1(n8457), .A2(n9762), .ZN(n8146) );
  OAI211_X1 U10490 ( .C1(n6449), .C2(n9468), .A(n8147), .B(n8146), .ZN(n12769)
         );
  INV_X1 U10491 ( .A(n12769), .ZN(n10036) );
  NAND2_X1 U10492 ( .A1(n8148), .A2(n10036), .ZN(n8791) );
  NAND2_X1 U10493 ( .A1(n9262), .A2(n9267), .ZN(n10180) );
  NAND2_X1 U10494 ( .A1(n8513), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U10495 ( .A1(n6448), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8152) );
  INV_X1 U10496 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10194) );
  OR2_X1 U10497 ( .A1(n8182), .A2(n10194), .ZN(n8151) );
  INV_X1 U10498 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8149) );
  OR2_X1 U10499 ( .A1(n8163), .A2(n8149), .ZN(n8150) );
  NAND2_X1 U10500 ( .A1(n9478), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8156) );
  XNOR2_X1 U10501 ( .A(n8169), .B(n8171), .ZN(n9489) );
  NAND2_X1 U10502 ( .A1(n8144), .A2(SI_2_), .ZN(n8162) );
  NAND2_X1 U10503 ( .A1(n8457), .A2(n6450), .ZN(n8161) );
  NAND2_X1 U10504 ( .A1(n12760), .A2(n10183), .ZN(n8794) );
  NAND2_X1 U10505 ( .A1(n12383), .A2(n10078), .ZN(n8795) );
  INV_X1 U10506 ( .A(n10186), .ZN(n10179) );
  NAND2_X1 U10507 ( .A1(n10180), .A2(n10179), .ZN(n10182) );
  NAND2_X1 U10508 ( .A1(n10182), .A2(n8794), .ZN(n10083) );
  NAND2_X1 U10509 ( .A1(n8513), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10510 ( .A1(n8198), .A2(n10384), .ZN(n8167) );
  INV_X1 U10511 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8164) );
  OR2_X1 U10512 ( .A1(n8753), .A2(n8164), .ZN(n8166) );
  INV_X1 U10513 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9998) );
  OR2_X1 U10514 ( .A1(n8182), .A2(n9998), .ZN(n8165) );
  INV_X1 U10515 ( .A(SI_3_), .ZN(n9481) );
  NAND2_X1 U10516 ( .A1(n8144), .A2(n9481), .ZN(n8180) );
  NAND2_X1 U10517 ( .A1(n9505), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8172) );
  XNOR2_X1 U10518 ( .A(n8190), .B(n8188), .ZN(n9482) );
  NAND2_X1 U10519 ( .A1(n8243), .A2(n9482), .ZN(n8179) );
  MUX2_X1 U10520 ( .A(n8361), .B(n8174), .S(P3_IR_REG_3__SCAN_IN), .Z(n8175)
         );
  INV_X1 U10521 ( .A(n8175), .ZN(n8177) );
  NAND2_X1 U10522 ( .A1(n8177), .A2(n8212), .ZN(n10015) );
  NAND2_X1 U10523 ( .A1(n8457), .A2(n10015), .ZN(n8178) );
  NAND2_X1 U10524 ( .A1(n10466), .A2(n10091), .ZN(n8802) );
  INV_X1 U10525 ( .A(n10091), .ZN(n10385) );
  NAND2_X1 U10526 ( .A1(n8513), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U10527 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8181) );
  NAND2_X1 U10528 ( .A1(n8200), .A2(n8181), .ZN(n10460) );
  NAND2_X1 U10529 ( .A1(n8604), .A2(n10460), .ZN(n8186) );
  INV_X1 U10530 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10018) );
  OR2_X1 U10531 ( .A1(n8756), .A2(n10018), .ZN(n8185) );
  INV_X1 U10532 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8183) );
  OR2_X1 U10533 ( .A1(n8753), .A2(n8183), .ZN(n8184) );
  AND4_X2 U10534 ( .A1(n8187), .A2(n8186), .A3(n8185), .A4(n8184), .ZN(n10638)
         );
  INV_X1 U10535 ( .A(SI_4_), .ZN(n9479) );
  NAND2_X1 U10536 ( .A1(n8762), .A2(n9479), .ZN(n8197) );
  XNOR2_X1 U10537 ( .A(n8209), .B(n8207), .ZN(n9480) );
  NAND2_X1 U10538 ( .A1(n8243), .A2(n9480), .ZN(n8196) );
  NAND2_X1 U10539 ( .A1(n8212), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8194) );
  INV_X1 U10540 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8193) );
  XNOR2_X1 U10541 ( .A(n8194), .B(n8193), .ZN(n15033) );
  NAND2_X1 U10542 ( .A1(n8457), .A2(n15033), .ZN(n8195) );
  INV_X1 U10543 ( .A(n10199), .ZN(n10467) );
  NAND2_X1 U10544 ( .A1(n12381), .A2(n10467), .ZN(n8805) );
  NAND2_X1 U10545 ( .A1(n8606), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U10546 ( .A1(n8200), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8201) );
  NAND2_X1 U10547 ( .A1(n8219), .A2(n8201), .ZN(n10641) );
  NAND2_X1 U10548 ( .A1(n8604), .A2(n10641), .ZN(n8205) );
  INV_X1 U10549 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10474) );
  OR2_X1 U10550 ( .A1(n8756), .A2(n10474), .ZN(n8204) );
  INV_X1 U10551 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8202) );
  OR2_X1 U10552 ( .A1(n8753), .A2(n8202), .ZN(n8203) );
  AND4_X2 U10553 ( .A1(n8206), .A2(n8205), .A3(n8204), .A4(n8203), .ZN(n10776)
         );
  NAND2_X1 U10554 ( .A1(n9504), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8210) );
  XNOR2_X1 U10555 ( .A(n8228), .B(n8226), .ZN(n9500) );
  NAND2_X1 U10556 ( .A1(n8762), .A2(SI_5_), .ZN(n8218) );
  NAND2_X1 U10557 ( .A1(n8214), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8213) );
  MUX2_X1 U10558 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8213), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8216) );
  INV_X1 U10559 ( .A(n8248), .ZN(n8215) );
  NAND2_X1 U10560 ( .A1(n8457), .A2(n10010), .ZN(n8217) );
  NAND2_X1 U10561 ( .A1(n10776), .A2(n10475), .ZN(n8809) );
  NAND2_X1 U10562 ( .A1(n12380), .A2(n10639), .ZN(n8810) );
  AND2_X2 U10563 ( .A1(n8809), .A2(n8810), .ZN(n10424) );
  NAND2_X1 U10564 ( .A1(n8606), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U10565 ( .A1(n8219), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U10566 ( .A1(n8235), .A2(n8220), .ZN(n10772) );
  NAND2_X1 U10567 ( .A1(n8604), .A2(n10772), .ZN(n8224) );
  INV_X1 U10568 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10570) );
  OR2_X1 U10569 ( .A1(n8756), .A2(n10570), .ZN(n8223) );
  INV_X1 U10570 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8221) );
  OR2_X1 U10571 ( .A1(n8753), .A2(n8221), .ZN(n8222) );
  NAND2_X1 U10572 ( .A1(n9503), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8229) );
  XNOR2_X1 U10573 ( .A(n9501), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8230) );
  XNOR2_X1 U10574 ( .A(n8245), .B(n8230), .ZN(n9498) );
  NAND2_X1 U10575 ( .A1(n8762), .A2(SI_6_), .ZN(n8233) );
  OR2_X1 U10576 ( .A1(n8248), .A2(n8361), .ZN(n8231) );
  NAND2_X1 U10577 ( .A1(n8457), .A2(n10060), .ZN(n8232) );
  OAI211_X1 U10578 ( .C1(n6449), .C2(n9498), .A(n8233), .B(n8232), .ZN(n10681)
         );
  NAND2_X1 U10579 ( .A1(n10862), .A2(n10681), .ZN(n8817) );
  INV_X1 U10580 ( .A(n10862), .ZN(n12379) );
  INV_X1 U10581 ( .A(n10681), .ZN(n10777) );
  NAND2_X1 U10582 ( .A1(n12379), .A2(n10777), .ZN(n8816) );
  NAND2_X1 U10583 ( .A1(n10564), .A2(n10565), .ZN(n10563) );
  NAND2_X1 U10584 ( .A1(n10563), .A2(n8817), .ZN(n10813) );
  NAND2_X1 U10585 ( .A1(n8606), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U10586 ( .A1(n8235), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U10587 ( .A1(n8254), .A2(n8236), .ZN(n10858) );
  NAND2_X1 U10588 ( .A1(n8604), .A2(n10858), .ZN(n8241) );
  INV_X1 U10589 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8237) );
  OR2_X1 U10590 ( .A1(n8753), .A2(n8237), .ZN(n8240) );
  INV_X1 U10591 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8238) );
  OR2_X1 U10592 ( .A1(n8756), .A2(n8238), .ZN(n8239) );
  NAND2_X1 U10593 ( .A1(n9496), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8246) );
  XNOR2_X1 U10594 ( .A(n8262), .B(n8261), .ZN(n9471) );
  NAND2_X1 U10595 ( .A1(n8243), .A2(n9471), .ZN(n8253) );
  INV_X1 U10596 ( .A(SI_7_), .ZN(n9470) );
  NAND2_X1 U10597 ( .A1(n8762), .A2(n9470), .ZN(n8252) );
  NAND2_X1 U10598 ( .A1(n8248), .A2(n8247), .ZN(n8265) );
  NAND2_X1 U10599 ( .A1(n8265), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8250) );
  INV_X1 U10600 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8249) );
  XNOR2_X1 U10601 ( .A(n8250), .B(n8249), .ZN(n10298) );
  NAND2_X1 U10602 ( .A1(n8457), .A2(n10298), .ZN(n8251) );
  NAND2_X1 U10603 ( .A1(n10960), .A2(n10820), .ZN(n8820) );
  NAND2_X1 U10604 ( .A1(n12378), .A2(n10988), .ZN(n8821) );
  INV_X1 U10605 ( .A(n10815), .ZN(n10812) );
  NAND2_X1 U10606 ( .A1(n8606), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U10607 ( .A1(n8254), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8255) );
  NAND2_X1 U10608 ( .A1(n8274), .A2(n8255), .ZN(n11046) );
  NAND2_X1 U10609 ( .A1(n8604), .A2(n11046), .ZN(n8259) );
  INV_X1 U10610 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8256) );
  OR2_X1 U10611 ( .A1(n8753), .A2(n8256), .ZN(n8258) );
  INV_X1 U10612 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11045) );
  OR2_X1 U10613 ( .A1(n8756), .A2(n11045), .ZN(n8257) );
  NAND2_X1 U10614 ( .A1(n9522), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8263) );
  XNOR2_X1 U10615 ( .A(n8281), .B(n8280), .ZN(n9475) );
  NAND2_X1 U10616 ( .A1(n8762), .A2(SI_8_), .ZN(n8272) );
  NAND2_X1 U10617 ( .A1(n8268), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8267) );
  MUX2_X1 U10618 ( .A(n8267), .B(P3_IR_REG_31__SCAN_IN), .S(n8266), .Z(n8270)
         );
  INV_X1 U10619 ( .A(n8284), .ZN(n8269) );
  NAND2_X1 U10620 ( .A1(n8457), .A2(n10906), .ZN(n8271) );
  OAI211_X1 U10621 ( .C1(n6449), .C2(n9475), .A(n8272), .B(n8271), .ZN(n11092)
         );
  NAND2_X1 U10622 ( .A1(n11205), .A2(n11092), .ZN(n8825) );
  INV_X1 U10623 ( .A(n11205), .ZN(n12377) );
  NAND2_X1 U10624 ( .A1(n12377), .A2(n11094), .ZN(n8824) );
  NAND2_X1 U10625 ( .A1(n8825), .A2(n8824), .ZN(n11042) );
  INV_X1 U10626 ( .A(n11042), .ZN(n11039) );
  NAND2_X1 U10627 ( .A1(n8673), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8279) );
  INV_X1 U10628 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15065) );
  OR2_X1 U10629 ( .A1(n8756), .A2(n15065), .ZN(n8278) );
  NAND2_X1 U10630 ( .A1(n8606), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U10631 ( .A1(n8274), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U10632 ( .A1(n8289), .A2(n8275), .ZN(n11208) );
  NAND2_X1 U10633 ( .A1(n8604), .A2(n11208), .ZN(n8276) );
  NAND2_X1 U10634 ( .A1(n9529), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8282) );
  XNOR2_X1 U10635 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8297) );
  XNOR2_X1 U10636 ( .A(n8298), .B(n8297), .ZN(n9473) );
  NAND2_X1 U10637 ( .A1(n8243), .A2(n9473), .ZN(n8287) );
  OR2_X1 U10638 ( .A1(n8284), .A2(n8361), .ZN(n8283) );
  MUX2_X1 U10639 ( .A(n8283), .B(P3_IR_REG_31__SCAN_IN), .S(n7030), .Z(n8285)
         );
  NAND2_X1 U10640 ( .A1(n8284), .A2(n7030), .ZN(n8317) );
  NAND2_X1 U10641 ( .A1(n8285), .A2(n8317), .ZN(n15071) );
  NAND2_X1 U10642 ( .A1(n8457), .A2(n15071), .ZN(n8286) );
  NAND2_X1 U10643 ( .A1(n12376), .A2(n11206), .ZN(n8829) );
  INV_X1 U10644 ( .A(n11206), .ZN(n11083) );
  NAND2_X1 U10645 ( .A1(n11341), .A2(n11083), .ZN(n8828) );
  NAND2_X1 U10646 ( .A1(n8606), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U10647 ( .A1(n8289), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10648 ( .A1(n8304), .A2(n8290), .ZN(n11336) );
  NAND2_X1 U10649 ( .A1(n8604), .A2(n11336), .ZN(n8294) );
  INV_X1 U10650 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8291) );
  OR2_X1 U10651 ( .A1(n8753), .A2(n8291), .ZN(n8293) );
  INV_X1 U10652 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10897) );
  OR2_X1 U10653 ( .A1(n8756), .A2(n10897), .ZN(n8292) );
  NAND2_X1 U10654 ( .A1(n8317), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8296) );
  XNOR2_X1 U10655 ( .A(n8296), .B(P3_IR_REG_10__SCAN_IN), .ZN(n15101) );
  INV_X1 U10656 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U10657 ( .A1(n8299), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8300) );
  XNOR2_X1 U10658 ( .A(n9599), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n8311) );
  XNOR2_X1 U10659 ( .A(n8313), .B(n8311), .ZN(n9483) );
  NAND2_X1 U10660 ( .A1(n9483), .A2(n8243), .ZN(n8302) );
  NAND2_X1 U10661 ( .A1(n8762), .A2(SI_10_), .ZN(n8301) );
  OAI211_X1 U10662 ( .C1(n9734), .C2(n10904), .A(n8302), .B(n8301), .ZN(n11196) );
  INV_X1 U10663 ( .A(n11196), .ZN(n11367) );
  NAND2_X1 U10664 ( .A1(n12375), .A2(n11367), .ZN(n8833) );
  NAND2_X1 U10665 ( .A1(n11195), .A2(n8833), .ZN(n8303) );
  NAND2_X1 U10666 ( .A1(n11405), .A2(n11196), .ZN(n8832) );
  NAND2_X1 U10667 ( .A1(n8303), .A2(n8832), .ZN(n11408) );
  NAND2_X1 U10668 ( .A1(n8606), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U10669 ( .A1(n8304), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U10670 ( .A1(n8333), .A2(n8305), .ZN(n11562) );
  NAND2_X1 U10671 ( .A1(n8604), .A2(n11562), .ZN(n8309) );
  INV_X1 U10672 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11411) );
  OR2_X1 U10673 ( .A1(n8756), .A2(n11411), .ZN(n8308) );
  INV_X1 U10674 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8306) );
  OR2_X1 U10675 ( .A1(n8753), .A2(n8306), .ZN(n8307) );
  INV_X1 U10676 ( .A(n8311), .ZN(n8312) );
  NAND2_X1 U10677 ( .A1(n9599), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8314) );
  XNOR2_X1 U10678 ( .A(n9692), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8316) );
  XNOR2_X1 U10679 ( .A(n8322), .B(n8316), .ZN(n9486) );
  NAND2_X1 U10680 ( .A1(n9486), .A2(n8243), .ZN(n8320) );
  OAI21_X1 U10681 ( .B1(n8317), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8318) );
  XNOR2_X1 U10682 ( .A(n8318), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U10683 ( .A1(n8762), .A2(SI_11_), .B1(n8457), .B2(n11143), .ZN(
        n8319) );
  NAND2_X1 U10684 ( .A1(n11646), .A2(n11409), .ZN(n8837) );
  NAND2_X1 U10685 ( .A1(n11560), .A2(n12374), .ZN(n8838) );
  NAND2_X1 U10686 ( .A1(n11408), .A2(n11407), .ZN(n11406) );
  NAND2_X1 U10687 ( .A1(n9692), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10688 ( .A1(n9842), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10689 ( .A1(n9840), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10690 ( .A1(n8341), .A2(n8324), .ZN(n8339) );
  XNOR2_X1 U10691 ( .A(n8340), .B(n8339), .ZN(n14403) );
  NAND2_X1 U10692 ( .A1(n14403), .A2(n8243), .ZN(n8329) );
  NAND2_X1 U10693 ( .A1(n8325), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8326) );
  XNOR2_X1 U10694 ( .A(n8326), .B(n8106), .ZN(n14406) );
  AOI22_X1 U10695 ( .A1(n8762), .A2(n8327), .B1(n8457), .B2(n14406), .ZN(n8328) );
  NAND2_X1 U10696 ( .A1(n8329), .A2(n8328), .ZN(n14471) );
  NAND2_X1 U10697 ( .A1(n8673), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8338) );
  INV_X1 U10698 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n8330) );
  OR2_X1 U10699 ( .A1(n8756), .A2(n8330), .ZN(n8337) );
  NAND2_X1 U10700 ( .A1(n8606), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8336) );
  INV_X1 U10701 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10702 ( .A1(n8333), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U10703 ( .A1(n8350), .A2(n8334), .ZN(n11642) );
  NAND2_X1 U10704 ( .A1(n8604), .A2(n11642), .ZN(n8335) );
  NAND4_X1 U10705 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(n12373) );
  OR2_X1 U10706 ( .A1(n14471), .A2(n12373), .ZN(n8843) );
  NAND2_X1 U10707 ( .A1(n14471), .A2(n12373), .ZN(n8842) );
  XNOR2_X1 U10708 ( .A(n8357), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n14407) );
  NAND2_X1 U10709 ( .A1(n14407), .A2(n8243), .ZN(n8348) );
  NAND2_X1 U10710 ( .A1(n8343), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8344) );
  MUX2_X1 U10711 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8344), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8345) );
  INV_X1 U10712 ( .A(n8345), .ZN(n8346) );
  NOR2_X1 U10713 ( .A1(n8346), .A2(n8396), .ZN(n12405) );
  AOI22_X1 U10714 ( .A1(n8762), .A2(SI_13_), .B1(n8457), .B2(n12405), .ZN(
        n8347) );
  NAND2_X1 U10715 ( .A1(n8348), .A2(n8347), .ZN(n11519) );
  NAND2_X1 U10716 ( .A1(n8606), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8356) );
  INV_X1 U10717 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U10718 ( .A1(n8350), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U10719 ( .A1(n8365), .A2(n8351), .ZN(n11514) );
  NAND2_X1 U10720 ( .A1(n8604), .A2(n11514), .ZN(n8355) );
  INV_X1 U10721 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n11653) );
  OR2_X1 U10722 ( .A1(n8753), .A2(n11653), .ZN(n8354) );
  INV_X1 U10723 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8352) );
  OR2_X1 U10724 ( .A1(n8756), .A2(n8352), .ZN(n8353) );
  OR2_X1 U10725 ( .A1(n11519), .A2(n11328), .ZN(n8848) );
  NAND2_X1 U10726 ( .A1(n11519), .A2(n11328), .ZN(n8847) );
  INV_X1 U10727 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U10728 ( .A1(n10100), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8374) );
  INV_X1 U10729 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10102) );
  NAND2_X1 U10730 ( .A1(n10102), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8360) );
  AND2_X1 U10731 ( .A1(n8374), .A2(n8360), .ZN(n8372) );
  XNOR2_X1 U10732 ( .A(n8373), .B(n8372), .ZN(n9535) );
  NAND2_X1 U10733 ( .A1(n9535), .A2(n8243), .ZN(n8364) );
  OR2_X1 U10734 ( .A1(n8396), .A2(n8361), .ZN(n8362) );
  XNOR2_X1 U10735 ( .A(n8362), .B(n12100), .ZN(n12440) );
  AOI22_X1 U10736 ( .A1(n8762), .A2(n7261), .B1(n8457), .B2(n12440), .ZN(n8363) );
  NAND2_X1 U10737 ( .A1(n8606), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8370) );
  INV_X1 U10738 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12407) );
  OR2_X1 U10739 ( .A1(n8756), .A2(n12407), .ZN(n8369) );
  NAND2_X1 U10740 ( .A1(n8673), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10741 ( .A1(n8365), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U10742 ( .A1(n8383), .A2(n8366), .ZN(n11633) );
  NAND2_X1 U10743 ( .A1(n8604), .A2(n11633), .ZN(n8367) );
  NAND4_X1 U10744 ( .A1(n8370), .A2(n8369), .A3(n8368), .A4(n8367), .ZN(n12371) );
  NAND2_X1 U10745 ( .A1(n11630), .A2(n12371), .ZN(n8852) );
  NAND2_X1 U10746 ( .A1(n11445), .A2(n11446), .ZN(n8371) );
  NAND2_X1 U10747 ( .A1(n8371), .A2(n8853), .ZN(n11664) );
  NAND2_X1 U10748 ( .A1(n10176), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10749 ( .A1(n10178), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U10750 ( .A1(n8393), .A2(n8376), .ZN(n8390) );
  XNOR2_X1 U10751 ( .A(n8392), .B(n8390), .ZN(n14413) );
  NAND2_X1 U10752 ( .A1(n14413), .A2(n8243), .ZN(n8380) );
  NAND2_X1 U10753 ( .A1(n8396), .A2(n12100), .ZN(n8377) );
  NAND2_X1 U10754 ( .A1(n8377), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8378) );
  XNOR2_X1 U10755 ( .A(n8378), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U10756 ( .A1(n8762), .A2(SI_15_), .B1(n8457), .B2(n12462), .ZN(
        n8379) );
  NAND2_X1 U10757 ( .A1(n8673), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8388) );
  INV_X1 U10758 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12434) );
  OR2_X1 U10759 ( .A1(n8756), .A2(n12434), .ZN(n8387) );
  NAND2_X1 U10760 ( .A1(n8606), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8386) );
  INV_X1 U10761 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U10762 ( .A1(n8383), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U10763 ( .A1(n8400), .A2(n8384), .ZN(n12357) );
  NAND2_X1 U10764 ( .A1(n8604), .A2(n12357), .ZN(n8385) );
  NAND4_X1 U10765 ( .A1(n8388), .A2(n8387), .A3(n8386), .A4(n8385), .ZN(n12370) );
  OR2_X1 U10766 ( .A1(n11666), .A2(n11629), .ZN(n8857) );
  NAND2_X1 U10767 ( .A1(n11666), .A2(n11629), .ZN(n8856) );
  NAND2_X1 U10768 ( .A1(n11664), .A2(n11665), .ZN(n8389) );
  NAND2_X1 U10769 ( .A1(n8389), .A2(n8856), .ZN(n11605) );
  INV_X1 U10770 ( .A(n8390), .ZN(n8391) );
  NAND2_X1 U10771 ( .A1(n10436), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10772 ( .A1(n10459), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10773 ( .A1(n8410), .A2(n8394), .ZN(n8407) );
  XNOR2_X1 U10774 ( .A(n8409), .B(n8407), .ZN(n14416) );
  NAND2_X1 U10775 ( .A1(n14416), .A2(n8243), .ZN(n8399) );
  NOR2_X1 U10776 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n8395) );
  OR2_X1 U10777 ( .A1(n8413), .A2(n8361), .ZN(n8397) );
  XNOR2_X1 U10778 ( .A(n8397), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U10779 ( .A1(n8762), .A2(SI_16_), .B1(n8457), .B2(n12494), .ZN(
        n8398) );
  NAND2_X1 U10780 ( .A1(n8673), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8405) );
  INV_X1 U10781 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12464) );
  OR2_X1 U10782 ( .A1(n8756), .A2(n12464), .ZN(n8404) );
  NAND2_X1 U10783 ( .A1(n8606), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10784 ( .A1(n8400), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10785 ( .A1(n8424), .A2(n8401), .ZN(n12293) );
  NAND2_X1 U10786 ( .A1(n8604), .A2(n12293), .ZN(n8402) );
  NAND4_X1 U10787 ( .A1(n8405), .A2(n8404), .A3(n8403), .A4(n8402), .ZN(n12369) );
  XNOR2_X1 U10788 ( .A(n12747), .B(n12369), .ZN(n11604) );
  NAND2_X1 U10789 ( .A1(n11605), .A2(n11604), .ZN(n8406) );
  INV_X1 U10790 ( .A(n12369), .ZN(n12682) );
  NAND2_X1 U10791 ( .A1(n12747), .A2(n12682), .ZN(n8863) );
  NAND2_X1 U10792 ( .A1(n8406), .A2(n8863), .ZN(n12684) );
  INV_X1 U10793 ( .A(n8407), .ZN(n8408) );
  AOI22_X1 U10794 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10472), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n10496), .ZN(n8411) );
  XNOR2_X1 U10795 ( .A(n8433), .B(n8411), .ZN(n14395) );
  NAND2_X1 U10796 ( .A1(n14395), .A2(n8243), .ZN(n8421) );
  INV_X1 U10797 ( .A(SI_17_), .ZN(n8419) );
  INV_X1 U10798 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8412) );
  NOR2_X1 U10799 ( .A1(n8417), .A2(n8361), .ZN(n8414) );
  MUX2_X1 U10800 ( .A(n8361), .B(n8414), .S(P3_IR_REG_17__SCAN_IN), .Z(n8415)
         );
  INV_X1 U10801 ( .A(n8415), .ZN(n8418) );
  INV_X1 U10802 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U10803 ( .A1(n8418), .A2(n8455), .ZN(n14398) );
  AOI22_X1 U10804 ( .A1(n8762), .A2(n8419), .B1(n8457), .B2(n14398), .ZN(n8420) );
  NAND2_X1 U10805 ( .A1(n8673), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8430) );
  INV_X1 U10806 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U10807 ( .A1(n8424), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10808 ( .A1(n8444), .A2(n8425), .ZN(n12686) );
  NAND2_X1 U10809 ( .A1(n12686), .A2(n8604), .ZN(n8429) );
  NAND2_X1 U10810 ( .A1(n8606), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10811 ( .A1(n8426), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8427) );
  NAND4_X1 U10812 ( .A1(n8430), .A2(n8429), .A3(n8428), .A4(n8427), .ZN(n12668) );
  NAND2_X1 U10813 ( .A1(n12813), .A2(n12668), .ZN(n8868) );
  NAND2_X1 U10814 ( .A1(n12684), .A2(n12685), .ZN(n8431) );
  NAND2_X1 U10815 ( .A1(n8431), .A2(n8870), .ZN(n12672) );
  INV_X1 U10816 ( .A(n12672), .ZN(n8451) );
  NAND2_X1 U10817 ( .A1(n10472), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U10818 ( .A1(n10496), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8434) );
  INV_X1 U10819 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10884) );
  NAND2_X1 U10820 ( .A1(n10884), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8452) );
  INV_X1 U10821 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U10822 ( .A1(n10882), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10823 ( .A1(n8452), .A2(n8436), .ZN(n8437) );
  NAND2_X1 U10824 ( .A1(n8438), .A2(n8437), .ZN(n8439) );
  NAND2_X1 U10825 ( .A1(n8453), .A2(n8439), .ZN(n14423) );
  NAND2_X1 U10826 ( .A1(n14423), .A2(n8243), .ZN(n8443) );
  NAND2_X1 U10827 ( .A1(n8455), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8441) );
  XNOR2_X1 U10828 ( .A(n8441), .B(n8440), .ZN(n14425) );
  INV_X1 U10829 ( .A(n14425), .ZN(n12509) );
  AOI22_X1 U10830 ( .A1(n8762), .A2(SI_18_), .B1(n8457), .B2(n12509), .ZN(
        n8442) );
  NAND2_X1 U10831 ( .A1(n8444), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10832 ( .A1(n8461), .A2(n8445), .ZN(n12673) );
  NAND2_X1 U10833 ( .A1(n12673), .A2(n8604), .ZN(n8450) );
  NAND2_X1 U10834 ( .A1(n8673), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10835 ( .A1(n8606), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8446) );
  AND2_X1 U10836 ( .A1(n8447), .A2(n8446), .ZN(n8449) );
  NAND2_X1 U10837 ( .A1(n8426), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U10838 ( .A1(n12739), .A2(n12681), .ZN(n8872) );
  INV_X1 U10839 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12129) );
  INV_X1 U10840 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U10841 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(
        P1_DATAO_REG_19__SCAN_IN), .B1(n12129), .B2(n10986), .ZN(n8454) );
  XNOR2_X1 U10842 ( .A(n8467), .B(n8454), .ZN(n10074) );
  NAND2_X1 U10843 ( .A1(n10074), .A2(n8243), .ZN(n8459) );
  INV_X1 U10844 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8456) );
  AOI22_X1 U10845 ( .A1(n8762), .A2(n10073), .B1(n8457), .B2(n12517), .ZN(
        n8458) );
  INV_X1 U10846 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n8465) );
  INV_X1 U10847 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12262) );
  NAND2_X1 U10848 ( .A1(n8461), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U10849 ( .A1(n8470), .A2(n8462), .ZN(n12660) );
  NAND2_X1 U10850 ( .A1(n12660), .A2(n8604), .ZN(n8464) );
  AOI22_X1 U10851 ( .A1(n8673), .A2(P3_REG0_REG_19__SCAN_IN), .B1(n8606), .B2(
        P3_REG1_REG_19__SCAN_IN), .ZN(n8463) );
  OAI211_X1 U10852 ( .C1(n8756), .C2(n8465), .A(n8464), .B(n8463), .ZN(n12667)
         );
  NAND2_X1 U10853 ( .A1(n12808), .A2(n12667), .ZN(n8877) );
  OR2_X1 U10854 ( .A1(n12808), .A2(n12667), .ZN(n8876) );
  NAND2_X1 U10855 ( .A1(n8466), .A2(n8876), .ZN(n12644) );
  INV_X1 U10856 ( .A(n12644), .ZN(n8475) );
  XNOR2_X1 U10857 ( .A(n8476), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U10858 ( .A1(n10368), .A2(n8243), .ZN(n8469) );
  NAND2_X1 U10859 ( .A1(n8762), .A2(SI_20_), .ZN(n8468) );
  NAND2_X1 U10860 ( .A1(n8470), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U10861 ( .A1(n8485), .A2(n8471), .ZN(n12647) );
  NAND2_X1 U10862 ( .A1(n12647), .A2(n8604), .ZN(n8474) );
  AOI22_X1 U10863 ( .A1(n8673), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n8513), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10864 ( .A1(n8426), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U10865 ( .A1(n12646), .A2(n12654), .ZN(n8882) );
  NAND2_X1 U10866 ( .A1(n8477), .A2(n11037), .ZN(n8478) );
  INV_X1 U10867 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U10868 ( .A1(n11186), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10869 ( .A1(n11189), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8480) );
  AND2_X1 U10870 ( .A1(n8495), .A2(n8480), .ZN(n8492) );
  XNOR2_X1 U10871 ( .A(n8494), .B(n8492), .ZN(n10497) );
  NAND2_X1 U10872 ( .A1(n10497), .A2(n8243), .ZN(n8482) );
  NAND2_X1 U10873 ( .A1(n8762), .A2(SI_21_), .ZN(n8481) );
  INV_X1 U10874 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U10875 ( .A1(n8485), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10876 ( .A1(n8498), .A2(n8486), .ZN(n12632) );
  INV_X1 U10877 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10878 ( .A1(n8673), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10879 ( .A1(n8606), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8487) );
  OAI211_X1 U10880 ( .C1(n8489), .C2(n8756), .A(n8488), .B(n8487), .ZN(n8490)
         );
  AOI21_X1 U10881 ( .B1(n12632), .B2(n8604), .A(n8490), .ZN(n12641) );
  OR2_X1 U10882 ( .A1(n12631), .A2(n12641), .ZN(n8784) );
  NAND2_X1 U10883 ( .A1(n12631), .A2(n12641), .ZN(n8785) );
  INV_X1 U10884 ( .A(n8492), .ZN(n8493) );
  XNOR2_X1 U10885 ( .A(n11371), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8506) );
  XNOR2_X1 U10886 ( .A(n8507), .B(n8506), .ZN(n10559) );
  NAND2_X1 U10887 ( .A1(n10559), .A2(n8243), .ZN(n8497) );
  NAND2_X1 U10888 ( .A1(n8762), .A2(SI_22_), .ZN(n8496) );
  NAND2_X1 U10889 ( .A1(n8498), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U10890 ( .A1(n8511), .A2(n8499), .ZN(n12621) );
  NAND2_X1 U10891 ( .A1(n12621), .A2(n8604), .ZN(n8505) );
  INV_X1 U10892 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U10893 ( .A1(n8673), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U10894 ( .A1(n8513), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8500) );
  OAI211_X1 U10895 ( .C1(n8502), .C2(n8756), .A(n8501), .B(n8500), .ZN(n8503)
         );
  INV_X1 U10896 ( .A(n8503), .ZN(n8504) );
  NAND2_X1 U10897 ( .A1(n8505), .A2(n8504), .ZN(n12365) );
  AND2_X1 U10898 ( .A1(n12324), .A2(n12628), .ZN(n8783) );
  OR2_X1 U10899 ( .A1(n12324), .A2(n12628), .ZN(n8888) );
  NAND2_X1 U10900 ( .A1(n11371), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8508) );
  XNOR2_X1 U10901 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8520) );
  XNOR2_X1 U10902 ( .A(n8521), .B(n8520), .ZN(n10827) );
  NAND2_X1 U10903 ( .A1(n10827), .A2(n8243), .ZN(n8510) );
  NAND2_X1 U10904 ( .A1(n8762), .A2(SI_23_), .ZN(n8509) );
  NAND2_X1 U10905 ( .A1(n8511), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U10906 ( .A1(n8530), .A2(n8512), .ZN(n12611) );
  NAND2_X1 U10907 ( .A1(n12611), .A2(n8604), .ZN(n8518) );
  INV_X1 U10908 ( .A(n8513), .ZN(n8676) );
  INV_X1 U10909 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12720) );
  NAND2_X1 U10910 ( .A1(n8673), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10911 ( .A1(n8426), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8514) );
  OAI211_X1 U10912 ( .C1(n8676), .C2(n12720), .A(n8515), .B(n8514), .ZN(n8516)
         );
  INV_X1 U10913 ( .A(n8516), .ZN(n8517) );
  NAND2_X1 U10914 ( .A1(n12610), .A2(n12618), .ZN(n8519) );
  INV_X1 U10915 ( .A(n12608), .ZN(n8891) );
  NAND2_X1 U10916 ( .A1(n11420), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U10917 ( .A1(n8524), .A2(n13468), .ZN(n8525) );
  INV_X1 U10918 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14287) );
  XNOR2_X1 U10919 ( .A(n8537), .B(n14287), .ZN(n11128) );
  NAND2_X1 U10920 ( .A1(n11128), .A2(n8243), .ZN(n8527) );
  NAND2_X1 U10921 ( .A1(n8762), .A2(SI_24_), .ZN(n8526) );
  INV_X1 U10922 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10923 ( .A1(n8530), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8531) );
  NAND2_X1 U10924 ( .A1(n8543), .A2(n8531), .ZN(n12599) );
  NAND2_X1 U10925 ( .A1(n12599), .A2(n8604), .ZN(n8536) );
  INV_X1 U10926 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12121) );
  NAND2_X1 U10927 ( .A1(n8673), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10928 ( .A1(n8513), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8532) );
  OAI211_X1 U10929 ( .C1(n12121), .C2(n8756), .A(n8533), .B(n8532), .ZN(n8534)
         );
  INV_X1 U10930 ( .A(n8534), .ZN(n8535) );
  INV_X1 U10931 ( .A(n12592), .ZN(n8938) );
  NAND2_X1 U10932 ( .A1(n12591), .A2(n12579), .ZN(n8551) );
  XNOR2_X1 U10933 ( .A(n13464), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8538) );
  XNOR2_X1 U10934 ( .A(n8553), .B(n8538), .ZN(n12252) );
  NAND2_X1 U10935 ( .A1(n12252), .A2(n8243), .ZN(n8540) );
  NAND2_X1 U10936 ( .A1(n8762), .A2(SI_25_), .ZN(n8539) );
  INV_X1 U10937 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U10938 ( .A1(n8543), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10939 ( .A1(n8560), .A2(n8544), .ZN(n12583) );
  NAND2_X1 U10940 ( .A1(n12583), .A2(n8604), .ZN(n8550) );
  INV_X1 U10941 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10942 ( .A1(n8673), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U10943 ( .A1(n8513), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8545) );
  OAI211_X1 U10944 ( .C1(n8547), .C2(n8756), .A(n8546), .B(n8545), .ZN(n8548)
         );
  INV_X1 U10945 ( .A(n8548), .ZN(n8549) );
  XNOR2_X1 U10946 ( .A(n12709), .B(n12594), .ZN(n12580) );
  INV_X1 U10947 ( .A(n12580), .ZN(n8939) );
  NAND2_X1 U10948 ( .A1(n8551), .A2(n8939), .ZN(n12582) );
  NAND2_X1 U10949 ( .A1(n12709), .A2(n12594), .ZN(n8897) );
  NAND2_X1 U10950 ( .A1(n13464), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U10951 ( .A1(n14283), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8554) );
  AOI22_X1 U10952 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13459), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14278), .ZN(n8556) );
  XNOR2_X1 U10953 ( .A(n8570), .B(n8556), .ZN(n11324) );
  NAND2_X1 U10954 ( .A1(n8762), .A2(SI_26_), .ZN(n8558) );
  INV_X2 U10955 ( .A(n9340), .ZN(n12783) );
  NAND2_X1 U10956 ( .A1(n8560), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10957 ( .A1(n8578), .A2(n8561), .ZN(n12567) );
  NAND2_X1 U10958 ( .A1(n12567), .A2(n8604), .ZN(n8567) );
  INV_X1 U10959 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U10960 ( .A1(n8673), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U10961 ( .A1(n8513), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8562) );
  OAI211_X1 U10962 ( .C1(n8564), .C2(n8756), .A(n8563), .B(n8562), .ZN(n8565)
         );
  INV_X1 U10963 ( .A(n8565), .ZN(n8566) );
  NAND2_X1 U10964 ( .A1(n12783), .A2(n12578), .ZN(n8902) );
  INV_X1 U10965 ( .A(n12578), .ZN(n12283) );
  NAND2_X1 U10966 ( .A1(n9340), .A2(n12283), .ZN(n8903) );
  AND2_X1 U10967 ( .A1(n14278), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10968 ( .A1(n13459), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8571) );
  AOI22_X1 U10969 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13454), .B2(n11774), .ZN(n8572) );
  INV_X1 U10970 ( .A(n8572), .ZN(n8573) );
  NAND2_X1 U10971 ( .A1(n11450), .A2(n8243), .ZN(n8575) );
  NAND2_X1 U10972 ( .A1(n8762), .A2(SI_27_), .ZN(n8574) );
  INV_X1 U10973 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U10974 ( .A1(n8578), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U10975 ( .A1(n8593), .A2(n8579), .ZN(n12557) );
  NAND2_X1 U10976 ( .A1(n12557), .A2(n8604), .ZN(n8585) );
  INV_X1 U10977 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U10978 ( .A1(n8606), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U10979 ( .A1(n8673), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8580) );
  OAI211_X1 U10980 ( .C1(n8756), .C2(n8582), .A(n8581), .B(n8580), .ZN(n8583)
         );
  INV_X1 U10981 ( .A(n8583), .ZN(n8584) );
  NAND2_X1 U10982 ( .A1(n12701), .A2(n12564), .ZN(n8908) );
  AND2_X1 U10983 ( .A1(n13454), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U10984 ( .A1(n11774), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8586) );
  OAI21_X2 U10985 ( .B1(n8588), .B2(n8587), .A(n8586), .ZN(n8599) );
  AOI22_X1 U10986 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8600), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n11773), .ZN(n8589) );
  INV_X1 U10987 ( .A(n8589), .ZN(n8590) );
  XNOR2_X1 U10988 ( .A(n8599), .B(n8590), .ZN(n12828) );
  NAND2_X1 U10989 ( .A1(n12828), .A2(n8243), .ZN(n8592) );
  NAND2_X1 U10990 ( .A1(n8762), .A2(SI_28_), .ZN(n8591) );
  NAND2_X1 U10991 ( .A1(n8593), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10992 ( .A1(n12526), .A2(n8594), .ZN(n12545) );
  INV_X1 U10993 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12187) );
  NAND2_X1 U10994 ( .A1(n8513), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8596) );
  INV_X1 U10995 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12776) );
  OR2_X1 U10996 ( .A1(n8753), .A2(n12776), .ZN(n8595) );
  OAI211_X1 U10997 ( .C1(n12187), .C2(n8756), .A(n8596), .B(n8595), .ZN(n8597)
         );
  AOI21_X1 U10998 ( .B1(n12545), .B2(n8604), .A(n8597), .ZN(n9368) );
  AND2_X1 U10999 ( .A1(n11773), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U11000 ( .A1(n8600), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8601) );
  XNOR2_X1 U11001 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n8745) );
  XNOR2_X1 U11002 ( .A(n8747), .B(n8745), .ZN(n12002) );
  NAND2_X1 U11003 ( .A1(n12002), .A2(n8243), .ZN(n8603) );
  NAND2_X1 U11004 ( .A1(n8762), .A2(SI_29_), .ZN(n8602) );
  INV_X1 U11005 ( .A(n12526), .ZN(n8605) );
  NAND2_X1 U11006 ( .A1(n8605), .A2(n8198), .ZN(n8759) );
  INV_X1 U11007 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n8609) );
  NAND2_X1 U11008 ( .A1(n8606), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U11009 ( .A1(n8673), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8607) );
  OAI211_X1 U11010 ( .C1(n8756), .C2(n8609), .A(n8608), .B(n8607), .ZN(n8610)
         );
  INV_X1 U11011 ( .A(n8610), .ZN(n8611) );
  NAND2_X1 U11012 ( .A1(n8759), .A2(n8611), .ZN(n12539) );
  INV_X1 U11013 ( .A(n8686), .ZN(n8615) );
  NAND2_X1 U11014 ( .A1(n8615), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8612) );
  INV_X1 U11015 ( .A(n10560), .ZN(n8732) );
  NAND2_X1 U11016 ( .A1(n8613), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8614) );
  MUX2_X1 U11017 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8614), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8616) );
  INV_X1 U11018 ( .A(n8617), .ZN(n8618) );
  NAND2_X1 U11019 ( .A1(n8618), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8619) );
  MUX2_X1 U11020 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8619), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8620) );
  NAND2_X1 U11021 ( .A1(n8620), .A2(n8613), .ZN(n10371) );
  NAND2_X1 U11022 ( .A1(n10500), .A2(n10371), .ZN(n8731) );
  XNOR2_X1 U11023 ( .A(n8731), .B(n10560), .ZN(n8622) );
  NAND2_X1 U11024 ( .A1(n12517), .A2(n10500), .ZN(n8621) );
  AND2_X1 U11025 ( .A1(n8622), .A2(n8621), .ZN(n8714) );
  INV_X1 U11026 ( .A(n8714), .ZN(n9349) );
  NAND2_X1 U11027 ( .A1(n8732), .A2(n10500), .ZN(n14470) );
  NAND2_X1 U11028 ( .A1(n9349), .A2(n14470), .ZN(n9979) );
  MUX2_X1 U11029 ( .A(n8732), .B(n9979), .S(n10371), .Z(n8623) );
  INV_X1 U11030 ( .A(n8623), .ZN(n8624) );
  NAND2_X1 U11031 ( .A1(n8624), .A2(n12517), .ZN(n12766) );
  NAND2_X1 U11032 ( .A1(n8947), .A2(n10371), .ZN(n15109) );
  OR2_X1 U11033 ( .A1(n15109), .A2(n10560), .ZN(n12713) );
  NAND2_X2 U11034 ( .A1(n12766), .A2(n12713), .ZN(n14475) );
  INV_X1 U11035 ( .A(n9368), .ZN(n12552) );
  NAND2_X1 U11036 ( .A1(n12757), .A2(n10114), .ZN(n9263) );
  NAND2_X1 U11037 ( .A1(n12765), .A2(n9263), .ZN(n8626) );
  NAND2_X1 U11038 ( .A1(n9265), .A2(n10036), .ZN(n8625) );
  NAND2_X1 U11039 ( .A1(n10185), .A2(n10186), .ZN(n8628) );
  NAND2_X1 U11040 ( .A1(n12760), .A2(n10078), .ZN(n8627) );
  NAND2_X1 U11041 ( .A1(n8628), .A2(n8627), .ZN(n10085) );
  INV_X1 U11042 ( .A(n10085), .ZN(n8630) );
  NAND2_X1 U11043 ( .A1(n8630), .A2(n8629), .ZN(n10087) );
  NAND2_X1 U11044 ( .A1(n12382), .A2(n10091), .ZN(n8631) );
  NAND2_X1 U11045 ( .A1(n10087), .A2(n8631), .ZN(n10132) );
  NAND2_X1 U11046 ( .A1(n12381), .A2(n10199), .ZN(n8632) );
  NAND2_X1 U11047 ( .A1(n10776), .A2(n10639), .ZN(n8634) );
  INV_X1 U11048 ( .A(n10566), .ZN(n8636) );
  INV_X1 U11049 ( .A(n10565), .ZN(n8635) );
  NAND2_X1 U11050 ( .A1(n8636), .A2(n8635), .ZN(n10568) );
  NAND2_X1 U11051 ( .A1(n12379), .A2(n10681), .ZN(n8637) );
  NAND2_X1 U11052 ( .A1(n10568), .A2(n8637), .ZN(n10816) );
  NAND2_X1 U11053 ( .A1(n12378), .A2(n10820), .ZN(n8638) );
  NAND2_X1 U11054 ( .A1(n11205), .A2(n11094), .ZN(n8639) );
  XNOR2_X1 U11055 ( .A(n12376), .B(n11206), .ZN(n11071) );
  NAND2_X1 U11056 ( .A1(n12376), .A2(n11083), .ZN(n8640) );
  NAND2_X1 U11057 ( .A1(n8832), .A2(n8833), .ZN(n11190) );
  NAND2_X1 U11058 ( .A1(n11646), .A2(n11560), .ZN(n8649) );
  AND2_X1 U11059 ( .A1(n11190), .A2(n8649), .ZN(n8641) );
  NAND2_X1 U11060 ( .A1(n11191), .A2(n8641), .ZN(n8645) );
  INV_X1 U11061 ( .A(n8649), .ZN(n8643) );
  NAND2_X1 U11062 ( .A1(n12375), .A2(n11196), .ZN(n11401) );
  NAND2_X1 U11063 ( .A1(n12374), .A2(n11409), .ZN(n8642) );
  AND2_X1 U11064 ( .A1(n11401), .A2(n8642), .ZN(n8647) );
  OR2_X1 U11065 ( .A1(n8643), .A2(n8647), .ZN(n8644) );
  NAND2_X1 U11066 ( .A1(n11326), .A2(n12373), .ZN(n8646) );
  NAND2_X1 U11067 ( .A1(n8646), .A2(n14471), .ZN(n8653) );
  INV_X1 U11068 ( .A(n12373), .ZN(n11556) );
  AND2_X1 U11069 ( .A1(n8647), .A2(n11556), .ZN(n8648) );
  NAND2_X1 U11070 ( .A1(n11402), .A2(n8648), .ZN(n8651) );
  OR2_X1 U11071 ( .A1(n12373), .A2(n8649), .ZN(n8650) );
  NAND2_X1 U11072 ( .A1(n8653), .A2(n8652), .ZN(n11487) );
  NAND2_X1 U11073 ( .A1(n8848), .A2(n8847), .ZN(n8841) );
  NAND2_X1 U11074 ( .A1(n11487), .A2(n8841), .ZN(n8655) );
  OR2_X1 U11075 ( .A1(n11519), .A2(n12372), .ZN(n8654) );
  INV_X1 U11076 ( .A(n12371), .ZN(n11663) );
  OR2_X1 U11077 ( .A1(n11630), .A2(n11663), .ZN(n11659) );
  NAND2_X1 U11078 ( .A1(n11666), .A2(n12370), .ZN(n8656) );
  AND2_X1 U11079 ( .A1(n11659), .A2(n8656), .ZN(n8657) );
  OR2_X1 U11080 ( .A1(n7434), .A2(n8657), .ZN(n8658) );
  AND2_X1 U11081 ( .A1(n12747), .A2(n12369), .ZN(n8659) );
  INV_X1 U11082 ( .A(n12668), .ZN(n12291) );
  INV_X1 U11083 ( .A(n8660), .ZN(n12665) );
  NAND2_X1 U11084 ( .A1(n12665), .A2(n8661), .ZN(n12664) );
  INV_X1 U11085 ( .A(n12681), .ZN(n12368) );
  OR2_X1 U11086 ( .A1(n12739), .A2(n12368), .ZN(n8662) );
  NAND2_X1 U11087 ( .A1(n8876), .A2(n8877), .ZN(n12658) );
  INV_X1 U11088 ( .A(n12667), .ZN(n12332) );
  OR2_X1 U11089 ( .A1(n12808), .A2(n12332), .ZN(n8663) );
  NAND2_X1 U11090 ( .A1(n12646), .A2(n12367), .ZN(n8664) );
  INV_X1 U11091 ( .A(n12641), .ZN(n12366) );
  NOR2_X1 U11092 ( .A1(n12324), .A2(n12365), .ZN(n8665) );
  NAND2_X1 U11093 ( .A1(n12605), .A2(n12608), .ZN(n8667) );
  NAND2_X1 U11094 ( .A1(n12610), .A2(n12364), .ZN(n8666) );
  INV_X1 U11095 ( .A(n12607), .ZN(n12363) );
  OR2_X1 U11096 ( .A1(n12297), .A2(n12363), .ZN(n12573) );
  AND2_X1 U11097 ( .A1(n12580), .A2(n12573), .ZN(n8668) );
  NAND2_X1 U11098 ( .A1(n12709), .A2(n12362), .ZN(n8669) );
  NAND2_X1 U11099 ( .A1(n12572), .A2(n8669), .ZN(n12562) );
  AND2_X1 U11100 ( .A1(n9340), .A2(n12578), .ZN(n8671) );
  NAND2_X1 U11101 ( .A1(n12783), .A2(n12283), .ZN(n8670) );
  NAND2_X1 U11102 ( .A1(n8947), .A2(n10560), .ZN(n8734) );
  INV_X1 U11103 ( .A(n10371), .ZN(n8736) );
  NAND2_X1 U11104 ( .A1(n9258), .A2(n8736), .ZN(n8776) );
  INV_X1 U11105 ( .A(n12833), .ZN(n9755) );
  INV_X1 U11106 ( .A(n6622), .ZN(n12511) );
  NAND2_X1 U11107 ( .A1(n9755), .A2(n12511), .ZN(n9737) );
  NAND2_X1 U11108 ( .A1(n9737), .A2(n9734), .ZN(n8679) );
  INV_X1 U11109 ( .A(n8679), .ZN(n8672) );
  INV_X1 U11110 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14469) );
  NAND2_X1 U11111 ( .A1(n8673), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11112 ( .A1(n8426), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8674) );
  OAI211_X1 U11113 ( .C1(n8676), .C2(n14469), .A(n8675), .B(n8674), .ZN(n8677)
         );
  INV_X1 U11114 ( .A(n8677), .ZN(n8678) );
  AND2_X1 U11115 ( .A1(n8759), .A2(n8678), .ZN(n10826) );
  NAND2_X1 U11116 ( .A1(n9755), .A2(P3_B_REG_SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11117 ( .A1(n12666), .A2(n8680), .ZN(n12524) );
  NOR2_X1 U11118 ( .A1(n10826), .A2(n12524), .ZN(n8681) );
  INV_X1 U11119 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8685) );
  INV_X1 U11120 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U11121 ( .A1(n8720), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8688) );
  MUX2_X1 U11122 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8688), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8689) );
  NAND2_X1 U11123 ( .A1(n8689), .A2(n8692), .ZN(n11130) );
  XNOR2_X1 U11124 ( .A(n11130), .B(P3_B_REG_SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11125 ( .A1(n8692), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8690) );
  XNOR2_X1 U11126 ( .A(n8690), .B(n12094), .ZN(n12255) );
  NAND2_X1 U11127 ( .A1(n8691), .A2(n12255), .ZN(n8694) );
  OR2_X1 U11128 ( .A1(n8697), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U11129 ( .A1(n11325), .A2(n12255), .ZN(n8695) );
  INV_X1 U11130 ( .A(n8697), .ZN(n8699) );
  INV_X1 U11131 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U11132 ( .A1(n11325), .A2(n11130), .ZN(n8700) );
  NOR4_X1 U11133 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8710) );
  OR4_X1 U11134 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n8707) );
  NOR4_X1 U11135 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8705) );
  NOR4_X1 U11136 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8704) );
  NOR4_X1 U11137 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8703) );
  NOR4_X1 U11138 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8702) );
  NAND4_X1 U11139 ( .A1(n8705), .A2(n8704), .A3(n8703), .A4(n8702), .ZN(n8706)
         );
  NOR4_X1 U11140 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n8707), .A4(n8706), .ZN(n8709) );
  NOR4_X1 U11141 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8708) );
  AND3_X1 U11142 ( .A1(n8710), .A2(n8709), .A3(n8708), .ZN(n8711) );
  OR2_X1 U11143 ( .A1(n8697), .A2(n8711), .ZN(n8728) );
  NAND3_X1 U11144 ( .A1(n12820), .A2(n12822), .A3(n8728), .ZN(n9350) );
  NAND2_X1 U11145 ( .A1(n10500), .A2(n8736), .ZN(n8949) );
  OR2_X1 U11146 ( .A1(n8949), .A2(n8734), .ZN(n9351) );
  INV_X1 U11147 ( .A(n12820), .ZN(n8713) );
  INV_X1 U11148 ( .A(n12822), .ZN(n8712) );
  NAND3_X1 U11149 ( .A1(n8713), .A2(n8712), .A3(n8728), .ZN(n9366) );
  OAI22_X1 U11150 ( .A1(n9350), .A2(n9351), .B1(n9366), .B2(n8714), .ZN(n8722)
         );
  INV_X1 U11151 ( .A(n12255), .ZN(n8716) );
  INV_X1 U11152 ( .A(n11130), .ZN(n8715) );
  AND2_X1 U11153 ( .A1(n8716), .A2(n8715), .ZN(n8718) );
  NAND2_X1 U11154 ( .A1(n8718), .A2(n8717), .ZN(n9376) );
  NAND2_X1 U11155 ( .A1(n6599), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8719) );
  MUX2_X1 U11156 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8719), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8721) );
  NAND2_X1 U11157 ( .A1(n8721), .A2(n8720), .ZN(n9732) );
  NAND2_X1 U11158 ( .A1(n8722), .A2(n9731), .ZN(n8725) );
  INV_X1 U11159 ( .A(n9350), .ZN(n9346) );
  INV_X1 U11160 ( .A(n9731), .ZN(n8723) );
  OR2_X1 U11161 ( .A1(n8723), .A2(n9353), .ZN(n9361) );
  NOR2_X1 U11162 ( .A1(n9361), .A2(n9970), .ZN(n9358) );
  NAND2_X1 U11163 ( .A1(n9346), .A2(n9358), .ZN(n8724) );
  INV_X2 U11164 ( .A(n15127), .ZN(n15129) );
  INV_X1 U11165 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8742) );
  XNOR2_X1 U11166 ( .A(n12822), .B(n12820), .ZN(n8730) );
  NAND2_X1 U11167 ( .A1(n9731), .A2(n8728), .ZN(n8729) );
  NOR2_X1 U11168 ( .A1(n8730), .A2(n8729), .ZN(n9977) );
  NAND2_X1 U11169 ( .A1(n8732), .A2(n8731), .ZN(n8733) );
  NAND3_X1 U11170 ( .A1(n9353), .A2(n8734), .A3(n8733), .ZN(n8735) );
  AND2_X1 U11171 ( .A1(n8735), .A2(n9970), .ZN(n8738) );
  NAND3_X1 U11172 ( .A1(n12517), .A2(n8736), .A3(n10560), .ZN(n9971) );
  MUX2_X1 U11173 ( .A(n9353), .B(n9971), .S(n9970), .Z(n9969) );
  NAND2_X1 U11174 ( .A1(n12820), .A2(n9969), .ZN(n8737) );
  OAI21_X1 U11175 ( .B1(n12820), .B2(n8738), .A(n8737), .ZN(n8739) );
  INV_X1 U11176 ( .A(n8739), .ZN(n8740) );
  AND2_X2 U11177 ( .A1(n9977), .A2(n8740), .ZN(n15133) );
  INV_X1 U11178 ( .A(n12539), .ZN(n12246) );
  OR2_X1 U11179 ( .A1(n8767), .A2(n12246), .ZN(n8919) );
  INV_X1 U11180 ( .A(n8745), .ZN(n8746) );
  INV_X1 U11181 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12214) );
  XNOR2_X1 U11182 ( .A(n12214), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n8760) );
  INV_X1 U11183 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12234) );
  XNOR2_X1 U11184 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n8748) );
  XNOR2_X1 U11185 ( .A(n8749), .B(n8748), .ZN(n12823) );
  NAND2_X1 U11186 ( .A1(n12823), .A2(n8243), .ZN(n8751) );
  NAND2_X1 U11187 ( .A1(n8762), .A2(SI_31_), .ZN(n8750) );
  NAND2_X2 U11188 ( .A1(n8751), .A2(n8750), .ZN(n12773) );
  INV_X1 U11189 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U11190 ( .A1(n8513), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8755) );
  INV_X1 U11191 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n8752) );
  OR2_X1 U11192 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  OAI211_X1 U11193 ( .C1(n12528), .C2(n8756), .A(n8755), .B(n8754), .ZN(n8757)
         );
  INV_X1 U11194 ( .A(n8757), .ZN(n8758) );
  XNOR2_X1 U11195 ( .A(n8761), .B(n8760), .ZN(n12236) );
  NAND2_X1 U11196 ( .A1(n12236), .A2(n8243), .ZN(n8764) );
  NAND2_X1 U11197 ( .A1(n8762), .A2(SI_30_), .ZN(n8763) );
  NAND2_X2 U11198 ( .A1(n8764), .A2(n8763), .ZN(n14468) );
  NAND2_X1 U11199 ( .A1(n14468), .A2(n10826), .ZN(n8765) );
  NAND2_X1 U11200 ( .A1(n8766), .A2(n8765), .ZN(n8778) );
  INV_X1 U11201 ( .A(n14468), .ZN(n8768) );
  INV_X1 U11202 ( .A(n12525), .ZN(n12361) );
  NAND2_X1 U11203 ( .A1(n8767), .A2(n12246), .ZN(n8916) );
  OAI21_X1 U11204 ( .B1(n8768), .B2(n12361), .A(n8916), .ZN(n8769) );
  NOR2_X1 U11205 ( .A1(n8778), .A2(n8769), .ZN(n8773) );
  NOR2_X1 U11206 ( .A1(n14468), .A2(n10826), .ZN(n8942) );
  NAND2_X1 U11207 ( .A1(n8942), .A2(n12773), .ZN(n8770) );
  AOI21_X2 U11208 ( .B1(n8774), .B2(n8773), .A(n8772), .ZN(n8775) );
  XNOR2_X1 U11209 ( .A(n8775), .B(n8947), .ZN(n8777) );
  NOR2_X1 U11210 ( .A1(n8777), .A2(n8776), .ZN(n8952) );
  INV_X1 U11211 ( .A(n15109), .ZN(n10184) );
  INV_X1 U11212 ( .A(n9353), .ZN(n8923) );
  INV_X1 U11213 ( .A(n8778), .ZN(n8945) );
  INV_X1 U11214 ( .A(n12542), .ZN(n8914) );
  AND2_X2 U11215 ( .A1(n8902), .A2(n8903), .ZN(n12565) );
  NAND2_X1 U11216 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  NAND2_X1 U11217 ( .A1(n8781), .A2(n12579), .ZN(n8782) );
  INV_X1 U11218 ( .A(n8783), .ZN(n8887) );
  MUX2_X1 U11219 ( .A(n8785), .B(n8784), .S(n9970), .Z(n8886) );
  NAND2_X1 U11220 ( .A1(n12757), .A2(n12001), .ZN(n8925) );
  NAND2_X1 U11221 ( .A1(n8925), .A2(n10560), .ZN(n8788) );
  NAND2_X1 U11222 ( .A1(n8925), .A2(n9258), .ZN(n8786) );
  NAND3_X1 U11223 ( .A1(n9267), .A2(n8786), .A3(n9970), .ZN(n8787) );
  OAI21_X1 U11224 ( .B1(n12765), .B2(n8788), .A(n8787), .ZN(n8790) );
  NAND2_X1 U11225 ( .A1(n12764), .A2(n10500), .ZN(n8789) );
  NAND2_X1 U11226 ( .A1(n8790), .A2(n8789), .ZN(n8793) );
  MUX2_X1 U11227 ( .A(n9267), .B(n8791), .S(n9970), .Z(n8792) );
  NAND3_X1 U11228 ( .A1(n8793), .A2(n10179), .A3(n8792), .ZN(n8800) );
  NAND2_X1 U11229 ( .A1(n8802), .A2(n8794), .ZN(n8797) );
  NAND2_X1 U11230 ( .A1(n8801), .A2(n8795), .ZN(n8796) );
  MUX2_X1 U11231 ( .A(n8797), .B(n8796), .S(n9733), .Z(n8798) );
  INV_X1 U11232 ( .A(n8798), .ZN(n8799) );
  NAND2_X1 U11233 ( .A1(n8800), .A2(n8799), .ZN(n8804) );
  MUX2_X1 U11234 ( .A(n8802), .B(n8801), .S(n9970), .Z(n8803) );
  NAND3_X1 U11235 ( .A1(n8804), .A2(n10138), .A3(n8803), .ZN(n8808) );
  MUX2_X1 U11236 ( .A(n8806), .B(n8805), .S(n9733), .Z(n8807) );
  NAND3_X1 U11237 ( .A1(n8808), .A2(n10424), .A3(n8807), .ZN(n8815) );
  NAND2_X1 U11238 ( .A1(n8817), .A2(n8809), .ZN(n8812) );
  NAND2_X1 U11239 ( .A1(n8816), .A2(n8810), .ZN(n8811) );
  MUX2_X1 U11240 ( .A(n8812), .B(n8811), .S(n9970), .Z(n8813) );
  INV_X1 U11241 ( .A(n8813), .ZN(n8814) );
  NAND2_X1 U11242 ( .A1(n8815), .A2(n8814), .ZN(n8819) );
  MUX2_X1 U11243 ( .A(n8817), .B(n8816), .S(n9733), .Z(n8818) );
  NAND3_X1 U11244 ( .A1(n8819), .A2(n10812), .A3(n8818), .ZN(n8823) );
  MUX2_X1 U11245 ( .A(n8821), .B(n8820), .S(n9733), .Z(n8822) );
  NAND3_X1 U11246 ( .A1(n8823), .A2(n11039), .A3(n8822), .ZN(n8827) );
  INV_X1 U11247 ( .A(n11071), .ZN(n11068) );
  MUX2_X1 U11248 ( .A(n8825), .B(n8824), .S(n9733), .Z(n8826) );
  NAND3_X1 U11249 ( .A1(n8827), .A2(n11068), .A3(n8826), .ZN(n8831) );
  MUX2_X1 U11250 ( .A(n8829), .B(n8828), .S(n9733), .Z(n8830) );
  NAND2_X1 U11251 ( .A1(n8831), .A2(n8830), .ZN(n8836) );
  INV_X1 U11252 ( .A(n11190), .ZN(n11194) );
  MUX2_X1 U11253 ( .A(n8833), .B(n8832), .S(n9733), .Z(n8834) );
  NAND2_X1 U11254 ( .A1(n8834), .A2(n11407), .ZN(n8835) );
  AOI21_X1 U11255 ( .B1(n8836), .B2(n11194), .A(n8835), .ZN(n8846) );
  NAND2_X1 U11256 ( .A1(n8843), .A2(n8837), .ZN(n8840) );
  NAND2_X1 U11257 ( .A1(n8842), .A2(n8838), .ZN(n8839) );
  MUX2_X1 U11258 ( .A(n8840), .B(n8839), .S(n9733), .Z(n8845) );
  INV_X1 U11259 ( .A(n8841), .ZN(n11489) );
  MUX2_X1 U11260 ( .A(n8843), .B(n8842), .S(n9970), .Z(n8844) );
  OAI211_X1 U11261 ( .C1(n8846), .C2(n8845), .A(n11489), .B(n8844), .ZN(n8850)
         );
  MUX2_X1 U11262 ( .A(n8848), .B(n8847), .S(n9970), .Z(n8849) );
  NAND2_X1 U11263 ( .A1(n8850), .A2(n8849), .ZN(n8851) );
  NAND2_X1 U11264 ( .A1(n8851), .A2(n11446), .ZN(n8855) );
  MUX2_X1 U11265 ( .A(n8853), .B(n8852), .S(n9733), .Z(n8854) );
  NAND3_X1 U11266 ( .A1(n8855), .A2(n11665), .A3(n8854), .ZN(n8861) );
  AND2_X1 U11267 ( .A1(n8863), .A2(n8856), .ZN(n8859) );
  OR2_X1 U11268 ( .A1(n12747), .A2(n12682), .ZN(n8862) );
  AND2_X1 U11269 ( .A1(n8862), .A2(n8857), .ZN(n8858) );
  MUX2_X1 U11270 ( .A(n8859), .B(n8858), .S(n9970), .Z(n8860) );
  NAND2_X1 U11271 ( .A1(n8861), .A2(n8860), .ZN(n8866) );
  MUX2_X1 U11272 ( .A(n8863), .B(n8862), .S(n9733), .Z(n8865) );
  NAND2_X1 U11273 ( .A1(n8933), .A2(n12685), .ZN(n8864) );
  AOI21_X1 U11274 ( .B1(n8866), .B2(n8865), .A(n8864), .ZN(n8880) );
  INV_X1 U11275 ( .A(n8872), .ZN(n8869) );
  OAI211_X1 U11276 ( .C1(n8869), .C2(n8868), .A(n8877), .B(n8867), .ZN(n8875)
         );
  INV_X1 U11277 ( .A(n8870), .ZN(n8871) );
  NAND2_X1 U11278 ( .A1(n8933), .A2(n8871), .ZN(n8873) );
  NAND3_X1 U11279 ( .A1(n8876), .A2(n8873), .A3(n8872), .ZN(n8874) );
  MUX2_X1 U11280 ( .A(n8875), .B(n8874), .S(n9970), .Z(n8879) );
  MUX2_X1 U11281 ( .A(n8877), .B(n8876), .S(n9733), .Z(n8878) );
  OAI21_X1 U11282 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8884) );
  MUX2_X1 U11283 ( .A(n8882), .B(n8881), .S(n9733), .Z(n8883) );
  OAI211_X1 U11284 ( .C1(n12645), .C2(n8884), .A(n12629), .B(n8883), .ZN(n8885) );
  NAND3_X1 U11285 ( .A1(n12619), .A2(n8886), .A3(n8885), .ZN(n8890) );
  MUX2_X1 U11286 ( .A(n8888), .B(n8887), .S(n9970), .Z(n8889) );
  NAND3_X1 U11287 ( .A1(n8891), .A2(n8890), .A3(n8889), .ZN(n8893) );
  NAND3_X1 U11288 ( .A1(n12610), .A2(n12618), .A3(n9733), .ZN(n8892) );
  NAND2_X1 U11289 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  NAND2_X1 U11290 ( .A1(n12592), .A2(n8894), .ZN(n8895) );
  NAND2_X1 U11291 ( .A1(n8896), .A2(n8895), .ZN(n8900) );
  OR2_X1 U11292 ( .A1(n12709), .A2(n12594), .ZN(n8898) );
  MUX2_X1 U11293 ( .A(n8898), .B(n8897), .S(n9970), .Z(n8899) );
  OAI21_X1 U11294 ( .B1(n8900), .B2(n12580), .A(n8899), .ZN(n8901) );
  AND2_X1 U11295 ( .A1(n8905), .A2(n8904), .ZN(n8906) );
  OAI21_X1 U11296 ( .B1(n12564), .B2(n12701), .A(n8912), .ZN(n8907) );
  NAND3_X1 U11297 ( .A1(n8909), .A2(n9733), .A3(n8908), .ZN(n8910) );
  INV_X1 U11298 ( .A(n8912), .ZN(n8913) );
  NAND3_X1 U11299 ( .A1(n8914), .A2(n9733), .A3(n8913), .ZN(n8915) );
  NAND3_X1 U11300 ( .A1(n8917), .A2(n8916), .A3(n8915), .ZN(n8920) );
  INV_X1 U11301 ( .A(n8942), .ZN(n8918) );
  NAND3_X1 U11302 ( .A1(n8920), .A2(n8919), .A3(n8918), .ZN(n8921) );
  INV_X1 U11303 ( .A(n12619), .ZN(n8937) );
  NOR2_X1 U11304 ( .A1(n10815), .A2(n10186), .ZN(n8924) );
  NAND4_X1 U11305 ( .A1(n8924), .A2(n10138), .A3(n10424), .A4(n11039), .ZN(
        n8928) );
  INV_X1 U11306 ( .A(n8925), .ZN(n8926) );
  NOR2_X1 U11307 ( .A1(n12764), .A2(n8926), .ZN(n10116) );
  INV_X1 U11308 ( .A(n12765), .ZN(n10030) );
  NAND4_X1 U11309 ( .A1(n10116), .A2(n10084), .A3(n10565), .A4(n10030), .ZN(
        n8927) );
  NOR2_X1 U11310 ( .A1(n8928), .A2(n8927), .ZN(n8929) );
  NAND4_X1 U11311 ( .A1(n8929), .A2(n11407), .A3(n11194), .A4(n11068), .ZN(
        n8930) );
  NOR2_X1 U11312 ( .A1(n8930), .A2(n7043), .ZN(n8931) );
  AND4_X1 U11313 ( .A1(n11665), .A2(n11446), .A3(n11489), .A4(n8931), .ZN(
        n8932) );
  NAND4_X1 U11314 ( .A1(n8933), .A2(n12685), .A3(n8932), .A4(n11604), .ZN(
        n8934) );
  NOR2_X1 U11315 ( .A1(n12658), .A2(n8934), .ZN(n8935) );
  NAND3_X1 U11316 ( .A1(n12629), .A2(n7187), .A3(n8935), .ZN(n8936) );
  NOR4_X1 U11317 ( .A1(n8938), .A2(n12608), .A3(n8937), .A4(n8936), .ZN(n8940)
         );
  NAND3_X1 U11318 ( .A1(n12565), .A2(n8940), .A3(n8939), .ZN(n8941) );
  NOR4_X1 U11319 ( .A1(n8942), .A2(n12550), .A3(n12542), .A4(n8941), .ZN(n8946) );
  NAND4_X1 U11320 ( .A1(n8945), .A2(n8946), .A3(n8944), .A4(n8771), .ZN(n8948)
         );
  XNOR2_X1 U11321 ( .A(n8948), .B(n8947), .ZN(n8950) );
  INV_X1 U11322 ( .A(n8949), .ZN(n9257) );
  NOR2_X1 U11323 ( .A1(n9732), .A2(P3_U3151), .ZN(n9730) );
  INV_X1 U11324 ( .A(n9730), .ZN(n10828) );
  INV_X1 U11325 ( .A(n9361), .ZN(n9364) );
  NAND3_X1 U11326 ( .A1(n9364), .A2(n12756), .A3(n6622), .ZN(n8953) );
  OAI211_X1 U11327 ( .C1(n10560), .C2(n10828), .A(n8953), .B(P3_B_REG_SCAN_IN), 
        .ZN(n8954) );
  NAND2_X1 U11328 ( .A1(n8955), .A2(n8954), .ZN(P3_U3296) );
  NAND2_X1 U11329 ( .A1(n8959), .A2(n8958), .ZN(n8961) );
  NAND2_X1 U11330 ( .A1(n8960), .A2(n8981), .ZN(n8963) );
  NAND2_X1 U11331 ( .A1(n8961), .A2(n8963), .ZN(n8965) );
  AOI21_X1 U11332 ( .B1(n6463), .B2(n11369), .A(n10120), .ZN(n8962) );
  OAI21_X1 U11333 ( .B1(n8963), .B2(n10165), .A(n8962), .ZN(n8964) );
  NAND2_X1 U11334 ( .A1(n8965), .A2(n8964), .ZN(n8970) );
  NAND2_X1 U11335 ( .A1(n9126), .A2(n10121), .ZN(n8966) );
  NAND2_X1 U11336 ( .A1(n8967), .A2(n8966), .ZN(n8968) );
  NAND2_X1 U11337 ( .A1(n8970), .A2(n8969), .ZN(n8971) );
  NAND2_X1 U11338 ( .A1(n8973), .A2(n6462), .ZN(n8975) );
  NAND2_X1 U11339 ( .A1(n9204), .A2(n10321), .ZN(n8974) );
  NAND2_X1 U11340 ( .A1(n8975), .A2(n8974), .ZN(n8978) );
  AOI22_X1 U11341 ( .A1(n8973), .A2(n9126), .B1(n6461), .B2(n10321), .ZN(n8976) );
  INV_X1 U11342 ( .A(n8977), .ZN(n8980) );
  NAND2_X1 U11343 ( .A1(n8980), .A2(n7430), .ZN(n8987) );
  NAND2_X1 U11344 ( .A1(n13047), .A2(n9204), .ZN(n8983) );
  NAND2_X1 U11345 ( .A1(n6461), .A2(n14939), .ZN(n8982) );
  NAND2_X1 U11346 ( .A1(n8983), .A2(n8982), .ZN(n8986) );
  AOI22_X1 U11347 ( .A1(n13047), .A2(n6462), .B1(n9204), .B2(n14939), .ZN(
        n8984) );
  AOI21_X1 U11348 ( .B1(n8987), .B2(n8986), .A(n8984), .ZN(n8985) );
  NAND2_X1 U11349 ( .A1(n13046), .A2(n6461), .ZN(n8989) );
  NAND2_X1 U11350 ( .A1(n9192), .A2(n10743), .ZN(n8988) );
  NAND2_X1 U11351 ( .A1(n8989), .A2(n8988), .ZN(n8995) );
  NAND2_X1 U11352 ( .A1(n13046), .A2(n9204), .ZN(n8991) );
  NAND2_X1 U11353 ( .A1(n6461), .A2(n10743), .ZN(n8990) );
  NAND2_X1 U11354 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  NAND2_X1 U11355 ( .A1(n8993), .A2(n8992), .ZN(n8999) );
  INV_X1 U11356 ( .A(n8994), .ZN(n8997) );
  INV_X1 U11357 ( .A(n8995), .ZN(n8996) );
  NAND2_X1 U11358 ( .A1(n8997), .A2(n8996), .ZN(n8998) );
  NAND2_X1 U11359 ( .A1(n13045), .A2(n9204), .ZN(n9001) );
  NAND2_X1 U11360 ( .A1(n6462), .A2(n10831), .ZN(n9000) );
  AOI22_X1 U11361 ( .A1(n13045), .A2(n6461), .B1(n9192), .B2(n10831), .ZN(
        n9002) );
  NAND2_X1 U11362 ( .A1(n13044), .A2(n6462), .ZN(n9005) );
  NAND2_X1 U11363 ( .A1(n9192), .A2(n10855), .ZN(n9004) );
  NAND2_X1 U11364 ( .A1(n9005), .A2(n9004), .ZN(n9011) );
  NAND2_X1 U11365 ( .A1(n13044), .A2(n9204), .ZN(n9007) );
  NAND2_X1 U11366 ( .A1(n6462), .A2(n10855), .ZN(n9006) );
  NAND2_X1 U11367 ( .A1(n9007), .A2(n9006), .ZN(n9008) );
  NAND2_X1 U11368 ( .A1(n9009), .A2(n9008), .ZN(n9013) );
  NAND2_X1 U11369 ( .A1(n13043), .A2(n9204), .ZN(n9015) );
  NAND2_X1 U11370 ( .A1(n6461), .A2(n10954), .ZN(n9014) );
  NAND2_X1 U11371 ( .A1(n9015), .A2(n9014), .ZN(n9017) );
  AOI22_X1 U11372 ( .A1(n13043), .A2(n6462), .B1(n9204), .B2(n10954), .ZN(
        n9016) );
  NAND2_X1 U11373 ( .A1(n13042), .A2(n6461), .ZN(n9019) );
  NAND2_X1 U11374 ( .A1(n11173), .A2(n9204), .ZN(n9018) );
  NAND2_X1 U11375 ( .A1(n9019), .A2(n9018), .ZN(n9025) );
  NAND2_X1 U11376 ( .A1(n9024), .A2(n9025), .ZN(n9023) );
  NAND2_X1 U11377 ( .A1(n13042), .A2(n9204), .ZN(n9021) );
  NAND2_X1 U11378 ( .A1(n11173), .A2(n6462), .ZN(n9020) );
  NAND2_X1 U11379 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  NAND2_X1 U11380 ( .A1(n9023), .A2(n9022), .ZN(n9029) );
  NAND2_X1 U11381 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  NAND2_X1 U11382 ( .A1(n11316), .A2(n6462), .ZN(n9031) );
  NAND2_X1 U11383 ( .A1(n13041), .A2(n9204), .ZN(n9030) );
  AOI22_X1 U11384 ( .A1(n11316), .A2(n9204), .B1(n6461), .B2(n13041), .ZN(
        n9032) );
  NAND2_X1 U11385 ( .A1(n11308), .A2(n9204), .ZN(n9034) );
  NAND2_X1 U11386 ( .A1(n13040), .A2(n6462), .ZN(n9033) );
  NAND2_X1 U11387 ( .A1(n9034), .A2(n9033), .ZN(n9037) );
  AOI22_X1 U11388 ( .A1(n11308), .A2(n6461), .B1(n9192), .B2(n13040), .ZN(
        n9035) );
  INV_X1 U11389 ( .A(n9036), .ZN(n9039) );
  NAND2_X1 U11390 ( .A1(n11467), .A2(n6462), .ZN(n9041) );
  NAND2_X1 U11391 ( .A1(n13039), .A2(n9204), .ZN(n9040) );
  NAND2_X1 U11392 ( .A1(n9041), .A2(n9040), .ZN(n9043) );
  INV_X1 U11393 ( .A(n9043), .ZN(n9042) );
  NAND2_X1 U11394 ( .A1(n11467), .A2(n9204), .ZN(n9045) );
  NAND2_X1 U11395 ( .A1(n13039), .A2(n6461), .ZN(n9044) );
  NAND2_X1 U11396 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U11397 ( .A1(n11565), .A2(n9204), .ZN(n9048) );
  NAND2_X1 U11398 ( .A1(n13038), .A2(n6461), .ZN(n9047) );
  NAND2_X1 U11399 ( .A1(n9048), .A2(n9047), .ZN(n9051) );
  AOI22_X1 U11400 ( .A1(n11565), .A2(n6462), .B1(n9204), .B2(n13038), .ZN(
        n9049) );
  INV_X1 U11401 ( .A(n9050), .ZN(n9053) );
  NAND2_X1 U11402 ( .A1(n9053), .A2(n7419), .ZN(n9058) );
  NAND2_X1 U11403 ( .A1(n14527), .A2(n6461), .ZN(n9055) );
  NAND2_X1 U11404 ( .A1(n14483), .A2(n9204), .ZN(n9054) );
  NAND2_X1 U11405 ( .A1(n14527), .A2(n9204), .ZN(n9057) );
  NAND2_X1 U11406 ( .A1(n14483), .A2(n6462), .ZN(n9056) );
  NAND2_X1 U11407 ( .A1(n14503), .A2(n9192), .ZN(n9060) );
  NAND2_X1 U11408 ( .A1(n13037), .A2(n6461), .ZN(n9059) );
  AOI22_X1 U11409 ( .A1(n14503), .A2(n6462), .B1(n9204), .B2(n13037), .ZN(
        n9061) );
  NAND2_X1 U11410 ( .A1(n11767), .A2(n6461), .ZN(n9063) );
  NAND2_X1 U11411 ( .A1(n14482), .A2(n9192), .ZN(n9062) );
  NAND2_X1 U11412 ( .A1(n9063), .A2(n9062), .ZN(n9068) );
  AND2_X1 U11413 ( .A1(n13036), .A2(n6462), .ZN(n9064) );
  AOI21_X1 U11414 ( .B1(n13399), .B2(n9126), .A(n9064), .ZN(n9073) );
  NAND2_X1 U11415 ( .A1(n13399), .A2(n6461), .ZN(n9066) );
  NAND2_X1 U11416 ( .A1(n13036), .A2(n9192), .ZN(n9065) );
  NAND2_X1 U11417 ( .A1(n9066), .A2(n9065), .ZN(n9072) );
  AOI22_X1 U11418 ( .A1(n11767), .A2(n9204), .B1(n6462), .B2(n14482), .ZN(
        n9067) );
  AOI21_X1 U11419 ( .B1(n9069), .B2(n9068), .A(n9067), .ZN(n9076) );
  AOI22_X1 U11420 ( .A1(n13439), .A2(n9126), .B1(n6462), .B2(n13035), .ZN(
        n9074) );
  NAND2_X1 U11421 ( .A1(n13439), .A2(n6462), .ZN(n9071) );
  NAND2_X1 U11422 ( .A1(n13035), .A2(n9192), .ZN(n9070) );
  NAND2_X1 U11423 ( .A1(n9071), .A2(n9070), .ZN(n9078) );
  AOI22_X1 U11424 ( .A1(n9074), .A2(n9078), .B1(n9073), .B2(n9072), .ZN(n9075)
         );
  INV_X1 U11425 ( .A(n9078), .ZN(n9079) );
  NAND2_X1 U11426 ( .A1(n9079), .A2(n9221), .ZN(n9080) );
  NAND2_X1 U11427 ( .A1(n13435), .A2(n9192), .ZN(n9083) );
  NAND2_X1 U11428 ( .A1(n13034), .A2(n6462), .ZN(n9082) );
  NAND2_X1 U11429 ( .A1(n9083), .A2(n9082), .ZN(n9085) );
  INV_X1 U11430 ( .A(n9085), .ZN(n9084) );
  AOI22_X1 U11431 ( .A1(n13435), .A2(n6461), .B1(n9192), .B2(n13034), .ZN(
        n9086) );
  NAND2_X1 U11432 ( .A1(n13277), .A2(n6461), .ZN(n9090) );
  NAND2_X1 U11433 ( .A1(n13033), .A2(n9192), .ZN(n9089) );
  NAND2_X1 U11434 ( .A1(n9090), .A2(n9089), .ZN(n9092) );
  AOI22_X1 U11435 ( .A1(n13277), .A2(n9126), .B1(n6462), .B2(n13033), .ZN(
        n9091) );
  AOI21_X1 U11436 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9095) );
  NOR2_X1 U11437 ( .A1(n9093), .A2(n9092), .ZN(n9094) );
  NAND2_X1 U11438 ( .A1(n13367), .A2(n9192), .ZN(n9097) );
  NAND2_X1 U11439 ( .A1(n13032), .A2(n6462), .ZN(n9096) );
  NAND2_X1 U11440 ( .A1(n9097), .A2(n9096), .ZN(n9099) );
  AOI22_X1 U11441 ( .A1(n13367), .A2(n6461), .B1(n9204), .B2(n13032), .ZN(
        n9098) );
  NAND2_X1 U11442 ( .A1(n13425), .A2(n6461), .ZN(n9101) );
  NAND2_X1 U11443 ( .A1(n13031), .A2(n9192), .ZN(n9100) );
  NAND2_X1 U11444 ( .A1(n9101), .A2(n9100), .ZN(n9103) );
  AOI22_X1 U11445 ( .A1(n13425), .A2(n9126), .B1(n6462), .B2(n13031), .ZN(
        n9102) );
  NAND2_X1 U11446 ( .A1(n13421), .A2(n9192), .ZN(n9106) );
  NAND2_X1 U11447 ( .A1(n13030), .A2(n6462), .ZN(n9105) );
  NAND2_X1 U11448 ( .A1(n9106), .A2(n9105), .ZN(n9108) );
  AOI22_X1 U11449 ( .A1(n13421), .A2(n6461), .B1(n9204), .B2(n13030), .ZN(
        n9107) );
  NOR2_X1 U11450 ( .A1(n9109), .A2(n9108), .ZN(n9113) );
  AND2_X1 U11451 ( .A1(n13029), .A2(n6461), .ZN(n9110) );
  AOI21_X1 U11452 ( .B1(n13345), .B2(n9126), .A(n9110), .ZN(n9130) );
  NAND2_X1 U11453 ( .A1(n13345), .A2(n6461), .ZN(n9112) );
  NAND2_X1 U11454 ( .A1(n13029), .A2(n9192), .ZN(n9111) );
  NAND2_X1 U11455 ( .A1(n9112), .A2(n9111), .ZN(n9129) );
  OAI22_X1 U11456 ( .A1(n9114), .A2(n9113), .B1(n9130), .B2(n9129), .ZN(n9115)
         );
  AND2_X1 U11457 ( .A1(n13025), .A2(n6462), .ZN(n9116) );
  AOI21_X1 U11458 ( .B1(n13320), .B2(n9126), .A(n9116), .ZN(n9174) );
  NAND2_X1 U11459 ( .A1(n13320), .A2(n6462), .ZN(n9118) );
  NAND2_X1 U11460 ( .A1(n13025), .A2(n9192), .ZN(n9117) );
  NAND2_X1 U11461 ( .A1(n9118), .A2(n9117), .ZN(n9173) );
  NAND2_X1 U11462 ( .A1(n9174), .A2(n9173), .ZN(n9179) );
  AND2_X1 U11463 ( .A1(n13026), .A2(n6462), .ZN(n9119) );
  AOI21_X1 U11464 ( .B1(n13176), .B2(n9126), .A(n9119), .ZN(n9168) );
  NAND2_X1 U11465 ( .A1(n13176), .A2(n6461), .ZN(n9121) );
  NAND2_X1 U11466 ( .A1(n13026), .A2(n9192), .ZN(n9120) );
  NAND2_X1 U11467 ( .A1(n9121), .A2(n9120), .ZN(n9165) );
  AND2_X1 U11468 ( .A1(n13027), .A2(n6461), .ZN(n9122) );
  AOI21_X1 U11469 ( .B1(n13193), .B2(n9204), .A(n9122), .ZN(n9160) );
  NAND2_X1 U11470 ( .A1(n13193), .A2(n6461), .ZN(n9124) );
  NAND2_X1 U11471 ( .A1(n13027), .A2(n9192), .ZN(n9123) );
  NAND2_X1 U11472 ( .A1(n9160), .A2(n9164), .ZN(n9132) );
  AND2_X1 U11473 ( .A1(n13028), .A2(n6461), .ZN(n9125) );
  AOI21_X1 U11474 ( .B1(n13339), .B2(n9126), .A(n9125), .ZN(n9157) );
  NAND2_X1 U11475 ( .A1(n13339), .A2(n6462), .ZN(n9128) );
  NAND2_X1 U11476 ( .A1(n13028), .A2(n9192), .ZN(n9127) );
  NAND2_X1 U11477 ( .A1(n9128), .A2(n9127), .ZN(n9156) );
  AOI22_X1 U11478 ( .A1(n9157), .A2(n9156), .B1(n9130), .B2(n9129), .ZN(n9131)
         );
  NAND2_X1 U11479 ( .A1(n9132), .A2(n9131), .ZN(n9133) );
  AOI21_X1 U11480 ( .B1(n9168), .B2(n9165), .A(n9133), .ZN(n9134) );
  INV_X1 U11481 ( .A(SI_29_), .ZN(n12005) );
  NAND2_X1 U11482 ( .A1(n9137), .A2(n12005), .ZN(n9138) );
  MUX2_X1 U11483 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9139), .Z(n9140) );
  NAND2_X1 U11484 ( .A1(n9140), .A2(SI_30_), .ZN(n9141) );
  OAI21_X1 U11485 ( .B1(n9140), .B2(SI_30_), .A(n9141), .ZN(n9187) );
  MUX2_X1 U11486 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9139), .Z(n9142) );
  XNOR2_X1 U11487 ( .A(n9142), .B(SI_31_), .ZN(n9143) );
  NAND2_X1 U11488 ( .A1(n13757), .A2(n7612), .ZN(n9147) );
  INV_X1 U11489 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9145) );
  OR2_X1 U11490 ( .A1(n7919), .A2(n9145), .ZN(n9146) );
  INV_X1 U11491 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U11492 ( .A1(n7506), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U11493 ( .A1(n9148), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9149) );
  OAI211_X1 U11494 ( .C1(n9152), .C2(n9151), .A(n9150), .B(n9149), .ZN(n13021)
         );
  AND2_X1 U11495 ( .A1(n13023), .A2(n9192), .ZN(n9153) );
  AOI21_X1 U11496 ( .B1(n13313), .B2(n6461), .A(n9153), .ZN(n9199) );
  NAND2_X1 U11497 ( .A1(n13313), .A2(n9192), .ZN(n9155) );
  NAND2_X1 U11498 ( .A1(n13023), .A2(n6462), .ZN(n9154) );
  INV_X1 U11499 ( .A(n9156), .ZN(n9159) );
  INV_X1 U11500 ( .A(n9157), .ZN(n9158) );
  NAND2_X1 U11501 ( .A1(n9159), .A2(n9158), .ZN(n9163) );
  NAND2_X1 U11502 ( .A1(n9164), .A2(n9163), .ZN(n9162) );
  INV_X1 U11503 ( .A(n9160), .ZN(n9161) );
  OR2_X1 U11504 ( .A1(n9164), .A2(n9163), .ZN(n9166) );
  NAND3_X1 U11505 ( .A1(n9168), .A2(n9167), .A3(n9166), .ZN(n9172) );
  INV_X1 U11506 ( .A(n9165), .ZN(n9171) );
  NAND2_X1 U11507 ( .A1(n9167), .A2(n9166), .ZN(n9170) );
  INV_X1 U11508 ( .A(n9168), .ZN(n9169) );
  AND2_X1 U11509 ( .A1(n13024), .A2(n9192), .ZN(n9175) );
  AOI21_X1 U11510 ( .B1(n12924), .B2(n6461), .A(n9175), .ZN(n9182) );
  NAND2_X1 U11511 ( .A1(n12924), .A2(n9192), .ZN(n9177) );
  NAND2_X1 U11512 ( .A1(n13024), .A2(n6462), .ZN(n9176) );
  NAND2_X1 U11513 ( .A1(n9177), .A2(n9176), .ZN(n9181) );
  AOI22_X1 U11514 ( .A1(n9179), .A2(n9178), .B1(n9182), .B2(n9181), .ZN(n9180)
         );
  INV_X1 U11515 ( .A(n9181), .ZN(n9185) );
  INV_X1 U11516 ( .A(n9182), .ZN(n9183) );
  NAND2_X1 U11517 ( .A1(n13021), .A2(n6461), .ZN(n9186) );
  OR2_X1 U11518 ( .A1(n7919), .A2(n12214), .ZN(n9190) );
  AND2_X1 U11519 ( .A1(n9249), .A2(n9897), .ZN(n9191) );
  OR2_X1 U11520 ( .A1(n8054), .A2(n11369), .ZN(n9211) );
  AND2_X1 U11521 ( .A1(n9191), .A2(n9211), .ZN(n9194) );
  NAND2_X1 U11522 ( .A1(n13021), .A2(n9192), .ZN(n9205) );
  AOI21_X1 U11523 ( .B1(n9194), .B2(n9205), .A(n9193), .ZN(n9195) );
  AOI21_X1 U11524 ( .B1(n13408), .B2(n6461), .A(n9195), .ZN(n9202) );
  NAND2_X1 U11525 ( .A1(n13408), .A2(n9192), .ZN(n9197) );
  NAND2_X1 U11526 ( .A1(n13022), .A2(n6462), .ZN(n9196) );
  NAND2_X1 U11527 ( .A1(n9202), .A2(n9201), .ZN(n9209) );
  AND2_X1 U11528 ( .A1(n6461), .A2(n13021), .ZN(n9207) );
  AND2_X1 U11529 ( .A1(n9205), .A2(n9204), .ZN(n9206) );
  MUX2_X1 U11530 ( .A(n9207), .B(n9206), .S(n13138), .Z(n9208) );
  AOI21_X2 U11531 ( .B1(n9210), .B2(n9209), .A(n9208), .ZN(n9250) );
  OAI21_X1 U11532 ( .B1(n9212), .B2(n10984), .A(n9211), .ZN(n9213) );
  INV_X1 U11533 ( .A(n10120), .ZN(n9214) );
  NAND2_X1 U11534 ( .A1(n11369), .A2(n9214), .ZN(n9215) );
  OAI211_X1 U11535 ( .C1(n6463), .C2(n11187), .A(n9897), .B(n9215), .ZN(n9216)
         );
  NAND2_X1 U11536 ( .A1(n9250), .A2(n9216), .ZN(n9217) );
  OAI21_X1 U11537 ( .B1(n9250), .B2(n9218), .A(n9217), .ZN(n9252) );
  XNOR2_X1 U11538 ( .A(n13408), .B(n13022), .ZN(n9246) );
  XNOR2_X1 U11539 ( .A(n13367), .B(n9219), .ZN(n13270) );
  XNOR2_X1 U11540 ( .A(n13277), .B(n13033), .ZN(n13278) );
  AND2_X1 U11541 ( .A1(n9221), .A2(n9220), .ZN(n11741) );
  OR2_X1 U11542 ( .A1(n8960), .A2(n10165), .ZN(n9222) );
  NAND2_X1 U11543 ( .A1(n10158), .A2(n9222), .ZN(n10444) );
  AND2_X1 U11544 ( .A1(n10444), .A2(n9223), .ZN(n9226) );
  NAND4_X1 U11545 ( .A1(n9226), .A2(n9225), .A3(n10162), .A4(n9224), .ZN(n9227) );
  NOR2_X1 U11546 ( .A1(n9227), .A2(n10668), .ZN(n9230) );
  NAND4_X1 U11547 ( .A1(n9230), .A2(n9229), .A3(n10648), .A4(n9228), .ZN(n9231) );
  NOR4_X1 U11548 ( .A1(n11254), .A2(n11156), .A3(n9231), .A4(n10970), .ZN(
        n9235) );
  AND2_X1 U11549 ( .A1(n9233), .A2(n9232), .ZN(n11473) );
  NAND4_X1 U11550 ( .A1(n9235), .A2(n11473), .A3(n9234), .A4(n11241), .ZN(
        n9236) );
  NOR4_X1 U11551 ( .A1(n11741), .A2(n9237), .A3(n14505), .A4(n9236), .ZN(n9239) );
  NAND4_X1 U11552 ( .A1(n13278), .A2(n9239), .A3(n9238), .A4(n11691), .ZN(
        n9240) );
  NOR4_X1 U11553 ( .A1(n13228), .A2(n13255), .A3(n13270), .A4(n9240), .ZN(
        n9241) );
  NAND4_X1 U11554 ( .A1(n13186), .A2(n9241), .A3(n13197), .A4(n13223), .ZN(
        n9242) );
  NOR4_X1 U11555 ( .A1(n9243), .A2(n13158), .A3(n13173), .A4(n9242), .ZN(n9245) );
  OR2_X1 U11556 ( .A1(n9801), .A2(P2_U3088), .ZN(n11418) );
  NOR4_X1 U11557 ( .A1(n14961), .A2(n9897), .A3(n13455), .A4(n12900), .ZN(
        n9255) );
  OAI21_X1 U11558 ( .B1(n11418), .B2(n9253), .A(P2_B_REG_SCAN_IN), .ZN(n9254)
         );
  NAND2_X1 U11559 ( .A1(n9258), .A2(n10371), .ZN(n9259) );
  XNOR2_X1 U11560 ( .A(n11666), .B(n12240), .ZN(n9301) );
  INV_X4 U11561 ( .A(n9261), .ZN(n9302) );
  XNOR2_X1 U11562 ( .A(n9302), .B(n11083), .ZN(n9288) );
  INV_X1 U11563 ( .A(n9288), .ZN(n9289) );
  XNOR2_X1 U11564 ( .A(n9302), .B(n11094), .ZN(n9286) );
  INV_X1 U11565 ( .A(n9286), .ZN(n9287) );
  XNOR2_X1 U11566 ( .A(n9302), .B(n10777), .ZN(n9281) );
  INV_X1 U11567 ( .A(n9281), .ZN(n9282) );
  NAND2_X1 U11568 ( .A1(n9262), .A2(n9302), .ZN(n9264) );
  INV_X1 U11569 ( .A(n9263), .ZN(n10034) );
  INV_X1 U11570 ( .A(n9265), .ZN(n12384) );
  OAI21_X1 U11571 ( .B1(n9283), .B2(n12384), .A(n9267), .ZN(n9269) );
  NAND2_X1 U11572 ( .A1(n9269), .A2(n9268), .ZN(n9272) );
  INV_X1 U11573 ( .A(n9272), .ZN(n9273) );
  NOR2_X1 U11574 ( .A1(n10031), .A2(n9273), .ZN(n10075) );
  XNOR2_X1 U11575 ( .A(n9302), .B(n10078), .ZN(n9274) );
  XNOR2_X1 U11576 ( .A(n9274), .B(n12383), .ZN(n10076) );
  XNOR2_X1 U11577 ( .A(n9302), .B(n10091), .ZN(n9275) );
  XNOR2_X1 U11578 ( .A(n9275), .B(n10466), .ZN(n10382) );
  INV_X1 U11579 ( .A(n9275), .ZN(n9276) );
  XNOR2_X1 U11580 ( .A(n9302), .B(n10199), .ZN(n9277) );
  XNOR2_X1 U11581 ( .A(n9277), .B(n12381), .ZN(n10463) );
  XNOR2_X1 U11582 ( .A(n9302), .B(n10639), .ZN(n9279) );
  XNOR2_X1 U11583 ( .A(n9279), .B(n10776), .ZN(n10635) );
  INV_X1 U11584 ( .A(n9279), .ZN(n9280) );
  XNOR2_X1 U11585 ( .A(n9281), .B(n10862), .ZN(n10774) );
  NAND2_X1 U11586 ( .A1(n10775), .A2(n10774), .ZN(n10773) );
  OAI21_X1 U11587 ( .B1(n10862), .B2(n9282), .A(n10773), .ZN(n10861) );
  XNOR2_X1 U11588 ( .A(n9261), .B(n10815), .ZN(n10860) );
  INV_X1 U11589 ( .A(n10860), .ZN(n9284) );
  NAND2_X1 U11590 ( .A1(n9284), .A2(n12378), .ZN(n9285) );
  XNOR2_X1 U11591 ( .A(n9286), .B(n11205), .ZN(n10958) );
  NAND2_X1 U11592 ( .A1(n10959), .A2(n10958), .ZN(n10957) );
  OAI21_X1 U11593 ( .B1(n11205), .B2(n9287), .A(n10957), .ZN(n11203) );
  XNOR2_X1 U11594 ( .A(n9288), .B(n11341), .ZN(n11204) );
  OAI21_X1 U11595 ( .B1(n9289), .B2(n12376), .A(n11201), .ZN(n11338) );
  XNOR2_X1 U11596 ( .A(n9302), .B(n11367), .ZN(n9290) );
  XNOR2_X1 U11597 ( .A(n9290), .B(n12375), .ZN(n11337) );
  NAND2_X1 U11598 ( .A1(n9290), .A2(n12375), .ZN(n9291) );
  XNOR2_X1 U11599 ( .A(n9302), .B(n11560), .ZN(n11637) );
  INV_X1 U11600 ( .A(n11637), .ZN(n9292) );
  XNOR2_X1 U11601 ( .A(n9302), .B(n14471), .ZN(n11639) );
  NAND2_X1 U11602 ( .A1(n11639), .A2(n12373), .ZN(n9294) );
  OAI21_X1 U11603 ( .B1(n9292), .B2(n11646), .A(n9294), .ZN(n9297) );
  NOR2_X1 U11604 ( .A1(n11637), .A2(n12374), .ZN(n9295) );
  INV_X1 U11605 ( .A(n11639), .ZN(n9293) );
  AOI22_X1 U11606 ( .A1(n9295), .A2(n9294), .B1(n11556), .B2(n9293), .ZN(n9296) );
  XOR2_X1 U11607 ( .A(n9302), .B(n11519), .Z(n11511) );
  NOR2_X1 U11608 ( .A1(n11511), .A2(n12372), .ZN(n9298) );
  XNOR2_X1 U11609 ( .A(n11630), .B(n9261), .ZN(n11625) );
  NOR2_X1 U11610 ( .A1(n11625), .A2(n11663), .ZN(n9300) );
  INV_X1 U11611 ( .A(n11625), .ZN(n9299) );
  XNOR2_X1 U11612 ( .A(n9301), .B(n11629), .ZN(n12348) );
  XOR2_X1 U11613 ( .A(n12240), .B(n12747), .Z(n12287) );
  XNOR2_X1 U11614 ( .A(n12813), .B(n12240), .ZN(n9303) );
  XNOR2_X1 U11615 ( .A(n9303), .B(n12668), .ZN(n11989) );
  NAND2_X1 U11616 ( .A1(n9303), .A2(n12668), .ZN(n12327) );
  XNOR2_X1 U11617 ( .A(n12739), .B(n12240), .ZN(n9306) );
  INV_X1 U11618 ( .A(n9306), .ZN(n9304) );
  NAND2_X1 U11619 ( .A1(n9304), .A2(n12368), .ZN(n9305) );
  AND2_X1 U11620 ( .A1(n12327), .A2(n9305), .ZN(n9308) );
  INV_X1 U11621 ( .A(n9305), .ZN(n9307) );
  XNOR2_X1 U11622 ( .A(n9306), .B(n12368), .ZN(n12329) );
  XNOR2_X1 U11623 ( .A(n12808), .B(n12240), .ZN(n9311) );
  XNOR2_X1 U11624 ( .A(n9311), .B(n12332), .ZN(n12305) );
  XNOR2_X1 U11625 ( .A(n12646), .B(n12240), .ZN(n9313) );
  XNOR2_X1 U11626 ( .A(n9313), .B(n12367), .ZN(n12309) );
  AND2_X1 U11627 ( .A1(n12305), .A2(n12309), .ZN(n9309) );
  XNOR2_X1 U11628 ( .A(n12631), .B(n12240), .ZN(n9310) );
  NAND2_X1 U11629 ( .A1(n9310), .A2(n12641), .ZN(n9319) );
  OAI21_X1 U11630 ( .B1(n9310), .B2(n12641), .A(n9319), .ZN(n12271) );
  INV_X1 U11631 ( .A(n12271), .ZN(n9317) );
  INV_X1 U11632 ( .A(n12309), .ZN(n9312) );
  NAND2_X1 U11633 ( .A1(n9311), .A2(n12667), .ZN(n12307) );
  INV_X1 U11634 ( .A(n9313), .ZN(n9314) );
  NAND2_X1 U11635 ( .A1(n9314), .A2(n12367), .ZN(n9315) );
  XNOR2_X1 U11636 ( .A(n12796), .B(n12240), .ZN(n9321) );
  NAND2_X1 U11637 ( .A1(n9320), .A2(n9321), .ZN(n9324) );
  INV_X1 U11638 ( .A(n9321), .ZN(n9322) );
  OR2_X2 U11639 ( .A1(n12320), .A2(n12365), .ZN(n12318) );
  NAND2_X1 U11640 ( .A1(n12318), .A2(n9326), .ZN(n9331) );
  XNOR2_X1 U11641 ( .A(n12610), .B(n12240), .ZN(n9330) );
  INV_X1 U11642 ( .A(n12320), .ZN(n9325) );
  INV_X1 U11643 ( .A(n9330), .ZN(n9327) );
  AND2_X2 U11644 ( .A1(n9329), .A2(n9328), .ZN(n12298) );
  OAI21_X1 U11645 ( .B1(n9331), .B2(n9330), .A(n12298), .ZN(n12256) );
  XNOR2_X1 U11646 ( .A(n12297), .B(n12240), .ZN(n9332) );
  NAND2_X1 U11647 ( .A1(n9332), .A2(n12607), .ZN(n12277) );
  INV_X1 U11648 ( .A(n9332), .ZN(n9333) );
  NAND2_X1 U11649 ( .A1(n9333), .A2(n12363), .ZN(n9334) );
  XNOR2_X1 U11650 ( .A(n12709), .B(n12240), .ZN(n9335) );
  NAND2_X1 U11651 ( .A1(n9335), .A2(n12594), .ZN(n9339) );
  INV_X1 U11652 ( .A(n9335), .ZN(n9336) );
  NAND2_X1 U11653 ( .A1(n9336), .A2(n12362), .ZN(n9337) );
  NAND2_X1 U11654 ( .A1(n9338), .A2(n12278), .ZN(n12279) );
  XNOR2_X1 U11655 ( .A(n9340), .B(n9261), .ZN(n9341) );
  AOI21_X1 U11656 ( .B1(n9341), .B2(n12578), .A(n9342), .ZN(n12340) );
  XNOR2_X1 U11657 ( .A(n12701), .B(n9261), .ZN(n12247) );
  NOR2_X1 U11658 ( .A1(n12247), .A2(n7018), .ZN(n12242) );
  OAI22_X1 U11659 ( .A1(n9350), .A2(n9979), .B1(n9366), .B2(n9351), .ZN(n9344)
         );
  INV_X1 U11660 ( .A(n12701), .ZN(n12559) );
  AND2_X1 U11661 ( .A1(n9731), .A2(n14467), .ZN(n9345) );
  NAND2_X1 U11662 ( .A1(n9346), .A2(n9345), .ZN(n9348) );
  NOR2_X1 U11663 ( .A1(n15109), .A2(n14470), .ZN(n9347) );
  NAND2_X1 U11664 ( .A1(n9731), .A2(n9347), .ZN(n15111) );
  NAND2_X1 U11665 ( .A1(n9350), .A2(n9349), .ZN(n9356) );
  INV_X1 U11666 ( .A(n9351), .ZN(n9352) );
  NAND2_X1 U11667 ( .A1(n9366), .A2(n9352), .ZN(n9355) );
  NAND2_X1 U11668 ( .A1(n9353), .A2(n9733), .ZN(n9354) );
  NAND4_X1 U11669 ( .A1(n9356), .A2(n9376), .A3(n9355), .A4(n9354), .ZN(n9357)
         );
  NAND2_X1 U11670 ( .A1(n9357), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9360) );
  AOI21_X1 U11671 ( .B1(n9358), .B2(n9366), .A(n9730), .ZN(n9359) );
  INV_X1 U11672 ( .A(n9366), .ZN(n9363) );
  NOR2_X1 U11673 ( .A1(n9361), .A2(n12759), .ZN(n9362) );
  NAND2_X1 U11674 ( .A1(n9363), .A2(n9362), .ZN(n12354) );
  NAND2_X1 U11675 ( .A1(n9364), .A2(n12756), .ZN(n9365) );
  NOR2_X2 U11676 ( .A1(n9366), .A2(n9365), .ZN(n12352) );
  AOI22_X1 U11677 ( .A1(n12578), .A2(n12352), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9367) );
  OAI21_X1 U11678 ( .B1(n9368), .B2(n12354), .A(n9367), .ZN(n9369) );
  AOI21_X1 U11679 ( .B1(n12557), .B2(n12356), .A(n9369), .ZN(n9370) );
  OAI21_X1 U11680 ( .B1(n12559), .B2(n12360), .A(n9370), .ZN(n9371) );
  NAND2_X1 U11681 ( .A1(n9373), .A2(n9372), .ZN(P3_U3154) );
  INV_X1 U11682 ( .A(n9801), .ZN(n9374) );
  NOR2_X1 U11683 ( .A1(n9375), .A2(n9374), .ZN(n9804) );
  AND2_X1 U11684 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9804), .ZN(P2_U3947) );
  INV_X1 U11685 ( .A(n9490), .ZN(n12821) );
  OR2_X2 U11686 ( .A1(n9376), .A2(n12821), .ZN(n12385) );
  NOR2_X2 U11687 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9377) );
  NAND4_X1 U11688 ( .A1(n9378), .A2(n9377), .A3(n9532), .A4(n9905), .ZN(n9381)
         );
  NAND4_X1 U11689 ( .A1(n9595), .A2(n10096), .A3(n9379), .A4(n9402), .ZN(n9380) );
  NOR3_X1 U11690 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .A3(P1_IR_REG_15__SCAN_IN), .ZN(n9382) );
  OAI21_X1 U11691 ( .B1(n9430), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9387) );
  XNOR2_X1 U11692 ( .A(n9387), .B(n9388), .ZN(n9668) );
  NAND2_X1 U11693 ( .A1(n9668), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9518) );
  NAND4_X1 U11694 ( .A1(n9390), .A2(n9389), .A3(n9431), .A4(n9388), .ZN(n9392)
         );
  NAND2_X1 U11695 ( .A1(n9386), .A2(n9538), .ZN(n9391) );
  INV_X1 U11696 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9398) );
  OAI21_X1 U11697 ( .B1(n9395), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9394) );
  XNOR2_X1 U11698 ( .A(n9394), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9515) );
  INV_X1 U11699 ( .A(n9515), .ZN(n14280) );
  NAND2_X1 U11700 ( .A1(n9395), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9397) );
  INV_X1 U11701 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U11702 ( .A1(n9427), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9399) );
  XNOR2_X1 U11703 ( .A(n9399), .B(n9398), .ZN(n14284) );
  OR2_X2 U11704 ( .A1(n9518), .A2(n9667), .ZN(n13847) );
  INV_X1 U11705 ( .A(n13847), .ZN(P1_U4016) );
  INV_X1 U11706 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10271) );
  INV_X1 U11707 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14272) );
  NOR2_X1 U11708 ( .A1(n10173), .A2(n14272), .ZN(n9401) );
  MUX2_X1 U11709 ( .A(n14272), .B(n9401), .S(P1_IR_REG_5__SCAN_IN), .Z(n9404)
         );
  NAND2_X1 U11710 ( .A1(n10173), .A2(n9402), .ZN(n9520) );
  INV_X1 U11711 ( .A(n9520), .ZN(n9403) );
  OR2_X1 U11712 ( .A1(n9404), .A2(n9403), .ZN(n10252) );
  MUX2_X1 U11713 ( .A(n10271), .B(P1_REG1_REG_5__SCAN_IN), .S(n10252), .Z(
        n9604) );
  INV_X1 U11714 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9407) );
  OR2_X1 U11715 ( .A1(n9405), .A2(n14272), .ZN(n9406) );
  XNOR2_X1 U11716 ( .A(n9406), .B(P1_IR_REG_2__SCAN_IN), .ZN(n13868) );
  MUX2_X1 U11717 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9407), .S(n13868), .Z(n9411) );
  INV_X1 U11718 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U11719 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9408) );
  XNOR2_X1 U11720 ( .A(n9408), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13852) );
  MUX2_X1 U11721 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9409), .S(n13852), .Z(
        n13850) );
  AND2_X1 U11722 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13851) );
  NAND2_X1 U11723 ( .A1(n13850), .A2(n13851), .ZN(n13870) );
  NAND2_X1 U11724 ( .A1(n13852), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n13869) );
  NAND2_X1 U11725 ( .A1(n13870), .A2(n13869), .ZN(n9410) );
  NAND2_X1 U11726 ( .A1(n9411), .A2(n9410), .ZN(n13883) );
  NAND2_X1 U11727 ( .A1(n13868), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13881) );
  NAND2_X1 U11728 ( .A1(n13883), .A2(n13881), .ZN(n9416) );
  INV_X1 U11729 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11730 ( .A1(n9412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9413) );
  XNOR2_X1 U11731 ( .A(n9413), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13885) );
  MUX2_X1 U11732 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9414), .S(n13885), .Z(n9415) );
  NAND2_X1 U11733 ( .A1(n9416), .A2(n9415), .ZN(n14668) );
  NAND2_X1 U11734 ( .A1(n13885), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14667) );
  NAND2_X1 U11735 ( .A1(n14668), .A2(n14667), .ZN(n9421) );
  NAND2_X1 U11736 ( .A1(n9417), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9419) );
  INV_X1 U11737 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9418) );
  XNOR2_X1 U11738 ( .A(n9419), .B(n9418), .ZN(n14665) );
  MUX2_X1 U11739 ( .A(n14811), .B(P1_REG1_REG_4__SCAN_IN), .S(n14665), .Z(
        n9420) );
  NAND2_X1 U11740 ( .A1(n9421), .A2(n9420), .ZN(n14670) );
  INV_X1 U11741 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14811) );
  OR2_X1 U11742 ( .A1(n14665), .A2(n14811), .ZN(n9422) );
  AND2_X1 U11743 ( .A1(n14670), .A2(n9422), .ZN(n9603) );
  NAND2_X1 U11744 ( .A1(n9604), .A2(n9603), .ZN(n9602) );
  NAND2_X1 U11745 ( .A1(n10252), .A2(n10271), .ZN(n9423) );
  NAND2_X1 U11746 ( .A1(n9602), .A2(n9423), .ZN(n9445) );
  INV_X1 U11747 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10788) );
  NAND2_X1 U11748 ( .A1(n9520), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9424) );
  XNOR2_X1 U11749 ( .A(n9424), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10522) );
  MUX2_X1 U11750 ( .A(n10788), .B(P1_REG1_REG_6__SCAN_IN), .S(n10522), .Z(
        n9444) );
  NOR2_X1 U11751 ( .A1(n9445), .A2(n9444), .ZN(n13902) );
  NOR2_X1 U11752 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9438) );
  INV_X1 U11753 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U11754 ( .A1(n9438), .A2(n9425), .ZN(n9426) );
  INV_X1 U11755 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9428) );
  INV_X1 U11756 ( .A(n9667), .ZN(n9661) );
  OR2_X1 U11757 ( .A1(n9668), .A2(P1_U3086), .ZN(n13817) );
  NAND2_X1 U11758 ( .A1(n10353), .A2(n13817), .ZN(n9463) );
  INV_X1 U11759 ( .A(n9433), .ZN(n9434) );
  NAND2_X1 U11760 ( .A1(n9565), .A2(n9564), .ZN(n13762) );
  INV_X1 U11761 ( .A(n13762), .ZN(n9436) );
  NAND2_X1 U11762 ( .A1(n9436), .A2(n9668), .ZN(n9442) );
  NOR2_X1 U11763 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n9437) );
  INV_X1 U11764 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U11765 ( .A1(n9442), .A2(n11895), .ZN(n9462) );
  INV_X1 U11766 ( .A(n9462), .ZN(n9443) );
  NAND2_X1 U11767 ( .A1(n9463), .A2(n9443), .ZN(n9447) );
  INV_X1 U11768 ( .A(n9447), .ZN(n9509) );
  AND2_X1 U11769 ( .A1(n6455), .A2(n9509), .ZN(n14689) );
  INV_X1 U11770 ( .A(n14689), .ZN(n13913) );
  AOI211_X1 U11771 ( .C1(n9445), .C2(n9444), .A(n13902), .B(n13913), .ZN(n9467) );
  INV_X1 U11772 ( .A(n11772), .ZN(n13860) );
  OR2_X1 U11773 ( .A1(n9447), .A2(n13860), .ZN(n13955) );
  INV_X1 U11774 ( .A(n10522), .ZN(n9615) );
  NOR2_X1 U11775 ( .A1(n13955), .A2(n9615), .ZN(n9466) );
  INV_X1 U11776 ( .A(n6455), .ZN(n13857) );
  NAND2_X1 U11777 ( .A1(n13860), .A2(n13857), .ZN(n9446) );
  OR2_X1 U11778 ( .A1(n9447), .A2(n9446), .ZN(n13956) );
  INV_X1 U11779 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9448) );
  MUX2_X1 U11780 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9448), .S(n13868), .Z(n9451) );
  INV_X1 U11781 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9449) );
  MUX2_X1 U11782 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9449), .S(n13852), .Z(
        n13849) );
  AND2_X1 U11783 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13858) );
  NAND2_X1 U11784 ( .A1(n13849), .A2(n13858), .ZN(n13865) );
  NAND2_X1 U11785 ( .A1(n13852), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n13864) );
  NAND2_X1 U11786 ( .A1(n13865), .A2(n13864), .ZN(n9450) );
  NAND2_X1 U11787 ( .A1(n9451), .A2(n9450), .ZN(n13888) );
  NAND2_X1 U11788 ( .A1(n13868), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13886) );
  NAND2_X1 U11789 ( .A1(n13888), .A2(n13886), .ZN(n9454) );
  INV_X1 U11790 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9452) );
  MUX2_X1 U11791 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9452), .S(n13885), .Z(n9453) );
  NAND2_X1 U11792 ( .A1(n9454), .A2(n9453), .ZN(n14662) );
  NAND2_X1 U11793 ( .A1(n13885), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14661) );
  NAND2_X1 U11794 ( .A1(n14662), .A2(n14661), .ZN(n9456) );
  INV_X1 U11795 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10485) );
  MUX2_X1 U11796 ( .A(n10485), .B(P1_REG2_REG_4__SCAN_IN), .S(n14665), .Z(
        n9455) );
  NAND2_X1 U11797 ( .A1(n9456), .A2(n9455), .ZN(n14664) );
  INV_X1 U11798 ( .A(n14665), .ZN(n14671) );
  NAND2_X1 U11799 ( .A1(n14671), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9605) );
  INV_X1 U11800 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9457) );
  MUX2_X1 U11801 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9457), .S(n10252), .Z(n9606) );
  AOI21_X1 U11802 ( .B1(n14664), .B2(n9605), .A(n9606), .ZN(n9608) );
  NOR2_X1 U11803 ( .A1(n10252), .A2(n9457), .ZN(n9459) );
  INV_X1 U11804 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10719) );
  MUX2_X1 U11805 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10719), .S(n10522), .Z(
        n9458) );
  OAI21_X1 U11806 ( .B1(n9608), .B2(n9459), .A(n9458), .ZN(n13905) );
  INV_X1 U11807 ( .A(n13905), .ZN(n9461) );
  NOR3_X1 U11808 ( .A1(n9608), .A2(n9459), .A3(n9458), .ZN(n9460) );
  NOR3_X1 U11809 ( .A1(n13956), .A2(n9461), .A3(n9460), .ZN(n9465) );
  AND2_X1 U11810 ( .A1(n9463), .A2(n9462), .ZN(n14673) );
  INV_X1 U11811 ( .A(n14673), .ZN(n14694) );
  INV_X1 U11812 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14347) );
  INV_X1 U11813 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n12158) );
  OAI22_X1 U11814 ( .A1(n14694), .A2(n14347), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12158), .ZN(n9464) );
  OR4_X1 U11815 ( .A1(n9467), .A2(n9466), .A3(n9465), .A4(n9464), .ZN(P1_U3249) );
  INV_X1 U11816 ( .A(n9762), .ZN(n9790) );
  NAND2_X1 U11817 ( .A1(n8134), .A2(P3_U3151), .ZN(n12832) );
  OAI222_X1 U11818 ( .A1(P3_U3151), .A2(n9790), .B1(n12829), .B2(n9469), .C1(
        n12832), .C2(n9468), .ZN(P3_U3294) );
  OAI222_X1 U11819 ( .A1(n12832), .A2(n9471), .B1(n12829), .B2(n9470), .C1(
        n10298), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U11820 ( .A(SI_9_), .ZN(n9472) );
  OAI222_X1 U11821 ( .A1(n12832), .A2(n9473), .B1(n12829), .B2(n9472), .C1(
        n15071), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U11822 ( .A(SI_8_), .ZN(n9474) );
  INV_X1 U11823 ( .A(n10906), .ZN(n10886) );
  OAI222_X1 U11824 ( .A1(n12832), .A2(n9475), .B1(n12829), .B2(n9474), .C1(
        n10886), .C2(P3_U3151), .ZN(P3_U3287) );
  AND2_X1 U11825 ( .A1(n9139), .A2(P1_U3086), .ZN(n14275) );
  INV_X1 U11826 ( .A(n13852), .ZN(n9476) );
  OAI222_X1 U11827 ( .A1(n6454), .A2(n9477), .B1(n14286), .B2(n9712), .C1(
        P1_U3086), .C2(n9476), .ZN(P1_U3354) );
  NOR2_X1 U11828 ( .A1(n9139), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13451) );
  NAND2_X1 U11829 ( .A1(n9139), .A2(P2_U3088), .ZN(n13467) );
  OAI222_X1 U11830 ( .A1(n13458), .A2(n9478), .B1(n13467), .B2(n9712), .C1(
        P2_U3088), .C2(n9815), .ZN(P2_U3326) );
  OAI222_X1 U11831 ( .A1(n15033), .A2(P3_U3151), .B1(n12832), .B2(n9480), .C1(
        n9479), .C2(n12829), .ZN(P3_U3291) );
  OAI222_X1 U11832 ( .A1(n10015), .A2(P3_U3151), .B1(n12832), .B2(n9482), .C1(
        n9481), .C2(n12829), .ZN(P3_U3292) );
  INV_X1 U11833 ( .A(n9483), .ZN(n9485) );
  INV_X1 U11834 ( .A(SI_10_), .ZN(n9484) );
  OAI222_X1 U11835 ( .A1(n12832), .A2(n9485), .B1(n12829), .B2(n9484), .C1(
        n10904), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U11836 ( .A(n9486), .ZN(n9487) );
  INV_X1 U11837 ( .A(n11143), .ZN(n11137) );
  OAI222_X1 U11838 ( .A1(n12832), .A2(n9487), .B1(n12829), .B2(n12095), .C1(
        n11137), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U11839 ( .A(n6450), .ZN(n9775) );
  INV_X1 U11840 ( .A(SI_2_), .ZN(n9488) );
  OAI222_X1 U11841 ( .A1(n9775), .A2(P3_U3151), .B1(n12832), .B2(n9489), .C1(
        n9488), .C2(n12829), .ZN(P3_U3293) );
  AND2_X1 U11842 ( .A1(n8697), .A2(n9490), .ZN(n9512) );
  INV_X1 U11843 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n12164) );
  NOR2_X1 U11844 ( .A1(n9512), .A2(n12164), .ZN(P3_U3238) );
  INV_X1 U11845 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n12199) );
  NOR2_X1 U11846 ( .A1(n9512), .A2(n12199), .ZN(P3_U3263) );
  OAI222_X1 U11847 ( .A1(n6454), .A2(n10232), .B1(n14286), .B2(n10231), .C1(
        P1_U3086), .C2(n14665), .ZN(P1_U3351) );
  INV_X1 U11848 ( .A(n13885), .ZN(n9491) );
  OAI222_X1 U11849 ( .A1(n6454), .A2(n9492), .B1(n14286), .B2(n10228), .C1(
        P1_U3086), .C2(n9491), .ZN(P1_U3352) );
  OAI222_X1 U11850 ( .A1(n6454), .A2(n9493), .B1(n14286), .B2(n10251), .C1(
        P1_U3086), .C2(n10252), .ZN(P1_U3350) );
  INV_X1 U11851 ( .A(n13868), .ZN(n13875) );
  OAI222_X1 U11852 ( .A1(n6454), .A2(n6699), .B1(n14286), .B2(n9913), .C1(
        P1_U3086), .C2(n13875), .ZN(P1_U3353) );
  INV_X1 U11853 ( .A(n12832), .ZN(n14422) );
  AOI22_X1 U11854 ( .A1(n14422), .A2(n9494), .B1(P3_STATE_REG_SCAN_IN), .B2(
        P3_IR_REG_0__SCAN_IN), .ZN(n9495) );
  OAI21_X1 U11855 ( .B1(n9581), .B2(n12829), .A(n9495), .ZN(P3_U3295) );
  OAI222_X1 U11856 ( .A1(n6454), .A2(n9496), .B1(n14286), .B2(n10521), .C1(
        P1_U3086), .C2(n9615), .ZN(P1_U3349) );
  INV_X1 U11857 ( .A(SI_6_), .ZN(n9497) );
  OAI222_X1 U11858 ( .A1(n10065), .A2(P3_U3151), .B1(n12832), .B2(n9498), .C1(
        n9497), .C2(n12829), .ZN(P3_U3289) );
  INV_X1 U11859 ( .A(SI_5_), .ZN(n9499) );
  OAI222_X1 U11860 ( .A1(n15053), .A2(P3_U3151), .B1(n12832), .B2(n9500), .C1(
        n9499), .C2(n12829), .ZN(P3_U3290) );
  INV_X1 U11861 ( .A(n13467), .ZN(n11417) );
  INV_X1 U11862 ( .A(n11417), .ZN(n13461) );
  OAI222_X1 U11863 ( .A1(n13458), .A2(n9501), .B1(n13461), .B2(n10521), .C1(
        P2_U3088), .C2(n13071), .ZN(P2_U3321) );
  OAI222_X1 U11864 ( .A1(n13458), .A2(n9502), .B1(n13461), .B2(n10228), .C1(
        P2_U3088), .C2(n13051), .ZN(P2_U3324) );
  OAI222_X1 U11865 ( .A1(n13458), .A2(n9503), .B1(n13461), .B2(n10251), .C1(
        P2_U3088), .C2(n14858), .ZN(P2_U3322) );
  OAI222_X1 U11866 ( .A1(n13458), .A2(n9504), .B1(n13461), .B2(n10231), .C1(
        P2_U3088), .C2(n9823), .ZN(P2_U3323) );
  OAI222_X1 U11867 ( .A1(n13458), .A2(n9505), .B1(n13461), .B2(n9913), .C1(
        P2_U3088), .C2(n9818), .ZN(P2_U3325) );
  NOR2_X1 U11868 ( .A1(n14673), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11869 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9511) );
  INV_X1 U11870 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9506) );
  AOI21_X1 U11871 ( .B1(n13857), .B2(n9506), .A(n11772), .ZN(n13863) );
  OAI21_X1 U11872 ( .B1(n13857), .B2(P1_REG1_REG_0__SCAN_IN), .A(n13863), .ZN(
        n9507) );
  XNOR2_X1 U11873 ( .A(n9507), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9508) );
  AOI22_X1 U11874 ( .A1(n9509), .A2(n9508), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9510) );
  OAI21_X1 U11875 ( .B1(n14694), .B2(n9511), .A(n9510), .ZN(P1_U3243) );
  AND2_X1 U11876 ( .A1(n9513), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11877 ( .A1(n9513), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11878 ( .A1(n9513), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11879 ( .A1(n9513), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11880 ( .A1(n9513), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11881 ( .A1(n9513), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11882 ( .A1(n9513), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11883 ( .A1(n9513), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11884 ( .A1(n9513), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U11885 ( .A1(n9513), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11886 ( .A1(n9513), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11887 ( .A1(n9513), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11888 ( .A1(n9513), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11889 ( .A1(n9513), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11890 ( .A1(n9513), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11891 ( .A1(n9513), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11892 ( .A1(n9513), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11893 ( .A1(n9513), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11894 ( .A1(n9513), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11895 ( .A1(n9513), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11896 ( .A1(n9513), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11897 ( .A1(n9513), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11898 ( .A1(n9513), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11899 ( .A1(n9513), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11900 ( .A1(n9513), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11901 ( .A1(n9513), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11902 ( .A1(n9513), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11903 ( .A1(n9513), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  NAND3_X1 U11904 ( .A1(n14281), .A2(P1_B_REG_SCAN_IN), .A3(n14284), .ZN(n9514) );
  OAI211_X1 U11905 ( .C1(P1_B_REG_SCAN_IN), .C2(n14284), .A(n9515), .B(n9514), 
        .ZN(n9557) );
  INV_X1 U11906 ( .A(n9557), .ZN(n9516) );
  INV_X1 U11907 ( .A(n14744), .ZN(n14743) );
  NAND2_X1 U11908 ( .A1(n14280), .A2(n14281), .ZN(n9554) );
  OAI22_X1 U11909 ( .A1(n14743), .A2(P1_D_REG_1__SCAN_IN), .B1(n9518), .B2(
        n9554), .ZN(n9517) );
  INV_X1 U11910 ( .A(n9517), .ZN(P1_U3446) );
  NAND2_X1 U11911 ( .A1(n14280), .A2(n14284), .ZN(n9558) );
  OAI22_X1 U11912 ( .A1(n14743), .A2(P1_D_REG_0__SCAN_IN), .B1(n9558), .B2(
        n9518), .ZN(n9519) );
  INV_X1 U11913 ( .A(n9519), .ZN(P1_U3445) );
  INV_X1 U11914 ( .A(n10591), .ZN(n9524) );
  NAND2_X1 U11915 ( .A1(n9526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U11916 ( .A(n9521), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13897) );
  INV_X1 U11917 ( .A(n13897), .ZN(n9620) );
  OAI222_X1 U11918 ( .A1(n6454), .A2(n9522), .B1(n14286), .B2(n9524), .C1(
        P1_U3086), .C2(n9620), .ZN(P1_U3348) );
  INV_X1 U11919 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9525) );
  INV_X1 U11920 ( .A(n14873), .ZN(n9523) );
  OAI222_X1 U11921 ( .A1(n13458), .A2(n9525), .B1(n13461), .B2(n9524), .C1(
        P2_U3088), .C2(n9523), .ZN(P2_U3320) );
  INV_X1 U11922 ( .A(n10595), .ZN(n9530) );
  INV_X1 U11923 ( .A(n9533), .ZN(n9527) );
  NAND2_X1 U11924 ( .A1(n9527), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9528) );
  XNOR2_X1 U11925 ( .A(n9528), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10596) );
  INV_X1 U11926 ( .A(n10596), .ZN(n9699) );
  OAI222_X1 U11927 ( .A1(n6454), .A2(n9529), .B1(n14286), .B2(n9530), .C1(
        P1_U3086), .C2(n9699), .ZN(P1_U3347) );
  INV_X1 U11928 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9531) );
  OAI222_X1 U11929 ( .A1(n13458), .A2(n9531), .B1(n13461), .B2(n9530), .C1(
        P2_U3088), .C2(n9829), .ZN(P2_U3319) );
  INV_X1 U11930 ( .A(n10996), .ZN(n9536) );
  NAND2_X1 U11931 ( .A1(n9533), .A2(n9532), .ZN(n9613) );
  NAND2_X1 U11932 ( .A1(n9613), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9596) );
  XNOR2_X1 U11933 ( .A(n9596), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U11934 ( .A1(n10997), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n14275), .ZN(n9534) );
  OAI21_X1 U11935 ( .B1(n9536), .B2(n14286), .A(n9534), .ZN(P1_U3346) );
  OAI222_X1 U11936 ( .A1(n12440), .A2(P3_U3151), .B1(n12832), .B2(n9535), .C1(
        n7261), .C2(n12829), .ZN(P3_U3281) );
  INV_X1 U11937 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9537) );
  INV_X1 U11938 ( .A(n9864), .ZN(n9832) );
  OAI222_X1 U11939 ( .A1(n13458), .A2(n9537), .B1(n13461), .B2(n9536), .C1(
        P2_U3088), .C2(n9832), .ZN(P2_U3318) );
  NAND2_X1 U11940 ( .A1(n9541), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9542) );
  XNOR2_X2 U11941 ( .A(n9542), .B(n9386), .ZN(n14155) );
  AND2_X1 U11942 ( .A1(n13738), .A2(n14155), .ZN(n9655) );
  OR2_X1 U11943 ( .A1(n13762), .A2(n9655), .ZN(n9670) );
  NOR4_X1 U11944 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n9551) );
  NOR4_X1 U11945 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9550) );
  OR4_X1 U11946 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9548) );
  NOR4_X1 U11947 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n9546) );
  NOR4_X1 U11948 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n9545) );
  NOR4_X1 U11949 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9544) );
  NOR4_X1 U11950 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9543) );
  NAND4_X1 U11951 ( .A1(n9546), .A2(n9545), .A3(n9544), .A4(n9543), .ZN(n9547)
         );
  NOR4_X1 U11952 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9548), .A4(n9547), .ZN(n9549) );
  AND3_X1 U11953 ( .A1(n9551), .A2(n9550), .A3(n9549), .ZN(n9552) );
  OR2_X1 U11954 ( .A1(n9557), .A2(n9552), .ZN(n9654) );
  NAND2_X1 U11955 ( .A1(n9670), .A2(n9654), .ZN(n9553) );
  NOR2_X1 U11956 ( .A1(n10353), .A2(n9553), .ZN(n10358) );
  OR2_X1 U11957 ( .A1(n9557), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9555) );
  AND2_X1 U11958 ( .A1(n9555), .A2(n9554), .ZN(n9653) );
  INV_X1 U11959 ( .A(n9653), .ZN(n10356) );
  AND2_X1 U11960 ( .A1(n10354), .A2(n10356), .ZN(n9556) );
  OR2_X1 U11961 ( .A1(n9557), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9559) );
  INV_X1 U11962 ( .A(n10355), .ZN(n9560) );
  AND2_X2 U11963 ( .A1(n10219), .A2(n9560), .ZN(n14807) );
  INV_X1 U11964 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9594) );
  OR2_X1 U11965 ( .A1(n13569), .A2(n14155), .ZN(n9563) );
  NAND2_X1 U11966 ( .A1(n9564), .A2(n6806), .ZN(n9562) );
  NAND2_X1 U11967 ( .A1(n9565), .A2(n14155), .ZN(n13571) );
  OR2_X1 U11968 ( .A1(n13584), .A2(n13571), .ZN(n9566) );
  NAND2_X1 U11969 ( .A1(n10364), .A2(n14155), .ZN(n14130) );
  OR2_X1 U11970 ( .A1(n13761), .A2(n14155), .ZN(n14745) );
  NAND2_X1 U11971 ( .A1(n14130), .A2(n14745), .ZN(n14803) );
  INV_X1 U11972 ( .A(n9569), .ZN(n9568) );
  NAND2_X1 U11973 ( .A1(n6446), .A2(n9567), .ZN(n14273) );
  NAND2_X1 U11974 ( .A1(n9569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U11975 ( .A1(n14273), .A2(n9571), .ZN(n11770) );
  INV_X1 U11976 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U11977 ( .A1(n11961), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9579) );
  AND2_X2 U11978 ( .A1(n12235), .A2(n11770), .ZN(n10236) );
  NAND2_X1 U11979 ( .A1(n10236), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9578) );
  AND2_X2 U11980 ( .A1(n12235), .A2(n9574), .ZN(n9925) );
  NAND2_X1 U11981 ( .A1(n9925), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U11982 ( .A1(n10235), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9576) );
  NAND4_X2 U11983 ( .A1(n9579), .A2(n9578), .A3(n9577), .A4(n9576), .ZN(n13848) );
  INV_X1 U11984 ( .A(n13848), .ZN(n9585) );
  INV_X1 U11985 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9664) );
  OAI21_X1 U11986 ( .B1(n9139), .B2(n9581), .A(n9580), .ZN(n9583) );
  NAND2_X1 U11987 ( .A1(n9584), .A2(n9583), .ZN(n14289) );
  MUX2_X1 U11988 ( .A(n9664), .B(n14289), .S(n6458), .Z(n14731) );
  INV_X1 U11989 ( .A(n14731), .ZN(n10257) );
  NAND2_X1 U11990 ( .A1(n13848), .A2(n14731), .ZN(n9586) );
  NAND2_X1 U11991 ( .A1(n14722), .A2(n9586), .ZN(n13776) );
  OAI21_X1 U11992 ( .B1(n14784), .B2(n14803), .A(n13776), .ZN(n9592) );
  NAND2_X1 U11993 ( .A1(n11961), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9590) );
  NAND2_X1 U11994 ( .A1(n10236), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9589) );
  NAND2_X1 U11995 ( .A1(n9925), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9588) );
  NAND2_X1 U11996 ( .A1(n10235), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9587) );
  OR2_X1 U11997 ( .A1(n13762), .A2(n13860), .ZN(n13544) );
  INV_X2 U11998 ( .A(n13544), .ZN(n14645) );
  NAND2_X1 U11999 ( .A1(n13846), .A2(n14645), .ZN(n10360) );
  INV_X1 U12000 ( .A(n9564), .ZN(n13572) );
  NAND3_X1 U12001 ( .A1(n10257), .A2(n13572), .A3(n13569), .ZN(n9591) );
  NAND3_X1 U12002 ( .A1(n9592), .A2(n10360), .A3(n9591), .ZN(n14254) );
  NAND2_X1 U12003 ( .A1(n14254), .A2(n14807), .ZN(n9593) );
  OAI21_X1 U12004 ( .B1(n14807), .B2(n9594), .A(n9593), .ZN(P1_U3459) );
  INV_X1 U12005 ( .A(n11001), .ZN(n9600) );
  NAND2_X1 U12006 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  NAND2_X1 U12007 ( .A1(n9597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9598) );
  XNOR2_X1 U12008 ( .A(n9598), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11002) );
  INV_X1 U12009 ( .A(n11002), .ZN(n9625) );
  OAI222_X1 U12010 ( .A1(n6454), .A2(n9599), .B1(n14286), .B2(n9600), .C1(
        P1_U3086), .C2(n9625), .ZN(P1_U3345) );
  INV_X1 U12011 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9601) );
  INV_X1 U12012 ( .A(n9955), .ZN(n9812) );
  OAI222_X1 U12013 ( .A1(n13458), .A2(n9601), .B1(n13461), .B2(n9600), .C1(
        P2_U3088), .C2(n9812), .ZN(P2_U3317) );
  OAI21_X1 U12014 ( .B1(n9604), .B2(n9603), .A(n9602), .ZN(n9610) );
  AND3_X1 U12015 ( .A1(n9606), .A2(n14664), .A3(n9605), .ZN(n9607) );
  NOR3_X1 U12016 ( .A1(n13956), .A2(n9608), .A3(n9607), .ZN(n9609) );
  AOI21_X1 U12017 ( .B1(n14689), .B2(n9610), .A(n9609), .ZN(n9612) );
  AND2_X1 U12018 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10396) );
  AOI21_X1 U12019 ( .B1(n14673), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10396), .ZN(
        n9611) );
  OAI211_X1 U12020 ( .C1(n10252), .C2(n13955), .A(n9612), .B(n9611), .ZN(
        P1_U3248) );
  INV_X1 U12021 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14612) );
  NAND2_X1 U12022 ( .A1(n9677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9614) );
  XNOR2_X1 U12023 ( .A(n9614), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11099) );
  MUX2_X1 U12024 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14612), .S(n11099), .Z(
        n9619) );
  INV_X1 U12025 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14813) );
  NOR2_X1 U12026 ( .A1(n9615), .A2(n10788), .ZN(n13896) );
  MUX2_X1 U12027 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14813), .S(n13897), .Z(
        n9616) );
  OAI21_X1 U12028 ( .B1(n13902), .B2(n13896), .A(n9616), .ZN(n13900) );
  OAI21_X1 U12029 ( .B1(n14813), .B2(n9620), .A(n13900), .ZN(n9697) );
  INV_X1 U12030 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9617) );
  MUX2_X1 U12031 ( .A(n9617), .B(P1_REG1_REG_8__SCAN_IN), .S(n10596), .Z(n9698) );
  NOR2_X1 U12032 ( .A1(n9697), .A2(n9698), .ZN(n9696) );
  NOR2_X1 U12033 ( .A1(n10596), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9645) );
  INV_X1 U12034 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11065) );
  MUX2_X1 U12035 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n11065), .S(n10997), .Z(
        n9646) );
  OAI21_X1 U12036 ( .B1(n9696), .B2(n9645), .A(n9646), .ZN(n9644) );
  OAI21_X1 U12037 ( .B1(n10997), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9644), .ZN(
        n9937) );
  INV_X1 U12038 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14817) );
  MUX2_X1 U12039 ( .A(n14817), .B(P1_REG1_REG_10__SCAN_IN), .S(n11002), .Z(
        n9936) );
  NOR2_X1 U12040 ( .A1(n9937), .A2(n9936), .ZN(n9935) );
  AOI21_X1 U12041 ( .B1(n11002), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9935), .ZN(
        n9618) );
  NAND2_X1 U12042 ( .A1(n9618), .A2(n9619), .ZN(n9687) );
  OAI21_X1 U12043 ( .B1(n9619), .B2(n9618), .A(n9687), .ZN(n9636) );
  INV_X1 U12044 ( .A(n11099), .ZN(n9693) );
  NAND2_X1 U12045 ( .A1(n10522), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n13904) );
  INV_X1 U12046 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n12112) );
  MUX2_X1 U12047 ( .A(n12112), .B(P1_REG2_REG_7__SCAN_IN), .S(n13897), .Z(
        n13903) );
  AOI21_X1 U12048 ( .B1(n13905), .B2(n13904), .A(n13903), .ZN(n9701) );
  NOR2_X1 U12049 ( .A1(n9620), .A2(n12112), .ZN(n9702) );
  INV_X1 U12050 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9621) );
  MUX2_X1 U12051 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9621), .S(n10596), .Z(n9622) );
  OAI21_X1 U12052 ( .B1(n9701), .B2(n9702), .A(n9622), .ZN(n9706) );
  NAND2_X1 U12053 ( .A1(n10596), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9639) );
  INV_X1 U12054 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9623) );
  MUX2_X1 U12055 ( .A(n9623), .B(P1_REG2_REG_9__SCAN_IN), .S(n10997), .Z(n9638) );
  AOI21_X1 U12056 ( .B1(n9706), .B2(n9639), .A(n9638), .ZN(n9652) );
  AOI21_X1 U12057 ( .B1(n10997), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9652), .ZN(
        n9941) );
  INV_X1 U12058 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9624) );
  MUX2_X1 U12059 ( .A(n9624), .B(P1_REG2_REG_10__SCAN_IN), .S(n11002), .Z(
        n9940) );
  NOR2_X1 U12060 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  NOR2_X1 U12061 ( .A1(n9625), .A2(n9624), .ZN(n9630) );
  INV_X1 U12062 ( .A(n9630), .ZN(n9627) );
  MUX2_X1 U12063 ( .A(n9628), .B(P1_REG2_REG_11__SCAN_IN), .S(n11099), .Z(
        n9626) );
  NAND2_X1 U12064 ( .A1(n9627), .A2(n9626), .ZN(n9631) );
  INV_X1 U12065 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9628) );
  MUX2_X1 U12066 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n9628), .S(n11099), .Z(
        n9629) );
  OAI21_X1 U12067 ( .B1(n9939), .B2(n9630), .A(n9629), .ZN(n9679) );
  OAI211_X1 U12068 ( .C1(n9939), .C2(n9631), .A(n9679), .B(n14690), .ZN(n9634)
         );
  NOR2_X1 U12069 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11504), .ZN(n9632) );
  AOI21_X1 U12070 ( .B1(n14673), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n9632), .ZN(
        n9633) );
  OAI211_X1 U12071 ( .C1(n13955), .C2(n9693), .A(n9634), .B(n9633), .ZN(n9635)
         );
  AOI21_X1 U12072 ( .B1(n14689), .B2(n9636), .A(n9635), .ZN(n9637) );
  INV_X1 U12073 ( .A(n9637), .ZN(P1_U3254) );
  NAND3_X1 U12074 ( .A1(n9706), .A2(n9639), .A3(n9638), .ZN(n9640) );
  NAND2_X1 U12075 ( .A1(n14690), .A2(n9640), .ZN(n9651) );
  NOR2_X1 U12076 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11294), .ZN(n9643) );
  INV_X1 U12077 ( .A(n10997), .ZN(n9641) );
  NOR2_X1 U12078 ( .A1(n13955), .A2(n9641), .ZN(n9642) );
  AOI211_X1 U12079 ( .C1(n14673), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9643), .B(
        n9642), .ZN(n9650) );
  INV_X1 U12080 ( .A(n9644), .ZN(n9648) );
  NOR3_X1 U12081 ( .A1(n9696), .A2(n9646), .A3(n9645), .ZN(n9647) );
  OAI21_X1 U12082 ( .B1(n9648), .B2(n9647), .A(n14689), .ZN(n9649) );
  OAI211_X1 U12083 ( .C1(n9652), .C2(n9651), .A(n9650), .B(n9649), .ZN(
        P1_U3252) );
  AND2_X1 U12084 ( .A1(n10355), .A2(n9653), .ZN(n9673) );
  NAND2_X1 U12085 ( .A1(n9673), .A2(n9654), .ZN(n9666) );
  INV_X1 U12086 ( .A(n9666), .ZN(n9660) );
  INV_X1 U12087 ( .A(n9655), .ZN(n9656) );
  NAND2_X1 U12088 ( .A1(n13572), .A2(n9656), .ZN(n9657) );
  NAND2_X1 U12089 ( .A1(n14799), .A2(n13762), .ZN(n9658) );
  NOR2_X1 U12090 ( .A1(n10353), .A2(n9658), .ZN(n9659) );
  NAND2_X1 U12091 ( .A1(n9660), .A2(n9659), .ZN(n14651) );
  AND2_X2 U12092 ( .A1(n10547), .A2(n9667), .ZN(n9910) );
  NAND2_X1 U12093 ( .A1(n13848), .A2(n11834), .ZN(n9663) );
  AOI22_X1 U12094 ( .A1(n10257), .A2(n12222), .B1(P1_REG1_REG_0__SCAN_IN), 
        .B2(n9661), .ZN(n9662) );
  NAND2_X1 U12095 ( .A1(n9663), .A2(n9662), .ZN(n9717) );
  OAI22_X1 U12096 ( .A1(n14731), .A2(n11904), .B1(n9664), .B2(n9667), .ZN(
        n9665) );
  AOI21_X1 U12097 ( .B1(n12223), .B2(n13848), .A(n9665), .ZN(n9718) );
  XOR2_X1 U12098 ( .A(n9717), .B(n9718), .Z(n13859) );
  NAND2_X1 U12099 ( .A1(n9666), .A2(n10354), .ZN(n9672) );
  AND2_X1 U12100 ( .A1(n9668), .A2(n9667), .ZN(n9669) );
  AND2_X1 U12101 ( .A1(n9670), .A2(n9669), .ZN(n13815) );
  NAND2_X1 U12102 ( .A1(n9672), .A2(n13815), .ZN(n10344) );
  NOR2_X1 U12103 ( .A1(n10344), .A2(P1_U3086), .ZN(n9934) );
  INV_X1 U12104 ( .A(n9934), .ZN(n9675) );
  NOR2_X1 U12105 ( .A1(n10353), .A2(n14799), .ZN(n9671) );
  AND2_X1 U12106 ( .A1(n10358), .A2(n9673), .ZN(n14578) );
  OAI22_X1 U12107 ( .A1(n13567), .A2(n14731), .B1(n14649), .B2(n10360), .ZN(
        n9674) );
  AOI21_X1 U12108 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9675), .A(n9674), .ZN(
        n9676) );
  OAI21_X1 U12109 ( .B1(n14651), .B2(n13859), .A(n9676), .ZN(P1_U3232) );
  INV_X1 U12110 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9678) );
  OAI21_X1 U12111 ( .B1(n9677), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9906) );
  XNOR2_X1 U12112 ( .A(n9906), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11216) );
  MUX2_X1 U12113 ( .A(n9678), .B(P1_REG2_REG_12__SCAN_IN), .S(n11216), .Z(
        n9681) );
  OAI21_X1 U12114 ( .B1(n9628), .B2(n9693), .A(n9679), .ZN(n9680) );
  NOR2_X1 U12115 ( .A1(n9680), .A2(n9681), .ZN(n10040) );
  AOI21_X1 U12116 ( .B1(n9681), .B2(n9680), .A(n10040), .ZN(n9691) );
  INV_X1 U12117 ( .A(n13955), .ZN(n14686) );
  INV_X1 U12118 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9682) );
  NAND2_X1 U12119 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14567)
         );
  OAI21_X1 U12120 ( .B1(n14694), .B2(n9682), .A(n14567), .ZN(n9683) );
  AOI21_X1 U12121 ( .B1(n11216), .B2(n14686), .A(n9683), .ZN(n9690) );
  NAND2_X1 U12122 ( .A1(n9693), .A2(n14612), .ZN(n9685) );
  INV_X1 U12123 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9684) );
  MUX2_X1 U12124 ( .A(n9684), .B(P1_REG1_REG_12__SCAN_IN), .S(n11216), .Z(
        n9686) );
  AOI21_X1 U12125 ( .B1(n9687), .B2(n9685), .A(n9686), .ZN(n10045) );
  AND3_X1 U12126 ( .A1(n9687), .A2(n9686), .A3(n9685), .ZN(n9688) );
  OAI21_X1 U12127 ( .B1(n10045), .B2(n9688), .A(n14689), .ZN(n9689) );
  OAI211_X1 U12128 ( .C1(n9691), .C2(n13956), .A(n9690), .B(n9689), .ZN(
        P1_U3255) );
  INV_X1 U12129 ( .A(n11098), .ZN(n9694) );
  INV_X1 U12130 ( .A(n14888), .ZN(n9957) );
  OAI222_X1 U12131 ( .A1(n13458), .A2(n9692), .B1(n13461), .B2(n9694), .C1(
        P2_U3088), .C2(n9957), .ZN(P2_U3316) );
  OAI222_X1 U12132 ( .A1(n6454), .A2(n9695), .B1(n14286), .B2(n9694), .C1(
        P1_U3086), .C2(n9693), .ZN(P1_U3344) );
  AOI21_X1 U12133 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9709) );
  NOR2_X1 U12134 ( .A1(n10599), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10938) );
  NOR2_X1 U12135 ( .A1(n13955), .A2(n9699), .ZN(n9700) );
  AOI211_X1 U12136 ( .C1(n14673), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10938), .B(
        n9700), .ZN(n9708) );
  INV_X1 U12137 ( .A(n9701), .ZN(n13907) );
  INV_X1 U12138 ( .A(n9702), .ZN(n9704) );
  MUX2_X1 U12139 ( .A(n9621), .B(P1_REG2_REG_8__SCAN_IN), .S(n10596), .Z(n9703) );
  NAND3_X1 U12140 ( .A1(n13907), .A2(n9704), .A3(n9703), .ZN(n9705) );
  NAND3_X1 U12141 ( .A1(n14690), .A2(n9706), .A3(n9705), .ZN(n9707) );
  OAI211_X1 U12142 ( .C1(n9709), .C2(n13913), .A(n9708), .B(n9707), .ZN(
        P1_U3251) );
  INV_X1 U12143 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9729) );
  AOI22_X1 U12144 ( .A1(n13846), .A2(n9910), .B1(n9713), .B2(n6656), .ZN(n9714) );
  XNOR2_X1 U12145 ( .A(n9714), .B(n10393), .ZN(n9917) );
  AND2_X1 U12146 ( .A1(n6656), .A2(n9910), .ZN(n9715) );
  INV_X1 U12147 ( .A(n9716), .ZN(n9919) );
  XNOR2_X1 U12148 ( .A(n9917), .B(n9919), .ZN(n9720) );
  NAND2_X1 U12149 ( .A1(n9719), .A2(n9720), .ZN(n9921) );
  OAI21_X1 U12150 ( .B1(n9720), .B2(n9719), .A(n9921), .ZN(n9721) );
  NAND2_X1 U12151 ( .A1(n9721), .A2(n14576), .ZN(n9728) );
  NAND2_X1 U12152 ( .A1(n10236), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U12153 ( .A1(n9925), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U12154 ( .A1(n10235), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U12155 ( .A1(n14647), .A2(n14645), .ZN(n14746) );
  OR2_X1 U12156 ( .A1(n13762), .A2(n11772), .ZN(n13542) );
  NAND2_X1 U12157 ( .A1(n13848), .A2(n13551), .ZN(n14724) );
  AOI21_X1 U12158 ( .B1(n14746), .B2(n14724), .A(n14649), .ZN(n9726) );
  AOI21_X1 U12159 ( .B1(n14657), .B2(n6656), .A(n9726), .ZN(n9727) );
  OAI211_X1 U12160 ( .C1(n9934), .C2(n9729), .A(n9728), .B(n9727), .ZN(
        P1_U3222) );
  OR2_X1 U12161 ( .A1(n9731), .A2(n9730), .ZN(n9768) );
  NAND2_X1 U12162 ( .A1(n9733), .A2(n9732), .ZN(n9735) );
  AND2_X1 U12163 ( .A1(n9735), .A2(n9734), .ZN(n9766) );
  NAND2_X1 U12164 ( .A1(n9768), .A2(n9766), .ZN(n9736) );
  MUX2_X1 U12165 ( .A(n9736), .B(n12385), .S(n9755), .Z(n15070) );
  INV_X1 U12166 ( .A(n9736), .ZN(n9759) );
  INV_X1 U12167 ( .A(n9737), .ZN(n9738) );
  NAND2_X1 U12168 ( .A1(n9759), .A2(n9738), .ZN(n15091) );
  INV_X1 U12169 ( .A(n15091), .ZN(n12487) );
  XNOR2_X1 U12170 ( .A(n10014), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n9742) );
  INV_X1 U12171 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9988) );
  OAI21_X1 U12172 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n9988), .A(n9762), .ZN(
        n9739) );
  NAND2_X1 U12173 ( .A1(n8158), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U12174 ( .A1(n9739), .A2(n9740), .ZN(n9784) );
  NAND2_X1 U12175 ( .A1(n9742), .A2(n9741), .ZN(n10013) );
  OAI21_X1 U12176 ( .B1(n9742), .B2(n9741), .A(n10013), .ZN(n9758) );
  INV_X1 U12177 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9743) );
  MUX2_X1 U12178 ( .A(n9744), .B(n9743), .S(n12476), .Z(n9745) );
  NAND2_X1 U12179 ( .A1(n9745), .A2(n9762), .ZN(n9753) );
  INV_X1 U12180 ( .A(n9745), .ZN(n9746) );
  NAND2_X1 U12181 ( .A1(n9746), .A2(n9790), .ZN(n9747) );
  AND2_X1 U12182 ( .A1(n9753), .A2(n9747), .ZN(n9779) );
  MUX2_X1 U12183 ( .A(n9988), .B(n11999), .S(n12476), .Z(n9987) );
  AND2_X1 U12184 ( .A1(n9987), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U12185 ( .A1(n9778), .A2(n9753), .ZN(n9751) );
  INV_X1 U12186 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9760) );
  MUX2_X1 U12187 ( .A(n10194), .B(n9760), .S(n12476), .Z(n9748) );
  NAND2_X1 U12188 ( .A1(n9748), .A2(n6450), .ZN(n15010) );
  INV_X1 U12189 ( .A(n9748), .ZN(n9749) );
  NAND2_X1 U12190 ( .A1(n9749), .A2(n9775), .ZN(n9750) );
  AND2_X1 U12191 ( .A1(n15010), .A2(n9750), .ZN(n9752) );
  NAND2_X1 U12192 ( .A1(n9751), .A2(n9752), .ZN(n15011) );
  INV_X1 U12193 ( .A(n9752), .ZN(n9754) );
  NAND3_X1 U12194 ( .A1(n9778), .A2(n9754), .A3(n9753), .ZN(n9756) );
  NOR2_X1 U12195 ( .A1(n12385), .A2(n9755), .ZN(n15055) );
  AOI21_X1 U12196 ( .B1(n15011), .B2(n9756), .A(n15096), .ZN(n9757) );
  AOI21_X1 U12197 ( .B1(n12487), .B2(n9758), .A(n9757), .ZN(n9774) );
  NAND2_X1 U12198 ( .A1(n9759), .A2(n6622), .ZN(n15040) );
  MUX2_X1 U12199 ( .A(n9760), .B(P3_REG1_REG_2__SCAN_IN), .S(n6450), .Z(n9765)
         );
  INV_X1 U12200 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11999) );
  NOR2_X1 U12201 ( .A1(n11999), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9993) );
  INV_X1 U12202 ( .A(n9993), .ZN(n9763) );
  NOR2_X1 U12203 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9763), .ZN(n9761) );
  AOI21_X1 U12204 ( .B1(n9762), .B2(n9763), .A(n9761), .ZN(n9777) );
  NAND2_X1 U12205 ( .A1(n9777), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9776) );
  OAI21_X1 U12206 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n9763), .A(n9776), .ZN(
        n9764) );
  NAND2_X1 U12207 ( .A1(n9765), .A2(n9764), .ZN(n10007) );
  OAI21_X1 U12208 ( .B1(n9765), .B2(n9764), .A(n10007), .ZN(n9772) );
  INV_X1 U12209 ( .A(n9766), .ZN(n9767) );
  NAND2_X1 U12210 ( .A1(n9768), .A2(n9767), .ZN(n15106) );
  INV_X1 U12211 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9770) );
  INV_X1 U12212 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n9769) );
  OAI22_X1 U12213 ( .A1(n15106), .A2(n9770), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9769), .ZN(n9771) );
  AOI21_X1 U12214 ( .B1(n15086), .B2(n9772), .A(n9771), .ZN(n9773) );
  OAI211_X1 U12215 ( .C1(n9775), .C2(n15070), .A(n9774), .B(n9773), .ZN(
        P3_U3184) );
  OAI21_X1 U12216 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n9777), .A(n9776), .ZN(
        n9788) );
  INV_X1 U12217 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n9782) );
  OAI21_X1 U12218 ( .B1(n9986), .B2(n9779), .A(n9778), .ZN(n9780) );
  AOI22_X1 U12219 ( .A1(n15055), .A2(n9780), .B1(P3_REG3_REG_1__SCAN_IN), .B2(
        P3_U3151), .ZN(n9781) );
  OAI21_X1 U12220 ( .B1(n15106), .B2(n9782), .A(n9781), .ZN(n9787) );
  AOI21_X1 U12221 ( .B1(n9744), .B2(n9784), .A(n9783), .ZN(n9785) );
  NOR2_X1 U12222 ( .A1(n15091), .A2(n9785), .ZN(n9786) );
  AOI211_X1 U12223 ( .C1(n15086), .C2(n9788), .A(n9787), .B(n9786), .ZN(n9789)
         );
  OAI21_X1 U12224 ( .B1(n9790), .B2(n15070), .A(n9789), .ZN(P3_U3183) );
  INV_X1 U12225 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n13072) );
  INV_X1 U12226 ( .A(n9823), .ZN(n14844) );
  INV_X1 U12227 ( .A(n13051), .ZN(n9820) );
  INV_X1 U12228 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9791) );
  MUX2_X1 U12229 ( .A(n9791), .B(P2_REG2_REG_2__SCAN_IN), .S(n9818), .Z(n14834) );
  INV_X1 U12230 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9792) );
  MUX2_X1 U12231 ( .A(n9792), .B(P2_REG2_REG_1__SCAN_IN), .S(n9815), .Z(n9870)
         );
  NAND3_X1 U12232 ( .A1(n9870), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n9882) );
  OAI21_X1 U12233 ( .B1(n9792), .B2(n9815), .A(n9882), .ZN(n14835) );
  NAND2_X1 U12234 ( .A1(n14834), .A2(n14835), .ZN(n14833) );
  INV_X1 U12235 ( .A(n9818), .ZN(n14831) );
  NAND2_X1 U12236 ( .A1(n14831), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13059) );
  INV_X1 U12237 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n14950) );
  MUX2_X1 U12238 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n14950), .S(n13051), .Z(
        n13058) );
  AOI21_X1 U12239 ( .B1(n14833), .B2(n13059), .A(n13058), .ZN(n13057) );
  INV_X1 U12240 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9793) );
  MUX2_X1 U12241 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9793), .S(n9823), .Z(n14848) );
  NOR2_X1 U12242 ( .A1(n14849), .A2(n14848), .ZN(n14847) );
  AOI21_X1 U12243 ( .B1(n14844), .B2(P2_REG2_REG_4__SCAN_IN), .A(n14847), .ZN(
        n14865) );
  INV_X1 U12244 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9794) );
  MUX2_X1 U12245 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9794), .S(n14858), .Z(
        n14864) );
  NOR2_X1 U12246 ( .A1(n14865), .A2(n14864), .ZN(n14863) );
  NOR2_X1 U12247 ( .A1(n14858), .A2(n9794), .ZN(n13073) );
  MUX2_X1 U12248 ( .A(n13072), .B(P2_REG2_REG_6__SCAN_IN), .S(n13071), .Z(
        n9795) );
  OAI21_X1 U12249 ( .B1(n13072), .B2(n13071), .A(n13076), .ZN(n14878) );
  INV_X1 U12250 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9796) );
  MUX2_X1 U12251 ( .A(n9796), .B(P2_REG2_REG_7__SCAN_IN), .S(n14873), .Z(n9797) );
  INV_X1 U12252 ( .A(n9797), .ZN(n14877) );
  NAND2_X1 U12253 ( .A1(n14878), .A2(n14877), .ZN(n14876) );
  NAND2_X1 U12254 ( .A1(n14873), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9844) );
  INV_X1 U12255 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9798) );
  MUX2_X1 U12256 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9798), .S(n9829), .Z(n9843)
         );
  AOI21_X1 U12257 ( .B1(n14876), .B2(n9844), .A(n9843), .ZN(n9855) );
  INV_X1 U12258 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9799) );
  MUX2_X1 U12259 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9799), .S(n9864), .Z(n9862)
         );
  NAND2_X1 U12260 ( .A1(n9863), .A2(n9862), .ZN(n9861) );
  OAI21_X1 U12261 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n9864), .A(n9861), .ZN(
        n9807) );
  INV_X1 U12262 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9800) );
  MUX2_X1 U12263 ( .A(n9800), .B(P2_REG2_REG_10__SCAN_IN), .S(n9955), .Z(n9806) );
  NAND2_X1 U12264 ( .A1(n9894), .A2(n9801), .ZN(n9802) );
  AND2_X1 U12265 ( .A1(n9803), .A2(n9802), .ZN(n9805) );
  NOR2_X1 U12266 ( .A1(n8027), .A2(P2_U3088), .ZN(n13450) );
  NAND2_X1 U12267 ( .A1(n9809), .A2(n13450), .ZN(n9835) );
  NOR2_X2 U12268 ( .A1(n9835), .A2(n13455), .ZN(n14931) );
  INV_X1 U12269 ( .A(n14931), .ZN(n14862) );
  NOR2_X1 U12270 ( .A1(n9807), .A2(n9806), .ZN(n9954) );
  AOI211_X1 U12271 ( .C1(n9807), .C2(n9806), .A(n14862), .B(n9954), .ZN(n9814)
         );
  AND2_X1 U12272 ( .A1(n8027), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9808) );
  NAND2_X1 U12273 ( .A1(n9809), .A2(n9808), .ZN(n14937) );
  NOR2_X2 U12274 ( .A1(n9809), .A2(P2_U3088), .ZN(n14929) );
  NAND2_X1 U12275 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11304)
         );
  INV_X1 U12276 ( .A(n11304), .ZN(n9810) );
  AOI21_X1 U12277 ( .B1(n14929), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9810), .ZN(
        n9811) );
  OAI21_X1 U12278 ( .B1(n9812), .B2(n14937), .A(n9811), .ZN(n9813) );
  NOR2_X1 U12279 ( .A1(n9814), .A2(n9813), .ZN(n9839) );
  XNOR2_X1 U12280 ( .A(n9818), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n14829) );
  MUX2_X1 U12281 ( .A(n7470), .B(P2_REG1_REG_1__SCAN_IN), .S(n9815), .Z(n9875)
         );
  AND2_X1 U12282 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9874) );
  NAND2_X1 U12283 ( .A1(n9875), .A2(n9874), .ZN(n9873) );
  INV_X1 U12284 ( .A(n9815), .ZN(n9876) );
  NAND2_X1 U12285 ( .A1(n9876), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9816) );
  NAND2_X1 U12286 ( .A1(n9873), .A2(n9816), .ZN(n14828) );
  NAND2_X1 U12287 ( .A1(n14829), .A2(n14828), .ZN(n14827) );
  INV_X1 U12288 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9817) );
  OR2_X1 U12289 ( .A1(n9818), .A2(n9817), .ZN(n9819) );
  NAND2_X1 U12290 ( .A1(n14827), .A2(n9819), .ZN(n13055) );
  INV_X1 U12291 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n12183) );
  MUX2_X1 U12292 ( .A(n12183), .B(P2_REG1_REG_3__SCAN_IN), .S(n13051), .Z(
        n13056) );
  NAND2_X1 U12293 ( .A1(n13055), .A2(n13056), .ZN(n13054) );
  NAND2_X1 U12294 ( .A1(n9820), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U12295 ( .A1(n13054), .A2(n9821), .ZN(n14840) );
  MUX2_X1 U12296 ( .A(n9822), .B(P2_REG1_REG_4__SCAN_IN), .S(n9823), .Z(n14841) );
  NAND2_X1 U12297 ( .A1(n14840), .A2(n14841), .ZN(n14839) );
  INV_X1 U12298 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9822) );
  OR2_X1 U12299 ( .A1(n9823), .A2(n9822), .ZN(n9824) );
  NAND2_X1 U12300 ( .A1(n14839), .A2(n9824), .ZN(n14855) );
  MUX2_X1 U12301 ( .A(n7539), .B(P2_REG1_REG_5__SCAN_IN), .S(n14858), .Z(
        n14856) );
  NAND2_X1 U12302 ( .A1(n14855), .A2(n14856), .ZN(n14854) );
  OR2_X1 U12303 ( .A1(n14858), .A2(n7539), .ZN(n9825) );
  NAND2_X1 U12304 ( .A1(n14854), .A2(n9825), .ZN(n13069) );
  INV_X1 U12305 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14993) );
  MUX2_X1 U12306 ( .A(n14993), .B(P2_REG1_REG_6__SCAN_IN), .S(n13071), .Z(
        n13070) );
  NAND2_X1 U12307 ( .A1(n13069), .A2(n13070), .ZN(n13068) );
  INV_X1 U12308 ( .A(n13071), .ZN(n9826) );
  NAND2_X1 U12309 ( .A1(n9826), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U12310 ( .A1(n13068), .A2(n9827), .ZN(n14870) );
  INV_X1 U12311 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10926) );
  MUX2_X1 U12312 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10926), .S(n14873), .Z(
        n14871) );
  NAND2_X1 U12313 ( .A1(n14870), .A2(n14871), .ZN(n14869) );
  NAND2_X1 U12314 ( .A1(n14873), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U12315 ( .A1(n14869), .A2(n9828), .ZN(n9850) );
  INV_X1 U12316 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14995) );
  MUX2_X1 U12317 ( .A(n14995), .B(P2_REG1_REG_8__SCAN_IN), .S(n9829), .Z(n9851) );
  NAND2_X1 U12318 ( .A1(n9850), .A2(n9851), .ZN(n9849) );
  NAND2_X1 U12319 ( .A1(n9848), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U12320 ( .A1(n9849), .A2(n9830), .ZN(n9859) );
  INV_X1 U12321 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9831) );
  MUX2_X1 U12322 ( .A(n9831), .B(P2_REG1_REG_9__SCAN_IN), .S(n9864), .Z(n9860)
         );
  OR2_X1 U12323 ( .A1(n9859), .A2(n9860), .ZN(n9857) );
  NAND2_X1 U12324 ( .A1(n9832), .A2(n9831), .ZN(n9833) );
  AND2_X1 U12325 ( .A1(n9857), .A2(n9833), .ZN(n9837) );
  INV_X1 U12326 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n14997) );
  MUX2_X1 U12327 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14997), .S(n9955), .Z(
        n9836) );
  NAND2_X1 U12328 ( .A1(n9837), .A2(n9836), .ZN(n9949) );
  NOR2_X2 U12329 ( .A1(n9835), .A2(n9834), .ZN(n14900) );
  OAI211_X1 U12330 ( .C1(n9837), .C2(n9836), .A(n9949), .B(n14900), .ZN(n9838)
         );
  NAND2_X1 U12331 ( .A1(n9839), .A2(n9838), .ZN(P2_U3224) );
  INV_X1 U12332 ( .A(n11215), .ZN(n9841) );
  INV_X1 U12333 ( .A(n9959), .ZN(n10276) );
  OAI222_X1 U12334 ( .A1(n13467), .A2(n9841), .B1(n10276), .B2(P2_U3088), .C1(
        n9840), .C2(n13458), .ZN(P2_U3315) );
  INV_X1 U12335 ( .A(n11216), .ZN(n10046) );
  OAI222_X1 U12336 ( .A1(n6454), .A2(n9842), .B1(n14286), .B2(n9841), .C1(
        n10046), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND3_X1 U12337 ( .A1(n14876), .A2(n9844), .A3(n9843), .ZN(n9845) );
  NAND2_X1 U12338 ( .A1(n9845), .A2(n14931), .ZN(n9854) );
  INV_X1 U12339 ( .A(n14937), .ZN(n14889) );
  INV_X1 U12340 ( .A(n14929), .ZN(n14897) );
  INV_X1 U12341 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U12342 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11179) );
  OAI21_X1 U12343 ( .B1(n14897), .B2(n9846), .A(n11179), .ZN(n9847) );
  AOI21_X1 U12344 ( .B1(n9848), .B2(n14889), .A(n9847), .ZN(n9853) );
  OAI211_X1 U12345 ( .C1(n9851), .C2(n9850), .A(n14900), .B(n9849), .ZN(n9852)
         );
  OAI211_X1 U12346 ( .C1(n9855), .C2(n9854), .A(n9853), .B(n9852), .ZN(
        P2_U3222) );
  INV_X1 U12347 ( .A(n11375), .ZN(n9908) );
  OAI222_X1 U12348 ( .A1(n13467), .A2(n9908), .B1(n14911), .B2(P2_U3088), .C1(
        n9856), .C2(n13458), .ZN(P2_U3314) );
  INV_X1 U12349 ( .A(n9857), .ZN(n9858) );
  AOI21_X1 U12350 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(n9869) );
  INV_X1 U12351 ( .A(n14900), .ZN(n14923) );
  OAI21_X1 U12352 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9867) );
  INV_X1 U12353 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U12354 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n11279) );
  NAND2_X1 U12355 ( .A1(n14889), .A2(n9864), .ZN(n9865) );
  OAI211_X1 U12356 ( .C1(n14897), .C2(n14428), .A(n11279), .B(n9865), .ZN(
        n9866) );
  AOI21_X1 U12357 ( .B1(n9867), .B2(n14931), .A(n9866), .ZN(n9868) );
  OAI21_X1 U12358 ( .B1(n9869), .B2(n14923), .A(n9868), .ZN(P2_U3223) );
  INV_X1 U12359 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U12360 ( .A1(n14931), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n14820) );
  INV_X1 U12361 ( .A(n9870), .ZN(n9871) );
  OAI22_X1 U12362 ( .A1(n9872), .A2(n14820), .B1(n14862), .B2(n9871), .ZN(
        n9881) );
  INV_X1 U12363 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10373) );
  OAI211_X1 U12364 ( .C1(n9875), .C2(n9874), .A(n14900), .B(n9873), .ZN(n9878)
         );
  NAND2_X1 U12365 ( .A1(n14889), .A2(n9876), .ZN(n9877) );
  OAI211_X1 U12366 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10373), .A(n9878), .B(
        n9877), .ZN(n9880) );
  INV_X1 U12367 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14334) );
  NOR2_X1 U12368 ( .A1(n14334), .A2(n14897), .ZN(n9879) );
  AOI211_X1 U12369 ( .C1(n9882), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9883)
         );
  INV_X1 U12370 ( .A(n9883), .ZN(P2_U3215) );
  OAI21_X1 U12371 ( .B1(n9885), .B2(n14958), .A(n9884), .ZN(n9890) );
  INV_X1 U12372 ( .A(n9886), .ZN(n9887) );
  AND2_X1 U12373 ( .A1(n9888), .A2(n9887), .ZN(n9889) );
  NAND2_X1 U12374 ( .A1(n9890), .A2(n9889), .ZN(n10748) );
  OR2_X1 U12375 ( .A1(n10748), .A2(P2_U3088), .ZN(n10328) );
  INV_X1 U12376 ( .A(n10328), .ZN(n9904) );
  INV_X1 U12377 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9903) );
  INV_X1 U12378 ( .A(n8960), .ZN(n10126) );
  NOR3_X1 U12379 ( .A1(n10126), .A2(n10165), .A3(n6452), .ZN(n9896) );
  INV_X1 U12380 ( .A(n14958), .ZN(n10103) );
  AND2_X1 U12381 ( .A1(n10103), .A2(n14959), .ZN(n9893) );
  NAND2_X1 U12382 ( .A1(n9893), .A2(n9892), .ZN(n9899) );
  OR2_X1 U12383 ( .A1(n13398), .A2(n9894), .ZN(n9895) );
  OAI21_X1 U12384 ( .B1(n10122), .B2(n9896), .A(n12957), .ZN(n9902) );
  AND2_X1 U12385 ( .A1(n13048), .A2(n14481), .ZN(n10106) );
  INV_X1 U12386 ( .A(n14491), .ZN(n12983) );
  OR2_X1 U12387 ( .A1(n9899), .A2(n9898), .ZN(n9900) );
  NAND2_X1 U12388 ( .A1(n9900), .A2(n13295), .ZN(n13014) );
  AOI22_X1 U12389 ( .A1(n10106), .A2(n12983), .B1(n10165), .B2(n13014), .ZN(
        n9901) );
  OAI211_X1 U12390 ( .C1(n9904), .C2(n9903), .A(n9902), .B(n9901), .ZN(
        P2_U3204) );
  NAND2_X1 U12391 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  NAND2_X1 U12392 ( .A1(n9907), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10097) );
  XNOR2_X1 U12393 ( .A(n10097), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11376) );
  INV_X1 U12394 ( .A(n11376), .ZN(n10150) );
  OAI222_X1 U12395 ( .A1(n6454), .A2(n9909), .B1(n14286), .B2(n9908), .C1(
        n10150), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12396 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U12397 ( .A1(n14647), .A2(n11966), .ZN(n9915) );
  NAND2_X1 U12398 ( .A1(n11842), .A2(n13868), .ZN(n9911) );
  NAND2_X1 U12399 ( .A1(n6453), .A2(n12222), .ZN(n9914) );
  NAND2_X1 U12400 ( .A1(n9915), .A2(n9914), .ZN(n9916) );
  XNOR2_X1 U12401 ( .A(n9916), .B(n10393), .ZN(n10333) );
  AOI22_X1 U12402 ( .A1(n12223), .A2(n14647), .B1(n11966), .B2(n6453), .ZN(
        n10331) );
  XNOR2_X1 U12403 ( .A(n10333), .B(n10331), .ZN(n9923) );
  INV_X1 U12404 ( .A(n9917), .ZN(n9918) );
  NAND2_X1 U12405 ( .A1(n9921), .A2(n9920), .ZN(n9922) );
  NAND2_X1 U12406 ( .A1(n9922), .A2(n9923), .ZN(n10332) );
  OAI21_X1 U12407 ( .B1(n9923), .B2(n9922), .A(n10332), .ZN(n9924) );
  NAND2_X1 U12408 ( .A1(n9924), .A2(n14576), .ZN(n9933) );
  NAND2_X1 U12409 ( .A1(n13846), .A2(n13551), .ZN(n9931) );
  NAND2_X1 U12410 ( .A1(n10236), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9929) );
  INV_X1 U12411 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14710) );
  NAND2_X1 U12412 ( .A1(n12050), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9927) );
  NAND2_X1 U12413 ( .A1(n10235), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9926) );
  NAND4_X2 U12414 ( .A1(n9929), .A2(n9928), .A3(n9927), .A4(n9926), .ZN(n13845) );
  NAND2_X1 U12415 ( .A1(n13845), .A2(n14645), .ZN(n9930) );
  NAND2_X1 U12416 ( .A1(n9931), .A2(n9930), .ZN(n10575) );
  AOI22_X1 U12417 ( .A1(n14657), .A2(n6453), .B1(n14578), .B2(n10575), .ZN(
        n9932) );
  OAI211_X1 U12418 ( .C1(n9934), .C2(n10583), .A(n9933), .B(n9932), .ZN(
        P1_U3237) );
  AOI211_X1 U12419 ( .C1(n9937), .C2(n9936), .A(n13913), .B(n9935), .ZN(n9938)
         );
  AOI21_X1 U12420 ( .B1(n14686), .B2(n11002), .A(n9938), .ZN(n9946) );
  AND2_X1 U12421 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11358) );
  AOI211_X1 U12422 ( .C1(n9941), .C2(n9940), .A(n13956), .B(n9939), .ZN(n9942)
         );
  INV_X1 U12423 ( .A(n9942), .ZN(n9943) );
  OAI21_X1 U12424 ( .B1(n6808), .B2(n14694), .A(n9943), .ZN(n9944) );
  NOR2_X1 U12425 ( .A1(n11358), .A2(n9944), .ZN(n9945) );
  NAND2_X1 U12426 ( .A1(n9946), .A2(n9945), .ZN(P1_U3253) );
  OR2_X1 U12427 ( .A1(n9959), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U12428 ( .A1(n9959), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U12429 ( .A1(n10282), .A2(n9947), .ZN(n9953) );
  NAND2_X1 U12430 ( .A1(n9955), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12431 ( .A1(n9949), .A2(n9948), .ZN(n14884) );
  INV_X1 U12432 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15000) );
  MUX2_X1 U12433 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n15000), .S(n14888), .Z(
        n14883) );
  NAND2_X1 U12434 ( .A1(n14884), .A2(n14883), .ZN(n14882) );
  NAND2_X1 U12435 ( .A1(n14888), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12436 ( .A1(n14882), .A2(n9950), .ZN(n9952) );
  INV_X1 U12437 ( .A(n10283), .ZN(n9951) );
  AOI21_X1 U12438 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9968) );
  INV_X1 U12439 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9956) );
  MUX2_X1 U12440 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9956), .S(n14888), .Z(
        n14892) );
  NAND2_X1 U12441 ( .A1(n14891), .A2(n14892), .ZN(n14890) );
  NAND2_X1 U12442 ( .A1(n9957), .A2(n9956), .ZN(n9962) );
  INV_X1 U12443 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9958) );
  OR2_X1 U12444 ( .A1(n9959), .A2(n9958), .ZN(n9961) );
  NAND2_X1 U12445 ( .A1(n9959), .A2(n9958), .ZN(n9960) );
  AND2_X1 U12446 ( .A1(n9961), .A2(n9960), .ZN(n9963) );
  AOI21_X1 U12447 ( .B1(n14890), .B2(n9962), .A(n9963), .ZN(n10275) );
  AND3_X1 U12448 ( .A1(n14890), .A2(n9963), .A3(n9962), .ZN(n9964) );
  OAI21_X1 U12449 ( .B1(n10275), .B2(n9964), .A(n14931), .ZN(n9967) );
  AND2_X1 U12450 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11576) );
  NOR2_X1 U12451 ( .A1(n14937), .A2(n10276), .ZN(n9965) );
  AOI211_X1 U12452 ( .C1(n14929), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n11576), 
        .B(n9965), .ZN(n9966) );
  OAI211_X1 U12453 ( .C1(n9968), .C2(n14923), .A(n9967), .B(n9966), .ZN(
        P2_U3226) );
  INV_X1 U12454 ( .A(n9969), .ZN(n9974) );
  NAND2_X1 U12455 ( .A1(n9971), .A2(n9970), .ZN(n9972) );
  NAND2_X1 U12456 ( .A1(n12820), .A2(n9972), .ZN(n9973) );
  OAI21_X1 U12457 ( .B1(n12820), .B2(n9974), .A(n9973), .ZN(n9975) );
  INV_X1 U12458 ( .A(n9975), .ZN(n9976) );
  NAND2_X1 U12459 ( .A1(n9977), .A2(n9976), .ZN(n9983) );
  NAND2_X1 U12460 ( .A1(n15109), .A2(n14467), .ZN(n9978) );
  AOI22_X1 U12461 ( .A1(n14463), .A2(n10114), .B1(n12687), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n9985) );
  AND2_X1 U12462 ( .A1(n9979), .A2(n12680), .ZN(n9980) );
  OR2_X1 U12463 ( .A1(n10116), .A2(n9980), .ZN(n9982) );
  NAND2_X1 U12464 ( .A1(n12384), .A2(n12666), .ZN(n9981) );
  AND2_X1 U12465 ( .A1(n9982), .A2(n9981), .ZN(n11998) );
  MUX2_X1 U12466 ( .A(n9988), .B(n11998), .S(n15117), .Z(n9984) );
  NAND2_X1 U12467 ( .A1(n9985), .A2(n9984), .ZN(P3_U3233) );
  NOR3_X1 U12468 ( .A1(n12487), .A2(n15086), .A3(n15055), .ZN(n9997) );
  INV_X1 U12469 ( .A(n9986), .ZN(n9996) );
  OAI22_X1 U12470 ( .A1(n15091), .A2(n9988), .B1(n9987), .B2(n15096), .ZN(
        n9989) );
  INV_X1 U12471 ( .A(n15070), .ZN(n15102) );
  MUX2_X1 U12472 ( .A(n9989), .B(n15102), .S(P3_IR_REG_0__SCAN_IN), .Z(n9990)
         );
  INV_X1 U12473 ( .A(n9990), .ZN(n9995) );
  INV_X1 U12474 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n9991) );
  INV_X1 U12475 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n12203) );
  OAI22_X1 U12476 ( .A1(n15106), .A2(n9991), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12203), .ZN(n9992) );
  AOI21_X1 U12477 ( .B1(n15086), .B2(n9993), .A(n9992), .ZN(n9994) );
  OAI211_X1 U12478 ( .C1(n9997), .C2(n9996), .A(n9995), .B(n9994), .ZN(
        P3_U3182) );
  MUX2_X1 U12479 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n6622), .Z(n10054) );
  XNOR2_X1 U12480 ( .A(n10054), .B(n10060), .ZN(n10056) );
  INV_X1 U12481 ( .A(n15033), .ZN(n10019) );
  MUX2_X1 U12482 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12476), .Z(n10004) );
  INV_X1 U12483 ( .A(n10004), .ZN(n10005) );
  NAND2_X1 U12484 ( .A1(n15011), .A2(n15010), .ZN(n10002) );
  MUX2_X1 U12485 ( .A(n9998), .B(n12154), .S(n12476), .Z(n9999) );
  NAND2_X1 U12486 ( .A1(n9999), .A2(n15016), .ZN(n10003) );
  INV_X1 U12487 ( .A(n9999), .ZN(n10000) );
  NAND2_X1 U12488 ( .A1(n10000), .A2(n10015), .ZN(n10001) );
  AND2_X1 U12489 ( .A1(n10003), .A2(n10001), .ZN(n15008) );
  NAND2_X1 U12490 ( .A1(n10002), .A2(n15008), .ZN(n15013) );
  NAND2_X1 U12491 ( .A1(n15013), .A2(n10003), .ZN(n15027) );
  XNOR2_X1 U12492 ( .A(n10004), .B(n10019), .ZN(n15026) );
  AND2_X1 U12493 ( .A1(n15027), .A2(n15026), .ZN(n15029) );
  INV_X1 U12494 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15057) );
  MUX2_X1 U12495 ( .A(n10474), .B(n15057), .S(n6622), .Z(n10006) );
  NOR2_X1 U12496 ( .A1(n10006), .A2(n10010), .ZN(n15046) );
  NAND2_X1 U12497 ( .A1(n10006), .A2(n10010), .ZN(n15047) );
  OAI21_X1 U12498 ( .B1(n15050), .B2(n15046), .A(n15047), .ZN(n10057) );
  XOR2_X1 U12499 ( .A(n10056), .B(n10057), .Z(n10029) );
  INV_X1 U12500 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10009) );
  OAI21_X1 U12501 ( .B1(n6450), .B2(n9760), .A(n10007), .ZN(n10008) );
  XNOR2_X1 U12502 ( .A(n10008), .B(n15016), .ZN(n15017) );
  AOI22_X1 U12503 ( .A1(n15017), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n10015), 
        .B2(n10008), .ZN(n15038) );
  MUX2_X1 U12504 ( .A(n10009), .B(P3_REG1_REG_4__SCAN_IN), .S(n15033), .Z(
        n15037) );
  INV_X1 U12505 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U12506 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n10065), .B1(n10060), 
        .B2(n10059), .ZN(n10011) );
  NAND2_X1 U12507 ( .A1(n10011), .A2(n10012), .ZN(n10058) );
  OAI21_X1 U12508 ( .B1(n10012), .B2(n10011), .A(n10058), .ZN(n10027) );
  OAI21_X1 U12509 ( .B1(n6450), .B2(n10194), .A(n10013), .ZN(n10016) );
  INV_X1 U12510 ( .A(n10016), .ZN(n10017) );
  XNOR2_X1 U12511 ( .A(n10016), .B(n10015), .ZN(n15005) );
  OAI21_X1 U12512 ( .B1(n10017), .B2(n15016), .A(n15003), .ZN(n15024) );
  MUX2_X1 U12513 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10018), .S(n15033), .Z(
        n15023) );
  XNOR2_X1 U12514 ( .A(n10020), .B(n15053), .ZN(n15045) );
  AOI22_X1 U12515 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10060), .B1(n10065), 
        .B2(n10570), .ZN(n10021) );
  AOI21_X1 U12516 ( .B1(n10022), .B2(n10021), .A(n10064), .ZN(n10025) );
  NAND2_X1 U12517 ( .A1(n15102), .A2(n10060), .ZN(n10024) );
  INV_X1 U12518 ( .A(n15106), .ZN(n15075) );
  AND2_X1 U12519 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10779) );
  AOI21_X1 U12520 ( .B1(n15075), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10779), .ZN(
        n10023) );
  OAI211_X1 U12521 ( .C1(n10025), .C2(n15091), .A(n10024), .B(n10023), .ZN(
        n10026) );
  AOI21_X1 U12522 ( .B1(n15086), .B2(n10027), .A(n10026), .ZN(n10028) );
  OAI21_X1 U12523 ( .B1(n10029), .B2(n15096), .A(n10028), .ZN(P3_U3188) );
  NOR3_X1 U12524 ( .A1(n10030), .A2(n9261), .A3(n12764), .ZN(n10032) );
  AOI211_X1 U12525 ( .C1(n10034), .C2(n10033), .A(n10032), .B(n10031), .ZN(
        n10039) );
  INV_X1 U12526 ( .A(n12356), .ZN(n11345) );
  NAND2_X1 U12527 ( .A1(n11345), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10111) );
  AOI22_X1 U12528 ( .A1(n12311), .A2(n12383), .B1(n12352), .B2(n12757), .ZN(
        n10035) );
  OAI21_X1 U12529 ( .B1(n10036), .B2(n12360), .A(n10035), .ZN(n10037) );
  AOI21_X1 U12530 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n10111), .A(n10037), .ZN(
        n10038) );
  OAI21_X1 U12531 ( .B1(n10039), .B2(n12347), .A(n10038), .ZN(P3_U3162) );
  AOI21_X1 U12532 ( .B1(n9678), .B2(n10046), .A(n10040), .ZN(n10044) );
  INV_X1 U12533 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11396) );
  MUX2_X1 U12534 ( .A(n11396), .B(P1_REG2_REG_13__SCAN_IN), .S(n11376), .Z(
        n10041) );
  INV_X1 U12535 ( .A(n10041), .ZN(n10043) );
  MUX2_X1 U12536 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11396), .S(n11376), .Z(
        n10042) );
  NAND2_X1 U12537 ( .A1(n10044), .A2(n10042), .ZN(n10144) );
  OAI211_X1 U12538 ( .C1(n10044), .C2(n10043), .A(n10144), .B(n14690), .ZN(
        n10053) );
  NAND2_X1 U12539 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11736)
         );
  AOI21_X1 U12540 ( .B1(n9684), .B2(n10046), .A(n10045), .ZN(n10049) );
  INV_X1 U12541 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10047) );
  MUX2_X1 U12542 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10047), .S(n11376), .Z(
        n10048) );
  NAND2_X1 U12543 ( .A1(n10049), .A2(n10048), .ZN(n10149) );
  OAI211_X1 U12544 ( .C1(n10049), .C2(n10048), .A(n14689), .B(n10149), .ZN(
        n10050) );
  NAND2_X1 U12545 ( .A1(n11736), .A2(n10050), .ZN(n10051) );
  AOI21_X1 U12546 ( .B1(n14673), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10051), 
        .ZN(n10052) );
  OAI211_X1 U12547 ( .C1(n13955), .C2(n10150), .A(n10053), .B(n10052), .ZN(
        P1_U3256) );
  MUX2_X1 U12548 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n6622), .Z(n10294) );
  XNOR2_X1 U12549 ( .A(n10294), .B(n10298), .ZN(n10295) );
  INV_X1 U12550 ( .A(n10054), .ZN(n10055) );
  AOI22_X1 U12551 ( .A1(n10057), .A2(n10056), .B1(n10060), .B2(n10055), .ZN(
        n10296) );
  XOR2_X1 U12552 ( .A(n10296), .B(n10295), .Z(n10072) );
  OAI21_X1 U12553 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10061), .A(n10299), .ZN(
        n10070) );
  NOR2_X1 U12554 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10062), .ZN(n10864) );
  AOI21_X1 U12555 ( .B1(n15075), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10864), .ZN(
        n10063) );
  OAI21_X1 U12556 ( .B1(n15070), .B2(n10298), .A(n10063), .ZN(n10069) );
  INV_X1 U12557 ( .A(n10298), .ZN(n10305) );
  NOR2_X1 U12558 ( .A1(n8238), .A2(n10066), .ZN(n10306) );
  AOI21_X1 U12559 ( .B1(n10066), .B2(n8238), .A(n10306), .ZN(n10067) );
  NOR2_X1 U12560 ( .A1(n10067), .A2(n15091), .ZN(n10068) );
  AOI211_X1 U12561 ( .C1(n15086), .C2(n10070), .A(n10069), .B(n10068), .ZN(
        n10071) );
  OAI21_X1 U12562 ( .B1(n10072), .B2(n15096), .A(n10071), .ZN(P3_U3189) );
  OAI222_X1 U12563 ( .A1(n12517), .A2(P3_U3151), .B1(n12832), .B2(n10074), 
        .C1(n10073), .C2(n12829), .ZN(P3_U3276) );
  XOR2_X1 U12564 ( .A(n10076), .B(n10075), .Z(n10081) );
  AOI22_X1 U12565 ( .A1(n12311), .A2(n12382), .B1(n12352), .B2(n12384), .ZN(
        n10077) );
  OAI21_X1 U12566 ( .B1(n10078), .B2(n12360), .A(n10077), .ZN(n10079) );
  AOI21_X1 U12567 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10111), .A(n10079), .ZN(
        n10080) );
  OAI21_X1 U12568 ( .B1(n10081), .B2(n12347), .A(n10080), .ZN(P3_U3177) );
  OAI21_X1 U12569 ( .B1(n10083), .B2(n10084), .A(n10082), .ZN(n10217) );
  NAND2_X1 U12570 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  NAND3_X1 U12571 ( .A1(n10087), .A2(n12762), .A3(n10086), .ZN(n10090) );
  OAI22_X1 U12572 ( .A1(n12760), .A2(n12683), .B1(n10638), .B2(n12759), .ZN(
        n10088) );
  INV_X1 U12573 ( .A(n10088), .ZN(n10089) );
  NAND2_X1 U12574 ( .A1(n10090), .A2(n10089), .ZN(n10214) );
  AOI21_X1 U12575 ( .B1(n14475), .B2(n10217), .A(n10214), .ZN(n10095) );
  INV_X1 U12576 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U12577 ( .A1(n8743), .A2(n10091), .B1(n15131), .B2(
        P3_REG1_REG_3__SCAN_IN), .ZN(n10092) );
  OAI21_X1 U12578 ( .B1(n10095), .B2(n15131), .A(n10092), .ZN(P3_U3462) );
  OAI22_X1 U12579 ( .A1(n10385), .A2(n12818), .B1(n15129), .B2(n8164), .ZN(
        n10093) );
  INV_X1 U12580 ( .A(n10093), .ZN(n10094) );
  OAI21_X1 U12581 ( .B1(n10095), .B2(n15127), .A(n10094), .ZN(P3_U3399) );
  INV_X1 U12582 ( .A(n11523), .ZN(n10101) );
  NAND2_X1 U12583 ( .A1(n10097), .A2(n10096), .ZN(n10098) );
  NAND2_X1 U12584 ( .A1(n10098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10099) );
  XNOR2_X1 U12585 ( .A(n10099), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11524) );
  INV_X1 U12586 ( .A(n11524), .ZN(n10157) );
  OAI222_X1 U12587 ( .A1(n6454), .A2(n10100), .B1(n14286), .B2(n10101), .C1(
        P1_U3086), .C2(n10157), .ZN(P1_U3341) );
  OAI222_X1 U12588 ( .A1(n13458), .A2(n10102), .B1(n13461), .B2(n10101), .C1(
        P2_U3088), .C2(n6659), .ZN(P2_U3313) );
  AOI21_X1 U12589 ( .B1(n13371), .B2(n11255), .A(n10444), .ZN(n10107) );
  NOR2_X1 U12590 ( .A1(n10107), .A2(n10106), .ZN(n10439) );
  NAND2_X1 U12591 ( .A1(n10165), .A2(n10108), .ZN(n10440) );
  OAI211_X1 U12592 ( .C1(n10444), .C2(n11311), .A(n10439), .B(n10440), .ZN(
        n10117) );
  NAND2_X1 U12593 ( .A1(n10117), .A2(n10105), .ZN(n10109) );
  OAI21_X1 U12594 ( .B1(n10105), .B2(n10110), .A(n10109), .ZN(P2_U3430) );
  NAND2_X1 U12595 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(n10111), .ZN(n10112) );
  OAI21_X1 U12596 ( .B1(n12354), .B2(n9265), .A(n10112), .ZN(n10113) );
  AOI21_X1 U12597 ( .B1(n12334), .B2(n10114), .A(n10113), .ZN(n10115) );
  OAI21_X1 U12598 ( .B1(n10116), .B2(n12347), .A(n10115), .ZN(P3_U3172) );
  NAND2_X1 U12599 ( .A1(n10117), .A2(n15002), .ZN(n10118) );
  OAI21_X1 U12600 ( .B1(n15002), .B2(n10119), .A(n10118), .ZN(P2_U3499) );
  XNOR2_X1 U12601 ( .A(n10121), .B(n12915), .ZN(n10317) );
  NAND2_X1 U12602 ( .A1(n13048), .A2(n12834), .ZN(n10319) );
  AOI21_X1 U12603 ( .B1(n10124), .B2(n10123), .A(n10318), .ZN(n10129) );
  INV_X1 U12604 ( .A(n8973), .ZN(n10125) );
  OAI22_X1 U12605 ( .A1(n10126), .A2(n12900), .B1(n10125), .B2(n12898), .ZN(
        n10163) );
  AOI22_X1 U12606 ( .A1(n10163), .A2(n12983), .B1(n10121), .B2(n13014), .ZN(
        n10128) );
  NAND2_X1 U12607 ( .A1(n10328), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n10127) );
  OAI211_X1 U12608 ( .C1(n10129), .C2(n14490), .A(n10128), .B(n10127), .ZN(
        P2_U3194) );
  OAI211_X1 U12609 ( .C1(n10132), .C2(n10131), .A(n10130), .B(n12762), .ZN(
        n10134) );
  AOI22_X1 U12610 ( .A1(n12666), .A2(n12380), .B1(n12382), .B2(n12756), .ZN(
        n10133) );
  NAND2_X1 U12611 ( .A1(n10134), .A2(n10133), .ZN(n10197) );
  INV_X1 U12612 ( .A(n10197), .ZN(n10143) );
  NOR2_X1 U12613 ( .A1(n15109), .A2(n10500), .ZN(n10135) );
  NAND2_X1 U12614 ( .A1(n15117), .A2(n10135), .ZN(n15114) );
  INV_X1 U12615 ( .A(n12766), .ZN(n12596) );
  NAND2_X1 U12616 ( .A1(n15117), .A2(n12596), .ZN(n10136) );
  OAI21_X1 U12617 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(n10198) );
  AOI22_X1 U12618 ( .A1(n14463), .A2(n10199), .B1(n12687), .B2(n10460), .ZN(
        n10140) );
  OAI21_X1 U12619 ( .B1(n10018), .B2(n15117), .A(n10140), .ZN(n10141) );
  AOI21_X1 U12620 ( .B1(n12691), .B2(n10198), .A(n10141), .ZN(n10142) );
  OAI21_X1 U12621 ( .B1(n15119), .B2(n10143), .A(n10142), .ZN(P3_U3229) );
  OAI21_X1 U12622 ( .B1(n11396), .B2(n10150), .A(n10144), .ZN(n10148) );
  INV_X1 U12623 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10145) );
  MUX2_X1 U12624 ( .A(n10145), .B(P1_REG2_REG_14__SCAN_IN), .S(n11524), .Z(
        n10146) );
  INV_X1 U12625 ( .A(n10146), .ZN(n10147) );
  NAND2_X1 U12626 ( .A1(n10147), .A2(n10148), .ZN(n10684) );
  OAI211_X1 U12627 ( .C1(n10148), .C2(n10147), .A(n14690), .B(n10684), .ZN(
        n10156) );
  NAND2_X1 U12628 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14559)
         );
  INV_X1 U12629 ( .A(n14559), .ZN(n10154) );
  INV_X1 U12630 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14606) );
  NOR2_X1 U12631 ( .A1(n10157), .A2(n14606), .ZN(n10692) );
  AOI21_X1 U12632 ( .B1(n14606), .B2(n10157), .A(n10692), .ZN(n10152) );
  OAI21_X1 U12633 ( .B1(n10047), .B2(n10150), .A(n10149), .ZN(n10691) );
  OAI21_X1 U12634 ( .B1(n10152), .B2(n10691), .A(n14689), .ZN(n10151) );
  AOI21_X1 U12635 ( .B1(n10152), .B2(n10691), .A(n10151), .ZN(n10153) );
  AOI211_X1 U12636 ( .C1(n14673), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n10154), 
        .B(n10153), .ZN(n10155) );
  OAI211_X1 U12637 ( .C1(n13955), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        P1_U3257) );
  INV_X1 U12638 ( .A(n10159), .ZN(n10160) );
  AOI21_X1 U12639 ( .B1(n7484), .B2(n10162), .A(n10160), .ZN(n10379) );
  XNOR2_X1 U12640 ( .A(n10162), .B(n10161), .ZN(n10164) );
  AOI21_X1 U12641 ( .B1(n10164), .B2(n14535), .A(n10163), .ZN(n10372) );
  AOI211_X1 U12642 ( .C1(n10165), .C2(n10121), .A(n13217), .B(n8035), .ZN(
        n10376) );
  INV_X1 U12643 ( .A(n10376), .ZN(n10166) );
  OAI211_X1 U12644 ( .C1(n10379), .C2(n14530), .A(n10372), .B(n10166), .ZN(
        n10171) );
  NAND2_X1 U12645 ( .A1(n10105), .A2(n13398), .ZN(n13431) );
  INV_X1 U12646 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10167) );
  OAI22_X1 U12647 ( .A1(n13431), .A2(n10374), .B1(n10105), .B2(n10167), .ZN(
        n10168) );
  AOI21_X1 U12648 ( .B1(n10171), .B2(n10105), .A(n10168), .ZN(n10169) );
  INV_X1 U12649 ( .A(n10169), .ZN(P2_U3433) );
  OAI22_X1 U12650 ( .A1(n13378), .A2(n10374), .B1(n15002), .B2(n7470), .ZN(
        n10170) );
  AOI21_X1 U12651 ( .B1(n10171), .B2(n15002), .A(n10170), .ZN(n10172) );
  INV_X1 U12652 ( .A(n10172), .ZN(P2_U3500) );
  INV_X1 U12653 ( .A(n11581), .ZN(n10177) );
  AND2_X1 U12654 ( .A1(n10174), .A2(n10173), .ZN(n10434) );
  OR2_X1 U12655 ( .A1(n10434), .A2(n14272), .ZN(n10175) );
  XNOR2_X1 U12656 ( .A(n10175), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14687) );
  INV_X1 U12657 ( .A(n14687), .ZN(n10693) );
  OAI222_X1 U12658 ( .A1(n6454), .A2(n10176), .B1(n14286), .B2(n10177), .C1(
        P1_U3086), .C2(n10693), .ZN(P1_U3340) );
  INV_X1 U12659 ( .A(n13096), .ZN(n14921) );
  OAI222_X1 U12660 ( .A1(n13458), .A2(n10178), .B1(n13467), .B2(n10177), .C1(
        P2_U3088), .C2(n14921), .ZN(P2_U3312) );
  OR2_X1 U12661 ( .A1(n10180), .A2(n10179), .ZN(n10181) );
  NAND2_X1 U12662 ( .A1(n10182), .A2(n10181), .ZN(n15122) );
  INV_X1 U12663 ( .A(n15122), .ZN(n10196) );
  NAND2_X1 U12664 ( .A1(n10183), .A2(n14467), .ZN(n15123) );
  NOR2_X1 U12665 ( .A1(n15123), .A2(n10184), .ZN(n10192) );
  XNOR2_X1 U12666 ( .A(n10186), .B(n10185), .ZN(n10187) );
  NAND2_X1 U12667 ( .A1(n10187), .A2(n12762), .ZN(n10191) );
  NAND2_X1 U12668 ( .A1(n15122), .A2(n12596), .ZN(n10190) );
  OAI22_X1 U12669 ( .A1(n9265), .A2(n12683), .B1(n10466), .B2(n12759), .ZN(
        n10188) );
  INV_X1 U12670 ( .A(n10188), .ZN(n10189) );
  NAND3_X1 U12671 ( .A1(n10191), .A2(n10190), .A3(n10189), .ZN(n15126) );
  AOI211_X1 U12672 ( .C1(n12687), .C2(P3_REG3_REG_2__SCAN_IN), .A(n10192), .B(
        n15126), .ZN(n10193) );
  MUX2_X1 U12673 ( .A(n10194), .B(n10193), .S(n15117), .Z(n10195) );
  OAI21_X1 U12674 ( .B1(n10196), .B2(n15114), .A(n10195), .ZN(P3_U3231) );
  AOI21_X1 U12675 ( .B1(n14475), .B2(n10198), .A(n10197), .ZN(n10203) );
  AOI22_X1 U12676 ( .A1(n8743), .A2(n10199), .B1(n15131), .B2(
        P3_REG1_REG_4__SCAN_IN), .ZN(n10200) );
  OAI21_X1 U12677 ( .B1(n10203), .B2(n15131), .A(n10200), .ZN(P3_U3463) );
  OAI22_X1 U12678 ( .A1(n10467), .A2(n12818), .B1(n15129), .B2(n8183), .ZN(
        n10201) );
  INV_X1 U12679 ( .A(n10201), .ZN(n10202) );
  OAI21_X1 U12680 ( .B1(n10203), .B2(n15127), .A(n10202), .ZN(P3_U3402) );
  OAI21_X1 U12681 ( .B1(n10205), .B2(n10207), .A(n10204), .ZN(n10448) );
  INV_X1 U12682 ( .A(n8035), .ZN(n10206) );
  AOI211_X1 U12683 ( .C1(n10321), .C2(n10206), .A(n13217), .B(n10405), .ZN(
        n10454) );
  XNOR2_X1 U12684 ( .A(n10208), .B(n10207), .ZN(n10209) );
  AOI22_X1 U12685 ( .A1(n14484), .A2(n13048), .B1(n13047), .B2(n14481), .ZN(
        n10326) );
  OAI21_X1 U12686 ( .B1(n10209), .B2(n13371), .A(n10326), .ZN(n10449) );
  AOI211_X1 U12687 ( .C1(n14983), .C2(n10448), .A(n10454), .B(n10449), .ZN(
        n10213) );
  AOI22_X1 U12688 ( .A1(n8070), .A2(n10321), .B1(P2_REG1_REG_2__SCAN_IN), .B2(
        n14999), .ZN(n10210) );
  OAI21_X1 U12689 ( .B1(n10213), .B2(n14999), .A(n10210), .ZN(P2_U3501) );
  OAI22_X1 U12690 ( .A1(n13431), .A2(n10450), .B1(n10105), .B2(n7488), .ZN(
        n10211) );
  INV_X1 U12691 ( .A(n10211), .ZN(n10212) );
  OAI21_X1 U12692 ( .B1(n10213), .B2(n14991), .A(n10212), .ZN(P2_U3436) );
  OAI22_X1 U12693 ( .A1(n12689), .A2(n10385), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15111), .ZN(n10216) );
  MUX2_X1 U12694 ( .A(n10214), .B(P3_REG2_REG_3__SCAN_IN), .S(n15119), .Z(
        n10215) );
  AOI211_X1 U12695 ( .C1(n12691), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10218) );
  INV_X1 U12696 ( .A(n10218), .ZN(P3_U3230) );
  AND2_X2 U12697 ( .A1(n10219), .A2(n10355), .ZN(n14819) );
  INV_X1 U12698 ( .A(n14722), .ZN(n10221) );
  NAND2_X1 U12699 ( .A1(n10256), .A2(n10221), .ZN(n10223) );
  NAND2_X1 U12700 ( .A1(n6665), .A2(n6656), .ZN(n10222) );
  NAND2_X1 U12701 ( .A1(n10223), .A2(n10222), .ZN(n10574) );
  NAND2_X1 U12702 ( .A1(n10574), .A2(n13777), .ZN(n10225) );
  INV_X1 U12703 ( .A(n14647), .ZN(n13580) );
  NAND2_X1 U12704 ( .A1(n13580), .A2(n6453), .ZN(n10224) );
  NAND2_X1 U12705 ( .A1(n10225), .A2(n10224), .ZN(n14705) );
  NAND2_X1 U12706 ( .A1(n6459), .A2(n13885), .ZN(n10226) );
  XNOR2_X2 U12707 ( .A(n13845), .B(n6457), .ZN(n14706) );
  INV_X1 U12708 ( .A(n13845), .ZN(n10336) );
  NAND2_X1 U12709 ( .A1(n10336), .A2(n6457), .ZN(n10230) );
  NOR2_X1 U12710 ( .A1(n10231), .A2(n6451), .ZN(n10234) );
  OAI22_X1 U12711 ( .A1(n13758), .A2(n10232), .B1(n11895), .B2(n14665), .ZN(
        n10233) );
  NAND2_X1 U12712 ( .A1(n10235), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10241) );
  NAND2_X1 U12713 ( .A1(n13730), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10240) );
  INV_X1 U12714 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n12111) );
  NAND2_X1 U12715 ( .A1(n14710), .A2(n12111), .ZN(n10237) );
  NAND2_X1 U12716 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10245) );
  AND2_X1 U12717 ( .A1(n10237), .A2(n10245), .ZN(n10345) );
  NAND2_X1 U12718 ( .A1(n12027), .A2(n10345), .ZN(n10239) );
  NAND2_X1 U12719 ( .A1(n12050), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10238) );
  NOR2_X1 U12720 ( .A1(n14768), .A2(n14646), .ZN(n10243) );
  NAND2_X1 U12721 ( .A1(n14768), .A2(n14646), .ZN(n10242) );
  NAND2_X1 U12722 ( .A1(n13730), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U12723 ( .A1(n12050), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10249) );
  INV_X1 U12724 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10244) );
  AND2_X1 U12725 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  NOR2_X1 U12726 ( .A1(n10260), .A2(n10246), .ZN(n10552) );
  NAND2_X1 U12727 ( .A1(n12027), .A2(n10552), .ZN(n10248) );
  NAND2_X1 U12728 ( .A1(n6456), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10247) );
  OR2_X1 U12729 ( .A1(n10251), .A2(n6451), .ZN(n10255) );
  INV_X4 U12730 ( .A(n13758), .ZN(n13728) );
  INV_X1 U12731 ( .A(n10252), .ZN(n10253) );
  AOI22_X1 U12732 ( .A1(n13728), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6459), 
        .B2(n10253), .ZN(n10254) );
  NAND2_X1 U12733 ( .A1(n10255), .A2(n10254), .ZN(n13608) );
  XNOR2_X1 U12734 ( .A(n10623), .B(n13608), .ZN(n13780) );
  XOR2_X1 U12735 ( .A(n10622), .B(n13780), .Z(n10558) );
  INV_X1 U12736 ( .A(n13777), .ZN(n10578) );
  INV_X1 U12737 ( .A(n6453), .ZN(n14753) );
  XNOR2_X1 U12738 ( .A(n14646), .B(n14768), .ZN(n13779) );
  INV_X1 U12739 ( .A(n13779), .ZN(n10480) );
  XNOR2_X1 U12740 ( .A(n10589), .B(n13780), .ZN(n10549) );
  NAND2_X1 U12741 ( .A1(n10549), .A2(n14803), .ZN(n10269) );
  INV_X1 U12742 ( .A(n14799), .ZN(n14786) );
  NAND2_X1 U12743 ( .A1(n14646), .A2(n13551), .ZN(n10267) );
  NAND2_X1 U12744 ( .A1(n6456), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U12745 ( .A1(n13730), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10264) );
  NAND2_X1 U12746 ( .A1(n10260), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10534) );
  OR2_X1 U12747 ( .A1(n10260), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10261) );
  AND2_X1 U12748 ( .A1(n10534), .A2(n10261), .ZN(n10531) );
  NAND2_X1 U12749 ( .A1(n12027), .A2(n10531), .ZN(n10263) );
  NAND2_X1 U12750 ( .A1(n12050), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10262) );
  NAND4_X1 U12751 ( .A1(n10265), .A2(n10264), .A3(n10263), .A4(n10262), .ZN(
        n13843) );
  NAND2_X1 U12752 ( .A1(n13843), .A2(n14645), .ZN(n10266) );
  NAND2_X1 U12753 ( .A1(n10267), .A2(n10266), .ZN(n10550) );
  NAND2_X1 U12754 ( .A1(n6664), .A2(n14731), .ZN(n14729) );
  NOR2_X1 U12755 ( .A1(n14729), .A2(n6453), .ZN(n14715) );
  INV_X1 U12756 ( .A(n14656), .ZN(n14760) );
  NAND2_X1 U12757 ( .A1(n14715), .A2(n14760), .ZN(n14714) );
  OR2_X1 U12758 ( .A1(n14714), .A2(n13601), .ZN(n10482) );
  AOI211_X1 U12759 ( .C1(n13608), .C2(n10482), .A(n14789), .B(n6849), .ZN(
        n10555) );
  AOI211_X1 U12760 ( .C1(n14786), .C2(n13608), .A(n10550), .B(n10555), .ZN(
        n10268) );
  OAI211_X1 U12761 ( .C1(n14795), .C2(n10558), .A(n10269), .B(n10268), .ZN(
        n10272) );
  NAND2_X1 U12762 ( .A1(n10272), .A2(n14819), .ZN(n10270) );
  OAI21_X1 U12763 ( .B1(n14819), .B2(n10271), .A(n10270), .ZN(P1_U3533) );
  INV_X1 U12764 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U12765 ( .A1(n10272), .A2(n14807), .ZN(n10273) );
  OAI21_X1 U12766 ( .B1(n14807), .B2(n10274), .A(n10273), .ZN(P1_U3474) );
  NAND2_X1 U12767 ( .A1(n10286), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10279) );
  AOI21_X1 U12768 ( .B1(n9958), .B2(n10276), .A(n10275), .ZN(n14908) );
  INV_X1 U12769 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11480) );
  NAND2_X1 U12770 ( .A1(n14911), .A2(n11480), .ZN(n10277) );
  OAI21_X1 U12771 ( .B1(n14911), .B2(n11480), .A(n10277), .ZN(n10278) );
  INV_X1 U12772 ( .A(n10278), .ZN(n14907) );
  NAND2_X1 U12773 ( .A1(n14908), .A2(n14907), .ZN(n14906) );
  NAND2_X1 U12774 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10280), .ZN(n13094) );
  OAI211_X1 U12775 ( .C1(n10280), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14931), 
        .B(n13094), .ZN(n10293) );
  OR2_X1 U12776 ( .A1(n10281), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14493) );
  OAI21_X1 U12777 ( .B1(n14937), .B2(n6659), .A(n14493), .ZN(n10291) );
  NAND2_X1 U12778 ( .A1(n10283), .A2(n10282), .ZN(n14899) );
  NAND2_X1 U12779 ( .A1(n14911), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10284) );
  OAI21_X1 U12780 ( .B1(n14911), .B2(P2_REG1_REG_13__SCAN_IN), .A(n10284), 
        .ZN(n10285) );
  INV_X1 U12781 ( .A(n10285), .ZN(n14898) );
  NOR2_X1 U12782 ( .A1(n14899), .A2(n14898), .ZN(n14903) );
  AOI21_X1 U12783 ( .B1(n10286), .B2(P2_REG1_REG_13__SCAN_IN), .A(n14903), 
        .ZN(n10289) );
  INV_X1 U12784 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14526) );
  NOR2_X1 U12785 ( .A1(n13093), .A2(n14526), .ZN(n10287) );
  AOI21_X1 U12786 ( .B1(n13093), .B2(n14526), .A(n10287), .ZN(n10288) );
  NOR2_X1 U12787 ( .A1(n10289), .A2(n10288), .ZN(n13081) );
  AOI211_X1 U12788 ( .C1(n10289), .C2(n10288), .A(n13081), .B(n14923), .ZN(
        n10290) );
  AOI211_X1 U12789 ( .C1(n14929), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n10291), 
        .B(n10290), .ZN(n10292) );
  NAND2_X1 U12790 ( .A1(n10293), .A2(n10292), .ZN(P2_U3228) );
  MUX2_X1 U12791 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n6622), .Z(n10890) );
  XNOR2_X1 U12792 ( .A(n10890), .B(n10906), .ZN(n10892) );
  OAI22_X1 U12793 ( .A1(n10296), .A2(n10295), .B1(n10294), .B2(n10298), .ZN(
        n10893) );
  XOR2_X1 U12794 ( .A(n10893), .B(n10892), .Z(n10316) );
  NAND2_X1 U12795 ( .A1(n10298), .A2(n10297), .ZN(n10300) );
  INV_X1 U12796 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10301) );
  MUX2_X1 U12797 ( .A(n10301), .B(P3_REG1_REG_8__SCAN_IN), .S(n10906), .Z(
        n10302) );
  NAND2_X1 U12798 ( .A1(n10303), .A2(n10302), .ZN(n10905) );
  OAI21_X1 U12799 ( .B1(n10303), .B2(n10302), .A(n10905), .ZN(n10314) );
  AND2_X1 U12800 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n10962) );
  NOR2_X1 U12801 ( .A1(n10305), .A2(n10304), .ZN(n10307) );
  MUX2_X1 U12802 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n11045), .S(n10906), .Z(
        n10308) );
  AOI21_X1 U12803 ( .B1(n10309), .B2(n10308), .A(n10885), .ZN(n10310) );
  NOR2_X1 U12804 ( .A1(n15091), .A2(n10310), .ZN(n10311) );
  AOI211_X1 U12805 ( .C1(n15075), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n10962), .B(
        n10311), .ZN(n10312) );
  OAI21_X1 U12806 ( .B1(n10886), .B2(n15070), .A(n10312), .ZN(n10313) );
  AOI21_X1 U12807 ( .B1(n15086), .B2(n10314), .A(n10313), .ZN(n10315) );
  OAI21_X1 U12808 ( .B1(n10316), .B2(n15096), .A(n10315), .ZN(P3_U3190) );
  INV_X1 U12809 ( .A(n10317), .ZN(n10320) );
  NAND2_X1 U12810 ( .A1(n8973), .A2(n12834), .ZN(n10323) );
  XNOR2_X1 U12811 ( .A(n10321), .B(n12873), .ZN(n10322) );
  NAND2_X1 U12812 ( .A1(n10323), .A2(n10322), .ZN(n10736) );
  OAI21_X1 U12813 ( .B1(n10323), .B2(n10322), .A(n10736), .ZN(n10324) );
  AOI21_X1 U12814 ( .B1(n10325), .B2(n10324), .A(n10738), .ZN(n10330) );
  OAI22_X1 U12815 ( .A1(n10326), .A2(n14491), .B1(n10450), .B2(n14488), .ZN(
        n10327) );
  AOI21_X1 U12816 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n10328), .A(n10327), .ZN(
        n10329) );
  OAI21_X1 U12817 ( .B1(n10330), .B2(n14490), .A(n10329), .ZN(P2_U3209) );
  INV_X1 U12818 ( .A(n10331), .ZN(n10334) );
  OAI21_X1 U12819 ( .B1(n10334), .B2(n10333), .A(n10332), .ZN(n14653) );
  AOI22_X1 U12820 ( .A1(n13845), .A2(n11966), .B1(n12222), .B2(n6457), .ZN(
        n10335) );
  XOR2_X1 U12821 ( .A(n10393), .B(n10335), .Z(n10338) );
  OAI22_X1 U12822 ( .A1(n10336), .A2(n11803), .B1(n14760), .B2(n11904), .ZN(
        n10337) );
  NAND2_X1 U12823 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  OAI21_X1 U12824 ( .B1(n10338), .B2(n10337), .A(n10339), .ZN(n14652) );
  INV_X1 U12825 ( .A(n10339), .ZN(n10340) );
  AOI22_X1 U12826 ( .A1(n12223), .A2(n14646), .B1(n11966), .B2(n13601), .ZN(
        n10341) );
  NAND2_X1 U12827 ( .A1(n7346), .A2(n10389), .ZN(n10343) );
  AOI22_X1 U12828 ( .A1(n14646), .A2(n11966), .B1(n13601), .B2(n12222), .ZN(
        n10342) );
  XOR2_X1 U12829 ( .A(n10393), .B(n10342), .Z(n10390) );
  XNOR2_X1 U12830 ( .A(n10343), .B(n10390), .ZN(n10351) );
  NAND2_X1 U12831 ( .A1(n10344), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14659) );
  INV_X1 U12832 ( .A(n10345), .ZN(n10487) );
  NAND2_X1 U12833 ( .A1(n13845), .A2(n13551), .ZN(n10347) );
  NAND2_X1 U12834 ( .A1(n13844), .A2(n14645), .ZN(n10346) );
  NAND2_X1 U12835 ( .A1(n10347), .A2(n10346), .ZN(n10484) );
  AND2_X1 U12836 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14672) );
  AOI21_X1 U12837 ( .B1(n14578), .B2(n10484), .A(n14672), .ZN(n10349) );
  NAND2_X1 U12838 ( .A1(n14657), .A2(n13601), .ZN(n10348) );
  OAI211_X1 U12839 ( .C1(n14659), .C2(n10487), .A(n10349), .B(n10348), .ZN(
        n10350) );
  AOI21_X1 U12840 ( .B1(n10351), .B2(n14576), .A(n10350), .ZN(n10352) );
  INV_X1 U12841 ( .A(n10352), .ZN(P1_U3230) );
  NOR2_X2 U12842 ( .A1(n10354), .A2(n10353), .ZN(n14728) );
  NOR2_X1 U12843 ( .A1(n10356), .A2(n10355), .ZN(n10357) );
  NAND2_X1 U12844 ( .A1(n10358), .A2(n10357), .ZN(n12057) );
  INV_X2 U12845 ( .A(n14120), .ZN(n14739) );
  INV_X1 U12846 ( .A(n14120), .ZN(n14697) );
  INV_X1 U12847 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10359) );
  OAI22_X1 U12848 ( .A1(n14697), .A2(n10360), .B1(n10359), .B2(n14116), .ZN(
        n10363) );
  OR2_X1 U12849 ( .A1(n9564), .A2(n13738), .ZN(n13765) );
  INV_X1 U12850 ( .A(n13765), .ZN(n13808) );
  NAND2_X1 U12851 ( .A1(n13808), .A2(n13569), .ZN(n10361) );
  NOR2_X1 U12852 ( .A1(n12057), .A2(n11394), .ZN(n12062) );
  INV_X1 U12853 ( .A(n12062), .ZN(n11124) );
  AOI21_X1 U12854 ( .B1(n14712), .B2(n11124), .A(n14731), .ZN(n10362) );
  AOI211_X1 U12855 ( .C1(n14739), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10363), .B(
        n10362), .ZN(n10367) );
  INV_X1 U12856 ( .A(n10364), .ZN(n10365) );
  INV_X1 U12857 ( .A(n14126), .ZN(n14093) );
  OAI21_X1 U12858 ( .B1(n14124), .B2(n14093), .A(n13776), .ZN(n10366) );
  NAND2_X1 U12859 ( .A1(n10367), .A2(n10366), .ZN(P1_U3293) );
  INV_X1 U12860 ( .A(n10368), .ZN(n10370) );
  INV_X1 U12861 ( .A(SI_20_), .ZN(n10369) );
  OAI222_X1 U12862 ( .A1(n10371), .A2(P3_U3151), .B1(n12832), .B2(n10370), 
        .C1(n10369), .C2(n12829), .ZN(P3_U3275) );
  MUX2_X1 U12863 ( .A(n10372), .B(n9792), .S(n14951), .Z(n10378) );
  OAI22_X1 U12864 ( .A1(n13205), .A2(n10374), .B1(n10373), .B2(n13295), .ZN(
        n10375) );
  AOI21_X1 U12865 ( .B1(n10376), .B2(n14509), .A(n10375), .ZN(n10377) );
  OAI211_X1 U12866 ( .C1(n10379), .C2(n13224), .A(n10378), .B(n10377), .ZN(
        P2_U3264) );
  AOI211_X1 U12867 ( .C1(n10382), .C2(n10381), .A(n12347), .B(n10380), .ZN(
        n10383) );
  INV_X1 U12868 ( .A(n10383), .ZN(n10388) );
  NOR2_X1 U12869 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10384), .ZN(n15006) );
  INV_X1 U12870 ( .A(n12352), .ZN(n12314) );
  OAI22_X1 U12871 ( .A1(n12360), .A2(n10385), .B1(n12314), .B2(n12760), .ZN(
        n10386) );
  AOI211_X1 U12872 ( .C1(n12311), .C2(n12381), .A(n15006), .B(n10386), .ZN(
        n10387) );
  OAI211_X1 U12873 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11345), .A(n10388), .B(
        n10387), .ZN(P3_U3158) );
  AOI22_X1 U12874 ( .A1(n12223), .A2(n13844), .B1(n13608), .B2(n11966), .ZN(
        n10518) );
  NAND2_X1 U12875 ( .A1(n13608), .A2(n12222), .ZN(n10392) );
  NAND2_X1 U12876 ( .A1(n13844), .A2(n11834), .ZN(n10391) );
  NAND2_X1 U12877 ( .A1(n10392), .A2(n10391), .ZN(n10394) );
  XNOR2_X1 U12878 ( .A(n10394), .B(n11810), .ZN(n10519) );
  XOR2_X1 U12879 ( .A(n10518), .B(n10519), .Z(n10395) );
  XNOR2_X1 U12880 ( .A(n10520), .B(n10395), .ZN(n10401) );
  INV_X1 U12881 ( .A(n10552), .ZN(n10399) );
  AOI21_X1 U12882 ( .B1(n14578), .B2(n10550), .A(n10396), .ZN(n10398) );
  NAND2_X1 U12883 ( .A1(n14657), .A2(n13608), .ZN(n10397) );
  OAI211_X1 U12884 ( .C1(n14659), .C2(n10399), .A(n10398), .B(n10397), .ZN(
        n10400) );
  AOI21_X1 U12885 ( .B1(n10401), .B2(n14576), .A(n10400), .ZN(n10402) );
  INV_X1 U12886 ( .A(n10402), .ZN(P1_U3227) );
  OAI21_X1 U12887 ( .B1(n10404), .B2(n10409), .A(n10403), .ZN(n14946) );
  INV_X1 U12888 ( .A(n10405), .ZN(n10406) );
  AOI211_X1 U12889 ( .C1(n14939), .C2(n10406), .A(n13217), .B(n6882), .ZN(
        n14938) );
  NAND2_X1 U12890 ( .A1(n10408), .A2(n10407), .ZN(n10410) );
  XNOR2_X1 U12891 ( .A(n10410), .B(n10409), .ZN(n10413) );
  NAND2_X1 U12892 ( .A1(n8973), .A2(n14484), .ZN(n10412) );
  NAND2_X1 U12893 ( .A1(n13046), .A2(n14481), .ZN(n10411) );
  AND2_X1 U12894 ( .A1(n10412), .A2(n10411), .ZN(n10792) );
  OAI21_X1 U12895 ( .B1(n10413), .B2(n13371), .A(n10792), .ZN(n14945) );
  AOI211_X1 U12896 ( .C1(n14983), .C2(n14946), .A(n14938), .B(n14945), .ZN(
        n10420) );
  OAI22_X1 U12897 ( .A1(n13378), .A2(n10417), .B1(n15002), .B2(n12183), .ZN(
        n10414) );
  INV_X1 U12898 ( .A(n10414), .ZN(n10415) );
  OAI21_X1 U12899 ( .B1(n10420), .B2(n14999), .A(n10415), .ZN(P2_U3502) );
  INV_X1 U12900 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10416) );
  OAI22_X1 U12901 ( .A1(n13431), .A2(n10417), .B1(n10105), .B2(n10416), .ZN(
        n10418) );
  INV_X1 U12902 ( .A(n10418), .ZN(n10419) );
  OAI21_X1 U12903 ( .B1(n10420), .B2(n14991), .A(n10419), .ZN(P2_U3439) );
  OAI21_X1 U12904 ( .B1(n10422), .B2(n10424), .A(n10421), .ZN(n10423) );
  INV_X1 U12905 ( .A(n10423), .ZN(n10478) );
  INV_X1 U12906 ( .A(n14475), .ZN(n10430) );
  NAND2_X1 U12907 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  NAND2_X1 U12908 ( .A1(n10427), .A2(n10426), .ZN(n10429) );
  OAI22_X1 U12909 ( .A1(n10638), .A2(n12683), .B1(n10862), .B2(n12759), .ZN(
        n10428) );
  AOI21_X1 U12910 ( .B1(n10429), .B2(n12762), .A(n10428), .ZN(n10473) );
  OAI21_X1 U12911 ( .B1(n10478), .B2(n10430), .A(n10473), .ZN(n10446) );
  OAI22_X1 U12912 ( .A1(n12755), .A2(n10639), .B1(n15133), .B2(n15057), .ZN(
        n10431) );
  AOI21_X1 U12913 ( .B1(n10446), .B2(n15133), .A(n10431), .ZN(n10432) );
  INV_X1 U12914 ( .A(n10432), .ZN(P3_U3464) );
  INV_X1 U12915 ( .A(n11695), .ZN(n10458) );
  INV_X1 U12916 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U12917 ( .A1(n10434), .A2(n10433), .ZN(n10493) );
  NAND2_X1 U12918 ( .A1(n10493), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10435) );
  XNOR2_X1 U12919 ( .A(n10435), .B(P1_IR_REG_16__SCAN_IN), .ZN(n13912) );
  INV_X1 U12920 ( .A(n13912), .ZN(n13922) );
  OAI222_X1 U12921 ( .A1(n6454), .A2(n10436), .B1(n14286), .B2(n10458), .C1(
        n13922), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12922 ( .A(n10437), .ZN(n10438) );
  NAND2_X1 U12923 ( .A1(n13298), .A2(n10438), .ZN(n11167) );
  OAI21_X1 U12924 ( .B1(n7968), .B2(n10440), .A(n10439), .ZN(n10441) );
  NAND2_X1 U12925 ( .A1(n10441), .A2(n13298), .ZN(n10443) );
  AOI22_X1 U12926 ( .A1(n14951), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n14941), .ZN(n10442) );
  OAI211_X1 U12927 ( .C1(n11167), .C2(n10444), .A(n10443), .B(n10442), .ZN(
        P2_U3265) );
  OAI22_X1 U12928 ( .A1(n10639), .A2(n12818), .B1(n15129), .B2(n8202), .ZN(
        n10445) );
  AOI21_X1 U12929 ( .B1(n10446), .B2(n15129), .A(n10445), .ZN(n10447) );
  INV_X1 U12930 ( .A(n10447), .ZN(P3_U3405) );
  INV_X1 U12931 ( .A(n10448), .ZN(n10457) );
  NAND2_X1 U12932 ( .A1(n10449), .A2(n14948), .ZN(n10456) );
  NOR2_X1 U12933 ( .A1(n13205), .A2(n10450), .ZN(n10453) );
  INV_X1 U12934 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10451) );
  OAI22_X1 U12935 ( .A1(n14948), .A2(n9791), .B1(n10451), .B2(n13295), .ZN(
        n10452) );
  AOI211_X1 U12936 ( .C1(n10454), .C2(n14509), .A(n10453), .B(n10452), .ZN(
        n10455) );
  OAI211_X1 U12937 ( .C1(n13224), .C2(n10457), .A(n10456), .B(n10455), .ZN(
        P2_U3263) );
  OAI222_X1 U12938 ( .A1(n13458), .A2(n10459), .B1(n14936), .B2(P2_U3088), 
        .C1(n13461), .C2(n10458), .ZN(P2_U3311) );
  INV_X1 U12939 ( .A(n10460), .ZN(n10471) );
  OAI21_X1 U12940 ( .B1(n10463), .B2(n10462), .A(n10461), .ZN(n10464) );
  NAND2_X1 U12941 ( .A1(n10464), .A2(n12341), .ZN(n10470) );
  NOR2_X1 U12942 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10465), .ZN(n15030) );
  OAI22_X1 U12943 ( .A1(n12360), .A2(n10467), .B1(n12314), .B2(n10466), .ZN(
        n10468) );
  AOI211_X1 U12944 ( .C1(n12311), .C2(n12380), .A(n15030), .B(n10468), .ZN(
        n10469) );
  OAI211_X1 U12945 ( .C1(n10471), .C2(n11345), .A(n10470), .B(n10469), .ZN(
        P3_U3170) );
  INV_X1 U12946 ( .A(n11816), .ZN(n10495) );
  INV_X1 U12947 ( .A(n13110), .ZN(n13106) );
  OAI222_X1 U12948 ( .A1(n13467), .A2(n10495), .B1(n13106), .B2(P2_U3088), 
        .C1(n10472), .C2(n13458), .ZN(P2_U3310) );
  INV_X1 U12949 ( .A(n12691), .ZN(n11080) );
  MUX2_X1 U12950 ( .A(n10474), .B(n10473), .S(n15117), .Z(n10477) );
  AOI22_X1 U12951 ( .A1(n14463), .A2(n10475), .B1(n12687), .B2(n10641), .ZN(
        n10476) );
  OAI211_X1 U12952 ( .C1(n11080), .C2(n10478), .A(n10477), .B(n10476), .ZN(
        P3_U3228) );
  XNOR2_X1 U12953 ( .A(n10480), .B(n10479), .ZN(n14774) );
  INV_X1 U12954 ( .A(n14774), .ZN(n10492) );
  AND2_X1 U12955 ( .A1(n10481), .A2(n10480), .ZN(n14770) );
  OR3_X1 U12956 ( .A1(n14771), .A2(n14770), .A3(n14160), .ZN(n10491) );
  AOI21_X1 U12957 ( .B1(n14714), .B2(n13601), .A(n14789), .ZN(n10483) );
  NAND2_X1 U12958 ( .A1(n10483), .A2(n10482), .ZN(n14767) );
  OR2_X1 U12959 ( .A1(n12057), .A2(n13568), .ZN(n14732) );
  NOR2_X1 U12960 ( .A1(n14767), .A2(n14732), .ZN(n10489) );
  INV_X1 U12961 ( .A(n10484), .ZN(n14766) );
  MUX2_X1 U12962 ( .A(n14766), .B(n10485), .S(n14739), .Z(n10486) );
  OAI21_X1 U12963 ( .B1(n14116), .B2(n10487), .A(n10486), .ZN(n10488) );
  AOI211_X1 U12964 ( .C1(n14735), .C2(n13601), .A(n10489), .B(n10488), .ZN(
        n10490) );
  OAI211_X1 U12965 ( .C1(n10492), .C2(n14126), .A(n10491), .B(n10490), .ZN(
        P1_U3289) );
  OAI21_X1 U12966 ( .B1(n10493), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10494) );
  XNOR2_X1 U12967 ( .A(n10494), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13936) );
  INV_X1 U12968 ( .A(n13936), .ZN(n13932) );
  OAI222_X1 U12969 ( .A1(n6454), .A2(n10496), .B1(n14286), .B2(n10495), .C1(
        n13932), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U12970 ( .A(SI_21_), .ZN(n10499) );
  INV_X1 U12971 ( .A(n10497), .ZN(n10498) );
  OAI222_X1 U12972 ( .A1(P3_U3151), .A2(n10500), .B1(n12829), .B2(n10499), 
        .C1(n12832), .C2(n10498), .ZN(P3_U3274) );
  NAND2_X1 U12973 ( .A1(n10501), .A2(n10502), .ZN(n10504) );
  NAND2_X1 U12974 ( .A1(n10504), .A2(n10503), .ZN(n10505) );
  XNOR2_X1 U12975 ( .A(n10505), .B(n10507), .ZN(n10729) );
  NAND2_X1 U12976 ( .A1(n13298), .A2(n14535), .ZN(n13305) );
  OAI21_X1 U12977 ( .B1(n10508), .B2(n10507), .A(n10506), .ZN(n10727) );
  AOI21_X1 U12978 ( .B1(n10665), .B2(n10831), .A(n13217), .ZN(n10509) );
  AND2_X1 U12979 ( .A1(n10656), .A2(n10509), .ZN(n10726) );
  NAND2_X1 U12980 ( .A1(n10726), .A2(n14509), .ZN(n10515) );
  NAND2_X1 U12981 ( .A1(n13046), .A2(n14484), .ZN(n10511) );
  NAND2_X1 U12982 ( .A1(n13044), .A2(n13013), .ZN(n10510) );
  NAND2_X1 U12983 ( .A1(n10511), .A2(n10510), .ZN(n10840) );
  MUX2_X1 U12984 ( .A(n10840), .B(P2_REG2_REG_5__SCAN_IN), .S(n14951), .Z(
        n10513) );
  OAI22_X1 U12985 ( .A1(n13205), .A2(n10839), .B1(n10842), .B2(n13295), .ZN(
        n10512) );
  NOR2_X1 U12986 ( .A1(n10513), .A2(n10512), .ZN(n10514) );
  NAND2_X1 U12987 ( .A1(n10515), .A2(n10514), .ZN(n10516) );
  AOI21_X1 U12988 ( .B1(n10727), .B2(n14510), .A(n10516), .ZN(n10517) );
  OAI21_X1 U12989 ( .B1(n10729), .B2(n13305), .A(n10517), .ZN(P2_U3260) );
  OR2_X1 U12990 ( .A1(n10521), .A2(n6451), .ZN(n10524) );
  AOI22_X1 U12991 ( .A1(n13728), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6459), 
        .B2(n10522), .ZN(n10523) );
  NAND2_X1 U12992 ( .A1(n10524), .A2(n10523), .ZN(n13616) );
  NAND2_X1 U12993 ( .A1(n13616), .A2(n12222), .ZN(n10526) );
  NAND2_X1 U12994 ( .A1(n13843), .A2(n11834), .ZN(n10525) );
  NAND2_X1 U12995 ( .A1(n10526), .A2(n10525), .ZN(n10527) );
  XNOR2_X1 U12996 ( .A(n10527), .B(n11810), .ZN(n10529) );
  AOI22_X1 U12997 ( .A1(n13616), .A2(n11966), .B1(n12223), .B2(n13843), .ZN(
        n10528) );
  NAND2_X1 U12998 ( .A1(n10529), .A2(n10528), .ZN(n10873) );
  NAND2_X1 U12999 ( .A1(n6592), .A2(n10873), .ZN(n10530) );
  XNOR2_X1 U13000 ( .A(n10874), .B(n10530), .ZN(n10545) );
  INV_X1 U13001 ( .A(n10531), .ZN(n10721) );
  NAND2_X1 U13002 ( .A1(n13844), .A2(n13551), .ZN(n10541) );
  NAND2_X1 U13003 ( .A1(n6456), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10539) );
  NAND2_X1 U13004 ( .A1(n12051), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U13005 ( .A1(n10534), .A2(n10533), .ZN(n10535) );
  AND2_X1 U13006 ( .A1(n10600), .A2(n10535), .ZN(n10867) );
  NAND2_X1 U13007 ( .A1(n12027), .A2(n10867), .ZN(n10537) );
  NAND2_X1 U13008 ( .A1(n12050), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10536) );
  NAND4_X1 U13009 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n13842) );
  NAND2_X1 U13010 ( .A1(n13842), .A2(n14645), .ZN(n10540) );
  NAND2_X1 U13011 ( .A1(n10541), .A2(n10540), .ZN(n10716) );
  AOI22_X1 U13012 ( .A1(n14578), .A2(n10716), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10543) );
  NAND2_X1 U13013 ( .A1(n14657), .A2(n13616), .ZN(n10542) );
  OAI211_X1 U13014 ( .C1(n14659), .C2(n10721), .A(n10543), .B(n10542), .ZN(
        n10544) );
  AOI21_X1 U13015 ( .B1(n10545), .B2(n14576), .A(n10544), .ZN(n10546) );
  INV_X1 U13016 ( .A(n10546), .ZN(P1_U3239) );
  NAND2_X1 U13017 ( .A1(n10547), .A2(n13568), .ZN(n13763) );
  INV_X1 U13018 ( .A(n13763), .ZN(n14727) );
  NAND2_X1 U13019 ( .A1(n14120), .A2(n14727), .ZN(n14139) );
  OAI21_X1 U13020 ( .B1(n14739), .B2(n14130), .A(n14139), .ZN(n10548) );
  NAND2_X1 U13021 ( .A1(n10549), .A2(n10548), .ZN(n10557) );
  INV_X1 U13022 ( .A(n14732), .ZN(n14717) );
  INV_X1 U13023 ( .A(n13608), .ZN(n10588) );
  MUX2_X1 U13024 ( .A(n10550), .B(P1_REG2_REG_5__SCAN_IN), .S(n14739), .Z(
        n10551) );
  AOI21_X1 U13025 ( .B1(n14728), .B2(n10552), .A(n10551), .ZN(n10553) );
  OAI21_X1 U13026 ( .B1(n10588), .B2(n14712), .A(n10553), .ZN(n10554) );
  AOI21_X1 U13027 ( .B1(n10555), .B2(n14717), .A(n10554), .ZN(n10556) );
  OAI211_X1 U13028 ( .C1(n10558), .C2(n14126), .A(n10557), .B(n10556), .ZN(
        P1_U3288) );
  INV_X1 U13029 ( .A(n10559), .ZN(n10562) );
  OAI22_X1 U13030 ( .A1(n10560), .A2(P3_U3151), .B1(SI_22_), .B2(n12829), .ZN(
        n10561) );
  AOI21_X1 U13031 ( .B1(n10562), .B2(n14422), .A(n10561), .ZN(P3_U3273) );
  OAI21_X1 U13032 ( .B1(n10564), .B2(n10565), .A(n10563), .ZN(n10678) );
  INV_X1 U13033 ( .A(n10678), .ZN(n10573) );
  AOI21_X1 U13034 ( .B1(n10566), .B2(n10565), .A(n12680), .ZN(n10569) );
  OAI22_X1 U13035 ( .A1(n10776), .A2(n12683), .B1(n10960), .B2(n12759), .ZN(
        n10567) );
  AOI21_X1 U13036 ( .B1(n10569), .B2(n10568), .A(n10567), .ZN(n10676) );
  MUX2_X1 U13037 ( .A(n10676), .B(n10570), .S(n15119), .Z(n10572) );
  AOI22_X1 U13038 ( .A1(n14463), .A2(n10681), .B1(n12687), .B2(n10772), .ZN(
        n10571) );
  OAI211_X1 U13039 ( .C1(n11080), .C2(n10573), .A(n10572), .B(n10571), .ZN(
        P3_U3227) );
  XNOR2_X1 U13040 ( .A(n13777), .B(n10574), .ZN(n10576) );
  AOI21_X1 U13041 ( .B1(n10576), .B2(n14784), .A(n10575), .ZN(n10580) );
  XNOR2_X1 U13042 ( .A(n10578), .B(n10577), .ZN(n14755) );
  INV_X1 U13043 ( .A(n14130), .ZN(n14723) );
  NAND2_X1 U13044 ( .A1(n14755), .A2(n14723), .ZN(n10579) );
  AND2_X1 U13045 ( .A1(n10580), .A2(n10579), .ZN(n14757) );
  INV_X1 U13046 ( .A(n14139), .ZN(n14718) );
  NAND2_X1 U13047 ( .A1(n14729), .A2(n6453), .ZN(n10581) );
  INV_X1 U13048 ( .A(n14789), .ZN(n14730) );
  NAND2_X1 U13049 ( .A1(n10581), .A2(n14730), .ZN(n10582) );
  OR2_X1 U13050 ( .A1(n14715), .A2(n10582), .ZN(n14752) );
  OAI22_X1 U13051 ( .A1(n14120), .A2(n9448), .B1(n10583), .B2(n14116), .ZN(
        n10584) );
  AOI21_X1 U13052 ( .B1(n14735), .B2(n6453), .A(n10584), .ZN(n10585) );
  OAI21_X1 U13053 ( .B1(n14732), .B2(n14752), .A(n10585), .ZN(n10586) );
  AOI21_X1 U13054 ( .B1(n14718), .B2(n14755), .A(n10586), .ZN(n10587) );
  OAI21_X1 U13055 ( .B1(n14739), .B2(n14757), .A(n10587), .ZN(P1_U3291) );
  INV_X1 U13056 ( .A(n13616), .ZN(n10722) );
  INV_X1 U13057 ( .A(n13843), .ZN(n10626) );
  NAND2_X1 U13058 ( .A1(n10722), .A2(n10626), .ZN(n10590) );
  NAND2_X1 U13059 ( .A1(n10591), .A2(n13756), .ZN(n10593) );
  AOI22_X1 U13060 ( .A1(n13728), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6459), 
        .B2(n13897), .ZN(n10592) );
  XNOR2_X1 U13061 ( .A(n13620), .B(n13842), .ZN(n13783) );
  NAND2_X1 U13062 ( .A1(n10595), .A2(n13756), .ZN(n10598) );
  AOI22_X1 U13063 ( .A1(n13728), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6459), 
        .B2(n10596), .ZN(n10597) );
  NAND2_X1 U13064 ( .A1(n6456), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U13065 ( .A1(n13730), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10605) );
  NAND2_X1 U13066 ( .A1(n10600), .A2(n10599), .ZN(n10601) );
  NAND2_X1 U13067 ( .A1(n10609), .A2(n10601), .ZN(n10941) );
  INV_X1 U13068 ( .A(n10941), .ZN(n10602) );
  NAND2_X1 U13069 ( .A1(n12027), .A2(n10602), .ZN(n10604) );
  NAND2_X1 U13070 ( .A1(n12050), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10603) );
  NAND4_X1 U13071 ( .A1(n10606), .A2(n10605), .A3(n10604), .A4(n10603), .ZN(
        n13841) );
  XNOR2_X1 U13072 ( .A(n14787), .B(n13841), .ZN(n13785) );
  OAI21_X1 U13073 ( .B1(n10607), .B2(n10630), .A(n10995), .ZN(n14793) );
  INV_X1 U13074 ( .A(n14793), .ZN(n10634) );
  INV_X1 U13075 ( .A(n13620), .ZN(n14776) );
  NAND2_X1 U13076 ( .A1(n10766), .A2(n14787), .ZN(n10608) );
  NAND2_X1 U13077 ( .A1(n11061), .A2(n10608), .ZN(n14790) );
  AND2_X1 U13078 ( .A1(n10609), .A2(n11294), .ZN(n10610) );
  NOR2_X1 U13079 ( .A1(n11005), .A2(n10610), .ZN(n14696) );
  NAND2_X1 U13080 ( .A1(n12027), .A2(n14696), .ZN(n10616) );
  NAND2_X1 U13081 ( .A1(n12050), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10615) );
  INV_X1 U13082 ( .A(n10235), .ZN(n10611) );
  OR2_X1 U13083 ( .A1(n10611), .A2(n9623), .ZN(n10614) );
  INV_X1 U13084 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10612) );
  OR2_X1 U13085 ( .A1(n10532), .A2(n10612), .ZN(n10613) );
  NAND2_X1 U13086 ( .A1(n13842), .A2(n13551), .ZN(n10617) );
  OAI21_X1 U13087 ( .B1(n11290), .B2(n13544), .A(n10617), .ZN(n14785) );
  INV_X1 U13088 ( .A(n14785), .ZN(n10618) );
  OAI21_X1 U13089 ( .B1(n14790), .B2(n11394), .A(n10618), .ZN(n10621) );
  NOR2_X1 U13090 ( .A1(n6847), .A2(n14712), .ZN(n10620) );
  OAI22_X1 U13091 ( .A1(n14120), .A2(n9621), .B1(n10941), .B2(n14116), .ZN(
        n10619) );
  AOI211_X1 U13092 ( .C1(n10621), .C2(n14120), .A(n10620), .B(n10619), .ZN(
        n10633) );
  NAND2_X1 U13093 ( .A1(n10623), .A2(n13608), .ZN(n10624) );
  INV_X1 U13094 ( .A(n13842), .ZN(n10628) );
  OR2_X1 U13095 ( .A1(n13620), .A2(n10628), .ZN(n10627) );
  INV_X1 U13096 ( .A(n10631), .ZN(n10629) );
  NAND2_X1 U13097 ( .A1(n10629), .A2(n13785), .ZN(n11015) );
  NAND2_X1 U13098 ( .A1(n10631), .A2(n10630), .ZN(n14783) );
  NAND3_X1 U13099 ( .A1(n11015), .A2(n14783), .A3(n14093), .ZN(n10632) );
  OAI211_X1 U13100 ( .C1(n10634), .C2(n14160), .A(n10633), .B(n10632), .ZN(
        P1_U3285) );
  XOR2_X1 U13101 ( .A(n10636), .B(n10635), .Z(n10644) );
  NOR2_X1 U13102 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10637), .ZN(n15051) );
  OAI22_X1 U13103 ( .A1(n12360), .A2(n10639), .B1(n12314), .B2(n10638), .ZN(
        n10640) );
  AOI211_X1 U13104 ( .C1(n12311), .C2(n12379), .A(n15051), .B(n10640), .ZN(
        n10643) );
  NAND2_X1 U13105 ( .A1(n12356), .A2(n10641), .ZN(n10642) );
  OAI211_X1 U13106 ( .C1(n10644), .C2(n12347), .A(n10643), .B(n10642), .ZN(
        P3_U3167) );
  NAND2_X1 U13107 ( .A1(n10501), .A2(n10645), .ZN(n10647) );
  NAND2_X1 U13108 ( .A1(n10647), .A2(n10646), .ZN(n10649) );
  OAI21_X1 U13109 ( .B1(n10649), .B2(n10648), .A(n6467), .ZN(n10652) );
  NAND2_X1 U13110 ( .A1(n13045), .A2(n14484), .ZN(n10651) );
  NAND2_X1 U13111 ( .A1(n13043), .A2(n14481), .ZN(n10650) );
  NAND2_X1 U13112 ( .A1(n10651), .A2(n10650), .ZN(n10851) );
  AOI21_X1 U13113 ( .B1(n10652), .B2(n14535), .A(n10851), .ZN(n14964) );
  OAI21_X1 U13114 ( .B1(n10655), .B2(n10654), .A(n10653), .ZN(n14967) );
  INV_X1 U13115 ( .A(n10656), .ZN(n10658) );
  INV_X1 U13116 ( .A(n10806), .ZN(n10657) );
  OAI211_X1 U13117 ( .C1(n14965), .C2(n10658), .A(n10657), .B(n6452), .ZN(
        n14963) );
  AOI22_X1 U13118 ( .A1(n14951), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n10850), 
        .B2(n14941), .ZN(n10660) );
  NAND2_X1 U13119 ( .A1(n14502), .A2(n10855), .ZN(n10659) );
  OAI211_X1 U13120 ( .C1(n14963), .C2(n13302), .A(n10660), .B(n10659), .ZN(
        n10661) );
  AOI21_X1 U13121 ( .B1(n14967), .B2(n14510), .A(n10661), .ZN(n10662) );
  OAI21_X1 U13122 ( .B1(n14964), .B2(n14951), .A(n10662), .ZN(P2_U3259) );
  OAI21_X1 U13123 ( .B1(n10664), .B2(n10668), .A(n10663), .ZN(n10705) );
  INV_X1 U13124 ( .A(n10665), .ZN(n10666) );
  AOI211_X1 U13125 ( .C1(n10743), .C2(n10667), .A(n13217), .B(n10666), .ZN(
        n10709) );
  XNOR2_X1 U13126 ( .A(n10501), .B(n10668), .ZN(n10669) );
  AOI22_X1 U13127 ( .A1(n14484), .A2(n13047), .B1(n13045), .B2(n14481), .ZN(
        n10750) );
  OAI21_X1 U13128 ( .B1(n10669), .B2(n13371), .A(n10750), .ZN(n10706) );
  AOI211_X1 U13129 ( .C1(n14983), .C2(n10705), .A(n10709), .B(n10706), .ZN(
        n10675) );
  INV_X1 U13130 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10670) );
  OAI22_X1 U13131 ( .A1(n13431), .A2(n6885), .B1(n10105), .B2(n10670), .ZN(
        n10671) );
  INV_X1 U13132 ( .A(n10671), .ZN(n10672) );
  OAI21_X1 U13133 ( .B1(n10675), .B2(n14991), .A(n10672), .ZN(P2_U3442) );
  OAI22_X1 U13134 ( .A1(n13378), .A2(n6885), .B1(n15002), .B2(n9822), .ZN(
        n10673) );
  INV_X1 U13135 ( .A(n10673), .ZN(n10674) );
  OAI21_X1 U13136 ( .B1(n10675), .B2(n14999), .A(n10674), .ZN(P2_U3503) );
  INV_X1 U13137 ( .A(n10676), .ZN(n10677) );
  AOI21_X1 U13138 ( .B1(n14475), .B2(n10678), .A(n10677), .ZN(n10683) );
  OAI22_X1 U13139 ( .A1(n10777), .A2(n12818), .B1(n15129), .B2(n8221), .ZN(
        n10679) );
  INV_X1 U13140 ( .A(n10679), .ZN(n10680) );
  OAI21_X1 U13141 ( .B1(n10683), .B2(n15127), .A(n10680), .ZN(P3_U3408) );
  AOI22_X1 U13142 ( .A1(n8743), .A2(n10681), .B1(n15131), .B2(
        P3_REG1_REG_6__SCAN_IN), .ZN(n10682) );
  OAI21_X1 U13143 ( .B1(n10683), .B2(n15131), .A(n10682), .ZN(P3_U3465) );
  NAND2_X1 U13144 ( .A1(n11524), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10685) );
  NAND2_X1 U13145 ( .A1(n10685), .A2(n10684), .ZN(n10686) );
  NOR2_X1 U13146 ( .A1(n14687), .A2(n10686), .ZN(n10687) );
  XOR2_X1 U13147 ( .A(n10686), .B(n10693), .Z(n14681) );
  NOR2_X1 U13148 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14681), .ZN(n14680) );
  NOR2_X1 U13149 ( .A1(n10687), .A2(n14680), .ZN(n10690) );
  INV_X1 U13150 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n13921) );
  NOR2_X1 U13151 ( .A1(n13922), .A2(n13921), .ZN(n10688) );
  AOI21_X1 U13152 ( .B1(n13921), .B2(n13922), .A(n10688), .ZN(n10689) );
  NAND2_X1 U13153 ( .A1(n10689), .A2(n10690), .ZN(n13920) );
  OAI211_X1 U13154 ( .C1(n10690), .C2(n10689), .A(n14690), .B(n13920), .ZN(
        n10704) );
  OAI22_X1 U13155 ( .A1(n10692), .A2(n10691), .B1(n11524), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n10694) );
  NAND2_X1 U13156 ( .A1(n10693), .A2(n10694), .ZN(n10695) );
  XNOR2_X1 U13157 ( .A(n14687), .B(n10694), .ZN(n14685) );
  INV_X1 U13158 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14684) );
  NAND2_X1 U13159 ( .A1(n14685), .A2(n14684), .ZN(n14683) );
  NAND2_X1 U13160 ( .A1(n10695), .A2(n14683), .ZN(n10698) );
  NOR2_X1 U13161 ( .A1(n13922), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n10696) );
  AOI21_X1 U13162 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n13922), .A(n10696), 
        .ZN(n10697) );
  NOR2_X1 U13163 ( .A1(n10697), .A2(n10698), .ZN(n13911) );
  AOI211_X1 U13164 ( .C1(n10698), .C2(n10697), .A(n13911), .B(n13913), .ZN(
        n10702) );
  NAND2_X1 U13165 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14579)
         );
  INV_X1 U13166 ( .A(n14579), .ZN(n10699) );
  AOI21_X1 U13167 ( .B1(n14673), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10699), 
        .ZN(n10700) );
  OAI21_X1 U13168 ( .B1(n13955), .B2(n13922), .A(n10700), .ZN(n10701) );
  NOR2_X1 U13169 ( .A1(n10702), .A2(n10701), .ZN(n10703) );
  NAND2_X1 U13170 ( .A1(n10704), .A2(n10703), .ZN(P1_U3259) );
  INV_X1 U13171 ( .A(n10705), .ZN(n10712) );
  INV_X1 U13172 ( .A(n10706), .ZN(n10707) );
  MUX2_X1 U13173 ( .A(n9793), .B(n10707), .S(n14948), .Z(n10711) );
  OAI22_X1 U13174 ( .A1(n13205), .A2(n6885), .B1(n13295), .B2(n10749), .ZN(
        n10708) );
  AOI21_X1 U13175 ( .B1(n10709), .B2(n14509), .A(n10708), .ZN(n10710) );
  OAI211_X1 U13176 ( .C1(n13224), .C2(n10712), .A(n10711), .B(n10710), .ZN(
        P2_U3261) );
  XNOR2_X1 U13177 ( .A(n13616), .B(n13843), .ZN(n13782) );
  XNOR2_X1 U13178 ( .A(n10713), .B(n13782), .ZN(n10718) );
  INV_X1 U13179 ( .A(n10718), .ZN(n10786) );
  XOR2_X1 U13180 ( .A(n13782), .B(n10714), .Z(n10715) );
  NOR2_X1 U13181 ( .A1(n10715), .A2(n14795), .ZN(n10717) );
  AOI211_X1 U13182 ( .C1(n10718), .C2(n14723), .A(n10717), .B(n10716), .ZN(
        n10785) );
  MUX2_X1 U13183 ( .A(n10719), .B(n10785), .S(n14120), .Z(n10725) );
  AOI21_X1 U13184 ( .B1(n13616), .B2(n10720), .A(n10764), .ZN(n10783) );
  OAI22_X1 U13185 ( .A1(n14712), .A2(n10722), .B1(n10721), .B2(n14116), .ZN(
        n10723) );
  AOI21_X1 U13186 ( .B1(n10783), .B2(n12062), .A(n10723), .ZN(n10724) );
  OAI211_X1 U13187 ( .C1(n10786), .C2(n14139), .A(n10725), .B(n10724), .ZN(
        P1_U3287) );
  AOI211_X1 U13188 ( .C1(n10727), .C2(n14983), .A(n10726), .B(n10840), .ZN(
        n10728) );
  OAI21_X1 U13189 ( .B1(n13371), .B2(n10729), .A(n10728), .ZN(n10734) );
  INV_X1 U13190 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10730) );
  OAI22_X1 U13191 ( .A1(n13431), .A2(n10839), .B1(n10105), .B2(n10730), .ZN(
        n10731) );
  AOI21_X1 U13192 ( .B1(n10734), .B2(n10105), .A(n10731), .ZN(n10732) );
  INV_X1 U13193 ( .A(n10732), .ZN(P2_U3445) );
  OAI22_X1 U13194 ( .A1(n13378), .A2(n10839), .B1(n15002), .B2(n7539), .ZN(
        n10733) );
  AOI21_X1 U13195 ( .B1(n10734), .B2(n15002), .A(n10733), .ZN(n10735) );
  INV_X1 U13196 ( .A(n10735), .ZN(P2_U3504) );
  INV_X1 U13197 ( .A(n10736), .ZN(n10737) );
  NAND2_X1 U13198 ( .A1(n13047), .A2(n12834), .ZN(n10739) );
  XNOR2_X1 U13199 ( .A(n14939), .B(n12915), .ZN(n10740) );
  XNOR2_X1 U13200 ( .A(n10739), .B(n10740), .ZN(n10793) );
  INV_X1 U13201 ( .A(n10739), .ZN(n10741) );
  AOI22_X1 U13202 ( .A1(n10794), .A2(n10793), .B1(n10741), .B2(n10740), .ZN(
        n10747) );
  NOR2_X1 U13203 ( .A1(n10742), .A2(n6452), .ZN(n10745) );
  XNOR2_X1 U13204 ( .A(n10743), .B(n12915), .ZN(n10744) );
  NOR2_X1 U13205 ( .A1(n10745), .A2(n10744), .ZN(n10834) );
  AOI21_X1 U13206 ( .B1(n10745), .B2(n10744), .A(n10834), .ZN(n10746) );
  NAND2_X1 U13207 ( .A1(n10747), .A2(n10746), .ZN(n10836) );
  OAI21_X1 U13208 ( .B1(n10747), .B2(n10746), .A(n10836), .ZN(n10753) );
  NAND2_X1 U13209 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14842) );
  OAI21_X1 U13210 ( .B1(n14488), .B2(n6885), .A(n14842), .ZN(n10752) );
  NAND2_X1 U13211 ( .A1(n10748), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14495) );
  OAI22_X1 U13212 ( .A1(n10750), .A2(n14491), .B1(n10749), .B2(n14495), .ZN(
        n10751) );
  AOI211_X1 U13213 ( .C1(n10753), .C2(n12957), .A(n10752), .B(n10751), .ZN(
        n10754) );
  INV_X1 U13214 ( .A(n10754), .ZN(P2_U3202) );
  OAI21_X1 U13215 ( .B1(n10756), .B2(n10757), .A(n10755), .ZN(n14780) );
  INV_X1 U13216 ( .A(n14780), .ZN(n10771) );
  XNOR2_X1 U13217 ( .A(n10758), .B(n10757), .ZN(n10762) );
  NAND2_X1 U13218 ( .A1(n14780), .A2(n14723), .ZN(n10761) );
  NAND2_X1 U13219 ( .A1(n13843), .A2(n13551), .ZN(n10760) );
  NAND2_X1 U13220 ( .A1(n13841), .A2(n14645), .ZN(n10759) );
  AND2_X1 U13221 ( .A1(n10760), .A2(n10759), .ZN(n10869) );
  OAI211_X1 U13222 ( .C1(n14795), .C2(n10762), .A(n10761), .B(n10869), .ZN(
        n14778) );
  NAND2_X1 U13223 ( .A1(n14778), .A2(n14120), .ZN(n10770) );
  INV_X1 U13224 ( .A(n10867), .ZN(n10763) );
  OAI22_X1 U13225 ( .A1(n14120), .A2(n12112), .B1(n10763), .B2(n14116), .ZN(
        n10768) );
  OR2_X1 U13226 ( .A1(n10764), .A2(n14776), .ZN(n10765) );
  NAND2_X1 U13227 ( .A1(n10766), .A2(n10765), .ZN(n14777) );
  NOR2_X1 U13228 ( .A1(n14777), .A2(n11124), .ZN(n10767) );
  AOI211_X1 U13229 ( .C1(n14735), .C2(n13620), .A(n10768), .B(n10767), .ZN(
        n10769) );
  OAI211_X1 U13230 ( .C1(n10771), .C2(n14139), .A(n10770), .B(n10769), .ZN(
        P1_U3286) );
  INV_X1 U13231 ( .A(n10772), .ZN(n10782) );
  OAI211_X1 U13232 ( .C1(n10775), .C2(n10774), .A(n10773), .B(n12341), .ZN(
        n10781) );
  OAI22_X1 U13233 ( .A1(n12360), .A2(n10777), .B1(n12314), .B2(n10776), .ZN(
        n10778) );
  AOI211_X1 U13234 ( .C1(n12311), .C2(n12378), .A(n10779), .B(n10778), .ZN(
        n10780) );
  OAI211_X1 U13235 ( .C1(n10782), .C2(n11345), .A(n10781), .B(n10780), .ZN(
        P3_U3179) );
  AOI22_X1 U13236 ( .A1(n10783), .A2(n14730), .B1(n14786), .B2(n13616), .ZN(
        n10784) );
  OAI211_X1 U13237 ( .C1(n14745), .C2(n10786), .A(n10785), .B(n10784), .ZN(
        n10789) );
  NAND2_X1 U13238 ( .A1(n10789), .A2(n14819), .ZN(n10787) );
  OAI21_X1 U13239 ( .B1(n14819), .B2(n10788), .A(n10787), .ZN(P1_U3534) );
  INV_X1 U13240 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n12137) );
  NAND2_X1 U13241 ( .A1(n10789), .A2(n14807), .ZN(n10790) );
  OAI21_X1 U13242 ( .B1(n14807), .B2(n12137), .A(n10790), .ZN(P1_U3477) );
  INV_X1 U13243 ( .A(n14495), .ZN(n13016) );
  INV_X1 U13244 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U13245 ( .A1(n13014), .A2(n14939), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10791) );
  OAI21_X1 U13246 ( .B1(n10792), .B2(n14491), .A(n10791), .ZN(n10797) );
  XNOR2_X1 U13247 ( .A(n10794), .B(n10793), .ZN(n10795) );
  NOR2_X1 U13248 ( .A1(n10795), .A2(n14490), .ZN(n10796) );
  AOI211_X1 U13249 ( .C1(n13016), .C2(n13050), .A(n10797), .B(n10796), .ZN(
        n10798) );
  INV_X1 U13250 ( .A(n10798), .ZN(P2_U3190) );
  AOI21_X1 U13251 ( .B1(n10799), .B2(n7088), .A(n13371), .ZN(n10803) );
  NAND2_X1 U13252 ( .A1(n13044), .A2(n14484), .ZN(n10801) );
  NAND2_X1 U13253 ( .A1(n13042), .A2(n13013), .ZN(n10800) );
  NAND2_X1 U13254 ( .A1(n10801), .A2(n10800), .ZN(n10949) );
  AOI21_X1 U13255 ( .B1(n10803), .B2(n10802), .A(n10949), .ZN(n10921) );
  OAI21_X1 U13256 ( .B1(n10805), .B2(n7088), .A(n10804), .ZN(n10919) );
  OAI211_X1 U13257 ( .C1(n10806), .C2(n10927), .A(n10978), .B(n6452), .ZN(
        n10920) );
  OAI22_X1 U13258 ( .A1(n14948), .A2(n9796), .B1(n10952), .B2(n13295), .ZN(
        n10807) );
  AOI21_X1 U13259 ( .B1(n14502), .B2(n10954), .A(n10807), .ZN(n10808) );
  OAI21_X1 U13260 ( .B1(n10920), .B2(n13302), .A(n10808), .ZN(n10809) );
  AOI21_X1 U13261 ( .B1(n10919), .B2(n14510), .A(n10809), .ZN(n10810) );
  OAI21_X1 U13262 ( .B1(n14951), .B2(n10921), .A(n10810), .ZN(P2_U3258) );
  OAI21_X1 U13263 ( .B1(n10813), .B2(n10812), .A(n10811), .ZN(n10992) );
  OAI211_X1 U13264 ( .C1(n10816), .C2(n10815), .A(n10814), .B(n12762), .ZN(
        n10819) );
  OAI22_X1 U13265 ( .A1(n10862), .A2(n12683), .B1(n11205), .B2(n12759), .ZN(
        n10817) );
  INV_X1 U13266 ( .A(n10817), .ZN(n10818) );
  NAND2_X1 U13267 ( .A1(n10819), .A2(n10818), .ZN(n10989) );
  AOI21_X1 U13268 ( .B1(n14475), .B2(n10992), .A(n10989), .ZN(n10824) );
  AOI22_X1 U13269 ( .A1(n8743), .A2(n10820), .B1(n15131), .B2(
        P3_REG1_REG_7__SCAN_IN), .ZN(n10821) );
  OAI21_X1 U13270 ( .B1(n10824), .B2(n15131), .A(n10821), .ZN(P3_U3466) );
  OAI22_X1 U13271 ( .A1(n10988), .A2(n12818), .B1(n15129), .B2(n8237), .ZN(
        n10822) );
  INV_X1 U13272 ( .A(n10822), .ZN(n10823) );
  OAI21_X1 U13273 ( .B1(n10824), .B2(n15127), .A(n10823), .ZN(P3_U3411) );
  NAND2_X1 U13274 ( .A1(n12385), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10825) );
  OAI21_X1 U13275 ( .B1(n10826), .B2(n12385), .A(n10825), .ZN(P3_U3521) );
  INV_X1 U13276 ( .A(SI_23_), .ZN(n10830) );
  NAND2_X1 U13277 ( .A1(n10827), .A2(n14422), .ZN(n10829) );
  OAI211_X1 U13278 ( .C1(n10830), .C2(n12829), .A(n10829), .B(n10828), .ZN(
        P3_U3272) );
  AND2_X1 U13279 ( .A1(n13045), .A2(n13217), .ZN(n10833) );
  XNOR2_X1 U13280 ( .A(n10831), .B(n12915), .ZN(n10832) );
  NOR2_X1 U13281 ( .A1(n10833), .A2(n10832), .ZN(n10847) );
  AOI21_X1 U13282 ( .B1(n10833), .B2(n10832), .A(n10847), .ZN(n10838) );
  INV_X1 U13283 ( .A(n10834), .ZN(n10835) );
  NAND2_X1 U13284 ( .A1(n10836), .A2(n10835), .ZN(n10837) );
  OAI21_X1 U13285 ( .B1(n10838), .B2(n10837), .A(n10849), .ZN(n10845) );
  NOR2_X1 U13286 ( .A1(n14488), .A2(n10839), .ZN(n10844) );
  NAND2_X1 U13287 ( .A1(n10840), .A2(n12983), .ZN(n10841) );
  NAND2_X1 U13288 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n14857) );
  OAI211_X1 U13289 ( .C1(n14495), .C2(n10842), .A(n10841), .B(n14857), .ZN(
        n10843) );
  AOI211_X1 U13290 ( .C1(n10845), .C2(n12957), .A(n10844), .B(n10843), .ZN(
        n10846) );
  INV_X1 U13291 ( .A(n10846), .ZN(P2_U3199) );
  INV_X1 U13292 ( .A(n10847), .ZN(n10848) );
  XNOR2_X1 U13293 ( .A(n10855), .B(n12915), .ZN(n10945) );
  NAND2_X1 U13294 ( .A1(n13044), .A2(n12834), .ZN(n10946) );
  XOR2_X1 U13295 ( .A(n10945), .B(n10946), .Z(n10947) );
  XNOR2_X1 U13296 ( .A(n10948), .B(n10947), .ZN(n10857) );
  INV_X1 U13297 ( .A(n10850), .ZN(n10853) );
  NAND2_X1 U13298 ( .A1(n10851), .A2(n12983), .ZN(n10852) );
  NAND2_X1 U13299 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13065) );
  OAI211_X1 U13300 ( .C1(n14495), .C2(n10853), .A(n10852), .B(n13065), .ZN(
        n10854) );
  AOI21_X1 U13301 ( .B1(n10855), .B2(n13014), .A(n10854), .ZN(n10856) );
  OAI21_X1 U13302 ( .B1(n10857), .B2(n14490), .A(n10856), .ZN(P2_U3211) );
  INV_X1 U13303 ( .A(n10858), .ZN(n10987) );
  OAI211_X1 U13304 ( .C1(n10861), .C2(n10860), .A(n10859), .B(n12341), .ZN(
        n10866) );
  OAI22_X1 U13305 ( .A1(n12360), .A2(n10988), .B1(n12314), .B2(n10862), .ZN(
        n10863) );
  AOI211_X1 U13306 ( .C1(n12311), .C2(n12377), .A(n10864), .B(n10863), .ZN(
        n10865) );
  OAI211_X1 U13307 ( .C1(n10987), .C2(n11345), .A(n10866), .B(n10865), .ZN(
        P3_U3153) );
  INV_X1 U13308 ( .A(n14659), .ZN(n13563) );
  NAND2_X1 U13309 ( .A1(n13563), .A2(n10867), .ZN(n10868) );
  NAND2_X1 U13310 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13893) );
  OAI211_X1 U13311 ( .C1(n10869), .C2(n14649), .A(n10868), .B(n13893), .ZN(
        n10878) );
  AOI22_X1 U13312 ( .A1(n13620), .A2(n11966), .B1(n12223), .B2(n13842), .ZN(
        n10932) );
  NAND2_X1 U13313 ( .A1(n13620), .A2(n12222), .ZN(n10871) );
  NAND2_X1 U13314 ( .A1(n13842), .A2(n11966), .ZN(n10870) );
  NAND2_X1 U13315 ( .A1(n10871), .A2(n10870), .ZN(n10872) );
  XNOR2_X1 U13316 ( .A(n10872), .B(n10393), .ZN(n10934) );
  XOR2_X1 U13317 ( .A(n10932), .B(n10934), .Z(n10876) );
  AOI211_X1 U13318 ( .C1(n10876), .C2(n10875), .A(n14651), .B(n10936), .ZN(
        n10877) );
  AOI211_X1 U13319 ( .C1(n14657), .C2(n13620), .A(n10878), .B(n10877), .ZN(
        n10879) );
  INV_X1 U13320 ( .A(n10879), .ZN(P1_U3213) );
  INV_X1 U13321 ( .A(n11826), .ZN(n10883) );
  NAND2_X1 U13322 ( .A1(n10880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10881) );
  XNOR2_X1 U13323 ( .A(n10881), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13951) );
  INV_X1 U13324 ( .A(n13951), .ZN(n13944) );
  OAI222_X1 U13325 ( .A1(n6454), .A2(n10882), .B1(n14286), .B2(n10883), .C1(
        P1_U3086), .C2(n13944), .ZN(P1_U3337) );
  INV_X1 U13326 ( .A(n13124), .ZN(n13118) );
  OAI222_X1 U13327 ( .A1(n13458), .A2(n10884), .B1(n13467), .B2(n10883), .C1(
        P2_U3088), .C2(n13118), .ZN(P2_U3309) );
  INV_X1 U13328 ( .A(n15071), .ZN(n10908) );
  NOR2_X1 U13329 ( .A1(n10908), .A2(n10887), .ZN(n10888) );
  NOR2_X1 U13330 ( .A1(n15065), .A2(n15064), .ZN(n15063) );
  AOI22_X1 U13331 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n15101), .B1(n10904), 
        .B2(n10897), .ZN(n15089) );
  AOI21_X1 U13332 ( .B1(n11411), .B2(n10889), .A(n11132), .ZN(n10918) );
  INV_X1 U13333 ( .A(n10890), .ZN(n10891) );
  AOI22_X1 U13334 ( .A1(n10893), .A2(n10892), .B1(n10906), .B2(n10891), .ZN(
        n15068) );
  INV_X1 U13335 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10894) );
  MUX2_X1 U13336 ( .A(n15065), .B(n10894), .S(n6622), .Z(n10895) );
  NOR2_X1 U13337 ( .A1(n10895), .A2(n10908), .ZN(n15066) );
  NOR2_X1 U13338 ( .A1(n15068), .A2(n15066), .ZN(n15095) );
  AND2_X1 U13339 ( .A1(n10895), .A2(n10908), .ZN(n15094) );
  INV_X1 U13340 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10896) );
  MUX2_X1 U13341 ( .A(n10897), .B(n10896), .S(n6622), .Z(n10898) );
  NAND2_X1 U13342 ( .A1(n10898), .A2(n15101), .ZN(n10901) );
  INV_X1 U13343 ( .A(n10898), .ZN(n10899) );
  NAND2_X1 U13344 ( .A1(n10899), .A2(n10904), .ZN(n10900) );
  AND2_X1 U13345 ( .A1(n10901), .A2(n10900), .ZN(n15093) );
  NAND2_X1 U13346 ( .A1(n15098), .A2(n10901), .ZN(n10903) );
  MUX2_X1 U13347 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6622), .Z(n11142) );
  XNOR2_X1 U13348 ( .A(n11142), .B(n11143), .ZN(n10902) );
  NAND2_X1 U13349 ( .A1(n10903), .A2(n10902), .ZN(n11146) );
  OAI21_X1 U13350 ( .B1(n10903), .B2(n10902), .A(n11146), .ZN(n10916) );
  AOI22_X1 U13351 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n10904), .B1(n15101), 
        .B2(n10896), .ZN(n15084) );
  OAI21_X1 U13352 ( .B1(n10906), .B2(n10301), .A(n10905), .ZN(n10907) );
  NAND2_X1 U13353 ( .A1(n15071), .A2(n10907), .ZN(n10909) );
  XNOR2_X1 U13354 ( .A(n10908), .B(n10907), .ZN(n15077) );
  NAND2_X1 U13355 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15077), .ZN(n15076) );
  NAND2_X1 U13356 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n10910), .ZN(n11138) );
  OAI21_X1 U13357 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n10910), .A(n11138), 
        .ZN(n10911) );
  NAND2_X1 U13358 ( .A1(n10911), .A2(n15086), .ZN(n10914) );
  INV_X1 U13359 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n10912) );
  NOR2_X1 U13360 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10912), .ZN(n11558) );
  AOI21_X1 U13361 ( .B1(n15075), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11558), 
        .ZN(n10913) );
  OAI211_X1 U13362 ( .C1(n15070), .C2(n11137), .A(n10914), .B(n10913), .ZN(
        n10915) );
  AOI21_X1 U13363 ( .B1(n10916), .B2(n15055), .A(n10915), .ZN(n10917) );
  OAI21_X1 U13364 ( .B1(n10918), .B2(n15091), .A(n10917), .ZN(P3_U3193) );
  INV_X1 U13365 ( .A(n10919), .ZN(n10922) );
  OAI211_X1 U13366 ( .C1(n10922), .C2(n14530), .A(n10921), .B(n10920), .ZN(
        n10929) );
  INV_X1 U13367 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10923) );
  OAI22_X1 U13368 ( .A1(n13431), .A2(n10927), .B1(n10105), .B2(n10923), .ZN(
        n10924) );
  AOI21_X1 U13369 ( .B1(n10929), .B2(n10105), .A(n10924), .ZN(n10925) );
  INV_X1 U13370 ( .A(n10925), .ZN(P2_U3451) );
  OAI22_X1 U13371 ( .A1(n13378), .A2(n10927), .B1(n15002), .B2(n10926), .ZN(
        n10928) );
  AOI21_X1 U13372 ( .B1(n10929), .B2(n15002), .A(n10928), .ZN(n10930) );
  INV_X1 U13373 ( .A(n10930), .ZN(P2_U3506) );
  AOI22_X1 U13374 ( .A1(n14787), .A2(n11966), .B1(n12223), .B2(n13841), .ZN(
        n11287) );
  AOI22_X1 U13375 ( .A1(n14787), .A2(n12222), .B1(n11966), .B2(n13841), .ZN(
        n10931) );
  XNOR2_X1 U13376 ( .A(n10931), .B(n10393), .ZN(n11286) );
  XOR2_X1 U13377 ( .A(n11287), .B(n11286), .Z(n10937) );
  INV_X1 U13378 ( .A(n10932), .ZN(n10933) );
  AND2_X1 U13379 ( .A1(n10934), .A2(n10933), .ZN(n10935) );
  OAI21_X1 U13380 ( .B1(n10937), .B2(n6600), .A(n11289), .ZN(n10943) );
  NAND2_X1 U13381 ( .A1(n14787), .A2(n14657), .ZN(n10940) );
  AOI21_X1 U13382 ( .B1(n14785), .B2(n14578), .A(n10938), .ZN(n10939) );
  OAI211_X1 U13383 ( .C1(n14659), .C2(n10941), .A(n10940), .B(n10939), .ZN(
        n10942) );
  AOI21_X1 U13384 ( .B1(n10943), .B2(n14576), .A(n10942), .ZN(n10944) );
  INV_X1 U13385 ( .A(n10944), .ZN(P1_U3221) );
  XNOR2_X1 U13386 ( .A(n10954), .B(n12915), .ZN(n11169) );
  NAND2_X1 U13387 ( .A1(n13043), .A2(n12834), .ZN(n11168) );
  XNOR2_X1 U13388 ( .A(n11169), .B(n11168), .ZN(n11171) );
  XNOR2_X1 U13389 ( .A(n11172), .B(n11171), .ZN(n10956) );
  NAND2_X1 U13390 ( .A1(n10949), .A2(n12983), .ZN(n10951) );
  AND2_X1 U13391 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14872) );
  INV_X1 U13392 ( .A(n14872), .ZN(n10950) );
  OAI211_X1 U13393 ( .C1(n14495), .C2(n10952), .A(n10951), .B(n10950), .ZN(
        n10953) );
  AOI21_X1 U13394 ( .B1(n10954), .B2(n13014), .A(n10953), .ZN(n10955) );
  OAI21_X1 U13395 ( .B1(n10956), .B2(n14490), .A(n10955), .ZN(P2_U3185) );
  INV_X1 U13396 ( .A(n11046), .ZN(n10965) );
  OAI211_X1 U13397 ( .C1(n10959), .C2(n10958), .A(n10957), .B(n12341), .ZN(
        n10964) );
  OAI22_X1 U13398 ( .A1(n12360), .A2(n11094), .B1(n12314), .B2(n10960), .ZN(
        n10961) );
  AOI211_X1 U13399 ( .C1(n12311), .C2(n12376), .A(n10962), .B(n10961), .ZN(
        n10963) );
  OAI211_X1 U13400 ( .C1(n10965), .C2(n11345), .A(n10964), .B(n10963), .ZN(
        P3_U3161) );
  NAND2_X1 U13401 ( .A1(n10967), .A2(n10966), .ZN(n10968) );
  NAND2_X1 U13402 ( .A1(n10969), .A2(n10968), .ZN(n10977) );
  OR2_X1 U13403 ( .A1(n10977), .A2(n11255), .ZN(n10976) );
  XNOR2_X1 U13404 ( .A(n10971), .B(n10970), .ZN(n10974) );
  NAND2_X1 U13405 ( .A1(n13043), .A2(n14484), .ZN(n10973) );
  NAND2_X1 U13406 ( .A1(n13041), .A2(n13013), .ZN(n10972) );
  NAND2_X1 U13407 ( .A1(n10973), .A2(n10972), .ZN(n11178) );
  AOI21_X1 U13408 ( .B1(n10974), .B2(n14535), .A(n11178), .ZN(n10975) );
  AND2_X1 U13409 ( .A1(n10976), .A2(n10975), .ZN(n14974) );
  INV_X1 U13410 ( .A(n10977), .ZN(n14972) );
  INV_X1 U13411 ( .A(n11167), .ZN(n11439) );
  AOI21_X1 U13412 ( .B1(n10978), .B2(n11173), .A(n13217), .ZN(n10979) );
  NAND2_X1 U13413 ( .A1(n10979), .A2(n11162), .ZN(n14969) );
  OAI22_X1 U13414 ( .A1(n14948), .A2(n9798), .B1(n11181), .B2(n13295), .ZN(
        n10980) );
  AOI21_X1 U13415 ( .B1(n14502), .B2(n11173), .A(n10980), .ZN(n10981) );
  OAI21_X1 U13416 ( .B1(n14969), .B2(n13302), .A(n10981), .ZN(n10982) );
  AOI21_X1 U13417 ( .B1(n14972), .B2(n11439), .A(n10982), .ZN(n10983) );
  OAI21_X1 U13418 ( .B1(n14974), .B2(n14951), .A(n10983), .ZN(P2_U3257) );
  INV_X1 U13419 ( .A(n11841), .ZN(n10985) );
  OAI222_X1 U13420 ( .A1(n13458), .A2(n12129), .B1(n13467), .B2(n10985), .C1(
        P2_U3088), .C2(n10984), .ZN(P2_U3308) );
  OAI222_X1 U13421 ( .A1(n6454), .A2(n10986), .B1(n14286), .B2(n10985), .C1(
        P1_U3086), .C2(n14155), .ZN(P1_U3336) );
  OAI22_X1 U13422 ( .A1(n12689), .A2(n10988), .B1(n10987), .B2(n15111), .ZN(
        n10991) );
  MUX2_X1 U13423 ( .A(n10989), .B(P3_REG2_REG_7__SCAN_IN), .S(n15119), .Z(
        n10990) );
  AOI211_X1 U13424 ( .C1(n12691), .C2(n10992), .A(n10991), .B(n10990), .ZN(
        n10993) );
  INV_X1 U13425 ( .A(n10993), .ZN(P3_U3226) );
  NAND2_X1 U13426 ( .A1(n10996), .A2(n13756), .ZN(n10999) );
  AOI22_X1 U13427 ( .A1(n13728), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6459), 
        .B2(n10997), .ZN(n10998) );
  XNOR2_X1 U13428 ( .A(n14698), .B(n13840), .ZN(n13788) );
  NAND2_X1 U13429 ( .A1(n11051), .A2(n11053), .ZN(n11050) );
  OR2_X1 U13430 ( .A1(n13840), .A2(n14698), .ZN(n11000) );
  NAND2_X1 U13431 ( .A1(n11050), .A2(n11000), .ZN(n11012) );
  NAND2_X1 U13432 ( .A1(n11001), .A2(n13756), .ZN(n11004) );
  AOI22_X1 U13433 ( .A1(n13728), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6459), 
        .B2(n11002), .ZN(n11003) );
  NAND2_X1 U13434 ( .A1(n6456), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U13435 ( .A1(n12051), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11009) );
  OR2_X1 U13436 ( .A1(n11005), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U13437 ( .A1(n11005), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11020) );
  AND2_X1 U13438 ( .A1(n11006), .A2(n11020), .ZN(n11359) );
  NAND2_X1 U13439 ( .A1(n12027), .A2(n11359), .ZN(n11008) );
  NAND2_X1 U13440 ( .A1(n12050), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11007) );
  NAND4_X1 U13441 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n13839) );
  INV_X1 U13442 ( .A(n13839), .ZN(n11351) );
  NAND2_X1 U13443 ( .A1(n13640), .A2(n11351), .ZN(n11011) );
  NAND2_X1 U13444 ( .A1(n11102), .A2(n11011), .ZN(n13787) );
  OAI21_X1 U13445 ( .B1(n11012), .B2(n13787), .A(n11118), .ZN(n14804) );
  INV_X1 U13446 ( .A(n13841), .ZN(n11013) );
  OR2_X1 U13447 ( .A1(n14787), .A2(n11013), .ZN(n11014) );
  NAND2_X1 U13448 ( .A1(n11015), .A2(n11014), .ZN(n11052) );
  INV_X1 U13449 ( .A(n11052), .ZN(n11016) );
  NAND2_X1 U13450 ( .A1(n14698), .A2(n11290), .ZN(n11017) );
  AND2_X1 U13451 ( .A1(n11018), .A2(n13787), .ZN(n14796) );
  NOR3_X1 U13452 ( .A1(n6479), .A2(n14796), .A3(n14126), .ZN(n11032) );
  INV_X1 U13453 ( .A(n13640), .ZN(n14800) );
  INV_X1 U13454 ( .A(n11121), .ZN(n11019) );
  OAI211_X1 U13455 ( .C1(n14800), .C2(n11060), .A(n11019), .B(n14730), .ZN(
        n11026) );
  NAND2_X1 U13456 ( .A1(n12051), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U13457 ( .A1(n11020), .A2(n11504), .ZN(n11021) );
  AND2_X1 U13458 ( .A1(n11105), .A2(n11021), .ZN(n11508) );
  NAND2_X1 U13459 ( .A1(n12027), .A2(n11508), .ZN(n11024) );
  NAND2_X1 U13460 ( .A1(n12050), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U13461 ( .A1(n6456), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11022) );
  NAND4_X1 U13462 ( .A1(n11025), .A2(n11024), .A3(n11023), .A4(n11022), .ZN(
        n13838) );
  NAND2_X1 U13463 ( .A1(n13838), .A2(n14645), .ZN(n11356) );
  AND2_X1 U13464 ( .A1(n11026), .A2(n11356), .ZN(n14798) );
  NAND2_X1 U13465 ( .A1(n13840), .A2(n13551), .ZN(n14797) );
  INV_X1 U13466 ( .A(n11359), .ZN(n11027) );
  OAI22_X1 U13467 ( .A1(n14697), .A2(n14797), .B1(n11027), .B2(n14116), .ZN(
        n11029) );
  NOR2_X1 U13468 ( .A1(n14800), .A2(n14712), .ZN(n11028) );
  AOI211_X1 U13469 ( .C1(n14697), .C2(P1_REG2_REG_10__SCAN_IN), .A(n11029), 
        .B(n11028), .ZN(n11030) );
  OAI21_X1 U13470 ( .B1(n14798), .B2(n14732), .A(n11030), .ZN(n11031) );
  AOI211_X1 U13471 ( .C1(n14804), .C2(n14124), .A(n11032), .B(n11031), .ZN(
        n11033) );
  INV_X1 U13472 ( .A(n11033), .ZN(P1_U3283) );
  INV_X1 U13473 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11034) );
  INV_X1 U13474 ( .A(n11861), .ZN(n11036) );
  OAI222_X1 U13475 ( .A1(n6454), .A2(n11034), .B1(n14286), .B2(n11036), .C1(
        P1_U3086), .C2(n13738), .ZN(P1_U3335) );
  OAI222_X1 U13476 ( .A1(n13458), .A2(n11037), .B1(n13467), .B2(n11036), .C1(
        P2_U3088), .C2(n11035), .ZN(P2_U3307) );
  OAI21_X1 U13477 ( .B1(n11040), .B2(n11039), .A(n11038), .ZN(n11091) );
  INV_X1 U13478 ( .A(n11091), .ZN(n11049) );
  OAI21_X1 U13479 ( .B1(n11043), .B2(n11042), .A(n11041), .ZN(n11044) );
  AOI222_X1 U13480 ( .A1(n12762), .A2(n11044), .B1(n12376), .B2(n12666), .C1(
        n12378), .C2(n12756), .ZN(n11089) );
  MUX2_X1 U13481 ( .A(n11045), .B(n11089), .S(n15117), .Z(n11048) );
  AOI22_X1 U13482 ( .A1(n14463), .A2(n11092), .B1(n12687), .B2(n11046), .ZN(
        n11047) );
  OAI211_X1 U13483 ( .C1(n11080), .C2(n11049), .A(n11048), .B(n11047), .ZN(
        P3_U3225) );
  OAI21_X1 U13484 ( .B1(n11051), .B2(n11053), .A(n11050), .ZN(n14700) );
  INV_X1 U13485 ( .A(n14700), .ZN(n11063) );
  NAND2_X1 U13486 ( .A1(n11052), .A2(n11053), .ZN(n11054) );
  AOI21_X1 U13487 ( .B1(n11055), .B2(n11054), .A(n14795), .ZN(n11059) );
  NAND2_X1 U13488 ( .A1(n13841), .A2(n13551), .ZN(n11057) );
  NAND2_X1 U13489 ( .A1(n13839), .A2(n14645), .ZN(n11056) );
  AND2_X1 U13490 ( .A1(n11057), .A2(n11056), .ZN(n11295) );
  INV_X1 U13491 ( .A(n11295), .ZN(n11058) );
  AOI211_X1 U13492 ( .C1(n14700), .C2(n14723), .A(n11059), .B(n11058), .ZN(
        n14703) );
  AOI211_X1 U13493 ( .C1(n14698), .C2(n11061), .A(n14789), .B(n11060), .ZN(
        n14699) );
  AOI21_X1 U13494 ( .B1(n14786), .B2(n14698), .A(n14699), .ZN(n11062) );
  OAI211_X1 U13495 ( .C1(n11063), .C2(n14745), .A(n14703), .B(n11062), .ZN(
        n11066) );
  NAND2_X1 U13496 ( .A1(n11066), .A2(n14819), .ZN(n11064) );
  OAI21_X1 U13497 ( .B1(n14819), .B2(n11065), .A(n11064), .ZN(P1_U3537) );
  NAND2_X1 U13498 ( .A1(n11066), .A2(n14807), .ZN(n11067) );
  OAI21_X1 U13499 ( .B1(n14807), .B2(n10612), .A(n11067), .ZN(P1_U3486) );
  XNOR2_X1 U13500 ( .A(n11069), .B(n11068), .ZN(n11082) );
  INV_X1 U13501 ( .A(n11082), .ZN(n11079) );
  OAI211_X1 U13502 ( .C1(n11072), .C2(n11071), .A(n11070), .B(n12762), .ZN(
        n11074) );
  AOI22_X1 U13503 ( .A1(n12756), .A2(n12377), .B1(n12375), .B2(n12666), .ZN(
        n11073) );
  NAND2_X1 U13504 ( .A1(n11074), .A2(n11073), .ZN(n11081) );
  NOR2_X1 U13505 ( .A1(n15117), .A2(n15065), .ZN(n11077) );
  INV_X1 U13506 ( .A(n11208), .ZN(n11075) );
  OAI22_X1 U13507 ( .A1(n12689), .A2(n11206), .B1(n11075), .B2(n15111), .ZN(
        n11076) );
  AOI211_X1 U13508 ( .C1(n11081), .C2(n15117), .A(n11077), .B(n11076), .ZN(
        n11078) );
  OAI21_X1 U13509 ( .B1(n11080), .B2(n11079), .A(n11078), .ZN(P3_U3224) );
  AOI21_X1 U13510 ( .B1(n11082), .B2(n14475), .A(n11081), .ZN(n11088) );
  AOI22_X1 U13511 ( .A1(n8743), .A2(n11083), .B1(P3_REG1_REG_9__SCAN_IN), .B2(
        n15131), .ZN(n11084) );
  OAI21_X1 U13512 ( .B1(n11088), .B2(n15131), .A(n11084), .ZN(P3_U3468) );
  INV_X1 U13513 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n11085) );
  OAI22_X1 U13514 ( .A1(n11206), .A2(n12818), .B1(n15129), .B2(n11085), .ZN(
        n11086) );
  INV_X1 U13515 ( .A(n11086), .ZN(n11087) );
  OAI21_X1 U13516 ( .B1(n11088), .B2(n15127), .A(n11087), .ZN(P3_U3417) );
  INV_X1 U13517 ( .A(n11089), .ZN(n11090) );
  AOI21_X1 U13518 ( .B1(n14475), .B2(n11091), .A(n11090), .ZN(n11097) );
  AOI22_X1 U13519 ( .A1(n8743), .A2(n11092), .B1(n15131), .B2(
        P3_REG1_REG_8__SCAN_IN), .ZN(n11093) );
  OAI21_X1 U13520 ( .B1(n11097), .B2(n15131), .A(n11093), .ZN(P3_U3467) );
  OAI22_X1 U13521 ( .A1(n11094), .A2(n12818), .B1(n15129), .B2(n8256), .ZN(
        n11095) );
  INV_X1 U13522 ( .A(n11095), .ZN(n11096) );
  OAI21_X1 U13523 ( .B1(n11097), .B2(n15127), .A(n11096), .ZN(P3_U3414) );
  NAND2_X1 U13524 ( .A1(n11098), .A2(n13756), .ZN(n11101) );
  AOI22_X1 U13525 ( .A1(n13728), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6459), 
        .B2(n11099), .ZN(n11100) );
  XNOR2_X1 U13526 ( .A(n13649), .B(n13838), .ZN(n13789) );
  INV_X1 U13527 ( .A(n13789), .ZN(n11119) );
  NAND2_X1 U13528 ( .A1(n11119), .A2(n11102), .ZN(n11103) );
  OAI211_X1 U13529 ( .C1(n6479), .C2(n11103), .A(n11214), .B(n14784), .ZN(
        n11116) );
  NAND2_X1 U13530 ( .A1(n13839), .A2(n13551), .ZN(n11115) );
  NAND2_X1 U13531 ( .A1(n12051), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11113) );
  INV_X1 U13532 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11104) );
  INV_X1 U13533 ( .A(n11226), .ZN(n11107) );
  NAND2_X1 U13534 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  NAND2_X1 U13535 ( .A1(n11107), .A2(n11106), .ZN(n14569) );
  INV_X1 U13536 ( .A(n14569), .ZN(n11108) );
  NAND2_X1 U13537 ( .A1(n12027), .A2(n11108), .ZN(n11112) );
  NAND2_X1 U13538 ( .A1(n11930), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U13539 ( .A1(n6456), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11110) );
  NAND4_X1 U13540 ( .A1(n11113), .A2(n11112), .A3(n11111), .A4(n11110), .ZN(
        n13837) );
  NAND2_X1 U13541 ( .A1(n13837), .A2(n14645), .ZN(n11114) );
  AND2_X1 U13542 ( .A1(n11115), .A2(n11114), .ZN(n11505) );
  NAND2_X1 U13543 ( .A1(n11116), .A2(n11505), .ZN(n14610) );
  INV_X1 U13544 ( .A(n14610), .ZN(n11127) );
  NAND2_X1 U13545 ( .A1(n11120), .A2(n11119), .ZN(n11221) );
  OAI21_X1 U13546 ( .B1(n11120), .B2(n11119), .A(n11221), .ZN(n14611) );
  INV_X1 U13547 ( .A(n13649), .ZN(n14607) );
  OAI21_X1 U13548 ( .B1(n11121), .B2(n14607), .A(n11224), .ZN(n14608) );
  AOI22_X1 U13549 ( .A1(n14697), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11508), 
        .B2(n14728), .ZN(n11123) );
  NAND2_X1 U13550 ( .A1(n13649), .A2(n14735), .ZN(n11122) );
  OAI211_X1 U13551 ( .C1(n14608), .C2(n11124), .A(n11123), .B(n11122), .ZN(
        n11125) );
  AOI21_X1 U13552 ( .B1(n14611), .B2(n14124), .A(n11125), .ZN(n11126) );
  OAI21_X1 U13553 ( .B1(n14739), .B2(n11127), .A(n11126), .ZN(P1_U3282) );
  INV_X1 U13554 ( .A(n11128), .ZN(n11129) );
  OAI222_X1 U13555 ( .A1(P3_U3151), .A2(n11130), .B1(n12832), .B2(n11129), 
        .C1(n12181), .C2(n12829), .ZN(P3_U3271) );
  NOR2_X1 U13556 ( .A1(n11143), .A2(n11131), .ZN(n11133) );
  INV_X1 U13557 ( .A(n14406), .ZN(n12393) );
  AOI22_X1 U13558 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12393), .B1(n14406), 
        .B2(n8330), .ZN(n11134) );
  AOI21_X1 U13559 ( .B1(n11135), .B2(n11134), .A(n12386), .ZN(n11154) );
  INV_X1 U13560 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14476) );
  AOI22_X1 U13561 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n14406), .B1(n12393), 
        .B2(n14476), .ZN(n11141) );
  NAND2_X1 U13562 ( .A1(n11137), .A2(n11136), .ZN(n11139) );
  OAI21_X1 U13563 ( .B1(n11141), .B2(n11140), .A(n12388), .ZN(n11152) );
  INV_X1 U13564 ( .A(n11142), .ZN(n11144) );
  NAND2_X1 U13565 ( .A1(n11144), .A2(n11143), .ZN(n11145) );
  AND2_X1 U13566 ( .A1(n11146), .A2(n11145), .ZN(n11148) );
  MUX2_X1 U13567 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6622), .Z(n12390) );
  XNOR2_X1 U13568 ( .A(n12390), .B(n12393), .ZN(n11147) );
  NAND3_X1 U13569 ( .A1(n11146), .A2(n11145), .A3(n11147), .ZN(n12391) );
  OAI211_X1 U13570 ( .C1(n11148), .C2(n11147), .A(n15055), .B(n12391), .ZN(
        n11150) );
  AND2_X1 U13571 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11643) );
  AOI21_X1 U13572 ( .B1(n15075), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11643), 
        .ZN(n11149) );
  OAI211_X1 U13573 ( .C1(n15070), .C2(n14406), .A(n11150), .B(n11149), .ZN(
        n11151) );
  AOI21_X1 U13574 ( .B1(n15086), .B2(n11152), .A(n11151), .ZN(n11153) );
  OAI21_X1 U13575 ( .B1(n11154), .B2(n15091), .A(n11153), .ZN(P3_U3194) );
  XNOR2_X1 U13576 ( .A(n11155), .B(n11156), .ZN(n11312) );
  XNOR2_X1 U13577 ( .A(n11157), .B(n11156), .ZN(n11160) );
  NAND2_X1 U13578 ( .A1(n13042), .A2(n14484), .ZN(n11159) );
  NAND2_X1 U13579 ( .A1(n13040), .A2(n14481), .ZN(n11158) );
  NAND2_X1 U13580 ( .A1(n11159), .A2(n11158), .ZN(n11278) );
  AOI21_X1 U13581 ( .B1(n11160), .B2(n14535), .A(n11278), .ZN(n11161) );
  OAI21_X1 U13582 ( .B1(n11312), .B2(n11255), .A(n11161), .ZN(n11313) );
  NAND2_X1 U13583 ( .A1(n11313), .A2(n13298), .ZN(n11166) );
  AOI211_X1 U13584 ( .C1(n11316), .C2(n11162), .A(n13217), .B(n11263), .ZN(
        n11314) );
  AOI22_X1 U13585 ( .A1(n14951), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11277), 
        .B2(n14941), .ZN(n11163) );
  OAI21_X1 U13586 ( .B1(n11319), .B2(n13205), .A(n11163), .ZN(n11164) );
  AOI21_X1 U13587 ( .B1(n11314), .B2(n14509), .A(n11164), .ZN(n11165) );
  OAI211_X1 U13588 ( .C1(n11312), .C2(n11167), .A(n11166), .B(n11165), .ZN(
        P2_U3256) );
  INV_X1 U13589 ( .A(n11168), .ZN(n11170) );
  AND2_X1 U13590 ( .A1(n13042), .A2(n13217), .ZN(n11175) );
  XNOR2_X1 U13591 ( .A(n11173), .B(n12915), .ZN(n11174) );
  NOR2_X1 U13592 ( .A1(n11174), .A2(n11175), .ZN(n11272) );
  AOI21_X1 U13593 ( .B1(n11175), .B2(n11174), .A(n11272), .ZN(n11176) );
  NAND2_X1 U13594 ( .A1(n11177), .A2(n11176), .ZN(n11274) );
  OAI21_X1 U13595 ( .B1(n11177), .B2(n11176), .A(n11274), .ZN(n11184) );
  NOR2_X1 U13596 ( .A1(n14488), .A2(n14970), .ZN(n11183) );
  NAND2_X1 U13597 ( .A1(n11178), .A2(n12983), .ZN(n11180) );
  OAI211_X1 U13598 ( .C1(n14495), .C2(n11181), .A(n11180), .B(n11179), .ZN(
        n11182) );
  AOI211_X1 U13599 ( .C1(n11184), .C2(n12957), .A(n11183), .B(n11182), .ZN(
        n11185) );
  INV_X1 U13600 ( .A(n11185), .ZN(P2_U3193) );
  INV_X1 U13601 ( .A(n11880), .ZN(n11188) );
  OAI222_X1 U13602 ( .A1(n6454), .A2(n11186), .B1(n14286), .B2(n11188), .C1(
        P1_U3086), .C2(n13572), .ZN(P1_U3334) );
  OAI222_X1 U13603 ( .A1(n13458), .A2(n11189), .B1(n13467), .B2(n11188), .C1(
        n11187), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI211_X1 U13604 ( .C1(n11191), .C2(n11190), .A(n11402), .B(n12762), .ZN(
        n11193) );
  AOI22_X1 U13605 ( .A1(n12374), .A2(n12666), .B1(n12756), .B2(n12376), .ZN(
        n11192) );
  NAND2_X1 U13606 ( .A1(n11193), .A2(n11192), .ZN(n11362) );
  INV_X1 U13607 ( .A(n11362), .ZN(n11200) );
  XNOR2_X1 U13608 ( .A(n11195), .B(n11194), .ZN(n11363) );
  AOI22_X1 U13609 ( .A1(n14463), .A2(n11196), .B1(n12687), .B2(n11336), .ZN(
        n11197) );
  OAI21_X1 U13610 ( .B1(n10897), .B2(n15117), .A(n11197), .ZN(n11198) );
  AOI21_X1 U13611 ( .B1(n11363), .B2(n12691), .A(n11198), .ZN(n11199) );
  OAI21_X1 U13612 ( .B1(n11200), .B2(n15119), .A(n11199), .ZN(P3_U3223) );
  INV_X1 U13613 ( .A(n11201), .ZN(n11202) );
  AOI21_X1 U13614 ( .B1(n11204), .B2(n11203), .A(n11202), .ZN(n11211) );
  NOR2_X1 U13615 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12142), .ZN(n15074) );
  OAI22_X1 U13616 ( .A1(n12360), .A2(n11206), .B1(n12314), .B2(n11205), .ZN(
        n11207) );
  AOI211_X1 U13617 ( .C1(n12311), .C2(n12375), .A(n15074), .B(n11207), .ZN(
        n11210) );
  NAND2_X1 U13618 ( .A1(n12356), .A2(n11208), .ZN(n11209) );
  OAI211_X1 U13619 ( .C1(n11211), .C2(n12347), .A(n11210), .B(n11209), .ZN(
        P3_U3171) );
  INV_X1 U13620 ( .A(n13838), .ZN(n11212) );
  OR2_X1 U13621 ( .A1(n13649), .A2(n11212), .ZN(n11213) );
  NAND2_X1 U13622 ( .A1(n11214), .A2(n11213), .ZN(n11219) );
  NAND2_X1 U13623 ( .A1(n11215), .A2(n13756), .ZN(n11218) );
  AOI22_X1 U13624 ( .A1(n13728), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11216), 
        .B2(n6459), .ZN(n11217) );
  XNOR2_X1 U13625 ( .A(n14564), .B(n13837), .ZN(n13791) );
  OAI21_X1 U13626 ( .B1(n11219), .B2(n13791), .A(n11374), .ZN(n14433) );
  INV_X1 U13627 ( .A(n13791), .ZN(n11222) );
  OAI21_X1 U13628 ( .B1(n11223), .B2(n11222), .A(n11381), .ZN(n14439) );
  AOI21_X1 U13629 ( .B1(n11224), .B2(n14564), .A(n14789), .ZN(n11225) );
  NAND2_X1 U13630 ( .A1(n11225), .A2(n11383), .ZN(n14435) );
  NOR2_X1 U13631 ( .A1(n14120), .A2(n9678), .ZN(n11235) );
  NAND2_X1 U13632 ( .A1(n13838), .A2(n13551), .ZN(n11233) );
  NAND2_X1 U13633 ( .A1(n6456), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11231) );
  NAND2_X1 U13634 ( .A1(n13730), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11230) );
  NAND2_X1 U13635 ( .A1(n11226), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11385) );
  OR2_X1 U13636 ( .A1(n11226), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11227) );
  AND2_X1 U13637 ( .A1(n11385), .A2(n11227), .ZN(n11738) );
  NAND2_X1 U13638 ( .A1(n12027), .A2(n11738), .ZN(n11229) );
  NAND2_X1 U13639 ( .A1(n11930), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11228) );
  NAND4_X1 U13640 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n13836) );
  NAND2_X1 U13641 ( .A1(n13836), .A2(n14645), .ZN(n11232) );
  NAND2_X1 U13642 ( .A1(n11233), .A2(n11232), .ZN(n14566) );
  INV_X1 U13643 ( .A(n14566), .ZN(n14434) );
  OAI22_X1 U13644 ( .A1(n14697), .A2(n14434), .B1(n14569), .B2(n14116), .ZN(
        n11234) );
  AOI211_X1 U13645 ( .C1(n14564), .C2(n14735), .A(n11235), .B(n11234), .ZN(
        n11236) );
  OAI21_X1 U13646 ( .B1(n14435), .B2(n14732), .A(n11236), .ZN(n11237) );
  AOI21_X1 U13647 ( .B1(n14439), .B2(n14124), .A(n11237), .ZN(n11238) );
  OAI21_X1 U13648 ( .B1(n14126), .B2(n14433), .A(n11238), .ZN(P1_U3281) );
  XNOR2_X1 U13649 ( .A(n11239), .B(n11241), .ZN(n14984) );
  INV_X1 U13650 ( .A(n14984), .ZN(n11252) );
  OAI21_X1 U13651 ( .B1(n11242), .B2(n11241), .A(n11240), .ZN(n11243) );
  NAND2_X1 U13652 ( .A1(n11243), .A2(n14535), .ZN(n11247) );
  NAND2_X1 U13653 ( .A1(n13040), .A2(n14484), .ZN(n11245) );
  NAND2_X1 U13654 ( .A1(n13038), .A2(n13013), .ZN(n11244) );
  NAND2_X1 U13655 ( .A1(n11245), .A2(n11244), .ZN(n11463) );
  INV_X1 U13656 ( .A(n11463), .ZN(n11246) );
  NAND2_X1 U13657 ( .A1(n11247), .A2(n11246), .ZN(n14990) );
  OAI211_X1 U13658 ( .C1(n11265), .C2(n14987), .A(n6452), .B(n11434), .ZN(
        n14985) );
  OAI22_X1 U13659 ( .A1(n14948), .A2(n9956), .B1(n11465), .B2(n13295), .ZN(
        n11248) );
  AOI21_X1 U13660 ( .B1(n11467), .B2(n14502), .A(n11248), .ZN(n11249) );
  OAI21_X1 U13661 ( .B1(n14985), .B2(n13302), .A(n11249), .ZN(n11250) );
  AOI21_X1 U13662 ( .B1(n14990), .B2(n14948), .A(n11250), .ZN(n11251) );
  OAI21_X1 U13663 ( .B1(n11252), .B2(n13224), .A(n11251), .ZN(P2_U3254) );
  INV_X1 U13664 ( .A(n11254), .ZN(n11256) );
  XNOR2_X1 U13665 ( .A(n11253), .B(n11256), .ZN(n14979) );
  INV_X1 U13666 ( .A(n11255), .ZN(n11425) );
  NAND2_X1 U13667 ( .A1(n14979), .A2(n11425), .ZN(n11262) );
  XNOR2_X1 U13668 ( .A(n11257), .B(n11256), .ZN(n11260) );
  NAND2_X1 U13669 ( .A1(n13041), .A2(n14484), .ZN(n11259) );
  NAND2_X1 U13670 ( .A1(n13039), .A2(n14481), .ZN(n11258) );
  NAND2_X1 U13671 ( .A1(n11259), .A2(n11258), .ZN(n11303) );
  AOI21_X1 U13672 ( .B1(n11260), .B2(n14535), .A(n11303), .ZN(n11261) );
  AND2_X1 U13673 ( .A1(n11262), .A2(n11261), .ZN(n14981) );
  OAI21_X1 U13674 ( .B1(n11263), .B2(n14977), .A(n6452), .ZN(n11264) );
  OR2_X1 U13675 ( .A1(n11265), .A2(n11264), .ZN(n14976) );
  OAI22_X1 U13676 ( .A1(n14948), .A2(n9800), .B1(n11306), .B2(n13295), .ZN(
        n11266) );
  AOI21_X1 U13677 ( .B1(n11308), .B2(n14502), .A(n11266), .ZN(n11267) );
  OAI21_X1 U13678 ( .B1(n14976), .B2(n13302), .A(n11267), .ZN(n11268) );
  AOI21_X1 U13679 ( .B1(n14979), .B2(n11439), .A(n11268), .ZN(n11269) );
  OAI21_X1 U13680 ( .B1(n14981), .B2(n14951), .A(n11269), .ZN(P2_U3255) );
  AND2_X1 U13681 ( .A1(n13041), .A2(n13217), .ZN(n11271) );
  XNOR2_X1 U13682 ( .A(n11316), .B(n12915), .ZN(n11270) );
  NOR2_X1 U13683 ( .A1(n11270), .A2(n11271), .ZN(n11300) );
  AOI21_X1 U13684 ( .B1(n11271), .B2(n11270), .A(n11300), .ZN(n11276) );
  INV_X1 U13685 ( .A(n11272), .ZN(n11273) );
  NAND2_X1 U13686 ( .A1(n11274), .A2(n11273), .ZN(n11275) );
  OAI21_X1 U13687 ( .B1(n11276), .B2(n11275), .A(n11302), .ZN(n11284) );
  NOR2_X1 U13688 ( .A1(n11319), .A2(n14488), .ZN(n11283) );
  INV_X1 U13689 ( .A(n11277), .ZN(n11281) );
  NAND2_X1 U13690 ( .A1(n11278), .A2(n12983), .ZN(n11280) );
  OAI211_X1 U13691 ( .C1(n14495), .C2(n11281), .A(n11280), .B(n11279), .ZN(
        n11282) );
  AOI211_X1 U13692 ( .C1(n11284), .C2(n12957), .A(n11283), .B(n11282), .ZN(
        n11285) );
  INV_X1 U13693 ( .A(n11285), .ZN(P2_U3203) );
  NOR2_X1 U13694 ( .A1(n11290), .A2(n11803), .ZN(n11291) );
  AOI21_X1 U13695 ( .B1(n14698), .B2(n11966), .A(n11291), .ZN(n11347) );
  INV_X1 U13696 ( .A(n11347), .ZN(n11292) );
  AOI22_X1 U13697 ( .A1(n14698), .A2(n12222), .B1(n11966), .B2(n13840), .ZN(
        n11293) );
  XNOR2_X1 U13698 ( .A(n11293), .B(n10393), .ZN(n11349) );
  XOR2_X1 U13699 ( .A(n11350), .B(n11349), .Z(n11299) );
  OAI22_X1 U13700 ( .A1(n14649), .A2(n11295), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11294), .ZN(n11296) );
  AOI21_X1 U13701 ( .B1(n14696), .B2(n13563), .A(n11296), .ZN(n11298) );
  NAND2_X1 U13702 ( .A1(n14698), .A2(n14657), .ZN(n11297) );
  OAI211_X1 U13703 ( .C1(n11299), .C2(n14651), .A(n11298), .B(n11297), .ZN(
        P1_U3231) );
  INV_X1 U13704 ( .A(n11300), .ZN(n11301) );
  NAND2_X1 U13705 ( .A1(n13040), .A2(n12834), .ZN(n11454) );
  XNOR2_X1 U13706 ( .A(n11308), .B(n12915), .ZN(n11453) );
  XOR2_X1 U13707 ( .A(n11454), .B(n11453), .Z(n11455) );
  XNOR2_X1 U13708 ( .A(n11456), .B(n11455), .ZN(n11310) );
  NAND2_X1 U13709 ( .A1(n11303), .A2(n12983), .ZN(n11305) );
  OAI211_X1 U13710 ( .C1(n14495), .C2(n11306), .A(n11305), .B(n11304), .ZN(
        n11307) );
  AOI21_X1 U13711 ( .B1(n11308), .B2(n13014), .A(n11307), .ZN(n11309) );
  OAI21_X1 U13712 ( .B1(n11310), .B2(n14490), .A(n11309), .ZN(P2_U3189) );
  INV_X1 U13713 ( .A(n11312), .ZN(n11315) );
  AOI211_X1 U13714 ( .C1(n8957), .C2(n11315), .A(n11314), .B(n11313), .ZN(
        n11322) );
  AOI22_X1 U13715 ( .A1(n8070), .A2(n11316), .B1(n14999), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11317) );
  OAI21_X1 U13716 ( .B1(n11322), .B2(n14999), .A(n11317), .ZN(P2_U3508) );
  INV_X1 U13717 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11318) );
  OAI22_X1 U13718 ( .A1(n11319), .A2(n13431), .B1(n10105), .B2(n11318), .ZN(
        n11320) );
  INV_X1 U13719 ( .A(n11320), .ZN(n11321) );
  OAI21_X1 U13720 ( .B1(n11322), .B2(n14991), .A(n11321), .ZN(P2_U3457) );
  OAI222_X1 U13721 ( .A1(P3_U3151), .A2(n11325), .B1(n12832), .B2(n11324), 
        .C1(n11323), .C2(n12829), .ZN(P3_U3269) );
  XNOR2_X1 U13722 ( .A(n11326), .B(n7043), .ZN(n11327) );
  OAI222_X1 U13723 ( .A1(n12759), .A2(n11328), .B1(n12683), .B2(n11646), .C1(
        n11327), .C2(n12680), .ZN(n14472) );
  INV_X1 U13724 ( .A(n14472), .ZN(n11335) );
  OAI21_X1 U13725 ( .B1(n11331), .B2(n11330), .A(n11329), .ZN(n14474) );
  INV_X1 U13726 ( .A(n14471), .ZN(n11648) );
  AOI22_X1 U13727 ( .A1(n14463), .A2(n11648), .B1(n12687), .B2(n11642), .ZN(
        n11332) );
  OAI21_X1 U13728 ( .B1(n8330), .B2(n15117), .A(n11332), .ZN(n11333) );
  AOI21_X1 U13729 ( .B1(n14474), .B2(n12691), .A(n11333), .ZN(n11334) );
  OAI21_X1 U13730 ( .B1(n11335), .B2(n15119), .A(n11334), .ZN(P3_U3221) );
  INV_X1 U13731 ( .A(n11336), .ZN(n11346) );
  AOI21_X1 U13732 ( .B1(n11338), .B2(n11337), .A(n12347), .ZN(n11340) );
  NAND2_X1 U13733 ( .A1(n11340), .A2(n11339), .ZN(n11344) );
  AND2_X1 U13734 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n15085) );
  OAI22_X1 U13735 ( .A1(n12360), .A2(n11367), .B1(n12314), .B2(n11341), .ZN(
        n11342) );
  AOI211_X1 U13736 ( .C1(n12311), .C2(n12374), .A(n15085), .B(n11342), .ZN(
        n11343) );
  OAI211_X1 U13737 ( .C1(n11346), .C2(n11345), .A(n11344), .B(n11343), .ZN(
        P3_U3157) );
  NOR2_X1 U13738 ( .A1(n11351), .A2(n11803), .ZN(n11352) );
  AOI21_X1 U13739 ( .B1(n13640), .B2(n11966), .A(n11352), .ZN(n11498) );
  AOI22_X1 U13740 ( .A1(n13640), .A2(n12222), .B1(n11966), .B2(n13839), .ZN(
        n11353) );
  XNOR2_X1 U13741 ( .A(n11353), .B(n10393), .ZN(n11497) );
  XOR2_X1 U13742 ( .A(n11498), .B(n11497), .Z(n11354) );
  OAI211_X1 U13743 ( .C1(n11355), .C2(n11354), .A(n11496), .B(n14576), .ZN(
        n11361) );
  AOI21_X1 U13744 ( .B1(n11356), .B2(n14797), .A(n14649), .ZN(n11357) );
  AOI211_X1 U13745 ( .C1(n13563), .C2(n11359), .A(n11358), .B(n11357), .ZN(
        n11360) );
  OAI211_X1 U13746 ( .C1(n14800), .C2(n13567), .A(n11361), .B(n11360), .ZN(
        P1_U3217) );
  AOI21_X1 U13747 ( .B1(n11363), .B2(n14475), .A(n11362), .ZN(n11365) );
  MUX2_X1 U13748 ( .A(n8291), .B(n11365), .S(n15129), .Z(n11364) );
  OAI21_X1 U13749 ( .B1(n11367), .B2(n12818), .A(n11364), .ZN(P3_U3420) );
  MUX2_X1 U13750 ( .A(n10896), .B(n11365), .S(n15133), .Z(n11366) );
  OAI21_X1 U13751 ( .B1(n11367), .B2(n12755), .A(n11366), .ZN(P3_U3469) );
  INV_X1 U13752 ( .A(n11368), .ZN(n11370) );
  OAI222_X1 U13753 ( .A1(n13458), .A2(n11371), .B1(n13467), .B2(n11370), .C1(
        n11369), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U13754 ( .A(n13837), .ZN(n11372) );
  NAND2_X1 U13755 ( .A1(n11375), .A2(n13756), .ZN(n11378) );
  AOI22_X1 U13756 ( .A1(n11376), .A2(n6459), .B1(n13728), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n11377) );
  INV_X1 U13757 ( .A(n13836), .ZN(n11732) );
  XNOR2_X1 U13758 ( .A(n13661), .B(n11732), .ZN(n13793) );
  OAI21_X1 U13759 ( .B1(n11379), .B2(n7214), .A(n11522), .ZN(n14253) );
  OAI21_X1 U13760 ( .B1(n11382), .B2(n13793), .A(n11529), .ZN(n14251) );
  NAND2_X1 U13761 ( .A1(n14251), .A2(n14124), .ZN(n11400) );
  AOI21_X1 U13762 ( .B1(n13661), .B2(n11383), .A(n11530), .ZN(n14247) );
  INV_X1 U13763 ( .A(n14247), .ZN(n11395) );
  INV_X1 U13764 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11384) );
  NAND2_X1 U13765 ( .A1(n11385), .A2(n11384), .ZN(n11386) );
  NAND2_X1 U13766 ( .A1(n11533), .A2(n11386), .ZN(n14561) );
  INV_X1 U13767 ( .A(n14561), .ZN(n11541) );
  NAND2_X1 U13768 ( .A1(n12027), .A2(n11541), .ZN(n11390) );
  NAND2_X1 U13769 ( .A1(n6456), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U13770 ( .A1(n11930), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11388) );
  NAND2_X1 U13771 ( .A1(n12051), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11387) );
  NAND4_X1 U13772 ( .A1(n11390), .A2(n11389), .A3(n11388), .A4(n11387), .ZN(
        n13835) );
  NAND2_X1 U13773 ( .A1(n13835), .A2(n14645), .ZN(n11392) );
  NAND2_X1 U13774 ( .A1(n13837), .A2(n13551), .ZN(n11391) );
  AND2_X1 U13775 ( .A1(n11392), .A2(n11391), .ZN(n14248) );
  NAND2_X1 U13776 ( .A1(n14728), .A2(n11738), .ZN(n11393) );
  OAI211_X1 U13777 ( .C1(n11395), .C2(n11394), .A(n14248), .B(n11393), .ZN(
        n11398) );
  OAI22_X1 U13778 ( .A1(n6857), .A2(n14712), .B1(n11396), .B2(n14120), .ZN(
        n11397) );
  AOI21_X1 U13779 ( .B1(n11398), .B2(n14120), .A(n11397), .ZN(n11399) );
  OAI211_X1 U13780 ( .C1(n14253), .C2(n14126), .A(n11400), .B(n11399), .ZN(
        P1_U3280) );
  NAND2_X1 U13781 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  XOR2_X1 U13782 ( .A(n11407), .B(n11403), .Z(n11404) );
  OAI222_X1 U13783 ( .A1(n12683), .A2(n11405), .B1(n12759), .B2(n11556), .C1(
        n11404), .C2(n12680), .ZN(n11550) );
  INV_X1 U13784 ( .A(n11550), .ZN(n11414) );
  OAI21_X1 U13785 ( .B1(n11408), .B2(n11407), .A(n11406), .ZN(n11551) );
  AOI22_X1 U13786 ( .A1(n14463), .A2(n11409), .B1(n12687), .B2(n11562), .ZN(
        n11410) );
  OAI21_X1 U13787 ( .B1(n11411), .B2(n15117), .A(n11410), .ZN(n11412) );
  AOI21_X1 U13788 ( .B1(n11551), .B2(n12691), .A(n11412), .ZN(n11413) );
  OAI21_X1 U13789 ( .B1(n11414), .B2(n15119), .A(n11413), .ZN(P3_U3222) );
  INV_X1 U13790 ( .A(n11911), .ZN(n11416) );
  NAND2_X1 U13791 ( .A1(n14275), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11415) );
  OAI211_X1 U13792 ( .C1(n11416), .C2(n14286), .A(n11415), .B(n13817), .ZN(
        P1_U3332) );
  NAND2_X1 U13793 ( .A1(n11911), .A2(n11417), .ZN(n11419) );
  OAI211_X1 U13794 ( .C1(n11420), .C2(n13458), .A(n11419), .B(n11418), .ZN(
        P2_U3304) );
  OR2_X1 U13795 ( .A1(n11239), .A2(n11421), .ZN(n11423) );
  NAND2_X1 U13796 ( .A1(n11423), .A2(n11422), .ZN(n11424) );
  XNOR2_X1 U13797 ( .A(n11424), .B(n11426), .ZN(n14540) );
  NAND2_X1 U13798 ( .A1(n14540), .A2(n11425), .ZN(n11433) );
  AOI21_X1 U13799 ( .B1(n11427), .B2(n11426), .A(n13371), .ZN(n11431) );
  NAND2_X1 U13800 ( .A1(n13039), .A2(n14484), .ZN(n11429) );
  NAND2_X1 U13801 ( .A1(n14483), .A2(n14481), .ZN(n11428) );
  NAND2_X1 U13802 ( .A1(n11429), .A2(n11428), .ZN(n11577) );
  AOI21_X1 U13803 ( .B1(n11431), .B2(n11430), .A(n11577), .ZN(n11432) );
  AOI21_X1 U13804 ( .B1(n11434), .B2(n11565), .A(n13217), .ZN(n11435) );
  NAND2_X1 U13805 ( .A1(n11435), .A2(n11475), .ZN(n14537) );
  AOI22_X1 U13806 ( .A1(n14951), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11573), 
        .B2(n14941), .ZN(n11437) );
  NAND2_X1 U13807 ( .A1(n11565), .A2(n14502), .ZN(n11436) );
  OAI211_X1 U13808 ( .C1(n14537), .C2(n13302), .A(n11437), .B(n11436), .ZN(
        n11438) );
  AOI21_X1 U13809 ( .B1(n14540), .B2(n11439), .A(n11438), .ZN(n11440) );
  OAI21_X1 U13810 ( .B1(n14542), .B2(n14951), .A(n11440), .ZN(P2_U3253) );
  OR2_X1 U13811 ( .A1(n11441), .A2(n11446), .ZN(n11660) );
  NAND2_X1 U13812 ( .A1(n11441), .A2(n11446), .ZN(n11442) );
  NAND3_X1 U13813 ( .A1(n11660), .A2(n12762), .A3(n11442), .ZN(n11444) );
  AOI22_X1 U13814 ( .A1(n12372), .A2(n12756), .B1(n12666), .B2(n12370), .ZN(
        n11443) );
  AND2_X1 U13815 ( .A1(n11444), .A2(n11443), .ZN(n11620) );
  XNOR2_X1 U13816 ( .A(n11445), .B(n11446), .ZN(n11618) );
  AOI22_X1 U13817 ( .A1(n15119), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n12687), 
        .B2(n11633), .ZN(n11447) );
  OAI21_X1 U13818 ( .B1(n11630), .B2(n12689), .A(n11447), .ZN(n11448) );
  AOI21_X1 U13819 ( .B1(n11618), .B2(n12691), .A(n11448), .ZN(n11449) );
  OAI21_X1 U13820 ( .B1(n11620), .B2(n15119), .A(n11449), .ZN(P3_U3219) );
  INV_X1 U13821 ( .A(n11450), .ZN(n11452) );
  INV_X1 U13822 ( .A(SI_27_), .ZN(n11451) );
  OAI222_X1 U13823 ( .A1(n6622), .A2(P3_U3151), .B1(n12832), .B2(n11452), .C1(
        n11451), .C2(n12829), .ZN(P3_U3268) );
  XNOR2_X1 U13824 ( .A(n11467), .B(n12873), .ZN(n11458) );
  NAND2_X1 U13825 ( .A1(n13039), .A2(n13217), .ZN(n11457) );
  NAND2_X1 U13826 ( .A1(n11458), .A2(n11457), .ZN(n11568) );
  OAI21_X1 U13827 ( .B1(n11458), .B2(n11457), .A(n11568), .ZN(n11460) );
  INV_X1 U13828 ( .A(n11569), .ZN(n11459) );
  AOI21_X1 U13829 ( .B1(n11461), .B2(n11460), .A(n11459), .ZN(n11469) );
  NOR2_X1 U13830 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11462), .ZN(n14887) );
  AOI21_X1 U13831 ( .B1(n11463), .B2(n12983), .A(n14887), .ZN(n11464) );
  OAI21_X1 U13832 ( .B1(n11465), .B2(n14495), .A(n11464), .ZN(n11466) );
  AOI21_X1 U13833 ( .B1(n11467), .B2(n13014), .A(n11466), .ZN(n11468) );
  OAI21_X1 U13834 ( .B1(n11469), .B2(n14490), .A(n11468), .ZN(P2_U3208) );
  NAND2_X1 U13835 ( .A1(n11471), .A2(n11470), .ZN(n11472) );
  XNOR2_X1 U13836 ( .A(n11472), .B(n11473), .ZN(n14531) );
  XOR2_X1 U13837 ( .A(n11474), .B(n11473), .Z(n14534) );
  INV_X1 U13838 ( .A(n13305), .ZN(n13212) );
  NAND2_X1 U13839 ( .A1(n11475), .A2(n14527), .ZN(n11476) );
  NAND2_X1 U13840 ( .A1(n11476), .A2(n6452), .ZN(n11477) );
  OR2_X1 U13841 ( .A1(n11477), .A2(n6590), .ZN(n14529) );
  NAND2_X1 U13842 ( .A1(n13037), .A2(n14481), .ZN(n11479) );
  NAND2_X1 U13843 ( .A1(n13038), .A2(n14484), .ZN(n11478) );
  AND2_X1 U13844 ( .A1(n11479), .A2(n11478), .ZN(n14528) );
  INV_X1 U13845 ( .A(n14528), .ZN(n11482) );
  OAI22_X1 U13846 ( .A1(n14948), .A2(n11480), .B1(n11613), .B2(n13295), .ZN(
        n11481) );
  AOI21_X1 U13847 ( .B1(n11482), .B2(n14948), .A(n11481), .ZN(n11484) );
  NAND2_X1 U13848 ( .A1(n14527), .A2(n14502), .ZN(n11483) );
  OAI211_X1 U13849 ( .C1(n14529), .C2(n13302), .A(n11484), .B(n11483), .ZN(
        n11485) );
  AOI21_X1 U13850 ( .B1(n14534), .B2(n13212), .A(n11485), .ZN(n11486) );
  OAI21_X1 U13851 ( .B1(n14531), .B2(n13224), .A(n11486), .ZN(P2_U3252) );
  XNOR2_X1 U13852 ( .A(n11487), .B(n11489), .ZN(n11488) );
  OAI222_X1 U13853 ( .A1(n12759), .A2(n11663), .B1(n12683), .B2(n11556), .C1(
        n12680), .C2(n11488), .ZN(n11651) );
  INV_X1 U13854 ( .A(n11651), .ZN(n11494) );
  XNOR2_X1 U13855 ( .A(n11490), .B(n11489), .ZN(n11652) );
  INV_X1 U13856 ( .A(n11519), .ZN(n11658) );
  AOI22_X1 U13857 ( .A1(n15119), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n12687), 
        .B2(n11514), .ZN(n11491) );
  OAI21_X1 U13858 ( .B1(n11658), .B2(n12689), .A(n11491), .ZN(n11492) );
  AOI21_X1 U13859 ( .B1(n11652), .B2(n12691), .A(n11492), .ZN(n11493) );
  OAI21_X1 U13860 ( .B1(n11494), .B2(n15119), .A(n11493), .ZN(P3_U3220) );
  AOI22_X1 U13861 ( .A1(n13649), .A2(n12222), .B1(n11966), .B2(n13838), .ZN(
        n11495) );
  XNOR2_X1 U13862 ( .A(n11495), .B(n10393), .ZN(n11718) );
  AOI22_X1 U13863 ( .A1(n13649), .A2(n11966), .B1(n12223), .B2(n13838), .ZN(
        n11719) );
  XNOR2_X1 U13864 ( .A(n11718), .B(n11719), .ZN(n11503) );
  INV_X1 U13865 ( .A(n11502), .ZN(n11500) );
  INV_X1 U13866 ( .A(n11503), .ZN(n11499) );
  INV_X1 U13867 ( .A(n11721), .ZN(n11501) );
  AOI21_X1 U13868 ( .B1(n11503), .B2(n11502), .A(n11501), .ZN(n11510) );
  OAI22_X1 U13869 ( .A1(n14649), .A2(n11505), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11504), .ZN(n11507) );
  NOR2_X1 U13870 ( .A1(n14607), .A2(n13567), .ZN(n11506) );
  AOI211_X1 U13871 ( .C1(n13563), .C2(n11508), .A(n11507), .B(n11506), .ZN(
        n11509) );
  OAI21_X1 U13872 ( .B1(n11510), .B2(n14651), .A(n11509), .ZN(P1_U3236) );
  XNOR2_X1 U13873 ( .A(n11511), .B(n12372), .ZN(n11512) );
  XNOR2_X1 U13874 ( .A(n11513), .B(n11512), .ZN(n11521) );
  NAND2_X1 U13875 ( .A1(n12356), .A2(n11514), .ZN(n11517) );
  NOR2_X1 U13876 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11515), .ZN(n12397) );
  AOI21_X1 U13877 ( .B1(n12311), .B2(n12371), .A(n12397), .ZN(n11516) );
  OAI211_X1 U13878 ( .C1(n11556), .C2(n12314), .A(n11517), .B(n11516), .ZN(
        n11518) );
  AOI21_X1 U13879 ( .B1(n11519), .B2(n12334), .A(n11518), .ZN(n11520) );
  OAI21_X1 U13880 ( .B1(n11521), .B2(n12347), .A(n11520), .ZN(P3_U3174) );
  NAND2_X1 U13881 ( .A1(n11523), .A2(n13756), .ZN(n11526) );
  AOI22_X1 U13882 ( .A1(n11524), .A2(n6459), .B1(n13728), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U13883 ( .A1(n14600), .A2(n11789), .ZN(n13665) );
  NAND2_X1 U13884 ( .A1(n11527), .A2(n13669), .ZN(n11580) );
  OAI21_X1 U13885 ( .B1(n11527), .B2(n13669), .A(n11580), .ZN(n14598) );
  OAI21_X1 U13886 ( .B1(n6588), .B2(n7217), .A(n7431), .ZN(n14603) );
  INV_X1 U13887 ( .A(n14603), .ZN(n11548) );
  INV_X1 U13888 ( .A(n14600), .ZN(n11585) );
  OAI21_X1 U13889 ( .B1(n11530), .B2(n11585), .A(n14730), .ZN(n11531) );
  OR2_X1 U13890 ( .A1(n11531), .A2(n11597), .ZN(n14601) );
  INV_X1 U13891 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11532) );
  AND2_X1 U13892 ( .A1(n11533), .A2(n11532), .ZN(n11534) );
  NOR2_X1 U13893 ( .A1(n11586), .A2(n11534), .ZN(n13564) );
  NAND2_X1 U13894 ( .A1(n13564), .A2(n12027), .ZN(n11538) );
  NAND2_X1 U13895 ( .A1(n6456), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U13896 ( .A1(n13730), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11536) );
  NAND2_X1 U13897 ( .A1(n11930), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11535) );
  NAND4_X1 U13898 ( .A1(n11538), .A2(n11537), .A3(n11536), .A4(n11535), .ZN(
        n13834) );
  NAND2_X1 U13899 ( .A1(n13834), .A2(n14645), .ZN(n11540) );
  NAND2_X1 U13900 ( .A1(n13836), .A2(n13551), .ZN(n11539) );
  NAND2_X1 U13901 ( .A1(n11540), .A2(n11539), .ZN(n14599) );
  INV_X1 U13902 ( .A(n14599), .ZN(n11544) );
  NAND2_X1 U13903 ( .A1(n14697), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11543) );
  NAND2_X1 U13904 ( .A1(n14728), .A2(n11541), .ZN(n11542) );
  OAI211_X1 U13905 ( .C1(n14739), .C2(n11544), .A(n11543), .B(n11542), .ZN(
        n11545) );
  AOI21_X1 U13906 ( .B1(n14600), .B2(n14735), .A(n11545), .ZN(n11546) );
  OAI21_X1 U13907 ( .B1(n14601), .B2(n14732), .A(n11546), .ZN(n11547) );
  AOI21_X1 U13908 ( .B1(n11548), .B2(n14124), .A(n11547), .ZN(n11549) );
  OAI21_X1 U13909 ( .B1(n14126), .B2(n14598), .A(n11549), .ZN(P1_U3279) );
  INV_X1 U13910 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11552) );
  AOI21_X1 U13911 ( .B1(n14475), .B2(n11551), .A(n11550), .ZN(n11554) );
  MUX2_X1 U13912 ( .A(n11552), .B(n11554), .S(n15133), .Z(n11553) );
  OAI21_X1 U13913 ( .B1(n11560), .B2(n12755), .A(n11553), .ZN(P3_U3470) );
  MUX2_X1 U13914 ( .A(n8306), .B(n11554), .S(n15129), .Z(n11555) );
  OAI21_X1 U13915 ( .B1(n11560), .B2(n12818), .A(n11555), .ZN(P3_U3423) );
  XNOR2_X1 U13916 ( .A(n11636), .B(n11637), .ZN(n11638) );
  XNOR2_X1 U13917 ( .A(n11638), .B(n11646), .ZN(n11564) );
  NOR2_X1 U13918 ( .A1(n12354), .A2(n11556), .ZN(n11557) );
  AOI211_X1 U13919 ( .C1(n12352), .C2(n12375), .A(n11558), .B(n11557), .ZN(
        n11559) );
  OAI21_X1 U13920 ( .B1(n11560), .B2(n12360), .A(n11559), .ZN(n11561) );
  AOI21_X1 U13921 ( .B1(n11562), .B2(n12356), .A(n11561), .ZN(n11563) );
  OAI21_X1 U13922 ( .B1(n11564), .B2(n12347), .A(n11563), .ZN(P3_U3176) );
  INV_X1 U13923 ( .A(n11565), .ZN(n14538) );
  AND2_X1 U13924 ( .A1(n13038), .A2(n13217), .ZN(n11567) );
  XNOR2_X1 U13925 ( .A(n11565), .B(n12915), .ZN(n11566) );
  NOR2_X1 U13926 ( .A1(n11566), .A2(n11567), .ZN(n11610) );
  AOI21_X1 U13927 ( .B1(n11567), .B2(n11566), .A(n11610), .ZN(n11571) );
  NAND2_X1 U13928 ( .A1(n11569), .A2(n11568), .ZN(n11570) );
  NAND2_X1 U13929 ( .A1(n11570), .A2(n11571), .ZN(n11612) );
  OAI21_X1 U13930 ( .B1(n11571), .B2(n11570), .A(n11612), .ZN(n11572) );
  NAND2_X1 U13931 ( .A1(n11572), .A2(n12957), .ZN(n11579) );
  INV_X1 U13932 ( .A(n11573), .ZN(n11574) );
  NOR2_X1 U13933 ( .A1(n14495), .A2(n11574), .ZN(n11575) );
  AOI211_X1 U13934 ( .C1(n12983), .C2(n11577), .A(n11576), .B(n11575), .ZN(
        n11578) );
  OAI211_X1 U13935 ( .C1(n14538), .C2(n14488), .A(n11579), .B(n11578), .ZN(
        P2_U3196) );
  NAND2_X1 U13936 ( .A1(n11580), .A2(n13664), .ZN(n11584) );
  NAND2_X1 U13937 ( .A1(n11581), .A2(n13756), .ZN(n11583) );
  AOI22_X1 U13938 ( .A1(n13728), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6459), 
        .B2(n14687), .ZN(n11582) );
  INV_X1 U13939 ( .A(n13834), .ZN(n11804) );
  NAND2_X1 U13940 ( .A1(n11799), .A2(n11804), .ZN(n13671) );
  NAND2_X1 U13941 ( .A1(n13672), .A2(n13671), .ZN(n13794) );
  OAI21_X1 U13942 ( .B1(n11584), .B2(n11700), .A(n11698), .ZN(n14591) );
  XNOR2_X1 U13943 ( .A(n11701), .B(n11700), .ZN(n14597) );
  NAND2_X1 U13944 ( .A1(n14597), .A2(n14124), .ZN(n11601) );
  INV_X1 U13945 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11596) );
  NOR2_X1 U13946 ( .A1(n11586), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11587) );
  OR2_X1 U13947 ( .A1(n11704), .A2(n11587), .ZN(n14581) );
  INV_X1 U13948 ( .A(n12027), .ZN(n11851) );
  NAND2_X1 U13949 ( .A1(n11930), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11589) );
  NAND2_X1 U13950 ( .A1(n6456), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11588) );
  AND2_X1 U13951 ( .A1(n11589), .A2(n11588), .ZN(n11591) );
  NAND2_X1 U13952 ( .A1(n12051), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11590) );
  OAI211_X1 U13953 ( .C1(n14581), .C2(n11851), .A(n11591), .B(n11590), .ZN(
        n13833) );
  NAND2_X1 U13954 ( .A1(n13833), .A2(n14645), .ZN(n11593) );
  NAND2_X1 U13955 ( .A1(n13835), .A2(n13551), .ZN(n11592) );
  AND2_X1 U13956 ( .A1(n11593), .A2(n11592), .ZN(n14592) );
  INV_X1 U13957 ( .A(n14592), .ZN(n11594) );
  AOI22_X1 U13958 ( .A1(n14120), .A2(n11594), .B1(n13564), .B2(n14728), .ZN(
        n11595) );
  OAI21_X1 U13959 ( .B1(n11596), .B2(n14120), .A(n11595), .ZN(n11599) );
  NAND2_X1 U13960 ( .A1(n11597), .A2(n14594), .ZN(n11710) );
  OAI211_X1 U13961 ( .C1(n11597), .C2(n14594), .A(n14730), .B(n11710), .ZN(
        n14593) );
  NOR2_X1 U13962 ( .A1(n14593), .A2(n14732), .ZN(n11598) );
  AOI211_X1 U13963 ( .C1(n14735), .C2(n11799), .A(n11599), .B(n11598), .ZN(
        n11600) );
  OAI211_X1 U13964 ( .C1(n14591), .C2(n14126), .A(n11601), .B(n11600), .ZN(
        P1_U3278) );
  XNOR2_X1 U13965 ( .A(n11602), .B(n11604), .ZN(n11603) );
  AOI222_X1 U13966 ( .A1(n12762), .A2(n11603), .B1(n12370), .B2(n12756), .C1(
        n12668), .C2(n12666), .ZN(n12750) );
  XNOR2_X1 U13967 ( .A(n11605), .B(n11604), .ZN(n12748) );
  INV_X1 U13968 ( .A(n12747), .ZN(n11607) );
  AOI22_X1 U13969 ( .A1(n15119), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12687), 
        .B2(n12293), .ZN(n11606) );
  OAI21_X1 U13970 ( .B1(n11607), .B2(n12689), .A(n11606), .ZN(n11608) );
  AOI21_X1 U13971 ( .B1(n12748), .B2(n12691), .A(n11608), .ZN(n11609) );
  OAI21_X1 U13972 ( .B1(n12750), .B2(n15119), .A(n11609), .ZN(P3_U3217) );
  INV_X1 U13973 ( .A(n11610), .ZN(n11611) );
  NAND2_X1 U13974 ( .A1(n14483), .A2(n13217), .ZN(n11755) );
  XNOR2_X1 U13975 ( .A(n14527), .B(n12915), .ZN(n11754) );
  XOR2_X1 U13976 ( .A(n11755), .B(n11754), .Z(n11757) );
  XNOR2_X1 U13977 ( .A(n11758), .B(n11757), .ZN(n11617) );
  NOR2_X1 U13978 ( .A1(n14495), .A2(n11613), .ZN(n11615) );
  OAI22_X1 U13979 ( .A1(n14528), .A2(n14491), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7688), .ZN(n11614) );
  AOI211_X1 U13980 ( .C1(n14527), .C2(n13014), .A(n11615), .B(n11614), .ZN(
        n11616) );
  OAI21_X1 U13981 ( .B1(n11617), .B2(n14490), .A(n11616), .ZN(P2_U3206) );
  NAND2_X1 U13982 ( .A1(n11618), .A2(n14475), .ZN(n11619) );
  AND2_X1 U13983 ( .A1(n11620), .A2(n11619), .ZN(n11623) );
  INV_X1 U13984 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11621) );
  MUX2_X1 U13985 ( .A(n11623), .B(n11621), .S(n15127), .Z(n11622) );
  OAI21_X1 U13986 ( .B1(n12818), .B2(n11630), .A(n11622), .ZN(P3_U3432) );
  INV_X1 U13987 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12413) );
  MUX2_X1 U13988 ( .A(n12413), .B(n11623), .S(n15133), .Z(n11624) );
  OAI21_X1 U13989 ( .B1(n12755), .B2(n11630), .A(n11624), .ZN(P3_U3473) );
  XNOR2_X1 U13990 ( .A(n11625), .B(n12371), .ZN(n11626) );
  XNOR2_X1 U13991 ( .A(n11627), .B(n11626), .ZN(n11635) );
  AND2_X1 U13992 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12417) );
  AOI21_X1 U13993 ( .B1(n12352), .B2(n12372), .A(n12417), .ZN(n11628) );
  OAI21_X1 U13994 ( .B1(n11629), .B2(n12354), .A(n11628), .ZN(n11632) );
  NOR2_X1 U13995 ( .A1(n11630), .A2(n12360), .ZN(n11631) );
  AOI211_X1 U13996 ( .C1(n11633), .C2(n12356), .A(n11632), .B(n11631), .ZN(
        n11634) );
  OAI21_X1 U13997 ( .B1(n11635), .B2(n12347), .A(n11634), .ZN(P3_U3155) );
  OAI22_X1 U13998 ( .A1(n11638), .A2(n12374), .B1(n11637), .B2(n11636), .ZN(
        n11641) );
  XNOR2_X1 U13999 ( .A(n11639), .B(n12373), .ZN(n11640) );
  XNOR2_X1 U14000 ( .A(n11641), .B(n11640), .ZN(n11650) );
  NAND2_X1 U14001 ( .A1(n12356), .A2(n11642), .ZN(n11645) );
  AOI21_X1 U14002 ( .B1(n12311), .B2(n12372), .A(n11643), .ZN(n11644) );
  OAI211_X1 U14003 ( .C1(n11646), .C2(n12314), .A(n11645), .B(n11644), .ZN(
        n11647) );
  AOI21_X1 U14004 ( .B1(n11648), .B2(n12334), .A(n11647), .ZN(n11649) );
  OAI21_X1 U14005 ( .B1(n11650), .B2(n12347), .A(n11649), .ZN(P3_U3164) );
  AOI21_X1 U14006 ( .B1(n11652), .B2(n14475), .A(n11651), .ZN(n11655) );
  MUX2_X1 U14007 ( .A(n11653), .B(n11655), .S(n15129), .Z(n11654) );
  OAI21_X1 U14008 ( .B1(n11658), .B2(n12818), .A(n11654), .ZN(P3_U3429) );
  INV_X1 U14009 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n11656) );
  MUX2_X1 U14010 ( .A(n11656), .B(n11655), .S(n15133), .Z(n11657) );
  OAI21_X1 U14011 ( .B1(n11658), .B2(n12755), .A(n11657), .ZN(P3_U3472) );
  NAND2_X1 U14012 ( .A1(n11660), .A2(n11659), .ZN(n11661) );
  XOR2_X1 U14013 ( .A(n11665), .B(n11661), .Z(n11662) );
  OAI222_X1 U14014 ( .A1(n12759), .A2(n12682), .B1(n12683), .B2(n11663), .C1(
        n11662), .C2(n12680), .ZN(n12751) );
  INV_X1 U14015 ( .A(n12751), .ZN(n11670) );
  XNOR2_X1 U14016 ( .A(n11664), .B(n11665), .ZN(n12752) );
  INV_X1 U14017 ( .A(n11666), .ZN(n12819) );
  AOI22_X1 U14018 ( .A1(n15119), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12687), 
        .B2(n12357), .ZN(n11667) );
  OAI21_X1 U14019 ( .B1(n12819), .B2(n12689), .A(n11667), .ZN(n11668) );
  AOI21_X1 U14020 ( .B1(n12752), .B2(n12691), .A(n11668), .ZN(n11669) );
  OAI21_X1 U14021 ( .B1(n11670), .B2(n15119), .A(n11669), .ZN(P3_U3218) );
  XNOR2_X1 U14022 ( .A(n11671), .B(n11672), .ZN(n14513) );
  XNOR2_X1 U14023 ( .A(n11673), .B(n11672), .ZN(n11674) );
  NAND2_X1 U14024 ( .A1(n11674), .A2(n14535), .ZN(n14517) );
  NAND2_X1 U14025 ( .A1(n13036), .A2(n13013), .ZN(n11676) );
  NAND2_X1 U14026 ( .A1(n13037), .A2(n14484), .ZN(n11675) );
  AND2_X1 U14027 ( .A1(n11676), .A2(n11675), .ZN(n14514) );
  OAI211_X1 U14028 ( .C1(n13295), .C2(n11764), .A(n14517), .B(n14514), .ZN(
        n11679) );
  OAI211_X1 U14029 ( .C1(n14506), .C2(n14516), .A(n6452), .B(n11686), .ZN(
        n14515) );
  AOI22_X1 U14030 ( .A1(n11767), .A2(n14502), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n14951), .ZN(n11677) );
  OAI21_X1 U14031 ( .B1(n14515), .B2(n13302), .A(n11677), .ZN(n11678) );
  AOI21_X1 U14032 ( .B1(n11679), .B2(n13298), .A(n11678), .ZN(n11680) );
  OAI21_X1 U14033 ( .B1(n13224), .B2(n14513), .A(n11680), .ZN(P2_U3250) );
  XNOR2_X1 U14034 ( .A(n11681), .B(n11691), .ZN(n13396) );
  INV_X1 U14035 ( .A(n13396), .ZN(n11694) );
  NAND2_X1 U14036 ( .A1(n13035), .A2(n13013), .ZN(n11683) );
  NAND2_X1 U14037 ( .A1(n14482), .A2(n14484), .ZN(n11682) );
  NAND2_X1 U14038 ( .A1(n11683), .A2(n11682), .ZN(n13397) );
  INV_X1 U14039 ( .A(n13397), .ZN(n11684) );
  OAI21_X1 U14040 ( .B1(n12948), .B2(n13295), .A(n11684), .ZN(n11685) );
  MUX2_X1 U14041 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n11685), .S(n14948), .Z(
        n11689) );
  AOI21_X1 U14042 ( .B1(n11686), .B2(n13399), .A(n13217), .ZN(n11687) );
  NAND2_X1 U14043 ( .A1(n11687), .A2(n11743), .ZN(n13402) );
  NOR2_X1 U14044 ( .A1(n13402), .A2(n13302), .ZN(n11688) );
  AOI211_X1 U14045 ( .C1(n14502), .C2(n13399), .A(n11689), .B(n11688), .ZN(
        n11693) );
  NAND2_X1 U14046 ( .A1(n11690), .A2(n11691), .ZN(n13400) );
  NAND3_X1 U14047 ( .A1(n13401), .A2(n13400), .A3(n14510), .ZN(n11692) );
  OAI211_X1 U14048 ( .C1(n11694), .C2(n13305), .A(n11693), .B(n11692), .ZN(
        P2_U3249) );
  NAND2_X1 U14049 ( .A1(n11695), .A2(n13756), .ZN(n11697) );
  AOI22_X1 U14050 ( .A1(n13728), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6459), 
        .B2(n13912), .ZN(n11696) );
  XNOR2_X1 U14051 ( .A(n14575), .B(n13833), .ZN(n13796) );
  NAND2_X1 U14052 ( .A1(n11698), .A2(n13672), .ZN(n11699) );
  AOI21_X1 U14053 ( .B1(n11702), .B2(n11699), .A(n12037), .ZN(n14586) );
  OAI21_X1 U14054 ( .B1(n11703), .B2(n11702), .A(n12007), .ZN(n14589) );
  INV_X1 U14055 ( .A(n14581), .ZN(n11713) );
  OR2_X1 U14056 ( .A1(n11704), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11705) );
  NAND2_X1 U14057 ( .A1(n11830), .A2(n11705), .ZN(n13512) );
  AOI22_X1 U14058 ( .A1(n6456), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n13730), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n11707) );
  NAND2_X1 U14059 ( .A1(n11930), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11706) );
  OAI211_X1 U14060 ( .C1(n13512), .C2(n11851), .A(n11707), .B(n11706), .ZN(
        n13832) );
  NAND2_X1 U14061 ( .A1(n13832), .A2(n14645), .ZN(n11709) );
  NAND2_X1 U14062 ( .A1(n13834), .A2(n13551), .ZN(n11708) );
  NAND2_X1 U14063 ( .A1(n11709), .A2(n11708), .ZN(n14582) );
  INV_X1 U14064 ( .A(n11710), .ZN(n11711) );
  INV_X1 U14065 ( .A(n14575), .ZN(n14585) );
  OAI211_X1 U14066 ( .C1(n11711), .C2(n14585), .A(n14730), .B(n14153), .ZN(
        n14584) );
  NOR2_X1 U14067 ( .A1(n14584), .A2(n13568), .ZN(n11712) );
  AOI211_X1 U14068 ( .C1(n14728), .C2(n11713), .A(n14582), .B(n11712), .ZN(
        n11715) );
  AOI22_X1 U14069 ( .A1(n14575), .A2(n14735), .B1(n14697), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n11714) );
  OAI21_X1 U14070 ( .B1(n11715), .B2(n14697), .A(n11714), .ZN(n11716) );
  AOI21_X1 U14071 ( .B1(n14589), .B2(n14124), .A(n11716), .ZN(n11717) );
  OAI21_X1 U14072 ( .B1(n14586), .B2(n14126), .A(n11717), .ZN(P1_U3277) );
  NAND2_X1 U14073 ( .A1(n14564), .A2(n12222), .ZN(n11723) );
  NAND2_X1 U14074 ( .A1(n13837), .A2(n11834), .ZN(n11722) );
  NAND2_X1 U14075 ( .A1(n11723), .A2(n11722), .ZN(n11724) );
  XNOR2_X1 U14076 ( .A(n11724), .B(n10393), .ZN(n11727) );
  AOI22_X1 U14077 ( .A1(n14564), .A2(n11966), .B1(n12223), .B2(n13837), .ZN(
        n11725) );
  XNOR2_X1 U14078 ( .A(n11727), .B(n11725), .ZN(n14562) );
  INV_X1 U14079 ( .A(n11725), .ZN(n11726) );
  NOR2_X1 U14080 ( .A1(n11727), .A2(n11726), .ZN(n11728) );
  NAND2_X1 U14081 ( .A1(n13661), .A2(n12222), .ZN(n11730) );
  NAND2_X1 U14082 ( .A1(n13836), .A2(n11834), .ZN(n11729) );
  NAND2_X1 U14083 ( .A1(n11730), .A2(n11729), .ZN(n11731) );
  XNOR2_X1 U14084 ( .A(n11731), .B(n10393), .ZN(n11793) );
  NOR2_X1 U14085 ( .A1(n11732), .A2(n11803), .ZN(n11733) );
  AOI21_X1 U14086 ( .B1(n13661), .B2(n11966), .A(n11733), .ZN(n11794) );
  XNOR2_X1 U14087 ( .A(n11793), .B(n11794), .ZN(n11734) );
  OAI211_X1 U14088 ( .C1(n11735), .C2(n11734), .A(n14552), .B(n14576), .ZN(
        n11740) );
  OAI21_X1 U14089 ( .B1(n14649), .B2(n14248), .A(n11736), .ZN(n11737) );
  AOI21_X1 U14090 ( .B1(n11738), .B2(n13563), .A(n11737), .ZN(n11739) );
  OAI211_X1 U14091 ( .C1(n6857), .C2(n13567), .A(n11740), .B(n11739), .ZN(
        P1_U3234) );
  XNOR2_X1 U14092 ( .A(n6568), .B(n11741), .ZN(n13387) );
  INV_X1 U14093 ( .A(n13387), .ZN(n11753) );
  XNOR2_X1 U14094 ( .A(n11742), .B(n11741), .ZN(n13388) );
  NAND2_X1 U14095 ( .A1(n11743), .A2(n13439), .ZN(n11744) );
  NAND2_X1 U14096 ( .A1(n11744), .A2(n6452), .ZN(n11745) );
  OR2_X1 U14097 ( .A1(n13292), .A2(n11745), .ZN(n13390) );
  NAND2_X1 U14098 ( .A1(n13034), .A2(n13013), .ZN(n11747) );
  NAND2_X1 U14099 ( .A1(n13036), .A2(n14484), .ZN(n11746) );
  AND2_X1 U14100 ( .A1(n11747), .A2(n11746), .ZN(n13389) );
  NOR2_X1 U14101 ( .A1(n13389), .A2(n14951), .ZN(n11749) );
  INV_X1 U14102 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13090) );
  OAI22_X1 U14103 ( .A1(n14948), .A2(n13090), .B1(n12959), .B2(n13295), .ZN(
        n11748) );
  AOI211_X1 U14104 ( .C1(n13439), .C2(n14502), .A(n11749), .B(n11748), .ZN(
        n11750) );
  OAI21_X1 U14105 ( .B1(n13390), .B2(n13302), .A(n11750), .ZN(n11751) );
  AOI21_X1 U14106 ( .B1(n13388), .B2(n13212), .A(n11751), .ZN(n11752) );
  OAI21_X1 U14107 ( .B1(n11753), .B2(n13224), .A(n11752), .ZN(P2_U3248) );
  INV_X1 U14108 ( .A(n11754), .ZN(n11756) );
  XNOR2_X1 U14109 ( .A(n14503), .B(n12873), .ZN(n11760) );
  NAND2_X1 U14110 ( .A1(n13037), .A2(n12834), .ZN(n11759) );
  NAND2_X1 U14111 ( .A1(n11760), .A2(n11759), .ZN(n12836) );
  OAI21_X1 U14112 ( .B1(n11760), .B2(n11759), .A(n12836), .ZN(n14487) );
  INV_X1 U14113 ( .A(n12836), .ZN(n11761) );
  NOR2_X1 U14114 ( .A1(n14485), .A2(n11761), .ZN(n11763) );
  XNOR2_X1 U14115 ( .A(n11767), .B(n12915), .ZN(n12838) );
  AND2_X1 U14116 ( .A1(n14482), .A2(n13217), .ZN(n12837) );
  INV_X1 U14117 ( .A(n12837), .ZN(n12839) );
  XNOR2_X1 U14118 ( .A(n12838), .B(n12839), .ZN(n11762) );
  XNOR2_X1 U14119 ( .A(n11763), .B(n11762), .ZN(n11769) );
  NOR2_X1 U14120 ( .A1(n14495), .A2(n11764), .ZN(n11766) );
  OAI22_X1 U14121 ( .A1(n14514), .A2(n14491), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7733), .ZN(n11765) );
  AOI211_X1 U14122 ( .C1(n11767), .C2(n13014), .A(n11766), .B(n11765), .ZN(
        n11768) );
  OAI21_X1 U14123 ( .B1(n11769), .B2(n14490), .A(n11768), .ZN(P2_U3213) );
  INV_X1 U14124 ( .A(n12034), .ZN(n13449) );
  OAI222_X1 U14125 ( .A1(n6454), .A2(n11771), .B1(n14286), .B2(n13449), .C1(
        n11770), .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U14126 ( .A(n12021), .ZN(n13453) );
  OAI222_X1 U14127 ( .A1(n6454), .A2(n11773), .B1(n14286), .B2(n13453), .C1(
        P1_U3086), .C2(n11772), .ZN(P1_U3327) );
  INV_X1 U14128 ( .A(n11775), .ZN(n13456) );
  OAI222_X1 U14129 ( .A1(n6454), .A2(n11774), .B1(n14286), .B2(n13456), .C1(
        n6455), .C2(P1_U3086), .ZN(P1_U3328) );
  NAND2_X1 U14130 ( .A1(n13728), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11776) );
  NAND2_X1 U14131 ( .A1(n13998), .A2(n12222), .ZN(n11784) );
  NAND2_X1 U14132 ( .A1(n12051), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11782) );
  NAND2_X1 U14133 ( .A1(n11930), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11781) );
  INV_X1 U14134 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11981) );
  INV_X1 U14135 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11829) );
  INV_X1 U14136 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13485) );
  INV_X1 U14137 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13494) );
  NAND2_X1 U14138 ( .A1(n11896), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11915) );
  NAND2_X1 U14139 ( .A1(n11943), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11778) );
  INV_X1 U14140 ( .A(n11778), .ZN(n11959) );
  NAND2_X1 U14141 ( .A1(n11959), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11974) );
  INV_X1 U14142 ( .A(n11974), .ZN(n12026) );
  AOI21_X1 U14143 ( .B1(n11981), .B2(n11778), .A(n12026), .ZN(n13999) );
  NAND2_X1 U14144 ( .A1(n12027), .A2(n13999), .ZN(n11780) );
  NAND2_X1 U14145 ( .A1(n6456), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11779) );
  NAND4_X1 U14146 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n13822) );
  NAND2_X1 U14147 ( .A1(n13822), .A2(n11834), .ZN(n11783) );
  NAND2_X1 U14148 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  XNOR2_X1 U14149 ( .A(n11785), .B(n10393), .ZN(n12218) );
  AOI22_X1 U14150 ( .A1(n13998), .A2(n9910), .B1(n12223), .B2(n13822), .ZN(
        n12219) );
  XNOR2_X1 U14151 ( .A(n12218), .B(n12219), .ZN(n12221) );
  NAND2_X1 U14152 ( .A1(n14600), .A2(n12222), .ZN(n11787) );
  NAND2_X1 U14153 ( .A1(n13835), .A2(n11834), .ZN(n11786) );
  NAND2_X1 U14154 ( .A1(n11787), .A2(n11786), .ZN(n11788) );
  XNOR2_X1 U14155 ( .A(n11788), .B(n11810), .ZN(n11792) );
  INV_X1 U14156 ( .A(n11792), .ZN(n11798) );
  NOR2_X1 U14157 ( .A1(n11789), .A2(n11803), .ZN(n11790) );
  AOI21_X1 U14158 ( .B1(n14600), .B2(n11966), .A(n11790), .ZN(n11791) );
  INV_X1 U14159 ( .A(n11791), .ZN(n11797) );
  XNOR2_X1 U14160 ( .A(n11792), .B(n11791), .ZN(n14553) );
  INV_X1 U14161 ( .A(n11793), .ZN(n11795) );
  NOR2_X1 U14162 ( .A1(n11795), .A2(n11794), .ZN(n14554) );
  NOR2_X1 U14163 ( .A1(n14553), .A2(n14554), .ZN(n11796) );
  NAND2_X1 U14164 ( .A1(n14552), .A2(n11796), .ZN(n14556) );
  OAI21_X1 U14165 ( .B1(n11798), .B2(n11797), .A(n14556), .ZN(n11805) );
  NAND2_X1 U14166 ( .A1(n11799), .A2(n12222), .ZN(n11801) );
  NAND2_X1 U14167 ( .A1(n13834), .A2(n11966), .ZN(n11800) );
  NAND2_X1 U14168 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  XNOR2_X1 U14169 ( .A(n11802), .B(n10393), .ZN(n11806) );
  XNOR2_X1 U14170 ( .A(n11805), .B(n11806), .ZN(n13561) );
  OAI22_X1 U14171 ( .A1(n14594), .A2(n11904), .B1(n11804), .B2(n11803), .ZN(
        n13560) );
  NAND2_X1 U14172 ( .A1(n13561), .A2(n13560), .ZN(n13559) );
  INV_X1 U14173 ( .A(n11805), .ZN(n11807) );
  NAND2_X1 U14174 ( .A1(n14575), .A2(n12222), .ZN(n11809) );
  NAND2_X1 U14175 ( .A1(n13833), .A2(n11966), .ZN(n11808) );
  NAND2_X1 U14176 ( .A1(n11809), .A2(n11808), .ZN(n11811) );
  XNOR2_X1 U14177 ( .A(n11811), .B(n11810), .ZN(n11814) );
  AOI22_X1 U14178 ( .A1(n14575), .A2(n11966), .B1(n12223), .B2(n13833), .ZN(
        n11813) );
  XNOR2_X1 U14179 ( .A(n11814), .B(n11813), .ZN(n14570) );
  NAND2_X1 U14180 ( .A1(n13559), .A2(n11812), .ZN(n14573) );
  NAND2_X1 U14181 ( .A1(n11814), .A2(n11813), .ZN(n11815) );
  NAND2_X1 U14182 ( .A1(n14573), .A2(n11815), .ZN(n13509) );
  NAND2_X1 U14183 ( .A1(n11816), .A2(n13756), .ZN(n11818) );
  AOI22_X1 U14184 ( .A1(n13728), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6459), 
        .B2(n13936), .ZN(n11817) );
  NAND2_X1 U14185 ( .A1(n14243), .A2(n12222), .ZN(n11820) );
  NAND2_X1 U14186 ( .A1(n13832), .A2(n11834), .ZN(n11819) );
  NAND2_X1 U14187 ( .A1(n11820), .A2(n11819), .ZN(n11821) );
  XNOR2_X1 U14188 ( .A(n11821), .B(n10393), .ZN(n11822) );
  AOI22_X1 U14189 ( .A1(n14243), .A2(n11966), .B1(n12223), .B2(n13832), .ZN(
        n11823) );
  XNOR2_X1 U14190 ( .A(n11822), .B(n11823), .ZN(n13510) );
  INV_X1 U14191 ( .A(n11822), .ZN(n11824) );
  NAND2_X1 U14192 ( .A1(n11824), .A2(n11823), .ZN(n11825) );
  NAND2_X1 U14193 ( .A1(n11826), .A2(n13756), .ZN(n11828) );
  AOI22_X1 U14194 ( .A1(n13728), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6459), 
        .B2(n13951), .ZN(n11827) );
  NAND2_X1 U14195 ( .A1(n14238), .A2(n12222), .ZN(n11836) );
  INV_X1 U14196 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n13938) );
  NAND2_X1 U14197 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  NAND2_X1 U14198 ( .A1(n11845), .A2(n11831), .ZN(n14135) );
  OR2_X1 U14199 ( .A1(n14135), .A2(n11851), .ZN(n11833) );
  AOI22_X1 U14200 ( .A1(n6456), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n12051), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n11832) );
  OAI211_X1 U14201 ( .C1(n11109), .C2(n13938), .A(n11833), .B(n11832), .ZN(
        n13831) );
  NAND2_X1 U14202 ( .A1(n13831), .A2(n11834), .ZN(n11835) );
  NAND2_X1 U14203 ( .A1(n11836), .A2(n11835), .ZN(n11837) );
  XNOR2_X1 U14204 ( .A(n11837), .B(n10393), .ZN(n11838) );
  AOI22_X1 U14205 ( .A1(n14238), .A2(n9910), .B1(n12223), .B2(n13831), .ZN(
        n11839) );
  XNOR2_X1 U14206 ( .A(n11838), .B(n11839), .ZN(n13540) );
  INV_X1 U14207 ( .A(n11838), .ZN(n11840) );
  NAND2_X1 U14208 ( .A1(n11841), .A2(n13756), .ZN(n11844) );
  AOI22_X1 U14209 ( .A1(n13728), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6459), 
        .B2(n13568), .ZN(n11843) );
  AND2_X1 U14210 ( .A1(n11845), .A2(n13485), .ZN(n11846) );
  OR2_X1 U14211 ( .A1(n11864), .A2(n11846), .ZN(n14117) );
  INV_X1 U14212 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13948) );
  NAND2_X1 U14213 ( .A1(n6456), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11848) );
  NAND2_X1 U14214 ( .A1(n13730), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11847) );
  OAI211_X1 U14215 ( .C1(n13948), .C2(n11109), .A(n11848), .B(n11847), .ZN(
        n11849) );
  INV_X1 U14216 ( .A(n11849), .ZN(n11850) );
  OAI21_X1 U14217 ( .B1(n14117), .B2(n11851), .A(n11850), .ZN(n13830) );
  AND2_X1 U14218 ( .A1(n13830), .A2(n12223), .ZN(n11852) );
  AOI21_X1 U14219 ( .B1(n14233), .B2(n9910), .A(n11852), .ZN(n11857) );
  NAND2_X1 U14220 ( .A1(n14233), .A2(n12222), .ZN(n11854) );
  NAND2_X1 U14221 ( .A1(n13830), .A2(n11966), .ZN(n11853) );
  NAND2_X1 U14222 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  XNOR2_X1 U14223 ( .A(n11855), .B(n10393), .ZN(n11859) );
  XOR2_X1 U14224 ( .A(n11857), .B(n11859), .Z(n13479) );
  INV_X1 U14225 ( .A(n11857), .ZN(n11858) );
  NAND2_X1 U14226 ( .A1(n11859), .A2(n11858), .ZN(n11860) );
  NAND2_X1 U14227 ( .A1(n13481), .A2(n11860), .ZN(n13525) );
  NAND2_X1 U14228 ( .A1(n11861), .A2(n13756), .ZN(n11863) );
  NAND2_X1 U14229 ( .A1(n13728), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n11862) );
  OR2_X1 U14230 ( .A1(n11864), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U14231 ( .A1(n11865), .A2(n11883), .ZN(n13526) );
  OR2_X1 U14232 ( .A1(n13526), .A2(n11851), .ZN(n11872) );
  INV_X1 U14233 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U14234 ( .A1(n11930), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11868) );
  NAND2_X1 U14235 ( .A1(n12051), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11867) );
  OAI211_X1 U14236 ( .C1(n10611), .C2(n11869), .A(n11868), .B(n11867), .ZN(
        n11870) );
  INV_X1 U14237 ( .A(n11870), .ZN(n11871) );
  NAND2_X1 U14238 ( .A1(n11872), .A2(n11871), .ZN(n13829) );
  AND2_X1 U14239 ( .A1(n13829), .A2(n12223), .ZN(n11873) );
  AOI21_X1 U14240 ( .B1(n14105), .B2(n11966), .A(n11873), .ZN(n11876) );
  AOI22_X1 U14241 ( .A1(n14105), .A2(n12222), .B1(n9910), .B2(n13829), .ZN(
        n11874) );
  XNOR2_X1 U14242 ( .A(n11874), .B(n10393), .ZN(n11875) );
  XOR2_X1 U14243 ( .A(n11876), .B(n11875), .Z(n13524) );
  INV_X1 U14244 ( .A(n11875), .ZN(n11878) );
  INV_X1 U14245 ( .A(n11876), .ZN(n11877) );
  NAND2_X1 U14246 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  NAND2_X1 U14247 ( .A1(n11880), .A2(n13756), .ZN(n11882) );
  NAND2_X1 U14248 ( .A1(n13728), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n11881) );
  NAND2_X1 U14249 ( .A1(n12051), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11887) );
  NAND2_X1 U14250 ( .A1(n11930), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11886) );
  AOI21_X1 U14251 ( .B1(n13494), .B2(n11883), .A(n11896), .ZN(n14087) );
  NAND2_X1 U14252 ( .A1(n12027), .A2(n14087), .ZN(n11885) );
  NAND2_X1 U14253 ( .A1(n6456), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11884) );
  NAND4_X1 U14254 ( .A1(n11887), .A2(n11886), .A3(n11885), .A4(n11884), .ZN(
        n13828) );
  AOI22_X1 U14255 ( .A1(n14090), .A2(n12222), .B1(n9910), .B2(n13828), .ZN(
        n11888) );
  XNOR2_X1 U14256 ( .A(n11888), .B(n10393), .ZN(n11891) );
  AOI22_X1 U14257 ( .A1(n14090), .A2(n11966), .B1(n12223), .B2(n13828), .ZN(
        n11890) );
  XNOR2_X1 U14258 ( .A(n11891), .B(n11890), .ZN(n13492) );
  INV_X1 U14259 ( .A(n13492), .ZN(n11889) );
  NAND2_X1 U14260 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  OR2_X1 U14261 ( .A1(n11893), .A2(n9139), .ZN(n11894) );
  XNOR2_X1 U14262 ( .A(n11894), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14288) );
  NAND2_X1 U14263 ( .A1(n12051), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11902) );
  NAND2_X1 U14264 ( .A1(n11930), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11901) );
  INV_X1 U14265 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13536) );
  INV_X1 U14266 ( .A(n11896), .ZN(n11898) );
  AOI21_X1 U14267 ( .B1(n13536), .B2(n11898), .A(n11897), .ZN(n14077) );
  NAND2_X1 U14268 ( .A1(n12027), .A2(n14077), .ZN(n11900) );
  NAND2_X1 U14269 ( .A1(n6456), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11899) );
  NAND4_X1 U14270 ( .A1(n11902), .A2(n11901), .A3(n11900), .A4(n11899), .ZN(
        n13827) );
  AOI22_X1 U14271 ( .A1(n14212), .A2(n12222), .B1(n9910), .B2(n13827), .ZN(
        n11903) );
  XNOR2_X1 U14272 ( .A(n11903), .B(n10393), .ZN(n11909) );
  OR2_X1 U14273 ( .A1(n14080), .A2(n11904), .ZN(n11906) );
  NAND2_X1 U14274 ( .A1(n12223), .A2(n13827), .ZN(n11905) );
  NAND2_X1 U14275 ( .A1(n11906), .A2(n11905), .ZN(n11907) );
  XNOR2_X1 U14276 ( .A(n11909), .B(n11907), .ZN(n13534) );
  INV_X1 U14277 ( .A(n11907), .ZN(n11908) );
  NAND2_X1 U14278 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  NAND2_X1 U14279 ( .A1(n11911), .A2(n13756), .ZN(n11913) );
  NAND2_X1 U14280 ( .A1(n13728), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U14281 ( .A1(n14059), .A2(n12222), .ZN(n11921) );
  NAND2_X1 U14282 ( .A1(n12051), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11919) );
  NAND2_X1 U14283 ( .A1(n6456), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11918) );
  INV_X1 U14284 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13474) );
  AOI21_X1 U14285 ( .B1(n13474), .B2(n11915), .A(n11914), .ZN(n14060) );
  NAND2_X1 U14286 ( .A1(n12027), .A2(n14060), .ZN(n11917) );
  NAND2_X1 U14287 ( .A1(n11930), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11916) );
  NAND4_X1 U14288 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n13826) );
  NAND2_X1 U14289 ( .A1(n13826), .A2(n11966), .ZN(n11920) );
  NAND2_X1 U14290 ( .A1(n11921), .A2(n11920), .ZN(n11922) );
  XNOR2_X1 U14291 ( .A(n11922), .B(n10393), .ZN(n11923) );
  AOI22_X1 U14292 ( .A1(n14059), .A2(n11966), .B1(n12223), .B2(n13826), .ZN(
        n11924) );
  XNOR2_X1 U14293 ( .A(n11923), .B(n11924), .ZN(n13471) );
  INV_X1 U14294 ( .A(n11923), .ZN(n11925) );
  NAND2_X1 U14295 ( .A1(n13728), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11926) );
  NAND2_X1 U14296 ( .A1(n14200), .A2(n12222), .ZN(n11936) );
  NAND2_X1 U14297 ( .A1(n6456), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11934) );
  NAND2_X1 U14298 ( .A1(n13730), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11933) );
  INV_X1 U14299 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13518) );
  AOI21_X1 U14300 ( .B1(n13518), .B2(n11929), .A(n11928), .ZN(n14046) );
  NAND2_X1 U14301 ( .A1(n12027), .A2(n14046), .ZN(n11932) );
  NAND2_X1 U14302 ( .A1(n11930), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11931) );
  NAND4_X1 U14303 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n13825) );
  NAND2_X1 U14304 ( .A1(n13825), .A2(n11966), .ZN(n11935) );
  NAND2_X1 U14305 ( .A1(n11936), .A2(n11935), .ZN(n11937) );
  XNOR2_X1 U14306 ( .A(n11937), .B(n10393), .ZN(n11938) );
  AOI22_X1 U14307 ( .A1(n14200), .A2(n11834), .B1(n12223), .B2(n13825), .ZN(
        n11939) );
  XNOR2_X1 U14308 ( .A(n11938), .B(n11939), .ZN(n13517) );
  INV_X1 U14309 ( .A(n11938), .ZN(n11940) );
  NAND2_X1 U14310 ( .A1(n13462), .A2(n13756), .ZN(n11942) );
  NAND2_X1 U14311 ( .A1(n13728), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U14312 ( .A1(n6693), .A2(n12222), .ZN(n11950) );
  NAND2_X1 U14313 ( .A1(n6456), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U14314 ( .A1(n12051), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11947) );
  INV_X1 U14315 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13503) );
  AOI21_X1 U14316 ( .B1(n13503), .B2(n11944), .A(n11943), .ZN(n14026) );
  NAND2_X1 U14317 ( .A1(n12027), .A2(n14026), .ZN(n11946) );
  NAND2_X1 U14318 ( .A1(n11930), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11945) );
  NAND4_X1 U14319 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n13824) );
  NAND2_X1 U14320 ( .A1(n13824), .A2(n11966), .ZN(n11949) );
  NAND2_X1 U14321 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  XNOR2_X1 U14322 ( .A(n11951), .B(n10393), .ZN(n11952) );
  AOI22_X1 U14323 ( .A1(n6693), .A2(n11966), .B1(n12223), .B2(n13824), .ZN(
        n11953) );
  XNOR2_X1 U14324 ( .A(n11952), .B(n11953), .ZN(n13500) );
  NAND2_X1 U14325 ( .A1(n13499), .A2(n13500), .ZN(n11956) );
  INV_X1 U14326 ( .A(n11952), .ZN(n11954) );
  NAND2_X1 U14327 ( .A1(n11954), .A2(n11953), .ZN(n11955) );
  NAND2_X1 U14328 ( .A1(n13728), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11957) );
  NAND2_X1 U14329 ( .A1(n13717), .A2(n12222), .ZN(n11968) );
  NAND2_X1 U14330 ( .A1(n12051), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11965) );
  NAND2_X1 U14331 ( .A1(n11930), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11964) );
  INV_X1 U14332 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13554) );
  AOI21_X1 U14333 ( .B1(n13554), .B2(n11960), .A(n11959), .ZN(n14014) );
  NAND2_X1 U14334 ( .A1(n12027), .A2(n14014), .ZN(n11963) );
  NAND2_X1 U14335 ( .A1(n6456), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11962) );
  NAND2_X1 U14336 ( .A1(n13823), .A2(n11966), .ZN(n11967) );
  NAND2_X1 U14337 ( .A1(n11968), .A2(n11967), .ZN(n11969) );
  XNOR2_X1 U14338 ( .A(n11969), .B(n10393), .ZN(n11970) );
  AOI22_X1 U14339 ( .A1(n13717), .A2(n11966), .B1(n12223), .B2(n13823), .ZN(
        n11971) );
  XNOR2_X1 U14340 ( .A(n11970), .B(n11971), .ZN(n13550) );
  INV_X1 U14341 ( .A(n11970), .ZN(n11972) );
  NAND2_X1 U14342 ( .A1(n11972), .A2(n11971), .ZN(n11973) );
  NAND2_X1 U14343 ( .A1(n13823), .A2(n13551), .ZN(n11980) );
  NAND2_X1 U14344 ( .A1(n6456), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U14345 ( .A1(n12051), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11977) );
  XNOR2_X1 U14346 ( .A(P1_REG3_REG_28__SCAN_IN), .B(n11974), .ZN(n13989) );
  NAND2_X1 U14347 ( .A1(n12027), .A2(n13989), .ZN(n11976) );
  NAND2_X1 U14348 ( .A1(n11930), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U14349 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n13821) );
  NAND2_X1 U14350 ( .A1(n13821), .A2(n14645), .ZN(n11979) );
  AND2_X1 U14351 ( .A1(n11980), .A2(n11979), .ZN(n14178) );
  OAI22_X1 U14352 ( .A1(n14649), .A2(n14178), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11981), .ZN(n11982) );
  AOI21_X1 U14353 ( .B1(n13999), .B2(n13563), .A(n11982), .ZN(n11984) );
  NAND2_X1 U14354 ( .A1(n13998), .A2(n14657), .ZN(n11983) );
  OAI211_X1 U14355 ( .C1(n11985), .C2(n14651), .A(n11984), .B(n11983), .ZN(
        P1_U3214) );
  NAND2_X1 U14356 ( .A1(n13021), .A2(n11987), .ZN(n13307) );
  NAND2_X1 U14357 ( .A1(n13141), .A2(n13307), .ZN(n12216) );
  XNOR2_X1 U14358 ( .A(n11990), .B(n11989), .ZN(n11995) );
  NAND2_X1 U14359 ( .A1(n12352), .A2(n12369), .ZN(n11991) );
  NAND2_X1 U14360 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14452)
         );
  OAI211_X1 U14361 ( .C1(n12681), .C2(n12354), .A(n11991), .B(n14452), .ZN(
        n11993) );
  NOR2_X1 U14362 ( .A1(n12813), .A2(n12360), .ZN(n11992) );
  AOI211_X1 U14363 ( .C1(n12686), .C2(n12356), .A(n11993), .B(n11992), .ZN(
        n11994) );
  OAI21_X1 U14364 ( .B1(n11995), .B2(n12347), .A(n11994), .ZN(P3_U3168) );
  INV_X1 U14365 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11996) );
  MUX2_X1 U14366 ( .A(n11998), .B(n11996), .S(n15127), .Z(n11997) );
  OAI21_X1 U14367 ( .B1(n12001), .B2(n12818), .A(n11997), .ZN(P3_U3390) );
  MUX2_X1 U14368 ( .A(n11999), .B(n11998), .S(n15133), .Z(n12000) );
  OAI21_X1 U14369 ( .B1(n12001), .B2(n12755), .A(n12000), .ZN(P3_U3459) );
  INV_X1 U14370 ( .A(n12002), .ZN(n12004) );
  OAI222_X1 U14371 ( .A1(n12829), .A2(n12005), .B1(n12832), .B2(n12004), .C1(
        P3_U3151), .C2(n12003), .ZN(P3_U3266) );
  INV_X1 U14372 ( .A(n13832), .ZN(n13543) );
  NAND2_X1 U14373 ( .A1(n14243), .A2(n13543), .ZN(n13683) );
  INV_X1 U14374 ( .A(n13831), .ZN(n12009) );
  NAND2_X1 U14375 ( .A1(n14238), .A2(n12009), .ZN(n12008) );
  INV_X1 U14376 ( .A(n14238), .ZN(n14138) );
  NAND2_X1 U14377 ( .A1(n14138), .A2(n12009), .ZN(n12010) );
  INV_X1 U14378 ( .A(n13830), .ZN(n13577) );
  INV_X1 U14379 ( .A(n13829), .ZN(n12012) );
  XNOR2_X1 U14380 ( .A(n14105), .B(n12012), .ZN(n13800) );
  INV_X1 U14381 ( .A(n13828), .ZN(n13693) );
  NOR2_X1 U14382 ( .A1(n14090), .A2(n13828), .ZN(n12013) );
  INV_X1 U14383 ( .A(n13827), .ZN(n12014) );
  NAND2_X1 U14384 ( .A1(n14212), .A2(n12014), .ZN(n13699) );
  NAND2_X1 U14385 ( .A1(n14080), .A2(n12014), .ZN(n12015) );
  XNOR2_X2 U14386 ( .A(n14200), .B(n13825), .ZN(n14038) );
  NAND2_X1 U14387 ( .A1(n14059), .A2(n13826), .ZN(n14035) );
  NAND2_X1 U14388 ( .A1(n6693), .A2(n13824), .ZN(n12017) );
  INV_X1 U14389 ( .A(n13823), .ZN(n12018) );
  NAND2_X1 U14390 ( .A1(n14009), .A2(n14008), .ZN(n12020) );
  NAND2_X1 U14391 ( .A1(n13717), .A2(n13823), .ZN(n12019) );
  NAND2_X1 U14392 ( .A1(n13728), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12022) );
  INV_X1 U14393 ( .A(n13821), .ZN(n12024) );
  NAND2_X1 U14394 ( .A1(n14174), .A2(n12024), .ZN(n12043) );
  AND2_X1 U14395 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n12026), .ZN(n12055) );
  NAND2_X1 U14396 ( .A1(n12027), .A2(n12055), .ZN(n12033) );
  NAND2_X1 U14397 ( .A1(n11930), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12032) );
  INV_X1 U14398 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n12028) );
  OR2_X1 U14399 ( .A1(n10611), .A2(n12028), .ZN(n12031) );
  INV_X1 U14400 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n12029) );
  OR2_X1 U14401 ( .A1(n10532), .A2(n12029), .ZN(n12030) );
  XNOR2_X1 U14402 ( .A(n12035), .B(n13804), .ZN(n14165) );
  NAND2_X1 U14403 ( .A1(n14165), .A2(n14124), .ZN(n12066) );
  INV_X1 U14404 ( .A(n13825), .ZN(n13574) );
  INV_X1 U14405 ( .A(n13833), .ZN(n13677) );
  NOR2_X1 U14406 ( .A1(n14109), .A2(n12040), .ZN(n14095) );
  OAI22_X1 U14407 ( .A1(n14084), .A2(n14085), .B1(n13693), .B2(n14090), .ZN(
        n14067) );
  INV_X1 U14408 ( .A(n13826), .ZN(n12041) );
  INV_X1 U14409 ( .A(n14029), .ZN(n14193) );
  INV_X1 U14410 ( .A(n14008), .ZN(n14011) );
  INV_X1 U14411 ( .A(n13804), .ZN(n12044) );
  INV_X1 U14412 ( .A(n14090), .ZN(n14218) );
  NAND2_X1 U14413 ( .A1(n14099), .A2(n14218), .ZN(n14086) );
  NOR2_X2 U14414 ( .A1(n14075), .A2(n14059), .ZN(n14043) );
  AOI21_X1 U14415 ( .B1(n13742), .B2(n13987), .A(n13974), .ZN(n14171) );
  INV_X1 U14416 ( .A(P1_B_REG_SCAN_IN), .ZN(n12048) );
  NOR2_X1 U14417 ( .A1(n6455), .A2(n12048), .ZN(n12049) );
  NOR2_X1 U14418 ( .A1(n13544), .A2(n12049), .ZN(n13969) );
  NAND2_X1 U14419 ( .A1(n12050), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12054) );
  NAND2_X1 U14420 ( .A1(n6456), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12053) );
  NAND2_X1 U14421 ( .A1(n12051), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12052) );
  NAND3_X1 U14422 ( .A1(n12054), .A2(n12053), .A3(n12052), .ZN(n13819) );
  NAND2_X1 U14423 ( .A1(n13969), .A2(n13819), .ZN(n14167) );
  NAND2_X1 U14424 ( .A1(n14728), .A2(n12055), .ZN(n12056) );
  OAI21_X1 U14425 ( .B1(n12057), .B2(n14167), .A(n12056), .ZN(n12059) );
  NAND2_X1 U14426 ( .A1(n13821), .A2(n13551), .ZN(n14168) );
  NOR2_X1 U14427 ( .A1(n14697), .A2(n14168), .ZN(n12058) );
  AOI211_X1 U14428 ( .C1(n14697), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12059), 
        .B(n12058), .ZN(n12060) );
  OAI21_X1 U14429 ( .B1(n14169), .B2(n14712), .A(n12060), .ZN(n12061) );
  AOI21_X1 U14430 ( .B1(n14171), .B2(n12062), .A(n12061), .ZN(n12063) );
  NAND2_X1 U14431 ( .A1(n12066), .A2(n12065), .ZN(n12213) );
  NOR3_X1 U14432 ( .A1(keyinput26), .A2(keyinput41), .A3(keyinput58), .ZN(
        n12079) );
  NAND2_X1 U14433 ( .A1(keyinput15), .A2(keyinput27), .ZN(n12070) );
  NOR4_X1 U14434 ( .A1(keyinput59), .A2(keyinput18), .A3(keyinput44), .A4(
        keyinput0), .ZN(n12068) );
  NOR2_X1 U14435 ( .A1(keyinput7), .A2(keyinput16), .ZN(n12067) );
  NAND4_X1 U14436 ( .A1(n12068), .A2(keyinput11), .A3(keyinput45), .A4(n12067), 
        .ZN(n12069) );
  NOR4_X1 U14437 ( .A1(keyinput8), .A2(keyinput34), .A3(n12070), .A4(n12069), 
        .ZN(n12078) );
  NAND2_X1 U14438 ( .A1(keyinput6), .A2(keyinput13), .ZN(n12076) );
  NOR2_X1 U14439 ( .A1(keyinput55), .A2(keyinput24), .ZN(n12074) );
  NAND3_X1 U14440 ( .A1(keyinput57), .A2(keyinput21), .A3(keyinput33), .ZN(
        n12072) );
  NAND3_X1 U14441 ( .A1(keyinput61), .A2(keyinput40), .A3(keyinput35), .ZN(
        n12071) );
  NOR4_X1 U14442 ( .A1(keyinput29), .A2(keyinput17), .A3(n12072), .A4(n12071), 
        .ZN(n12073) );
  NAND4_X1 U14443 ( .A1(keyinput48), .A2(keyinput49), .A3(n12074), .A4(n12073), 
        .ZN(n12075) );
  NOR4_X1 U14444 ( .A1(keyinput53), .A2(keyinput51), .A3(n12076), .A4(n12075), 
        .ZN(n12077) );
  NAND4_X1 U14445 ( .A1(keyinput63), .A2(n12079), .A3(n12078), .A4(n12077), 
        .ZN(n12211) );
  NAND3_X1 U14446 ( .A1(keyinput39), .A2(keyinput32), .A3(keyinput23), .ZN(
        n12081) );
  NAND3_X1 U14447 ( .A1(keyinput60), .A2(keyinput42), .A3(keyinput46), .ZN(
        n12080) );
  OR4_X1 U14448 ( .A1(n12081), .A2(n12080), .A3(keyinput19), .A4(keyinput2), 
        .ZN(n12093) );
  NOR3_X1 U14449 ( .A1(keyinput52), .A2(keyinput20), .A3(keyinput38), .ZN(
        n12086) );
  NAND2_X1 U14450 ( .A1(keyinput36), .A2(keyinput25), .ZN(n12082) );
  NOR3_X1 U14451 ( .A1(keyinput14), .A2(keyinput54), .A3(n12082), .ZN(n12085)
         );
  NAND2_X1 U14452 ( .A1(keyinput28), .A2(keyinput1), .ZN(n12083) );
  NOR3_X1 U14453 ( .A1(keyinput56), .A2(keyinput43), .A3(n12083), .ZN(n12084)
         );
  NAND4_X1 U14454 ( .A1(keyinput30), .A2(n12086), .A3(n12085), .A4(n12084), 
        .ZN(n12092) );
  NOR3_X1 U14455 ( .A1(keyinput3), .A2(keyinput50), .A3(keyinput5), .ZN(n12089) );
  INV_X1 U14456 ( .A(keyinput4), .ZN(n12087) );
  NOR3_X1 U14457 ( .A1(keyinput62), .A2(keyinput37), .A3(n12087), .ZN(n12088)
         );
  NAND4_X1 U14458 ( .A1(keyinput12), .A2(n12089), .A3(keyinput10), .A4(n12088), 
        .ZN(n12091) );
  INV_X1 U14459 ( .A(keyinput22), .ZN(n12136) );
  NAND4_X1 U14460 ( .A1(keyinput47), .A2(keyinput9), .A3(keyinput31), .A4(
        n12136), .ZN(n12090) );
  OR4_X1 U14461 ( .A1(n12093), .A2(n12092), .A3(n12091), .A4(n12090), .ZN(
        n12210) );
  XOR2_X1 U14462 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput35), .Z(n12099) );
  XOR2_X1 U14463 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput23), .Z(n12098) );
  XNOR2_X1 U14464 ( .A(n12094), .B(keyinput18), .ZN(n12097) );
  XNOR2_X1 U14465 ( .A(n12095), .B(keyinput43), .ZN(n12096) );
  NOR4_X1 U14466 ( .A1(n12099), .A2(n12098), .A3(n12097), .A4(n12096), .ZN(
        n12119) );
  XNOR2_X1 U14467 ( .A(n8266), .B(keyinput10), .ZN(n12105) );
  XOR2_X1 U14468 ( .A(P3_IR_REG_31__SCAN_IN), .B(keyinput32), .Z(n12104) );
  XNOR2_X1 U14469 ( .A(n12100), .B(keyinput28), .ZN(n12103) );
  XNOR2_X1 U14470 ( .A(n12101), .B(keyinput9), .ZN(n12102) );
  NOR4_X1 U14471 ( .A1(n12105), .A2(n12104), .A3(n12103), .A4(n12102), .ZN(
        n12118) );
  XNOR2_X1 U14472 ( .A(n12106), .B(keyinput6), .ZN(n12116) );
  XNOR2_X1 U14473 ( .A(P2_REG0_REG_21__SCAN_IN), .B(keyinput17), .ZN(n12110)
         );
  XNOR2_X1 U14474 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput40), .ZN(n12109) );
  XNOR2_X1 U14475 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput53), .ZN(n12108)
         );
  XNOR2_X1 U14476 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput8), .ZN(n12107) );
  NAND4_X1 U14477 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12115) );
  XNOR2_X1 U14478 ( .A(n12111), .B(keyinput13), .ZN(n12114) );
  XNOR2_X1 U14479 ( .A(keyinput59), .B(n12112), .ZN(n12113) );
  NOR4_X1 U14480 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12117) );
  NAND3_X1 U14481 ( .A1(n12119), .A2(n12118), .A3(n12117), .ZN(n12126) );
  INV_X1 U14482 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14590) );
  AOI22_X1 U14483 ( .A1(n14590), .A2(keyinput49), .B1(n12121), .B2(keyinput24), 
        .ZN(n12120) );
  OAI221_X1 U14484 ( .B1(n14590), .B2(keyinput49), .C1(n12121), .C2(keyinput24), .A(n12120), .ZN(n12125) );
  INV_X1 U14485 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14913) );
  AOI22_X1 U14486 ( .A1(n14913), .A2(keyinput3), .B1(keyinput50), .B2(n12407), 
        .ZN(n12122) );
  OAI221_X1 U14487 ( .B1(n14913), .B2(keyinput3), .C1(n12407), .C2(keyinput50), 
        .A(n12122), .ZN(n12124) );
  INV_X1 U14488 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14740) );
  XNOR2_X1 U14489 ( .A(n14740), .B(keyinput47), .ZN(n12123) );
  NOR4_X1 U14490 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n12123), .ZN(
        n12152) );
  INV_X1 U14491 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U14492 ( .A1(n12129), .A2(keyinput29), .B1(keyinput33), .B2(n12128), 
        .ZN(n12127) );
  OAI221_X1 U14493 ( .B1(n12129), .B2(keyinput29), .C1(n12128), .C2(keyinput33), .A(n12127), .ZN(n12130) );
  INV_X1 U14494 ( .A(n12130), .ZN(n12134) );
  XNOR2_X1 U14495 ( .A(keyinput61), .B(n12528), .ZN(n12132) );
  XNOR2_X1 U14496 ( .A(keyinput4), .B(n9449), .ZN(n12131) );
  NOR2_X1 U14497 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  NAND2_X1 U14498 ( .A1(n12134), .A2(n12133), .ZN(n12139) );
  AOI22_X1 U14499 ( .A1(n12137), .A2(keyinput31), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n12136), .ZN(n12135) );
  OAI221_X1 U14500 ( .B1(n12137), .B2(keyinput31), .C1(n12136), .C2(
        P3_ADDR_REG_15__SCAN_IN), .A(n12135), .ZN(n12138) );
  NOR2_X1 U14501 ( .A1(n12139), .A2(n12138), .ZN(n12151) );
  AOI22_X1 U14502 ( .A1(n8752), .A2(keyinput57), .B1(n12776), .B2(keyinput21), 
        .ZN(n12140) );
  OAI221_X1 U14503 ( .B1(n8752), .B2(keyinput57), .C1(n12776), .C2(keyinput21), 
        .A(n12140), .ZN(n12144) );
  AOI22_X1 U14504 ( .A1(n8698), .A2(keyinput34), .B1(keyinput27), .B2(n12142), 
        .ZN(n12141) );
  OAI221_X1 U14505 ( .B1(n8698), .B2(keyinput34), .C1(n12142), .C2(keyinput27), 
        .A(n12141), .ZN(n12143) );
  NOR2_X1 U14506 ( .A1(n12144), .A2(n12143), .ZN(n12150) );
  INV_X1 U14507 ( .A(keyinput51), .ZN(n12145) );
  XNOR2_X1 U14508 ( .A(n12145), .B(P3_DATAO_REG_12__SCAN_IN), .ZN(n12148) );
  INV_X1 U14509 ( .A(keyinput15), .ZN(n12146) );
  XNOR2_X1 U14510 ( .A(n12146), .B(P3_DATAO_REG_20__SCAN_IN), .ZN(n12147) );
  NOR2_X1 U14511 ( .A1(n12148), .A2(n12147), .ZN(n12149) );
  AND4_X1 U14512 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12195) );
  INV_X1 U14513 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14741) );
  AOI22_X1 U14514 ( .A1(n14741), .A2(keyinput11), .B1(n12154), .B2(keyinput45), 
        .ZN(n12153) );
  OAI221_X1 U14515 ( .B1(n14741), .B2(keyinput11), .C1(n12154), .C2(keyinput45), .A(n12153), .ZN(n12162) );
  INV_X1 U14516 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13127) );
  AOI22_X1 U14517 ( .A1(n13127), .A2(keyinput7), .B1(keyinput16), .B2(n12720), 
        .ZN(n12155) );
  OAI221_X1 U14518 ( .B1(n13127), .B2(keyinput7), .C1(n12720), .C2(keyinput16), 
        .A(n12155), .ZN(n12161) );
  INV_X1 U14519 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14544) );
  AOI22_X1 U14520 ( .A1(n14544), .A2(keyinput41), .B1(keyinput58), .B2(n13090), 
        .ZN(n12156) );
  OAI221_X1 U14521 ( .B1(n14544), .B2(keyinput41), .C1(n13090), .C2(keyinput58), .A(n12156), .ZN(n12160) );
  INV_X1 U14522 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n14954) );
  AOI22_X1 U14523 ( .A1(n12158), .A2(keyinput63), .B1(n14954), .B2(keyinput26), 
        .ZN(n12157) );
  OAI221_X1 U14524 ( .B1(n12158), .B2(keyinput63), .C1(n14954), .C2(keyinput26), .A(n12157), .ZN(n12159) );
  NOR4_X1 U14525 ( .A1(n12162), .A2(n12161), .A3(n12160), .A4(n12159), .ZN(
        n12194) );
  AOI22_X1 U14526 ( .A1(n12262), .A2(keyinput56), .B1(n12164), .B2(keyinput1), 
        .ZN(n12163) );
  OAI221_X1 U14527 ( .B1(n12262), .B2(keyinput56), .C1(n12164), .C2(keyinput1), 
        .A(n12163), .ZN(n12175) );
  INV_X1 U14528 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14742) );
  INV_X1 U14529 ( .A(keyinput0), .ZN(n12166) );
  AOI22_X1 U14530 ( .A1(n14742), .A2(keyinput44), .B1(P1_ADDR_REG_6__SCAN_IN), 
        .B2(n12166), .ZN(n12165) );
  OAI221_X1 U14531 ( .B1(n14742), .B2(keyinput44), .C1(n12166), .C2(
        P1_ADDR_REG_6__SCAN_IN), .A(n12165), .ZN(n12174) );
  INV_X1 U14532 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n12169) );
  INV_X1 U14533 ( .A(keyinput62), .ZN(n12168) );
  AOI22_X1 U14534 ( .A1(n12169), .A2(keyinput37), .B1(P3_DATAO_REG_28__SCAN_IN), .B2(n12168), .ZN(n12167) );
  OAI221_X1 U14535 ( .B1(n12169), .B2(keyinput37), .C1(n12168), .C2(
        P3_DATAO_REG_28__SCAN_IN), .A(n12167), .ZN(n12173) );
  INV_X1 U14536 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n12171) );
  INV_X1 U14537 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14953) );
  AOI22_X1 U14538 ( .A1(n12171), .A2(keyinput39), .B1(n14953), .B2(keyinput19), 
        .ZN(n12170) );
  OAI221_X1 U14539 ( .B1(n12171), .B2(keyinput39), .C1(n14953), .C2(keyinput19), .A(n12170), .ZN(n12172) );
  NOR4_X1 U14540 ( .A1(n12175), .A2(n12174), .A3(n12173), .A4(n12172), .ZN(
        n12193) );
  INV_X1 U14541 ( .A(keyinput5), .ZN(n12178) );
  INV_X1 U14542 ( .A(keyinput12), .ZN(n12177) );
  AOI22_X1 U14543 ( .A1(n12178), .A2(P3_DATAO_REG_1__SCAN_IN), .B1(
        P3_ADDR_REG_3__SCAN_IN), .B2(n12177), .ZN(n12176) );
  OAI221_X1 U14544 ( .B1(n12178), .B2(P3_DATAO_REG_1__SCAN_IN), .C1(n12177), 
        .C2(P3_ADDR_REG_3__SCAN_IN), .A(n12176), .ZN(n12191) );
  INV_X1 U14545 ( .A(keyinput46), .ZN(n12180) );
  AOI22_X1 U14546 ( .A1(n12181), .A2(keyinput42), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n12180), .ZN(n12179) );
  OAI221_X1 U14547 ( .B1(n12181), .B2(keyinput42), .C1(n12180), .C2(
        P1_ADDR_REG_16__SCAN_IN), .A(n12179), .ZN(n12190) );
  INV_X1 U14548 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U14549 ( .A1(n12184), .A2(keyinput48), .B1(n12183), .B2(keyinput55), 
        .ZN(n12182) );
  OAI221_X1 U14550 ( .B1(n12184), .B2(keyinput48), .C1(n12183), .C2(keyinput55), .A(n12182), .ZN(n12189) );
  INV_X1 U14551 ( .A(keyinput2), .ZN(n12186) );
  AOI22_X1 U14552 ( .A1(n12187), .A2(keyinput60), .B1(P1_ADDR_REG_2__SCAN_IN), 
        .B2(n12186), .ZN(n12185) );
  OAI221_X1 U14553 ( .B1(n12187), .B2(keyinput60), .C1(n12186), .C2(
        P1_ADDR_REG_2__SCAN_IN), .A(n12185), .ZN(n12188) );
  NOR4_X1 U14554 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12192) );
  AND4_X1 U14555 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n12209) );
  INV_X1 U14556 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14536) );
  INV_X1 U14557 ( .A(keyinput30), .ZN(n12197) );
  AOI22_X1 U14558 ( .A1(n14536), .A2(keyinput52), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n12197), .ZN(n12196) );
  OAI221_X1 U14559 ( .B1(n14536), .B2(keyinput52), .C1(n12197), .C2(
        P3_ADDR_REG_14__SCAN_IN), .A(n12196), .ZN(n12207) );
  AOI22_X1 U14560 ( .A1(n12199), .A2(keyinput20), .B1(keyinput38), .B2(n13494), 
        .ZN(n12198) );
  OAI221_X1 U14561 ( .B1(n12199), .B2(keyinput20), .C1(n13494), .C2(keyinput38), .A(n12198), .ZN(n12206) );
  INV_X1 U14562 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12201) );
  INV_X1 U14563 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U14564 ( .A1(n12201), .A2(keyinput14), .B1(keyinput25), .B2(n14448), 
        .ZN(n12200) );
  OAI221_X1 U14565 ( .B1(n12201), .B2(keyinput14), .C1(n14448), .C2(keyinput25), .A(n12200), .ZN(n12205) );
  INV_X1 U14566 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U14567 ( .A1(n12203), .A2(keyinput36), .B1(n12805), .B2(keyinput54), 
        .ZN(n12202) );
  OAI221_X1 U14568 ( .B1(n12203), .B2(keyinput36), .C1(n12805), .C2(keyinput54), .A(n12202), .ZN(n12204) );
  NOR4_X1 U14569 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12208) );
  OAI211_X1 U14570 ( .C1(n12211), .C2(n12210), .A(n12209), .B(n12208), .ZN(
        n12212) );
  XNOR2_X1 U14571 ( .A(n12213), .B(n12212), .ZN(P1_U3356) );
  OAI222_X1 U14572 ( .A1(n13461), .A2(n13727), .B1(n12215), .B2(P2_U3088), 
        .C1(n12214), .C2(n13458), .ZN(P2_U3297) );
  INV_X1 U14573 ( .A(n13431), .ZN(n13440) );
  INV_X1 U14574 ( .A(n12218), .ZN(n12220) );
  AOI22_X1 U14575 ( .A1(n14174), .A2(n12222), .B1(n9910), .B2(n13821), .ZN(
        n12226) );
  AOI22_X1 U14576 ( .A1(n14174), .A2(n11966), .B1(n12223), .B2(n13821), .ZN(
        n12224) );
  XNOR2_X1 U14577 ( .A(n12224), .B(n10393), .ZN(n12225) );
  XOR2_X1 U14578 ( .A(n12226), .B(n12225), .Z(n12227) );
  INV_X1 U14579 ( .A(n13989), .ZN(n12230) );
  OAI22_X1 U14580 ( .A1(n12228), .A2(n13542), .B1(n13741), .B2(n13544), .ZN(
        n13981) );
  AOI22_X1 U14581 ( .A1(n13981), .A2(n14578), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12229) );
  OAI21_X1 U14582 ( .B1(n12230), .B2(n14659), .A(n12229), .ZN(n12231) );
  AOI21_X1 U14583 ( .B1(n14174), .B2(n14657), .A(n12231), .ZN(n12232) );
  OAI21_X1 U14584 ( .B1(n12233), .B2(n14651), .A(n12232), .ZN(P1_U3220) );
  OAI222_X1 U14585 ( .A1(n12235), .A2(P1_U3086), .B1(n14286), .B2(n13727), 
        .C1(n12234), .C2(n6454), .ZN(P1_U3325) );
  INV_X1 U14586 ( .A(SI_30_), .ZN(n12238) );
  INV_X1 U14587 ( .A(n12236), .ZN(n12237) );
  OAI222_X1 U14588 ( .A1(P3_U3151), .A2(n12239), .B1(n12829), .B2(n12238), 
        .C1(n12832), .C2(n12237), .ZN(P3_U3265) );
  XNOR2_X1 U14589 ( .A(n12542), .B(n12240), .ZN(n12248) );
  INV_X1 U14590 ( .A(n12248), .ZN(n12241) );
  INV_X1 U14591 ( .A(n12242), .ZN(n12243) );
  AOI22_X1 U14592 ( .A1(n7018), .A2(n12352), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12245) );
  NAND2_X1 U14593 ( .A1(n12545), .A2(n12356), .ZN(n12244) );
  OAI211_X1 U14594 ( .C1(n12246), .C2(n12354), .A(n12245), .B(n12244), .ZN(
        n12250) );
  NOR4_X1 U14595 ( .A1(n12248), .A2(n12247), .A3(n7018), .A4(n12347), .ZN(
        n12249) );
  AOI211_X1 U14596 ( .C1(n12334), .C2(n12544), .A(n12250), .B(n12249), .ZN(
        n12251) );
  INV_X1 U14597 ( .A(n12252), .ZN(n12253) );
  OAI222_X1 U14598 ( .A1(n12255), .A2(P3_U3151), .B1(n12829), .B2(n12254), 
        .C1(n12832), .C2(n12253), .ZN(P3_U3270) );
  AOI21_X1 U14599 ( .B1(n12364), .B2(n12256), .A(n6466), .ZN(n12261) );
  AOI22_X1 U14600 ( .A1(n12365), .A2(n12352), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12258) );
  NAND2_X1 U14601 ( .A1(n12356), .A2(n12611), .ZN(n12257) );
  OAI211_X1 U14602 ( .C1(n12607), .C2(n12354), .A(n12258), .B(n12257), .ZN(
        n12259) );
  AOI21_X1 U14603 ( .B1(n12610), .B2(n12334), .A(n12259), .ZN(n12260) );
  OAI21_X1 U14604 ( .B1(n12261), .B2(n12347), .A(n12260), .ZN(P3_U3156) );
  XNOR2_X1 U14605 ( .A(n12306), .B(n12305), .ZN(n12267) );
  NOR2_X1 U14606 ( .A1(n12262), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12519) );
  AOI21_X1 U14607 ( .B1(n12367), .B2(n12311), .A(n12519), .ZN(n12263) );
  OAI21_X1 U14608 ( .B1(n12681), .B2(n12314), .A(n12263), .ZN(n12265) );
  NOR2_X1 U14609 ( .A1(n12808), .A2(n12360), .ZN(n12264) );
  AOI211_X1 U14610 ( .C1(n12660), .C2(n12356), .A(n12265), .B(n12264), .ZN(
        n12266) );
  OAI21_X1 U14611 ( .B1(n12267), .B2(n12347), .A(n12266), .ZN(P3_U3159) );
  NAND2_X1 U14612 ( .A1(n12269), .A2(n12268), .ZN(n12270) );
  AOI21_X1 U14613 ( .B1(n12271), .B2(n12270), .A(n6542), .ZN(n12276) );
  AOI22_X1 U14614 ( .A1(n12367), .A2(n12352), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12273) );
  NAND2_X1 U14615 ( .A1(n12356), .A2(n12632), .ZN(n12272) );
  OAI211_X1 U14616 ( .C1(n12628), .C2(n12354), .A(n12273), .B(n12272), .ZN(
        n12274) );
  AOI21_X1 U14617 ( .B1(n12631), .B2(n12334), .A(n12274), .ZN(n12275) );
  OAI21_X1 U14618 ( .B1(n12276), .B2(n12347), .A(n12275), .ZN(P3_U3163) );
  INV_X1 U14619 ( .A(n12709), .ZN(n12585) );
  NOR3_X1 U14620 ( .A1(n6482), .A2(n6756), .A3(n12278), .ZN(n12281) );
  INV_X1 U14621 ( .A(n12279), .ZN(n12280) );
  OAI21_X1 U14622 ( .B1(n12281), .B2(n12280), .A(n12341), .ZN(n12286) );
  AOI22_X1 U14623 ( .A1(n12363), .A2(n12352), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12282) );
  OAI21_X1 U14624 ( .B1(n12283), .B2(n12354), .A(n12282), .ZN(n12284) );
  AOI21_X1 U14625 ( .B1(n12583), .B2(n12356), .A(n12284), .ZN(n12285) );
  OAI211_X1 U14626 ( .C1(n12585), .C2(n12360), .A(n12286), .B(n12285), .ZN(
        P3_U3165) );
  XNOR2_X1 U14627 ( .A(n12287), .B(n12682), .ZN(n12288) );
  XNOR2_X1 U14628 ( .A(n12289), .B(n12288), .ZN(n12296) );
  NAND2_X1 U14629 ( .A1(n12352), .A2(n12370), .ZN(n12290) );
  NAND2_X1 U14630 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12468)
         );
  OAI211_X1 U14631 ( .C1(n12291), .C2(n12354), .A(n12290), .B(n12468), .ZN(
        n12292) );
  AOI21_X1 U14632 ( .B1(n12293), .B2(n12356), .A(n12292), .ZN(n12295) );
  NAND2_X1 U14633 ( .A1(n12747), .A2(n12334), .ZN(n12294) );
  OAI211_X1 U14634 ( .C1(n12296), .C2(n12347), .A(n12295), .B(n12294), .ZN(
        P3_U3166) );
  INV_X1 U14635 ( .A(n12297), .ZN(n12788) );
  NOR3_X1 U14636 ( .A1(n6466), .A2(n6761), .A3(n12299), .ZN(n12300) );
  OAI21_X1 U14637 ( .B1(n12300), .B2(n6482), .A(n12341), .ZN(n12304) );
  AOI22_X1 U14638 ( .A1(n12362), .A2(n12311), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12301) );
  OAI21_X1 U14639 ( .B1(n12618), .B2(n12314), .A(n12301), .ZN(n12302) );
  AOI21_X1 U14640 ( .B1(n12599), .B2(n12356), .A(n12302), .ZN(n12303) );
  OAI211_X1 U14641 ( .C1(n12788), .C2(n12360), .A(n12304), .B(n12303), .ZN(
        P3_U3169) );
  NAND2_X1 U14642 ( .A1(n12306), .A2(n12305), .ZN(n12308) );
  NAND2_X1 U14643 ( .A1(n12308), .A2(n12307), .ZN(n12310) );
  XNOR2_X1 U14644 ( .A(n12310), .B(n12309), .ZN(n12317) );
  AOI22_X1 U14645 ( .A1(n12366), .A2(n12311), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12313) );
  NAND2_X1 U14646 ( .A1(n12356), .A2(n12647), .ZN(n12312) );
  OAI211_X1 U14647 ( .C1(n12332), .C2(n12314), .A(n12313), .B(n12312), .ZN(
        n12315) );
  AOI21_X1 U14648 ( .B1(n12646), .B2(n12334), .A(n12315), .ZN(n12316) );
  OAI21_X1 U14649 ( .B1(n12317), .B2(n12347), .A(n12316), .ZN(P3_U3173) );
  INV_X1 U14650 ( .A(n12318), .ZN(n12319) );
  AOI21_X1 U14651 ( .B1(n12365), .B2(n12320), .A(n12319), .ZN(n12326) );
  AOI22_X1 U14652 ( .A1(n12366), .A2(n12352), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12322) );
  NAND2_X1 U14653 ( .A1(n12356), .A2(n12621), .ZN(n12321) );
  OAI211_X1 U14654 ( .C1(n12618), .C2(n12354), .A(n12322), .B(n12321), .ZN(
        n12323) );
  AOI21_X1 U14655 ( .B1(n12324), .B2(n12334), .A(n12323), .ZN(n12325) );
  OAI21_X1 U14656 ( .B1(n12326), .B2(n12347), .A(n12325), .ZN(P3_U3175) );
  NAND2_X1 U14657 ( .A1(n12328), .A2(n12327), .ZN(n12330) );
  XNOR2_X1 U14658 ( .A(n12330), .B(n12329), .ZN(n12337) );
  NAND2_X1 U14659 ( .A1(n12352), .A2(n12668), .ZN(n12331) );
  NAND2_X1 U14660 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12490)
         );
  OAI211_X1 U14661 ( .C1(n12332), .C2(n12354), .A(n12331), .B(n12490), .ZN(
        n12333) );
  AOI21_X1 U14662 ( .B1(n12673), .B2(n12356), .A(n12333), .ZN(n12336) );
  NAND2_X1 U14663 ( .A1(n12739), .A2(n12334), .ZN(n12335) );
  OAI211_X1 U14664 ( .C1(n12337), .C2(n12347), .A(n12336), .B(n12335), .ZN(
        P3_U3178) );
  NAND2_X1 U14665 ( .A1(n12342), .A2(n12341), .ZN(n12346) );
  AOI22_X1 U14666 ( .A1(n12362), .A2(n12352), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12343) );
  OAI21_X1 U14667 ( .B1(n12564), .B2(n12354), .A(n12343), .ZN(n12344) );
  AOI21_X1 U14668 ( .B1(n12567), .B2(n12356), .A(n12344), .ZN(n12345) );
  OAI211_X1 U14669 ( .C1(n12783), .C2(n12360), .A(n12346), .B(n12345), .ZN(
        P3_U3180) );
  AOI21_X1 U14670 ( .B1(n12349), .B2(n12348), .A(n12347), .ZN(n12351) );
  NAND2_X1 U14671 ( .A1(n12351), .A2(n12350), .ZN(n12359) );
  NAND2_X1 U14672 ( .A1(n12352), .A2(n12371), .ZN(n12353) );
  NAND2_X1 U14673 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12443)
         );
  OAI211_X1 U14674 ( .C1(n12682), .C2(n12354), .A(n12353), .B(n12443), .ZN(
        n12355) );
  AOI21_X1 U14675 ( .B1(n12357), .B2(n12356), .A(n12355), .ZN(n12358) );
  OAI211_X1 U14676 ( .C1(n12819), .C2(n12360), .A(n12359), .B(n12358), .ZN(
        P3_U3181) );
  MUX2_X1 U14677 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12361), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14678 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12539), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14679 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12552), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14680 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n7018), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14681 ( .A(n12578), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12385), .Z(
        P3_U3517) );
  MUX2_X1 U14682 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12362), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14683 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12363), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14684 ( .A(n12364), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12385), .Z(
        P3_U3514) );
  MUX2_X1 U14685 ( .A(n12365), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12385), .Z(
        P3_U3513) );
  MUX2_X1 U14686 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12366), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14687 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12367), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14688 ( .A(n12667), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12385), .Z(
        P3_U3510) );
  MUX2_X1 U14689 ( .A(n12368), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12385), .Z(
        P3_U3509) );
  MUX2_X1 U14690 ( .A(n12668), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12385), .Z(
        P3_U3508) );
  MUX2_X1 U14691 ( .A(n12369), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12385), .Z(
        P3_U3507) );
  MUX2_X1 U14692 ( .A(n12370), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12385), .Z(
        P3_U3506) );
  MUX2_X1 U14693 ( .A(n12371), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12385), .Z(
        P3_U3505) );
  MUX2_X1 U14694 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12372), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14695 ( .A(n12373), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12385), .Z(
        P3_U3503) );
  MUX2_X1 U14696 ( .A(n12374), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12385), .Z(
        P3_U3502) );
  MUX2_X1 U14697 ( .A(n12375), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12385), .Z(
        P3_U3501) );
  MUX2_X1 U14698 ( .A(n12376), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12385), .Z(
        P3_U3500) );
  MUX2_X1 U14699 ( .A(n12377), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12385), .Z(
        P3_U3499) );
  MUX2_X1 U14700 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12378), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14701 ( .A(n12379), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12385), .Z(
        P3_U3497) );
  MUX2_X1 U14702 ( .A(n12380), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12385), .Z(
        P3_U3496) );
  MUX2_X1 U14703 ( .A(n12381), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12385), .Z(
        P3_U3495) );
  MUX2_X1 U14704 ( .A(n12382), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12385), .Z(
        P3_U3494) );
  MUX2_X1 U14705 ( .A(n12383), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12385), .Z(
        P3_U3493) );
  MUX2_X1 U14706 ( .A(n12384), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12385), .Z(
        P3_U3492) );
  MUX2_X1 U14707 ( .A(n12757), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12385), .Z(
        P3_U3491) );
  INV_X1 U14708 ( .A(n12405), .ZN(n14409) );
  AOI21_X1 U14709 ( .B1(n8352), .B2(n12387), .A(n12406), .ZN(n12403) );
  NAND2_X1 U14710 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12389), .ZN(n12411) );
  OAI21_X1 U14711 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12389), .A(n12411), 
        .ZN(n12401) );
  MUX2_X1 U14712 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6622), .Z(n12419) );
  XNOR2_X1 U14713 ( .A(n12419), .B(n14409), .ZN(n12395) );
  INV_X1 U14714 ( .A(n12390), .ZN(n12392) );
  OAI21_X1 U14715 ( .B1(n12393), .B2(n12392), .A(n12391), .ZN(n12394) );
  NOR2_X1 U14716 ( .A1(n12394), .A2(n12395), .ZN(n12424) );
  AOI21_X1 U14717 ( .B1(n12395), .B2(n12394), .A(n12424), .ZN(n12399) );
  INV_X1 U14718 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14314) );
  NOR2_X1 U14719 ( .A1(n15106), .A2(n14314), .ZN(n12396) );
  AOI211_X1 U14720 ( .C1(n15102), .C2(n12405), .A(n12397), .B(n12396), .ZN(
        n12398) );
  OAI21_X1 U14721 ( .B1(n12399), .B2(n15096), .A(n12398), .ZN(n12400) );
  AOI21_X1 U14722 ( .B1(n15086), .B2(n12401), .A(n12400), .ZN(n12402) );
  OAI21_X1 U14723 ( .B1(n12403), .B2(n15091), .A(n12402), .ZN(P3_U3195) );
  INV_X1 U14724 ( .A(n12440), .ZN(n12414) );
  NAND2_X1 U14725 ( .A1(n12414), .A2(n12407), .ZN(n12408) );
  NAND2_X1 U14726 ( .A1(n6596), .A2(n12408), .ZN(n12422) );
  AOI21_X1 U14727 ( .B1(n12409), .B2(n12422), .A(n12432), .ZN(n12431) );
  NAND2_X1 U14728 ( .A1(n14409), .A2(n12410), .ZN(n12412) );
  NAND2_X1 U14729 ( .A1(n12414), .A2(n12413), .ZN(n12415) );
  NAND2_X1 U14730 ( .A1(n12440), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12436) );
  AND2_X1 U14731 ( .A1(n12415), .A2(n12436), .ZN(n12420) );
  OAI21_X1 U14732 ( .B1(n12416), .B2(n12420), .A(n12435), .ZN(n12429) );
  AOI21_X1 U14733 ( .B1(n15075), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12417), 
        .ZN(n12418) );
  OAI21_X1 U14734 ( .B1(n15070), .B2(n12440), .A(n12418), .ZN(n12428) );
  NOR2_X1 U14735 ( .A1(n12419), .A2(n14409), .ZN(n12423) );
  OR2_X1 U14736 ( .A1(n12424), .A2(n12423), .ZN(n12426) );
  INV_X1 U14737 ( .A(n12420), .ZN(n12421) );
  MUX2_X1 U14738 ( .A(n12422), .B(n12421), .S(n6622), .Z(n12425) );
  AOI211_X1 U14739 ( .C1(n12426), .C2(n12425), .A(n15096), .B(n12438), .ZN(
        n12427) );
  AOI211_X1 U14740 ( .C1(n15086), .C2(n12429), .A(n12428), .B(n12427), .ZN(
        n12430) );
  OAI21_X1 U14741 ( .B1(n12431), .B2(n15091), .A(n12430), .ZN(P3_U3196) );
  XNOR2_X1 U14742 ( .A(n12462), .B(n12451), .ZN(n12433) );
  NOR2_X1 U14743 ( .A1(n12434), .A2(n12433), .ZN(n12452) );
  AOI21_X1 U14744 ( .B1(n12434), .B2(n12433), .A(n12452), .ZN(n12450) );
  INV_X1 U14745 ( .A(n12462), .ZN(n14415) );
  NAND2_X1 U14746 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12437), .ZN(n12457) );
  OAI21_X1 U14747 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12437), .A(n12457), 
        .ZN(n12448) );
  MUX2_X1 U14748 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6622), .Z(n12442) );
  MUX2_X1 U14749 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n6622), .Z(n12439) );
  AOI21_X1 U14750 ( .B1(n12440), .B2(n12439), .A(n12438), .ZN(n12463) );
  XNOR2_X1 U14751 ( .A(n12463), .B(n12462), .ZN(n12441) );
  AOI21_X1 U14752 ( .B1(n12442), .B2(n12441), .A(n12461), .ZN(n12446) );
  INV_X1 U14753 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14318) );
  OAI21_X1 U14754 ( .B1(n15106), .B2(n14318), .A(n12443), .ZN(n12444) );
  AOI21_X1 U14755 ( .B1(n15102), .B2(n12462), .A(n12444), .ZN(n12445) );
  OAI21_X1 U14756 ( .B1(n12446), .B2(n15096), .A(n12445), .ZN(n12447) );
  AOI21_X1 U14757 ( .B1(n15086), .B2(n12448), .A(n12447), .ZN(n12449) );
  OAI21_X1 U14758 ( .B1(n12450), .B2(n15091), .A(n12449), .ZN(P3_U3197) );
  NOR2_X1 U14759 ( .A1(n12462), .A2(n12451), .ZN(n12453) );
  NOR2_X1 U14760 ( .A1(n12453), .A2(n12452), .ZN(n12455) );
  INV_X1 U14761 ( .A(n12494), .ZN(n14418) );
  AOI22_X1 U14762 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12494), .B1(n14418), 
        .B2(n12464), .ZN(n12454) );
  NOR2_X1 U14763 ( .A1(n12455), .A2(n12454), .ZN(n12483) );
  AOI21_X1 U14764 ( .B1(n12455), .B2(n12454), .A(n12483), .ZN(n12475) );
  INV_X1 U14765 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U14766 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n14418), .B1(n12494), 
        .B2(n12493), .ZN(n12460) );
  NAND2_X1 U14767 ( .A1(n14415), .A2(n12456), .ZN(n12458) );
  OAI21_X1 U14768 ( .B1(n12460), .B2(n12459), .A(n12492), .ZN(n12473) );
  AOI21_X1 U14769 ( .B1(n12463), .B2(n12462), .A(n12461), .ZN(n12479) );
  MUX2_X1 U14770 ( .A(n12464), .B(n12493), .S(n6622), .Z(n12465) );
  NOR2_X1 U14771 ( .A1(n12465), .A2(n12494), .ZN(n12478) );
  NAND2_X1 U14772 ( .A1(n12465), .A2(n12494), .ZN(n12477) );
  INV_X1 U14773 ( .A(n12477), .ZN(n12466) );
  NOR2_X1 U14774 ( .A1(n12478), .A2(n12466), .ZN(n12467) );
  XNOR2_X1 U14775 ( .A(n12479), .B(n12467), .ZN(n12471) );
  INV_X1 U14776 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14291) );
  OAI21_X1 U14777 ( .B1(n15106), .B2(n14291), .A(n12468), .ZN(n12469) );
  AOI21_X1 U14778 ( .B1(n15102), .B2(n12494), .A(n12469), .ZN(n12470) );
  OAI21_X1 U14779 ( .B1(n12471), .B2(n15096), .A(n12470), .ZN(n12472) );
  AOI21_X1 U14780 ( .B1(n15086), .B2(n12473), .A(n12472), .ZN(n12474) );
  OAI21_X1 U14781 ( .B1(n12475), .B2(n15091), .A(n12474), .ZN(P3_U3198) );
  MUX2_X1 U14782 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6622), .Z(n12482) );
  MUX2_X1 U14783 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6622), .Z(n12480) );
  OAI21_X1 U14784 ( .B1(n12479), .B2(n12478), .A(n12477), .ZN(n14456) );
  XNOR2_X1 U14785 ( .A(n12480), .B(n14398), .ZN(n14457) );
  NOR2_X1 U14786 ( .A1(n14456), .A2(n14457), .ZN(n14455) );
  XNOR2_X1 U14787 ( .A(n12510), .B(n12509), .ZN(n12481) );
  NOR2_X1 U14788 ( .A1(n12481), .A2(n12482), .ZN(n12508) );
  AOI21_X1 U14789 ( .B1(n12482), .B2(n12481), .A(n12508), .ZN(n12504) );
  INV_X1 U14790 ( .A(n14398), .ZN(n14451) );
  NAND2_X1 U14791 ( .A1(n14425), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12505) );
  OR2_X1 U14792 ( .A1(n14425), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12485) );
  AND2_X1 U14793 ( .A1(n12505), .A2(n12485), .ZN(n12486) );
  INV_X1 U14794 ( .A(n12506), .ZN(n12489) );
  NOR3_X1 U14795 ( .A1(n14446), .A2(n7432), .A3(n12486), .ZN(n12488) );
  OAI21_X1 U14796 ( .B1(n12489), .B2(n12488), .A(n12487), .ZN(n12503) );
  INV_X1 U14797 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12491) );
  OAI21_X1 U14798 ( .B1(n15106), .B2(n12491), .A(n12490), .ZN(n12501) );
  NAND2_X1 U14799 ( .A1(n12495), .A2(n14398), .ZN(n12497) );
  NAND2_X1 U14800 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14450), .ZN(n14449) );
  XNOR2_X1 U14801 ( .A(n14425), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12496) );
  AOI21_X1 U14802 ( .B1(n12497), .B2(n14449), .A(n12496), .ZN(n12515) );
  INV_X1 U14803 ( .A(n12515), .ZN(n12499) );
  NAND3_X1 U14804 ( .A1(n12497), .A2(n14449), .A3(n12496), .ZN(n12498) );
  AOI21_X1 U14805 ( .B1(n12499), .B2(n12498), .A(n15040), .ZN(n12500) );
  AOI211_X1 U14806 ( .C1(n15102), .C2(n12509), .A(n12501), .B(n12500), .ZN(
        n12502) );
  OAI211_X1 U14807 ( .C1(n12504), .C2(n15096), .A(n12503), .B(n12502), .ZN(
        P3_U3200) );
  NAND2_X1 U14808 ( .A1(n12506), .A2(n12505), .ZN(n12507) );
  XNOR2_X1 U14809 ( .A(n12517), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12512) );
  XNOR2_X1 U14810 ( .A(n12507), .B(n12512), .ZN(n12523) );
  AOI21_X1 U14811 ( .B1(n12510), .B2(n12509), .A(n12508), .ZN(n12514) );
  XNOR2_X1 U14812 ( .A(n12517), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12516) );
  MUX2_X1 U14813 ( .A(n12516), .B(n12512), .S(n12511), .Z(n12513) );
  XNOR2_X1 U14814 ( .A(n12514), .B(n12513), .ZN(n12521) );
  NOR2_X1 U14815 ( .A1(n15070), .A2(n12517), .ZN(n12518) );
  AOI211_X1 U14816 ( .C1(P3_ADDR_REG_19__SCAN_IN), .C2(n15075), .A(n12519), 
        .B(n12518), .ZN(n12520) );
  OAI21_X1 U14817 ( .B1(n12523), .B2(n15091), .A(n12522), .ZN(P3_U3201) );
  NAND2_X1 U14818 ( .A1(n12773), .A2(n14463), .ZN(n12527) );
  NOR2_X1 U14819 ( .A1(n12526), .A2(n15111), .ZN(n12530) );
  AOI21_X1 U14820 ( .B1(n14466), .B2(n15117), .A(n12530), .ZN(n14465) );
  OAI211_X1 U14821 ( .C1(n15117), .C2(n12528), .A(n12527), .B(n14465), .ZN(
        P3_U3202) );
  INV_X1 U14822 ( .A(n12529), .ZN(n12536) );
  AOI21_X1 U14823 ( .B1(n15119), .B2(P3_REG2_REG_29__SCAN_IN), .A(n12530), 
        .ZN(n12531) );
  OAI21_X1 U14824 ( .B1(n12532), .B2(n12689), .A(n12531), .ZN(n12533) );
  AOI21_X1 U14825 ( .B1(n12534), .B2(n12691), .A(n12533), .ZN(n12535) );
  OAI21_X1 U14826 ( .B1(n12536), .B2(n15119), .A(n12535), .ZN(P3_U3204) );
  AOI22_X1 U14827 ( .A1(n7018), .A2(n12756), .B1(n12539), .B2(n12666), .ZN(
        n12540) );
  INV_X1 U14828 ( .A(n12699), .ZN(n12549) );
  XNOR2_X1 U14829 ( .A(n12543), .B(n12542), .ZN(n12697) );
  INV_X1 U14830 ( .A(n12544), .ZN(n12778) );
  AOI22_X1 U14831 ( .A1(n12545), .A2(n12687), .B1(P3_REG2_REG_28__SCAN_IN), 
        .B2(n15119), .ZN(n12546) );
  OAI21_X1 U14832 ( .B1(n12778), .B2(n12689), .A(n12546), .ZN(n12547) );
  AOI21_X1 U14833 ( .B1(n12697), .B2(n12691), .A(n12547), .ZN(n12548) );
  OAI21_X1 U14834 ( .B1(n12549), .B2(n15119), .A(n12548), .ZN(P3_U3205) );
  XNOR2_X1 U14835 ( .A(n12551), .B(n12550), .ZN(n12553) );
  AOI222_X1 U14836 ( .A1(n12762), .A2(n12553), .B1(n12552), .B2(n12666), .C1(
        n12578), .C2(n12756), .ZN(n12704) );
  OAI21_X1 U14837 ( .B1(n12556), .B2(n12555), .A(n12554), .ZN(n12702) );
  AOI22_X1 U14838 ( .A1(n12557), .A2(n12687), .B1(n15119), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12558) );
  OAI21_X1 U14839 ( .B1(n12559), .B2(n12689), .A(n12558), .ZN(n12560) );
  AOI21_X1 U14840 ( .B1(n12702), .B2(n12691), .A(n12560), .ZN(n12561) );
  OAI21_X1 U14841 ( .B1(n12704), .B2(n15119), .A(n12561), .ZN(P3_U3206) );
  XOR2_X1 U14842 ( .A(n12562), .B(n12565), .Z(n12563) );
  OAI222_X1 U14843 ( .A1(n12683), .A2(n12594), .B1(n12759), .B2(n12564), .C1(
        n12563), .C2(n12680), .ZN(n12705) );
  INV_X1 U14844 ( .A(n12705), .ZN(n12571) );
  XNOR2_X1 U14845 ( .A(n12566), .B(n12565), .ZN(n12706) );
  AOI22_X1 U14846 ( .A1(n12567), .A2(n12687), .B1(n15119), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12568) );
  OAI21_X1 U14847 ( .B1(n12783), .B2(n12689), .A(n12568), .ZN(n12569) );
  AOI21_X1 U14848 ( .B1(n12706), .B2(n12691), .A(n12569), .ZN(n12570) );
  OAI21_X1 U14849 ( .B1(n12571), .B2(n15119), .A(n12570), .ZN(P3_U3207) );
  NOR2_X1 U14850 ( .A1(n12607), .A2(n12683), .ZN(n12577) );
  INV_X1 U14851 ( .A(n12572), .ZN(n12575) );
  AOI21_X1 U14852 ( .B1(n12588), .B2(n12573), .A(n12580), .ZN(n12574) );
  NOR3_X1 U14853 ( .A1(n12575), .A2(n12574), .A3(n12680), .ZN(n12576) );
  AOI211_X1 U14854 ( .C1(n12666), .C2(n12578), .A(n12577), .B(n12576), .ZN(
        n12712) );
  NAND3_X1 U14855 ( .A1(n12591), .A2(n12580), .A3(n12579), .ZN(n12581) );
  NAND2_X1 U14856 ( .A1(n12582), .A2(n12581), .ZN(n12710) );
  AOI22_X1 U14857 ( .A1(n12583), .A2(n12687), .B1(n15119), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12584) );
  OAI21_X1 U14858 ( .B1(n12585), .B2(n12689), .A(n12584), .ZN(n12586) );
  AOI21_X1 U14859 ( .B1(n12710), .B2(n12691), .A(n12586), .ZN(n12587) );
  OAI21_X1 U14860 ( .B1(n12712), .B2(n15119), .A(n12587), .ZN(P3_U3208) );
  INV_X1 U14861 ( .A(n12588), .ZN(n12589) );
  AOI21_X1 U14862 ( .B1(n12592), .B2(n12590), .A(n12589), .ZN(n12598) );
  OAI21_X1 U14863 ( .B1(n12593), .B2(n12592), .A(n12591), .ZN(n12715) );
  OAI22_X1 U14864 ( .A1(n12594), .A2(n12759), .B1(n12618), .B2(n12683), .ZN(
        n12595) );
  AOI21_X1 U14865 ( .B1(n12715), .B2(n12596), .A(n12595), .ZN(n12597) );
  OAI21_X1 U14866 ( .B1(n12598), .B2(n12680), .A(n12597), .ZN(n12714) );
  INV_X1 U14867 ( .A(n12714), .ZN(n12604) );
  INV_X1 U14868 ( .A(n15114), .ZN(n12602) );
  AOI22_X1 U14869 ( .A1(n15119), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12599), 
        .B2(n12687), .ZN(n12600) );
  OAI21_X1 U14870 ( .B1(n12788), .B2(n12689), .A(n12600), .ZN(n12601) );
  AOI21_X1 U14871 ( .B1(n12715), .B2(n12602), .A(n12601), .ZN(n12603) );
  OAI21_X1 U14872 ( .B1(n12604), .B2(n15119), .A(n12603), .ZN(P3_U3209) );
  XNOR2_X1 U14873 ( .A(n12605), .B(n12608), .ZN(n12606) );
  OAI222_X1 U14874 ( .A1(n12759), .A2(n12607), .B1(n12683), .B2(n12628), .C1(
        n12606), .C2(n12680), .ZN(n12718) );
  INV_X1 U14875 ( .A(n12718), .ZN(n12615) );
  XNOR2_X1 U14876 ( .A(n12609), .B(n12608), .ZN(n12719) );
  INV_X1 U14877 ( .A(n12610), .ZN(n12792) );
  AOI22_X1 U14878 ( .A1(n15119), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12687), 
        .B2(n12611), .ZN(n12612) );
  OAI21_X1 U14879 ( .B1(n12792), .B2(n12689), .A(n12612), .ZN(n12613) );
  AOI21_X1 U14880 ( .B1(n12719), .B2(n12691), .A(n12613), .ZN(n12614) );
  OAI21_X1 U14881 ( .B1(n12615), .B2(n15119), .A(n12614), .ZN(P3_U3210) );
  XNOR2_X1 U14882 ( .A(n12616), .B(n12619), .ZN(n12617) );
  OAI222_X1 U14883 ( .A1(n12683), .A2(n12641), .B1(n12759), .B2(n12618), .C1(
        n12680), .C2(n12617), .ZN(n12722) );
  INV_X1 U14884 ( .A(n12722), .ZN(n12625) );
  XNOR2_X1 U14885 ( .A(n12620), .B(n12619), .ZN(n12723) );
  AOI22_X1 U14886 ( .A1(n15119), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12687), 
        .B2(n12621), .ZN(n12622) );
  OAI21_X1 U14887 ( .B1(n12796), .B2(n12689), .A(n12622), .ZN(n12623) );
  AOI21_X1 U14888 ( .B1(n12723), .B2(n12691), .A(n12623), .ZN(n12624) );
  OAI21_X1 U14889 ( .B1(n12625), .B2(n15119), .A(n12624), .ZN(P3_U3211) );
  AOI21_X1 U14890 ( .B1(n12629), .B2(n12626), .A(n6524), .ZN(n12627) );
  OAI222_X1 U14891 ( .A1(n12683), .A2(n12654), .B1(n12759), .B2(n12628), .C1(
        n12680), .C2(n12627), .ZN(n12726) );
  INV_X1 U14892 ( .A(n12726), .ZN(n12636) );
  XOR2_X1 U14893 ( .A(n12630), .B(n12629), .Z(n12727) );
  INV_X1 U14894 ( .A(n12631), .ZN(n12800) );
  AOI22_X1 U14895 ( .A1(n15119), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12687), 
        .B2(n12632), .ZN(n12633) );
  OAI21_X1 U14896 ( .B1(n12800), .B2(n12689), .A(n12633), .ZN(n12634) );
  AOI21_X1 U14897 ( .B1(n12727), .B2(n12691), .A(n12634), .ZN(n12635) );
  OAI21_X1 U14898 ( .B1(n12636), .B2(n15119), .A(n12635), .ZN(P3_U3212) );
  OAI211_X1 U14899 ( .C1(n12638), .C2(n12645), .A(n12637), .B(n12762), .ZN(
        n12640) );
  NAND2_X1 U14900 ( .A1(n12667), .A2(n12756), .ZN(n12639) );
  OAI211_X1 U14901 ( .C1(n12641), .C2(n12759), .A(n12640), .B(n12639), .ZN(
        n12730) );
  INV_X1 U14902 ( .A(n12730), .ZN(n12651) );
  INV_X1 U14903 ( .A(n12642), .ZN(n12643) );
  AOI21_X1 U14904 ( .B1(n12645), .B2(n12644), .A(n12643), .ZN(n12731) );
  INV_X1 U14905 ( .A(n12646), .ZN(n12804) );
  AOI22_X1 U14906 ( .A1(n15119), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n12687), 
        .B2(n12647), .ZN(n12648) );
  OAI21_X1 U14907 ( .B1(n12804), .B2(n12689), .A(n12648), .ZN(n12649) );
  AOI21_X1 U14908 ( .B1(n12731), .B2(n12691), .A(n12649), .ZN(n12650) );
  OAI21_X1 U14909 ( .B1(n12651), .B2(n15119), .A(n12650), .ZN(P3_U3213) );
  OAI211_X1 U14910 ( .C1(n12653), .C2(n12658), .A(n12652), .B(n12762), .ZN(
        n12657) );
  OAI22_X1 U14911 ( .A1(n12654), .A2(n12759), .B1(n12681), .B2(n12683), .ZN(
        n12655) );
  INV_X1 U14912 ( .A(n12655), .ZN(n12656) );
  XNOR2_X1 U14913 ( .A(n12659), .B(n12658), .ZN(n12734) );
  AOI22_X1 U14914 ( .A1(n15119), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12687), 
        .B2(n12660), .ZN(n12661) );
  OAI21_X1 U14915 ( .B1(n12808), .B2(n12689), .A(n12661), .ZN(n12662) );
  AOI21_X1 U14916 ( .B1(n12734), .B2(n12691), .A(n12662), .ZN(n12663) );
  OAI21_X1 U14917 ( .B1(n12736), .B2(n15119), .A(n12663), .ZN(P3_U3214) );
  OAI21_X1 U14918 ( .B1(n12665), .B2(n8661), .A(n12664), .ZN(n12669) );
  AOI222_X1 U14919 ( .A1(n12762), .A2(n12669), .B1(n12668), .B2(n12756), .C1(
        n12667), .C2(n12666), .ZN(n12742) );
  INV_X1 U14920 ( .A(n12670), .ZN(n12671) );
  AOI21_X1 U14921 ( .B1(n8661), .B2(n12672), .A(n12671), .ZN(n12740) );
  INV_X1 U14922 ( .A(n12739), .ZN(n12675) );
  AOI22_X1 U14923 ( .A1(n15119), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n12687), 
        .B2(n12673), .ZN(n12674) );
  OAI21_X1 U14924 ( .B1(n12675), .B2(n12689), .A(n12674), .ZN(n12676) );
  AOI21_X1 U14925 ( .B1(n12740), .B2(n12691), .A(n12676), .ZN(n12677) );
  OAI21_X1 U14926 ( .B1(n12742), .B2(n15119), .A(n12677), .ZN(P3_U3215) );
  XNOR2_X1 U14927 ( .A(n12678), .B(n12685), .ZN(n12679) );
  OAI222_X1 U14928 ( .A1(n12683), .A2(n12682), .B1(n12759), .B2(n12681), .C1(
        n12680), .C2(n12679), .ZN(n12743) );
  INV_X1 U14929 ( .A(n12743), .ZN(n12693) );
  XNOR2_X1 U14930 ( .A(n12684), .B(n12685), .ZN(n12744) );
  AOI22_X1 U14931 ( .A1(n15119), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12687), 
        .B2(n12686), .ZN(n12688) );
  OAI21_X1 U14932 ( .B1(n12813), .B2(n12689), .A(n12688), .ZN(n12690) );
  AOI21_X1 U14933 ( .B1(n12744), .B2(n12691), .A(n12690), .ZN(n12692) );
  OAI21_X1 U14934 ( .B1(n12693), .B2(n15119), .A(n12692), .ZN(P3_U3216) );
  INV_X1 U14935 ( .A(n12773), .ZN(n12696) );
  NAND2_X1 U14936 ( .A1(n15131), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12695) );
  NAND2_X1 U14937 ( .A1(n14466), .A2(n15133), .ZN(n12694) );
  OAI211_X1 U14938 ( .C1(n12696), .C2(n12755), .A(n12695), .B(n12694), .ZN(
        P3_U3490) );
  INV_X1 U14939 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U14940 ( .A1(n12702), .A2(n14475), .B1(n14467), .B2(n12701), .ZN(
        n12703) );
  NAND2_X1 U14941 ( .A1(n12704), .A2(n12703), .ZN(n12779) );
  MUX2_X1 U14942 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12779), .S(n15133), .Z(
        P3_U3486) );
  INV_X1 U14943 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12707) );
  AOI21_X1 U14944 ( .B1(n12706), .B2(n14475), .A(n12705), .ZN(n12780) );
  MUX2_X1 U14945 ( .A(n12707), .B(n12780), .S(n15133), .Z(n12708) );
  OAI21_X1 U14946 ( .B1(n12783), .B2(n12755), .A(n12708), .ZN(P3_U3485) );
  AOI22_X1 U14947 ( .A1(n12710), .A2(n14475), .B1(n14467), .B2(n12709), .ZN(
        n12711) );
  NAND2_X1 U14948 ( .A1(n12712), .A2(n12711), .ZN(n12784) );
  MUX2_X1 U14949 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12784), .S(n15133), .Z(
        P3_U3484) );
  INV_X1 U14950 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12716) );
  INV_X1 U14951 ( .A(n12713), .ZN(n15121) );
  AOI21_X1 U14952 ( .B1(n15121), .B2(n12715), .A(n12714), .ZN(n12785) );
  MUX2_X1 U14953 ( .A(n12716), .B(n12785), .S(n15133), .Z(n12717) );
  OAI21_X1 U14954 ( .B1(n12788), .B2(n12755), .A(n12717), .ZN(P3_U3483) );
  AOI21_X1 U14955 ( .B1(n14475), .B2(n12719), .A(n12718), .ZN(n12789) );
  MUX2_X1 U14956 ( .A(n12720), .B(n12789), .S(n15133), .Z(n12721) );
  OAI21_X1 U14957 ( .B1(n12792), .B2(n12755), .A(n12721), .ZN(P3_U3482) );
  INV_X1 U14958 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12724) );
  AOI21_X1 U14959 ( .B1(n12723), .B2(n14475), .A(n12722), .ZN(n12793) );
  MUX2_X1 U14960 ( .A(n12724), .B(n12793), .S(n15133), .Z(n12725) );
  OAI21_X1 U14961 ( .B1(n12796), .B2(n12755), .A(n12725), .ZN(P3_U3481) );
  INV_X1 U14962 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12728) );
  AOI21_X1 U14963 ( .B1(n14475), .B2(n12727), .A(n12726), .ZN(n12797) );
  MUX2_X1 U14964 ( .A(n12728), .B(n12797), .S(n15133), .Z(n12729) );
  OAI21_X1 U14965 ( .B1(n12800), .B2(n12755), .A(n12729), .ZN(P3_U3480) );
  INV_X1 U14966 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12732) );
  AOI21_X1 U14967 ( .B1(n12731), .B2(n14475), .A(n12730), .ZN(n12801) );
  MUX2_X1 U14968 ( .A(n12732), .B(n12801), .S(n15133), .Z(n12733) );
  OAI21_X1 U14969 ( .B1(n12804), .B2(n12755), .A(n12733), .ZN(P3_U3479) );
  INV_X1 U14970 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12737) );
  NAND2_X1 U14971 ( .A1(n12734), .A2(n14475), .ZN(n12735) );
  MUX2_X1 U14972 ( .A(n12737), .B(n12806), .S(n15133), .Z(n12738) );
  OAI21_X1 U14973 ( .B1(n12755), .B2(n12808), .A(n12738), .ZN(P3_U3478) );
  AOI22_X1 U14974 ( .A1(n12740), .A2(n14475), .B1(n14467), .B2(n12739), .ZN(
        n12741) );
  NAND2_X1 U14975 ( .A1(n12742), .A2(n12741), .ZN(n12809) );
  MUX2_X1 U14976 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12809), .S(n15133), .Z(
        P3_U3477) );
  INV_X1 U14977 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12745) );
  AOI21_X1 U14978 ( .B1(n12744), .B2(n14475), .A(n12743), .ZN(n12810) );
  MUX2_X1 U14979 ( .A(n12745), .B(n12810), .S(n15133), .Z(n12746) );
  OAI21_X1 U14980 ( .B1(n12755), .B2(n12813), .A(n12746), .ZN(P3_U3476) );
  AOI22_X1 U14981 ( .A1(n12748), .A2(n14475), .B1(n14467), .B2(n12747), .ZN(
        n12749) );
  NAND2_X1 U14982 ( .A1(n12750), .A2(n12749), .ZN(n12814) );
  MUX2_X1 U14983 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12814), .S(n15133), .Z(
        P3_U3475) );
  INV_X1 U14984 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12753) );
  AOI21_X1 U14985 ( .B1(n12752), .B2(n14475), .A(n12751), .ZN(n12815) );
  MUX2_X1 U14986 ( .A(n12753), .B(n12815), .S(n15133), .Z(n12754) );
  OAI21_X1 U14987 ( .B1(n12819), .B2(n12755), .A(n12754), .ZN(P3_U3474) );
  XNOR2_X1 U14988 ( .A(n12765), .B(n9263), .ZN(n12763) );
  NAND2_X1 U14989 ( .A1(n12757), .A2(n12756), .ZN(n12758) );
  OAI21_X1 U14990 ( .B1(n12760), .B2(n12759), .A(n12758), .ZN(n12761) );
  AOI21_X1 U14991 ( .B1(n12763), .B2(n12762), .A(n12761), .ZN(n12768) );
  XNOR2_X1 U14992 ( .A(n12765), .B(n12764), .ZN(n15113) );
  OR2_X1 U14993 ( .A1(n15113), .A2(n12766), .ZN(n12767) );
  AND2_X1 U14994 ( .A1(n12768), .A2(n12767), .ZN(n15107) );
  INV_X1 U14995 ( .A(n15113), .ZN(n12770) );
  AND2_X1 U14996 ( .A1(n12769), .A2(n14467), .ZN(n15110) );
  AOI21_X1 U14997 ( .B1(n12770), .B2(n15121), .A(n15110), .ZN(n12771) );
  AND2_X1 U14998 ( .A1(n15107), .A2(n12771), .ZN(n15120) );
  INV_X1 U14999 ( .A(n15120), .ZN(n12772) );
  MUX2_X1 U15000 ( .A(n12772), .B(P3_REG1_REG_1__SCAN_IN), .S(n15131), .Z(
        P3_U3460) );
  NAND2_X1 U15001 ( .A1(n12773), .A2(n8727), .ZN(n12775) );
  NAND2_X1 U15002 ( .A1(n14466), .A2(n15129), .ZN(n12774) );
  OAI211_X1 U15003 ( .C1(n8752), .C2(n15129), .A(n12775), .B(n12774), .ZN(
        P3_U3458) );
  MUX2_X1 U15004 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12779), .S(n15129), .Z(
        P3_U3454) );
  INV_X1 U15005 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12781) );
  MUX2_X1 U15006 ( .A(n12781), .B(n12780), .S(n15129), .Z(n12782) );
  OAI21_X1 U15007 ( .B1(n12783), .B2(n12818), .A(n12782), .ZN(P3_U3453) );
  MUX2_X1 U15008 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12784), .S(n15129), .Z(
        P3_U3452) );
  INV_X1 U15009 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12786) );
  MUX2_X1 U15010 ( .A(n12786), .B(n12785), .S(n15129), .Z(n12787) );
  OAI21_X1 U15011 ( .B1(n12788), .B2(n12818), .A(n12787), .ZN(P3_U3451) );
  INV_X1 U15012 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12790) );
  MUX2_X1 U15013 ( .A(n12790), .B(n12789), .S(n15129), .Z(n12791) );
  OAI21_X1 U15014 ( .B1(n12792), .B2(n12818), .A(n12791), .ZN(P3_U3450) );
  INV_X1 U15015 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12794) );
  MUX2_X1 U15016 ( .A(n12794), .B(n12793), .S(n15129), .Z(n12795) );
  OAI21_X1 U15017 ( .B1(n12796), .B2(n12818), .A(n12795), .ZN(P3_U3449) );
  INV_X1 U15018 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12798) );
  MUX2_X1 U15019 ( .A(n12798), .B(n12797), .S(n15129), .Z(n12799) );
  OAI21_X1 U15020 ( .B1(n12800), .B2(n12818), .A(n12799), .ZN(P3_U3448) );
  INV_X1 U15021 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12802) );
  MUX2_X1 U15022 ( .A(n12802), .B(n12801), .S(n15129), .Z(n12803) );
  OAI21_X1 U15023 ( .B1(n12804), .B2(n12818), .A(n12803), .ZN(P3_U3447) );
  MUX2_X1 U15024 ( .A(n12806), .B(n12805), .S(n15127), .Z(n12807) );
  OAI21_X1 U15025 ( .B1(n12818), .B2(n12808), .A(n12807), .ZN(P3_U3446) );
  MUX2_X1 U15026 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n12809), .S(n15129), .Z(
        P3_U3444) );
  INV_X1 U15027 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12811) );
  MUX2_X1 U15028 ( .A(n12811), .B(n12810), .S(n15129), .Z(n12812) );
  OAI21_X1 U15029 ( .B1(n12818), .B2(n12813), .A(n12812), .ZN(P3_U3441) );
  MUX2_X1 U15030 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n12814), .S(n15129), .Z(
        P3_U3438) );
  INV_X1 U15031 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12816) );
  MUX2_X1 U15032 ( .A(n12816), .B(n12815), .S(n15129), .Z(n12817) );
  OAI21_X1 U15033 ( .B1(n12819), .B2(n12818), .A(n12817), .ZN(P3_U3435) );
  MUX2_X1 U15034 ( .A(n12820), .B(P3_D_REG_1__SCAN_IN), .S(n12821), .Z(
        P3_U3377) );
  MUX2_X1 U15035 ( .A(n12822), .B(P3_D_REG_0__SCAN_IN), .S(n12821), .Z(
        P3_U3376) );
  INV_X1 U15036 ( .A(n12823), .ZN(n12827) );
  INV_X1 U15037 ( .A(n12829), .ZN(n14421) );
  NOR4_X1 U15038 ( .A1(n12824), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), 
        .A4(n8361), .ZN(n12825) );
  AOI21_X1 U15039 ( .B1(n14421), .B2(SI_31_), .A(n12825), .ZN(n12826) );
  OAI21_X1 U15040 ( .B1(n12827), .B2(n12832), .A(n12826), .ZN(P3_U3264) );
  INV_X1 U15041 ( .A(n12828), .ZN(n12831) );
  OAI222_X1 U15042 ( .A1(n12833), .A2(P3_U3151), .B1(n12832), .B2(n12831), 
        .C1(n12830), .C2(n12829), .ZN(P3_U3267) );
  INV_X1 U15043 ( .A(n13320), .ZN(n13168) );
  XNOR2_X1 U15044 ( .A(n13435), .B(n12915), .ZN(n12852) );
  NOR2_X1 U15045 ( .A1(n12835), .A2(n6452), .ZN(n12851) );
  XNOR2_X1 U15046 ( .A(n12852), .B(n12851), .ZN(n13001) );
  OAI21_X1 U15047 ( .B1(n12838), .B2(n12837), .A(n12836), .ZN(n12841) );
  INV_X1 U15048 ( .A(n12838), .ZN(n12840) );
  XNOR2_X1 U15049 ( .A(n13399), .B(n12873), .ZN(n12843) );
  NAND2_X1 U15050 ( .A1(n13036), .A2(n13217), .ZN(n12842) );
  NAND2_X1 U15051 ( .A1(n12843), .A2(n12842), .ZN(n12952) );
  OAI21_X1 U15052 ( .B1(n12843), .B2(n12842), .A(n12952), .ZN(n12946) );
  AND2_X1 U15053 ( .A1(n13035), .A2(n13217), .ZN(n12845) );
  XNOR2_X1 U15054 ( .A(n13439), .B(n12915), .ZN(n12844) );
  NOR2_X1 U15055 ( .A1(n12844), .A2(n12845), .ZN(n12849) );
  AOI21_X1 U15056 ( .B1(n12845), .B2(n12844), .A(n12849), .ZN(n12956) );
  INV_X1 U15057 ( .A(n12956), .ZN(n12846) );
  OR2_X1 U15058 ( .A1(n12846), .A2(n12952), .ZN(n12847) );
  INV_X1 U15059 ( .A(n12849), .ZN(n12850) );
  NAND2_X1 U15060 ( .A1(n12954), .A2(n12850), .ZN(n13002) );
  AND2_X1 U15061 ( .A1(n13033), .A2(n13217), .ZN(n12854) );
  XNOR2_X1 U15062 ( .A(n13277), .B(n12915), .ZN(n12853) );
  NOR2_X1 U15063 ( .A1(n12853), .A2(n12854), .ZN(n12855) );
  AOI21_X1 U15064 ( .B1(n12854), .B2(n12853), .A(n12855), .ZN(n12907) );
  XNOR2_X1 U15065 ( .A(n13367), .B(n12915), .ZN(n12857) );
  AND2_X1 U15066 ( .A1(n13032), .A2(n13217), .ZN(n12856) );
  NOR2_X1 U15067 ( .A1(n12857), .A2(n12856), .ZN(n12976) );
  NAND2_X1 U15068 ( .A1(n12857), .A2(n12856), .ZN(n12977) );
  XNOR2_X1 U15069 ( .A(n13425), .B(n12915), .ZN(n12860) );
  NAND2_X1 U15070 ( .A1(n13031), .A2(n13217), .ZN(n12858) );
  XNOR2_X1 U15071 ( .A(n12860), .B(n12858), .ZN(n12927) );
  XNOR2_X1 U15072 ( .A(n13421), .B(n12873), .ZN(n12991) );
  NAND2_X1 U15073 ( .A1(n13030), .A2(n13217), .ZN(n12863) );
  INV_X1 U15074 ( .A(n12858), .ZN(n12859) );
  NAND2_X1 U15075 ( .A1(n12860), .A2(n12859), .ZN(n12988) );
  INV_X1 U15076 ( .A(n12991), .ZN(n12864) );
  INV_X1 U15077 ( .A(n12863), .ZN(n12990) );
  XNOR2_X1 U15078 ( .A(n13345), .B(n12915), .ZN(n12865) );
  NAND2_X1 U15079 ( .A1(n13029), .A2(n13217), .ZN(n12897) );
  NAND2_X1 U15080 ( .A1(n12896), .A2(n12897), .ZN(n12869) );
  INV_X1 U15081 ( .A(n12865), .ZN(n12866) );
  NAND2_X1 U15082 ( .A1(n12867), .A2(n12866), .ZN(n12868) );
  NAND2_X1 U15083 ( .A1(n12869), .A2(n12868), .ZN(n12966) );
  XNOR2_X1 U15084 ( .A(n6644), .B(n12915), .ZN(n12871) );
  AND2_X1 U15085 ( .A1(n13028), .A2(n13217), .ZN(n12870) );
  NAND2_X1 U15086 ( .A1(n12871), .A2(n12870), .ZN(n12872) );
  OAI21_X1 U15087 ( .B1(n12871), .B2(n12870), .A(n12872), .ZN(n12967) );
  XNOR2_X1 U15088 ( .A(n13193), .B(n12873), .ZN(n12875) );
  NAND2_X1 U15089 ( .A1(n13027), .A2(n12834), .ZN(n12874) );
  NOR2_X1 U15090 ( .A1(n12875), .A2(n12874), .ZN(n12876) );
  AOI21_X1 U15091 ( .B1(n12875), .B2(n12874), .A(n12876), .ZN(n12938) );
  INV_X1 U15092 ( .A(n12876), .ZN(n12877) );
  XNOR2_X1 U15093 ( .A(n13176), .B(n12915), .ZN(n12878) );
  NOR2_X1 U15094 ( .A1(n12890), .A2(n6452), .ZN(n12879) );
  XNOR2_X1 U15095 ( .A(n12878), .B(n12879), .ZN(n13009) );
  INV_X1 U15096 ( .A(n12878), .ZN(n12881) );
  INV_X1 U15097 ( .A(n12879), .ZN(n12880) );
  NAND2_X1 U15098 ( .A1(n12881), .A2(n12880), .ZN(n12886) );
  NAND2_X1 U15099 ( .A1(n13012), .A2(n12886), .ZN(n12884) );
  XNOR2_X1 U15100 ( .A(n13320), .B(n12915), .ZN(n12883) );
  AND2_X1 U15101 ( .A1(n13025), .A2(n13217), .ZN(n12882) );
  NAND2_X1 U15102 ( .A1(n12883), .A2(n12882), .ZN(n12913) );
  OAI21_X1 U15103 ( .B1(n12883), .B2(n12882), .A(n12913), .ZN(n12885) );
  AOI21_X1 U15104 ( .B1(n12884), .B2(n12885), .A(n14490), .ZN(n12889) );
  INV_X1 U15105 ( .A(n12885), .ZN(n12887) );
  AND2_X1 U15106 ( .A1(n12887), .A2(n12886), .ZN(n12888) );
  NAND2_X1 U15107 ( .A1(n12889), .A2(n12914), .ZN(n12895) );
  INV_X1 U15108 ( .A(n13024), .ZN(n12891) );
  OAI22_X1 U15109 ( .A1(n12891), .A2(n12898), .B1(n12890), .B2(n12900), .ZN(
        n13319) );
  OAI22_X1 U15110 ( .A1(n14495), .A2(n13164), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12892), .ZN(n12893) );
  AOI21_X1 U15111 ( .B1(n13319), .B2(n12983), .A(n12893), .ZN(n12894) );
  OAI211_X1 U15112 ( .C1(n13168), .C2(n14488), .A(n12895), .B(n12894), .ZN(
        P2_U3186) );
  XOR2_X1 U15113 ( .A(n12897), .B(n12896), .Z(n12905) );
  OAI22_X1 U15114 ( .A1(n12901), .A2(n12900), .B1(n12899), .B2(n12898), .ZN(
        n13215) );
  AOI22_X1 U15115 ( .A1(n13215), .A2(n12983), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12902) );
  OAI21_X1 U15116 ( .B1(n13222), .B2(n14495), .A(n12902), .ZN(n12903) );
  AOI21_X1 U15117 ( .B1(n13345), .B2(n13014), .A(n12903), .ZN(n12904) );
  OAI21_X1 U15118 ( .B1(n12905), .B2(n14490), .A(n12904), .ZN(P2_U3188) );
  OAI21_X1 U15119 ( .B1(n12908), .B2(n12907), .A(n12906), .ZN(n12909) );
  NAND2_X1 U15120 ( .A1(n12909), .A2(n12957), .ZN(n12912) );
  AOI22_X1 U15121 ( .A1(n14484), .A2(n13034), .B1(n13032), .B2(n14481), .ZN(
        n13280) );
  NAND2_X1 U15122 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13135)
         );
  OAI21_X1 U15123 ( .B1(n13280), .B2(n14491), .A(n13135), .ZN(n12910) );
  AOI21_X1 U15124 ( .B1(n13274), .B2(n13016), .A(n12910), .ZN(n12911) );
  OAI211_X1 U15125 ( .C1(n13432), .C2(n14488), .A(n12912), .B(n12911), .ZN(
        P2_U3191) );
  NAND2_X1 U15126 ( .A1(n12914), .A2(n12913), .ZN(n12919) );
  NAND2_X1 U15127 ( .A1(n13024), .A2(n13217), .ZN(n12916) );
  XNOR2_X1 U15128 ( .A(n12916), .B(n12915), .ZN(n12917) );
  XNOR2_X1 U15129 ( .A(n12919), .B(n12918), .ZN(n12926) );
  NOR2_X1 U15130 ( .A1(n13149), .A2(n14495), .ZN(n12923) );
  OAI22_X1 U15131 ( .A1(n12921), .A2(n14491), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12920), .ZN(n12922) );
  AOI211_X1 U15132 ( .C1(n12924), .C2(n13014), .A(n12923), .B(n12922), .ZN(
        n12925) );
  OAI21_X1 U15133 ( .B1(n12926), .B2(n14490), .A(n12925), .ZN(P2_U3192) );
  INV_X1 U15134 ( .A(n13425), .ZN(n12936) );
  OAI211_X1 U15135 ( .C1(n12928), .C2(n12927), .A(n12989), .B(n12957), .ZN(
        n12935) );
  INV_X1 U15136 ( .A(n13249), .ZN(n12933) );
  NAND2_X1 U15137 ( .A1(n13030), .A2(n13013), .ZN(n12930) );
  NAND2_X1 U15138 ( .A1(n13032), .A2(n14484), .ZN(n12929) );
  AND2_X1 U15139 ( .A1(n12930), .A2(n12929), .ZN(n13358) );
  OAI22_X1 U15140 ( .A1(n13358), .A2(n14491), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12931), .ZN(n12932) );
  AOI21_X1 U15141 ( .B1(n12933), .B2(n13016), .A(n12932), .ZN(n12934) );
  OAI211_X1 U15142 ( .C1(n12936), .C2(n14488), .A(n12935), .B(n12934), .ZN(
        P2_U3195) );
  OAI211_X1 U15143 ( .C1(n12939), .C2(n12938), .A(n12937), .B(n12957), .ZN(
        n12943) );
  AOI22_X1 U15144 ( .A1(n13026), .A2(n14481), .B1(n14484), .B2(n13028), .ZN(
        n13331) );
  OAI22_X1 U15145 ( .A1(n13331), .A2(n14491), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12940), .ZN(n12941) );
  AOI21_X1 U15146 ( .B1(n13190), .B2(n13016), .A(n12941), .ZN(n12942) );
  OAI211_X1 U15147 ( .C1(n8036), .C2(n14488), .A(n12943), .B(n12942), .ZN(
        P2_U3197) );
  OR2_X1 U15148 ( .A1(n12945), .A2(n12946), .ZN(n12953) );
  INV_X1 U15149 ( .A(n12953), .ZN(n12944) );
  AOI21_X1 U15150 ( .B1(n12946), .B2(n12945), .A(n12944), .ZN(n12951) );
  NAND2_X1 U15151 ( .A1(n13397), .A2(n12983), .ZN(n12947) );
  NAND2_X1 U15152 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14922)
         );
  OAI211_X1 U15153 ( .C1(n14495), .C2(n12948), .A(n12947), .B(n14922), .ZN(
        n12949) );
  AOI21_X1 U15154 ( .B1(n13399), .B2(n13014), .A(n12949), .ZN(n12950) );
  OAI21_X1 U15155 ( .B1(n12951), .B2(n14490), .A(n12950), .ZN(P2_U3198) );
  INV_X1 U15156 ( .A(n13439), .ZN(n12965) );
  NAND2_X1 U15157 ( .A1(n12953), .A2(n12952), .ZN(n12955) );
  OAI21_X1 U15158 ( .B1(n12956), .B2(n12955), .A(n12954), .ZN(n12958) );
  NAND2_X1 U15159 ( .A1(n12958), .A2(n12957), .ZN(n12964) );
  INV_X1 U15160 ( .A(n12959), .ZN(n12962) );
  OAI22_X1 U15161 ( .A1(n13389), .A2(n14491), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12960), .ZN(n12961) );
  AOI21_X1 U15162 ( .B1(n12962), .B2(n13016), .A(n12961), .ZN(n12963) );
  OAI211_X1 U15163 ( .C1(n12965), .C2(n14488), .A(n12964), .B(n12963), .ZN(
        P2_U3200) );
  INV_X1 U15164 ( .A(n6644), .ZN(n13206) );
  AOI21_X1 U15165 ( .B1(n12966), .B2(n12967), .A(n14490), .ZN(n12969) );
  NAND2_X1 U15166 ( .A1(n12969), .A2(n12968), .ZN(n12975) );
  NAND2_X1 U15167 ( .A1(n13027), .A2(n13013), .ZN(n12971) );
  NAND2_X1 U15168 ( .A1(n13029), .A2(n14484), .ZN(n12970) );
  NAND2_X1 U15169 ( .A1(n12971), .A2(n12970), .ZN(n13338) );
  OAI22_X1 U15170 ( .A1(n14495), .A2(n13200), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12972), .ZN(n12973) );
  AOI21_X1 U15171 ( .B1(n12983), .B2(n13338), .A(n12973), .ZN(n12974) );
  OAI211_X1 U15172 ( .C1(n13206), .C2(n14488), .A(n12975), .B(n12974), .ZN(
        P2_U3201) );
  INV_X1 U15173 ( .A(n12976), .ZN(n12978) );
  NAND2_X1 U15174 ( .A1(n12978), .A2(n12977), .ZN(n12979) );
  XNOR2_X1 U15175 ( .A(n12980), .B(n12979), .ZN(n12987) );
  NAND2_X1 U15176 ( .A1(n13033), .A2(n14484), .ZN(n12982) );
  NAND2_X1 U15177 ( .A1(n13031), .A2(n13013), .ZN(n12981) );
  NAND2_X1 U15178 ( .A1(n12982), .A2(n12981), .ZN(n13366) );
  AOI22_X1 U15179 ( .A1(n13366), .A2(n12983), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12984) );
  OAI21_X1 U15180 ( .B1(n13263), .B2(n14495), .A(n12984), .ZN(n12985) );
  AOI21_X1 U15181 ( .B1(n13367), .B2(n13014), .A(n12985), .ZN(n12986) );
  OAI21_X1 U15182 ( .B1(n12987), .B2(n14490), .A(n12986), .ZN(P2_U3205) );
  NAND2_X1 U15183 ( .A1(n12989), .A2(n12988), .ZN(n12993) );
  XNOR2_X1 U15184 ( .A(n12991), .B(n12990), .ZN(n12992) );
  XNOR2_X1 U15185 ( .A(n12993), .B(n12992), .ZN(n13000) );
  NAND2_X1 U15186 ( .A1(n13029), .A2(n14481), .ZN(n12995) );
  NAND2_X1 U15187 ( .A1(n13031), .A2(n14484), .ZN(n12994) );
  AND2_X1 U15188 ( .A1(n12995), .A2(n12994), .ZN(n13350) );
  OAI22_X1 U15189 ( .A1(n13350), .A2(n14491), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12996), .ZN(n12998) );
  NOR2_X1 U15190 ( .A1(n13235), .A2(n14488), .ZN(n12997) );
  AOI211_X1 U15191 ( .C1(n13016), .C2(n13236), .A(n12998), .B(n12997), .ZN(
        n12999) );
  OAI21_X1 U15192 ( .B1(n13000), .B2(n14490), .A(n12999), .ZN(P2_U3207) );
  XNOR2_X1 U15193 ( .A(n13002), .B(n13001), .ZN(n13008) );
  NOR2_X1 U15194 ( .A1(n14495), .A2(n13296), .ZN(n13006) );
  NAND2_X1 U15195 ( .A1(n13035), .A2(n14484), .ZN(n13004) );
  NAND2_X1 U15196 ( .A1(n13033), .A2(n14481), .ZN(n13003) );
  AND2_X1 U15197 ( .A1(n13004), .A2(n13003), .ZN(n13382) );
  NAND2_X1 U15198 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13108)
         );
  OAI21_X1 U15199 ( .B1(n13382), .B2(n14491), .A(n13108), .ZN(n13005) );
  AOI211_X1 U15200 ( .C1(n13435), .C2(n13014), .A(n13006), .B(n13005), .ZN(
        n13007) );
  OAI21_X1 U15201 ( .B1(n13008), .B2(n14490), .A(n13007), .ZN(P2_U3210) );
  NAND2_X1 U15202 ( .A1(n13010), .A2(n13009), .ZN(n13011) );
  AOI21_X1 U15203 ( .B1(n13012), .B2(n13011), .A(n14490), .ZN(n13020) );
  AOI22_X1 U15204 ( .A1(n13025), .A2(n13013), .B1(n14484), .B2(n13027), .ZN(
        n13324) );
  NAND2_X1 U15205 ( .A1(n13176), .A2(n13014), .ZN(n13018) );
  INV_X1 U15206 ( .A(n13015), .ZN(n13177) );
  AOI22_X1 U15207 ( .A1(n13016), .A2(n13177), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13017) );
  OAI211_X1 U15208 ( .C1(n13324), .C2(n14491), .A(n13018), .B(n13017), .ZN(
        n13019) );
  OR2_X1 U15209 ( .A1(n13020), .A2(n13019), .ZN(P2_U3212) );
  INV_X2 U15210 ( .A(P2_U3947), .ZN(n13049) );
  MUX2_X1 U15211 ( .A(n13021), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13049), .Z(
        P2_U3562) );
  MUX2_X1 U15212 ( .A(n13022), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13049), .Z(
        P2_U3561) );
  MUX2_X1 U15213 ( .A(n13023), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13049), .Z(
        P2_U3560) );
  MUX2_X1 U15214 ( .A(n13024), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13049), .Z(
        P2_U3559) );
  MUX2_X1 U15215 ( .A(n13025), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13049), .Z(
        P2_U3558) );
  MUX2_X1 U15216 ( .A(n13026), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13049), .Z(
        P2_U3557) );
  MUX2_X1 U15217 ( .A(n13027), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13049), .Z(
        P2_U3556) );
  MUX2_X1 U15218 ( .A(n13028), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13049), .Z(
        P2_U3555) );
  MUX2_X1 U15219 ( .A(n13029), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13049), .Z(
        P2_U3554) );
  MUX2_X1 U15220 ( .A(n13030), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13049), .Z(
        P2_U3553) );
  MUX2_X1 U15221 ( .A(n13031), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13049), .Z(
        P2_U3552) );
  MUX2_X1 U15222 ( .A(n13032), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13049), .Z(
        P2_U3551) );
  MUX2_X1 U15223 ( .A(n13033), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13049), .Z(
        P2_U3550) );
  MUX2_X1 U15224 ( .A(n13034), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13049), .Z(
        P2_U3549) );
  MUX2_X1 U15225 ( .A(n13035), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13049), .Z(
        P2_U3548) );
  MUX2_X1 U15226 ( .A(n13036), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13049), .Z(
        P2_U3547) );
  MUX2_X1 U15227 ( .A(n14482), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13049), .Z(
        P2_U3546) );
  MUX2_X1 U15228 ( .A(n13037), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13049), .Z(
        P2_U3545) );
  MUX2_X1 U15229 ( .A(n14483), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13049), .Z(
        P2_U3544) );
  MUX2_X1 U15230 ( .A(n13038), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13049), .Z(
        P2_U3543) );
  MUX2_X1 U15231 ( .A(n13039), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13049), .Z(
        P2_U3542) );
  MUX2_X1 U15232 ( .A(n13040), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13049), .Z(
        P2_U3541) );
  MUX2_X1 U15233 ( .A(n13041), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13049), .Z(
        P2_U3540) );
  MUX2_X1 U15234 ( .A(n13042), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13049), .Z(
        P2_U3539) );
  MUX2_X1 U15235 ( .A(n13043), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13049), .Z(
        P2_U3538) );
  MUX2_X1 U15236 ( .A(n13044), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13049), .Z(
        P2_U3537) );
  MUX2_X1 U15237 ( .A(n13045), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13049), .Z(
        P2_U3536) );
  MUX2_X1 U15238 ( .A(n13046), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13049), .Z(
        P2_U3535) );
  MUX2_X1 U15239 ( .A(n13047), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13049), .Z(
        P2_U3534) );
  MUX2_X1 U15240 ( .A(n8973), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13049), .Z(
        P2_U3533) );
  MUX2_X1 U15241 ( .A(n13048), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13049), .Z(
        P2_U3532) );
  MUX2_X1 U15242 ( .A(n8960), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13049), .Z(
        P2_U3531) );
  NOR2_X1 U15243 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13050), .ZN(n13053) );
  NOR2_X1 U15244 ( .A1(n14937), .A2(n13051), .ZN(n13052) );
  AOI211_X1 U15245 ( .C1(n14929), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n13053), .B(
        n13052), .ZN(n13064) );
  OAI211_X1 U15246 ( .C1(n13056), .C2(n13055), .A(n14900), .B(n13054), .ZN(
        n13063) );
  INV_X1 U15247 ( .A(n13057), .ZN(n13061) );
  NAND3_X1 U15248 ( .A1(n14833), .A2(n13059), .A3(n13058), .ZN(n13060) );
  NAND3_X1 U15249 ( .A1(n14931), .A2(n13061), .A3(n13060), .ZN(n13062) );
  NAND3_X1 U15250 ( .A1(n13064), .A2(n13063), .A3(n13062), .ZN(P2_U3217) );
  INV_X1 U15251 ( .A(n13065), .ZN(n13067) );
  NOR2_X1 U15252 ( .A1(n14937), .A2(n13071), .ZN(n13066) );
  AOI211_X1 U15253 ( .C1(n14929), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n13067), .B(
        n13066), .ZN(n13080) );
  OAI211_X1 U15254 ( .C1(n13070), .C2(n13069), .A(n14900), .B(n13068), .ZN(
        n13079) );
  MUX2_X1 U15255 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n13072), .S(n13071), .Z(
        n13075) );
  INV_X1 U15256 ( .A(n13073), .ZN(n13074) );
  NAND2_X1 U15257 ( .A1(n13075), .A2(n13074), .ZN(n13077) );
  OAI211_X1 U15258 ( .C1(n14863), .C2(n13077), .A(n14931), .B(n13076), .ZN(
        n13078) );
  NAND3_X1 U15259 ( .A1(n13080), .A2(n13079), .A3(n13078), .ZN(P2_U3220) );
  AOI21_X1 U15260 ( .B1(n13093), .B2(P2_REG1_REG_14__SCAN_IN), .A(n13081), 
        .ZN(n13082) );
  NOR2_X1 U15261 ( .A1(n13082), .A2(n14921), .ZN(n13083) );
  XNOR2_X1 U15262 ( .A(n14921), .B(n13082), .ZN(n14914) );
  NOR2_X1 U15263 ( .A1(n14913), .A2(n14914), .ZN(n14912) );
  NOR2_X1 U15264 ( .A1(n13083), .A2(n14912), .ZN(n14926) );
  XNOR2_X1 U15265 ( .A(n13084), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14925) );
  NOR2_X1 U15266 ( .A1(n14926), .A2(n14925), .ZN(n14924) );
  AOI21_X1 U15267 ( .B1(n13084), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14924), 
        .ZN(n13086) );
  XNOR2_X1 U15268 ( .A(n13110), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n13085) );
  NOR2_X1 U15269 ( .A1(n13086), .A2(n13085), .ZN(n13109) );
  AOI211_X1 U15270 ( .C1(n13086), .C2(n13085), .A(n13109), .B(n14923), .ZN(
        n13087) );
  INV_X1 U15271 ( .A(n13087), .ZN(n13104) );
  AND2_X1 U15272 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13089) );
  NOR2_X1 U15273 ( .A1(n14937), .A2(n13106), .ZN(n13088) );
  AOI211_X1 U15274 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n14929), .A(n13089), 
        .B(n13088), .ZN(n13103) );
  NOR2_X1 U15275 ( .A1(n13106), .A2(n13090), .ZN(n13091) );
  AOI21_X1 U15276 ( .B1(n13090), .B2(n13106), .A(n13091), .ZN(n13101) );
  INV_X1 U15277 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13099) );
  XNOR2_X1 U15278 ( .A(n14936), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n14932) );
  NAND2_X1 U15279 ( .A1(n13093), .A2(n13092), .ZN(n13095) );
  NAND2_X1 U15280 ( .A1(n13095), .A2(n13094), .ZN(n13097) );
  NAND2_X1 U15281 ( .A1(n13096), .A2(n13097), .ZN(n13098) );
  XNOR2_X1 U15282 ( .A(n13097), .B(n14921), .ZN(n14918) );
  NAND2_X1 U15283 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14918), .ZN(n14917) );
  NAND2_X1 U15284 ( .A1(n13098), .A2(n14917), .ZN(n14933) );
  NAND2_X1 U15285 ( .A1(n14932), .A2(n14933), .ZN(n14930) );
  OAI211_X1 U15286 ( .C1(n13101), .C2(n13100), .A(n14931), .B(n13105), .ZN(
        n13102) );
  NAND3_X1 U15287 ( .A1(n13104), .A2(n13103), .A3(n13102), .ZN(P2_U3231) );
  OAI21_X1 U15288 ( .B1(n13090), .B2(n13106), .A(n13105), .ZN(n13123) );
  XNOR2_X1 U15289 ( .A(n13124), .B(n13123), .ZN(n13107) );
  AOI21_X1 U15290 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13107), .A(n13126), 
        .ZN(n13117) );
  OAI21_X1 U15291 ( .B1(n14937), .B2(n13118), .A(n13108), .ZN(n13115) );
  AOI21_X1 U15292 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n13110), .A(n13109), 
        .ZN(n13119) );
  INV_X1 U15293 ( .A(n13119), .ZN(n13111) );
  XNOR2_X1 U15294 ( .A(n13124), .B(n13111), .ZN(n13113) );
  INV_X1 U15295 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13112) );
  NOR2_X1 U15296 ( .A1(n13112), .A2(n13113), .ZN(n13121) );
  AOI211_X1 U15297 ( .C1(n13113), .C2(n13112), .A(n13121), .B(n14923), .ZN(
        n13114) );
  AOI211_X1 U15298 ( .C1(n14929), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13115), 
        .B(n13114), .ZN(n13116) );
  OAI21_X1 U15299 ( .B1(n13117), .B2(n14862), .A(n13116), .ZN(P2_U3232) );
  NOR2_X1 U15300 ( .A1(n13119), .A2(n13118), .ZN(n13120) );
  NOR2_X1 U15301 ( .A1(n13121), .A2(n13120), .ZN(n13122) );
  XOR2_X1 U15302 ( .A(n13122), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13132) );
  NOR2_X1 U15303 ( .A1(n13124), .A2(n13123), .ZN(n13125) );
  NOR2_X1 U15304 ( .A1(n13126), .A2(n13125), .ZN(n13128) );
  XOR2_X1 U15305 ( .A(n13128), .B(n13127), .Z(n13130) );
  OAI22_X1 U15306 ( .A1(n13132), .A2(n14923), .B1(n13130), .B2(n14862), .ZN(
        n13129) );
  INV_X1 U15307 ( .A(n13129), .ZN(n13134) );
  AND2_X1 U15308 ( .A1(n13130), .A2(n14931), .ZN(n13131) );
  AOI211_X1 U15309 ( .C1(n13132), .C2(n14900), .A(n14889), .B(n13131), .ZN(
        n13133) );
  MUX2_X1 U15310 ( .A(n13134), .B(n13133), .S(n6463), .Z(n13136) );
  OAI211_X1 U15311 ( .C1(n13137), .C2(n14897), .A(n13136), .B(n13135), .ZN(
        P2_U3233) );
  NOR2_X1 U15312 ( .A1(n14951), .A2(n13307), .ZN(n13145) );
  AOI21_X1 U15313 ( .B1(n14951), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13145), 
        .ZN(n13140) );
  NAND2_X1 U15314 ( .A1(n13138), .A2(n14502), .ZN(n13139) );
  OAI211_X1 U15315 ( .C1(n13141), .C2(n13302), .A(n13140), .B(n13139), .ZN(
        P2_U3234) );
  NAND2_X1 U15316 ( .A1(n13408), .A2(n13142), .ZN(n13143) );
  NAND3_X1 U15317 ( .A1(n13144), .A2(n6452), .A3(n13143), .ZN(n13308) );
  AOI21_X1 U15318 ( .B1(n14951), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13145), 
        .ZN(n13147) );
  NAND2_X1 U15319 ( .A1(n13408), .A2(n14502), .ZN(n13146) );
  OAI211_X1 U15320 ( .C1(n13308), .C2(n13302), .A(n13147), .B(n13146), .ZN(
        P2_U3235) );
  OAI21_X1 U15321 ( .B1(n13149), .B2(n13295), .A(n13148), .ZN(n13150) );
  NAND2_X1 U15322 ( .A1(n13150), .A2(n14948), .ZN(n13156) );
  INV_X1 U15323 ( .A(n13151), .ZN(n13154) );
  INV_X1 U15324 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13152) );
  OAI22_X1 U15325 ( .A1(n13413), .A2(n13205), .B1(n14948), .B2(n13152), .ZN(
        n13153) );
  AOI21_X1 U15326 ( .B1(n13154), .B2(n14509), .A(n13153), .ZN(n13155) );
  OAI211_X1 U15327 ( .C1(n13157), .C2(n13224), .A(n13156), .B(n13155), .ZN(
        P2_U3237) );
  XNOR2_X1 U15328 ( .A(n13159), .B(n13158), .ZN(n13323) );
  NAND2_X1 U15329 ( .A1(n13160), .A2(n6908), .ZN(n13316) );
  NAND3_X1 U15330 ( .A1(n13317), .A2(n13316), .A3(n14510), .ZN(n13171) );
  NAND2_X1 U15331 ( .A1(n13320), .A2(n13174), .ZN(n13161) );
  NAND2_X1 U15332 ( .A1(n13161), .A2(n6452), .ZN(n13162) );
  NOR2_X1 U15333 ( .A1(n13163), .A2(n13162), .ZN(n13318) );
  INV_X1 U15334 ( .A(n13164), .ZN(n13165) );
  AOI22_X1 U15335 ( .A1(n13165), .A2(n14941), .B1(n14951), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n13167) );
  NAND2_X1 U15336 ( .A1(n13319), .A2(n14948), .ZN(n13166) );
  OAI211_X1 U15337 ( .C1(n13168), .C2(n13205), .A(n13167), .B(n13166), .ZN(
        n13169) );
  AOI21_X1 U15338 ( .B1(n13318), .B2(n14509), .A(n13169), .ZN(n13170) );
  OAI211_X1 U15339 ( .C1(n13323), .C2(n13305), .A(n13171), .B(n13170), .ZN(
        P2_U3238) );
  XNOR2_X1 U15340 ( .A(n13172), .B(n13173), .ZN(n13330) );
  INV_X1 U15341 ( .A(n13174), .ZN(n13175) );
  AOI211_X1 U15342 ( .C1(n13176), .C2(n13189), .A(n13217), .B(n13175), .ZN(
        n13327) );
  INV_X1 U15343 ( .A(n13176), .ZN(n13325) );
  NOR2_X1 U15344 ( .A1(n13325), .A2(n13205), .ZN(n13180) );
  AOI22_X1 U15345 ( .A1(n14951), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13177), 
        .B2(n14941), .ZN(n13178) );
  OAI21_X1 U15346 ( .B1(n13324), .B2(n14951), .A(n13178), .ZN(n13179) );
  AOI211_X1 U15347 ( .C1(n13327), .C2(n14509), .A(n13180), .B(n13179), .ZN(
        n13184) );
  XNOR2_X1 U15348 ( .A(n13182), .B(n13181), .ZN(n13328) );
  NAND2_X1 U15349 ( .A1(n13328), .A2(n13212), .ZN(n13183) );
  OAI211_X1 U15350 ( .C1(n13330), .C2(n13224), .A(n13184), .B(n13183), .ZN(
        P2_U3239) );
  XOR2_X1 U15351 ( .A(n13185), .B(n13186), .Z(n13336) );
  XNOR2_X1 U15352 ( .A(n13187), .B(n13186), .ZN(n13334) );
  OAI211_X1 U15353 ( .C1(n8036), .C2(n13188), .A(n6452), .B(n13189), .ZN(
        n13332) );
  AOI22_X1 U15354 ( .A1(n14951), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13190), 
        .B2(n14941), .ZN(n13191) );
  OAI21_X1 U15355 ( .B1(n13331), .B2(n14951), .A(n13191), .ZN(n13192) );
  AOI21_X1 U15356 ( .B1(n13193), .B2(n14502), .A(n13192), .ZN(n13194) );
  OAI21_X1 U15357 ( .B1(n13332), .B2(n13302), .A(n13194), .ZN(n13195) );
  AOI21_X1 U15358 ( .B1(n13334), .B2(n13212), .A(n13195), .ZN(n13196) );
  OAI21_X1 U15359 ( .B1(n13336), .B2(n13224), .A(n13196), .ZN(P2_U3240) );
  XNOR2_X1 U15360 ( .A(n13198), .B(n13197), .ZN(n13340) );
  AOI21_X1 U15361 ( .B1(n6644), .B2(n13218), .A(n13217), .ZN(n13199) );
  AND2_X1 U15362 ( .A1(n13199), .A2(n6871), .ZN(n13337) );
  NAND2_X1 U15363 ( .A1(n13337), .A2(n14509), .ZN(n13204) );
  INV_X1 U15364 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13201) );
  OAI22_X1 U15365 ( .A1(n14948), .A2(n13201), .B1(n13200), .B2(n13295), .ZN(
        n13202) );
  AOI21_X1 U15366 ( .B1(n13338), .B2(n13298), .A(n13202), .ZN(n13203) );
  OAI211_X1 U15367 ( .C1(n13206), .C2(n13205), .A(n13204), .B(n13203), .ZN(
        n13211) );
  OAI21_X1 U15368 ( .B1(n13209), .B2(n13208), .A(n13207), .ZN(n13343) );
  NOR2_X1 U15369 ( .A1(n13343), .A2(n13224), .ZN(n13210) );
  AOI211_X1 U15370 ( .C1(n13212), .C2(n13340), .A(n13211), .B(n13210), .ZN(
        n13213) );
  INV_X1 U15371 ( .A(n13213), .ZN(P2_U3241) );
  XNOR2_X1 U15372 ( .A(n13214), .B(n13223), .ZN(n13216) );
  AOI21_X1 U15373 ( .B1(n13216), .B2(n14535), .A(n13215), .ZN(n13347) );
  AOI21_X1 U15374 ( .B1(n13234), .B2(n13345), .A(n13217), .ZN(n13219) );
  AND2_X1 U15375 ( .A1(n13219), .A2(n13218), .ZN(n13344) );
  NAND2_X1 U15376 ( .A1(n13345), .A2(n14502), .ZN(n13221) );
  NAND2_X1 U15377 ( .A1(n14951), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n13220) );
  OAI211_X1 U15378 ( .C1(n13295), .C2(n13222), .A(n13221), .B(n13220), .ZN(
        n13226) );
  XNOR2_X1 U15379 ( .A(n6570), .B(n13223), .ZN(n13348) );
  NOR2_X1 U15380 ( .A1(n13348), .A2(n13224), .ZN(n13225) );
  AOI211_X1 U15381 ( .C1(n13344), .C2(n14509), .A(n13226), .B(n13225), .ZN(
        n13227) );
  OAI21_X1 U15382 ( .B1(n14951), .B2(n13347), .A(n13227), .ZN(P2_U3242) );
  XNOR2_X1 U15383 ( .A(n13229), .B(n13228), .ZN(n13354) );
  NAND2_X1 U15384 ( .A1(n13231), .A2(n13232), .ZN(n13233) );
  NAND2_X1 U15385 ( .A1(n13230), .A2(n13233), .ZN(n13349) );
  INV_X1 U15386 ( .A(n13349), .ZN(n13242) );
  OAI211_X1 U15387 ( .C1(n13235), .C2(n13248), .A(n6452), .B(n13234), .ZN(
        n13351) );
  NAND2_X1 U15388 ( .A1(n14941), .A2(n13236), .ZN(n13238) );
  NAND2_X1 U15389 ( .A1(n14951), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n13237) );
  OAI211_X1 U15390 ( .C1(n13350), .C2(n14951), .A(n13238), .B(n13237), .ZN(
        n13239) );
  AOI21_X1 U15391 ( .B1(n13421), .B2(n14502), .A(n13239), .ZN(n13240) );
  OAI21_X1 U15392 ( .B1(n13351), .B2(n13302), .A(n13240), .ZN(n13241) );
  AOI21_X1 U15393 ( .B1(n13242), .B2(n14510), .A(n13241), .ZN(n13243) );
  OAI21_X1 U15394 ( .B1(n13354), .B2(n13305), .A(n13243), .ZN(P2_U3243) );
  XNOR2_X1 U15395 ( .A(n13244), .B(n13245), .ZN(n13357) );
  NAND2_X1 U15396 ( .A1(n13261), .A2(n13425), .ZN(n13246) );
  NAND2_X1 U15397 ( .A1(n13246), .A2(n6452), .ZN(n13247) );
  OR2_X1 U15398 ( .A1(n13248), .A2(n13247), .ZN(n13359) );
  INV_X1 U15399 ( .A(n13358), .ZN(n13252) );
  INV_X1 U15400 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13250) );
  OAI22_X1 U15401 ( .A1(n14948), .A2(n13250), .B1(n13249), .B2(n13295), .ZN(
        n13251) );
  AOI21_X1 U15402 ( .B1(n13252), .B2(n13298), .A(n13251), .ZN(n13254) );
  NAND2_X1 U15403 ( .A1(n13425), .A2(n14502), .ZN(n13253) );
  OAI211_X1 U15404 ( .C1(n13359), .C2(n13302), .A(n13254), .B(n13253), .ZN(
        n13258) );
  XNOR2_X1 U15405 ( .A(n13256), .B(n13255), .ZN(n13362) );
  NOR2_X1 U15406 ( .A1(n13362), .A2(n13305), .ZN(n13257) );
  AOI211_X1 U15407 ( .C1(n14510), .C2(n13357), .A(n13258), .B(n13257), .ZN(
        n13259) );
  INV_X1 U15408 ( .A(n13259), .ZN(P2_U3244) );
  XOR2_X1 U15409 ( .A(n13260), .B(n13270), .Z(n13372) );
  AOI21_X1 U15410 ( .B1(n6587), .B2(n13367), .A(n13217), .ZN(n13262) );
  AND2_X1 U15411 ( .A1(n13262), .A2(n13261), .ZN(n13365) );
  NAND2_X1 U15412 ( .A1(n13367), .A2(n14502), .ZN(n13267) );
  INV_X1 U15413 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13264) );
  OAI22_X1 U15414 ( .A1(n13298), .A2(n13264), .B1(n13263), .B2(n13295), .ZN(
        n13265) );
  AOI21_X1 U15415 ( .B1(n13366), .B2(n13298), .A(n13265), .ZN(n13266) );
  NAND2_X1 U15416 ( .A1(n13267), .A2(n13266), .ZN(n13268) );
  AOI21_X1 U15417 ( .B1(n13365), .B2(n14509), .A(n13268), .ZN(n13272) );
  XNOR2_X1 U15418 ( .A(n13269), .B(n13270), .ZN(n13368) );
  NAND2_X1 U15419 ( .A1(n13368), .A2(n14510), .ZN(n13271) );
  OAI211_X1 U15420 ( .C1(n13372), .C2(n13305), .A(n13272), .B(n13271), .ZN(
        P2_U3245) );
  XOR2_X1 U15421 ( .A(n13273), .B(n13278), .Z(n13375) );
  NAND2_X1 U15422 ( .A1(n13375), .A2(n14510), .ZN(n13286) );
  INV_X1 U15423 ( .A(n13274), .ZN(n13275) );
  OAI22_X1 U15424 ( .A1(n14948), .A2(n13127), .B1(n13275), .B2(n13295), .ZN(
        n13276) );
  AOI21_X1 U15425 ( .B1(n13277), .B2(n14502), .A(n13276), .ZN(n13285) );
  XNOR2_X1 U15426 ( .A(n13279), .B(n13278), .ZN(n13281) );
  OAI21_X1 U15427 ( .B1(n13281), .B2(n13371), .A(n13280), .ZN(n13373) );
  NAND2_X1 U15428 ( .A1(n13373), .A2(n14948), .ZN(n13284) );
  OR2_X1 U15429 ( .A1(n13293), .A2(n13432), .ZN(n13282) );
  AND3_X1 U15430 ( .A1(n6587), .A2(n6452), .A3(n13282), .ZN(n13374) );
  NAND2_X1 U15431 ( .A1(n13374), .A2(n14509), .ZN(n13283) );
  NAND4_X1 U15432 ( .A1(n13286), .A2(n13285), .A3(n13284), .A4(n13283), .ZN(
        P2_U3246) );
  XNOR2_X1 U15433 ( .A(n13287), .B(n13289), .ZN(n13379) );
  INV_X1 U15434 ( .A(n13379), .ZN(n13306) );
  OAI21_X1 U15435 ( .B1(n13290), .B2(n13289), .A(n13288), .ZN(n13380) );
  OAI21_X1 U15436 ( .B1(n13292), .B2(n13291), .A(n6452), .ZN(n13294) );
  OR2_X1 U15437 ( .A1(n13294), .A2(n13293), .ZN(n13381) );
  NOR2_X1 U15438 ( .A1(n13382), .A2(n14951), .ZN(n13300) );
  INV_X1 U15439 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13297) );
  OAI22_X1 U15440 ( .A1(n13298), .A2(n13297), .B1(n13296), .B2(n13295), .ZN(
        n13299) );
  AOI211_X1 U15441 ( .C1(n13435), .C2(n14502), .A(n13300), .B(n13299), .ZN(
        n13301) );
  OAI21_X1 U15442 ( .B1(n13381), .B2(n13302), .A(n13301), .ZN(n13303) );
  AOI21_X1 U15443 ( .B1(n13380), .B2(n14510), .A(n13303), .ZN(n13304) );
  OAI21_X1 U15444 ( .B1(n13306), .B2(n13305), .A(n13304), .ZN(P2_U3247) );
  NAND2_X1 U15445 ( .A1(n13308), .A2(n13307), .ZN(n13406) );
  MUX2_X1 U15446 ( .A(n13406), .B(P2_REG1_REG_30__SCAN_IN), .S(n14999), .Z(
        n13309) );
  AOI21_X1 U15447 ( .B1(n8070), .B2(n13408), .A(n13309), .ZN(n13310) );
  INV_X1 U15448 ( .A(n13310), .ZN(P2_U3529) );
  NAND3_X1 U15449 ( .A1(n13317), .A2(n14983), .A3(n13316), .ZN(n13322) );
  AOI211_X1 U15450 ( .C1(n13398), .C2(n13320), .A(n13319), .B(n13318), .ZN(
        n13321) );
  OAI211_X1 U15451 ( .C1(n13371), .C2(n13323), .A(n13322), .B(n13321), .ZN(
        n13414) );
  MUX2_X1 U15452 ( .A(n13414), .B(P2_REG1_REG_27__SCAN_IN), .S(n14999), .Z(
        P2_U3526) );
  INV_X1 U15453 ( .A(n13398), .ZN(n14986) );
  OAI21_X1 U15454 ( .B1(n13325), .B2(n14986), .A(n13324), .ZN(n13326) );
  AOI211_X1 U15455 ( .C1(n13328), .C2(n14535), .A(n13327), .B(n13326), .ZN(
        n13329) );
  OAI21_X1 U15456 ( .B1(n13330), .B2(n14530), .A(n13329), .ZN(n13415) );
  MUX2_X1 U15457 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13415), .S(n15002), .Z(
        P2_U3525) );
  OAI211_X1 U15458 ( .C1(n8036), .C2(n14986), .A(n13332), .B(n13331), .ZN(
        n13333) );
  AOI21_X1 U15459 ( .B1(n13334), .B2(n14535), .A(n13333), .ZN(n13335) );
  OAI21_X1 U15460 ( .B1(n13336), .B2(n14530), .A(n13335), .ZN(n13416) );
  MUX2_X1 U15461 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13416), .S(n15002), .Z(
        P2_U3524) );
  AOI211_X1 U15462 ( .C1(n13398), .C2(n6644), .A(n13338), .B(n13337), .ZN(
        n13342) );
  NAND2_X1 U15463 ( .A1(n13340), .A2(n14535), .ZN(n13341) );
  OAI211_X1 U15464 ( .C1(n13343), .C2(n14530), .A(n13342), .B(n13341), .ZN(
        n13417) );
  MUX2_X1 U15465 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13417), .S(n15002), .Z(
        P2_U3523) );
  AOI21_X1 U15466 ( .B1(n13398), .B2(n13345), .A(n13344), .ZN(n13346) );
  OAI211_X1 U15467 ( .C1(n13348), .C2(n14530), .A(n13347), .B(n13346), .ZN(
        n13418) );
  MUX2_X1 U15468 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13418), .S(n15002), .Z(
        P2_U3522) );
  OR2_X1 U15469 ( .A1(n13349), .A2(n14530), .ZN(n13353) );
  AND2_X1 U15470 ( .A1(n13351), .A2(n13350), .ZN(n13352) );
  OAI211_X1 U15471 ( .C1(n13371), .C2(n13354), .A(n13353), .B(n13352), .ZN(
        n13419) );
  MUX2_X1 U15472 ( .A(n13419), .B(P2_REG1_REG_22__SCAN_IN), .S(n14999), .Z(
        n13355) );
  AOI21_X1 U15473 ( .B1(n8070), .B2(n13421), .A(n13355), .ZN(n13356) );
  INV_X1 U15474 ( .A(n13356), .ZN(P2_U3521) );
  NAND2_X1 U15475 ( .A1(n13357), .A2(n14983), .ZN(n13361) );
  AND2_X1 U15476 ( .A1(n13359), .A2(n13358), .ZN(n13360) );
  OAI211_X1 U15477 ( .C1(n13362), .C2(n13371), .A(n13361), .B(n13360), .ZN(
        n13423) );
  MUX2_X1 U15478 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13423), .S(n15002), .Z(
        n13363) );
  AOI21_X1 U15479 ( .B1(n8070), .B2(n13425), .A(n13363), .ZN(n13364) );
  INV_X1 U15480 ( .A(n13364), .ZN(P2_U3520) );
  AOI211_X1 U15481 ( .C1(n13398), .C2(n13367), .A(n13366), .B(n13365), .ZN(
        n13370) );
  NAND2_X1 U15482 ( .A1(n13368), .A2(n14983), .ZN(n13369) );
  OAI211_X1 U15483 ( .C1(n13372), .C2(n13371), .A(n13370), .B(n13369), .ZN(
        n13427) );
  MUX2_X1 U15484 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13427), .S(n15002), .Z(
        P2_U3519) );
  INV_X1 U15485 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13376) );
  AOI211_X1 U15486 ( .C1(n13375), .C2(n14983), .A(n13374), .B(n13373), .ZN(
        n13428) );
  MUX2_X1 U15487 ( .A(n13376), .B(n13428), .S(n15002), .Z(n13377) );
  OAI21_X1 U15488 ( .B1(n13432), .B2(n13378), .A(n13377), .ZN(P2_U3518) );
  NAND2_X1 U15489 ( .A1(n13379), .A2(n14535), .ZN(n13384) );
  NAND2_X1 U15490 ( .A1(n13380), .A2(n14983), .ZN(n13383) );
  NAND4_X1 U15491 ( .A1(n13384), .A2(n13383), .A3(n13382), .A4(n13381), .ZN(
        n13433) );
  MUX2_X1 U15492 ( .A(n13433), .B(P2_REG1_REG_18__SCAN_IN), .S(n14999), .Z(
        n13385) );
  AOI21_X1 U15493 ( .B1(n8070), .B2(n13435), .A(n13385), .ZN(n13386) );
  INV_X1 U15494 ( .A(n13386), .ZN(P2_U3517) );
  NAND2_X1 U15495 ( .A1(n13387), .A2(n14983), .ZN(n13393) );
  NAND2_X1 U15496 ( .A1(n13388), .A2(n14535), .ZN(n13392) );
  AND2_X1 U15497 ( .A1(n13390), .A2(n13389), .ZN(n13391) );
  NAND3_X1 U15498 ( .A1(n13393), .A2(n13392), .A3(n13391), .ZN(n13437) );
  MUX2_X1 U15499 ( .A(n13437), .B(P2_REG1_REG_17__SCAN_IN), .S(n14999), .Z(
        n13394) );
  AOI21_X1 U15500 ( .B1(n8070), .B2(n13439), .A(n13394), .ZN(n13395) );
  INV_X1 U15501 ( .A(n13395), .ZN(P2_U3516) );
  NAND2_X1 U15502 ( .A1(n13396), .A2(n14535), .ZN(n13405) );
  AOI21_X1 U15503 ( .B1(n13399), .B2(n13398), .A(n13397), .ZN(n13404) );
  NAND3_X1 U15504 ( .A1(n13401), .A2(n13400), .A3(n14983), .ZN(n13403) );
  NAND4_X1 U15505 ( .A1(n13405), .A2(n13404), .A3(n13403), .A4(n13402), .ZN(
        n13442) );
  MUX2_X1 U15506 ( .A(n13442), .B(P2_REG1_REG_16__SCAN_IN), .S(n14999), .Z(
        P2_U3515) );
  MUX2_X1 U15507 ( .A(n13406), .B(P2_REG0_REG_30__SCAN_IN), .S(n14991), .Z(
        n13407) );
  AOI21_X1 U15508 ( .B1(n13440), .B2(n13408), .A(n13407), .ZN(n13409) );
  INV_X1 U15509 ( .A(n13409), .ZN(P2_U3497) );
  OAI21_X1 U15510 ( .B1(n13413), .B2(n13431), .A(n13412), .ZN(P2_U3495) );
  MUX2_X1 U15511 ( .A(n13414), .B(P2_REG0_REG_27__SCAN_IN), .S(n14991), .Z(
        P2_U3494) );
  MUX2_X1 U15512 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13415), .S(n10105), .Z(
        P2_U3493) );
  MUX2_X1 U15513 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13416), .S(n10105), .Z(
        P2_U3492) );
  MUX2_X1 U15514 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13417), .S(n10105), .Z(
        P2_U3491) );
  MUX2_X1 U15515 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13418), .S(n10105), .Z(
        P2_U3490) );
  MUX2_X1 U15516 ( .A(n13419), .B(P2_REG0_REG_22__SCAN_IN), .S(n14991), .Z(
        n13420) );
  AOI21_X1 U15517 ( .B1(n13440), .B2(n13421), .A(n13420), .ZN(n13422) );
  INV_X1 U15518 ( .A(n13422), .ZN(P2_U3489) );
  MUX2_X1 U15519 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13423), .S(n10105), .Z(
        n13424) );
  AOI21_X1 U15520 ( .B1(n13440), .B2(n13425), .A(n13424), .ZN(n13426) );
  INV_X1 U15521 ( .A(n13426), .ZN(P2_U3488) );
  MUX2_X1 U15522 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13427), .S(n10105), .Z(
        P2_U3487) );
  INV_X1 U15523 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13429) );
  MUX2_X1 U15524 ( .A(n13429), .B(n13428), .S(n10105), .Z(n13430) );
  OAI21_X1 U15525 ( .B1(n13432), .B2(n13431), .A(n13430), .ZN(P2_U3486) );
  MUX2_X1 U15526 ( .A(n13433), .B(P2_REG0_REG_18__SCAN_IN), .S(n14991), .Z(
        n13434) );
  AOI21_X1 U15527 ( .B1(n13440), .B2(n13435), .A(n13434), .ZN(n13436) );
  INV_X1 U15528 ( .A(n13436), .ZN(P2_U3484) );
  MUX2_X1 U15529 ( .A(n13437), .B(P2_REG0_REG_17__SCAN_IN), .S(n14991), .Z(
        n13438) );
  AOI21_X1 U15530 ( .B1(n13440), .B2(n13439), .A(n13438), .ZN(n13441) );
  INV_X1 U15531 ( .A(n13441), .ZN(P2_U3481) );
  MUX2_X1 U15532 ( .A(n13442), .B(P2_REG0_REG_16__SCAN_IN), .S(n14991), .Z(
        P2_U3478) );
  INV_X1 U15533 ( .A(n13757), .ZN(n14277) );
  INV_X1 U15534 ( .A(n13443), .ZN(n13445) );
  NOR4_X1 U15535 ( .A1(n13445), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3088), 
        .A4(n13444), .ZN(n13446) );
  AOI21_X1 U15536 ( .B1(n13451), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13446), 
        .ZN(n13447) );
  OAI21_X1 U15537 ( .B1(n14277), .B2(n13461), .A(n13447), .ZN(P2_U3296) );
  OAI222_X1 U15538 ( .A1(n13461), .A2(n13449), .B1(n7468), .B2(P2_U3088), .C1(
        n13448), .C2(n13458), .ZN(P2_U3298) );
  AOI21_X1 U15539 ( .B1(n13451), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13450), 
        .ZN(n13452) );
  OAI21_X1 U15540 ( .B1(n13453), .B2(n13461), .A(n13452), .ZN(P2_U3299) );
  OAI222_X1 U15541 ( .A1(n13467), .A2(n13456), .B1(P2_U3088), .B2(n13455), 
        .C1(n13454), .C2(n13458), .ZN(P2_U3300) );
  INV_X1 U15542 ( .A(n13457), .ZN(n14279) );
  OAI222_X1 U15543 ( .A1(n13461), .A2(n14279), .B1(n13460), .B2(P2_U3088), 
        .C1(n13459), .C2(n13458), .ZN(P2_U3301) );
  INV_X1 U15544 ( .A(n13462), .ZN(n14282) );
  OAI222_X1 U15545 ( .A1(n13458), .A2(n13464), .B1(n13467), .B2(n14282), .C1(
        P2_U3088), .C2(n13463), .ZN(P2_U3302) );
  INV_X1 U15546 ( .A(n13465), .ZN(n14285) );
  OAI222_X1 U15547 ( .A1(n13458), .A2(n13468), .B1(n13467), .B2(n14285), .C1(
        P2_U3088), .C2(n13466), .ZN(P2_U3303) );
  MUX2_X1 U15548 ( .A(n13469), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15549 ( .A(n13471), .B(n13470), .Z(n13478) );
  NAND2_X1 U15550 ( .A1(n13827), .A2(n13551), .ZN(n13473) );
  NAND2_X1 U15551 ( .A1(n13825), .A2(n14645), .ZN(n13472) );
  AND2_X1 U15552 ( .A1(n13473), .A2(n13472), .ZN(n14204) );
  OAI22_X1 U15553 ( .A1(n14649), .A2(n14204), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13474), .ZN(n13475) );
  AOI21_X1 U15554 ( .B1(n14060), .B2(n13563), .A(n13475), .ZN(n13477) );
  NAND2_X1 U15555 ( .A1(n14059), .A2(n14657), .ZN(n13476) );
  OAI211_X1 U15556 ( .C1(n13478), .C2(n14651), .A(n13477), .B(n13476), .ZN(
        P1_U3216) );
  AOI21_X1 U15557 ( .B1(n13480), .B2(n13479), .A(n14651), .ZN(n13482) );
  NAND2_X1 U15558 ( .A1(n13482), .A2(n13481), .ZN(n13488) );
  NAND2_X1 U15559 ( .A1(n13829), .A2(n14645), .ZN(n13484) );
  NAND2_X1 U15560 ( .A1(n13831), .A2(n13551), .ZN(n13483) );
  NAND2_X1 U15561 ( .A1(n13484), .A2(n13483), .ZN(n14232) );
  NOR2_X1 U15562 ( .A1(n13485), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13963) );
  NOR2_X1 U15563 ( .A1(n14659), .A2(n14117), .ZN(n13486) );
  AOI211_X1 U15564 ( .C1(n14232), .C2(n14578), .A(n13963), .B(n13486), .ZN(
        n13487) );
  OAI211_X1 U15565 ( .C1(n6863), .C2(n13567), .A(n13488), .B(n13487), .ZN(
        P1_U3219) );
  INV_X1 U15566 ( .A(n13489), .ZN(n13490) );
  AOI21_X1 U15567 ( .B1(n13492), .B2(n13491), .A(n13490), .ZN(n13498) );
  AND2_X1 U15568 ( .A1(n13827), .A2(n14645), .ZN(n13493) );
  AOI21_X1 U15569 ( .B1(n13829), .B2(n13551), .A(n13493), .ZN(n14216) );
  OAI22_X1 U15570 ( .A1(n14216), .A2(n14649), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13494), .ZN(n13496) );
  NOR2_X1 U15571 ( .A1(n14218), .A2(n13567), .ZN(n13495) );
  AOI211_X1 U15572 ( .C1(n13563), .C2(n14087), .A(n13496), .B(n13495), .ZN(
        n13497) );
  OAI21_X1 U15573 ( .B1(n13498), .B2(n14651), .A(n13497), .ZN(P1_U3223) );
  XOR2_X1 U15574 ( .A(n13500), .B(n13499), .Z(n13507) );
  NAND2_X1 U15575 ( .A1(n13825), .A2(n13551), .ZN(n13502) );
  NAND2_X1 U15576 ( .A1(n13823), .A2(n14645), .ZN(n13501) );
  AND2_X1 U15577 ( .A1(n13502), .A2(n13501), .ZN(n14192) );
  OAI22_X1 U15578 ( .A1(n14649), .A2(n14192), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13503), .ZN(n13504) );
  AOI21_X1 U15579 ( .B1(n14026), .B2(n13563), .A(n13504), .ZN(n13506) );
  NAND2_X1 U15580 ( .A1(n6693), .A2(n14657), .ZN(n13505) );
  OAI211_X1 U15581 ( .C1(n13507), .C2(n14651), .A(n13506), .B(n13505), .ZN(
        P1_U3225) );
  OAI21_X1 U15582 ( .B1(n13510), .B2(n13509), .A(n13508), .ZN(n13511) );
  NAND2_X1 U15583 ( .A1(n13511), .A2(n14576), .ZN(n13515) );
  INV_X1 U15584 ( .A(n13512), .ZN(n14154) );
  AOI22_X1 U15585 ( .A1(n13831), .A2(n14645), .B1(n13551), .B2(n13833), .ZN(
        n14148) );
  NAND2_X1 U15586 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13917)
         );
  OAI21_X1 U15587 ( .B1(n14148), .B2(n14649), .A(n13917), .ZN(n13513) );
  AOI21_X1 U15588 ( .B1(n14154), .B2(n13563), .A(n13513), .ZN(n13514) );
  OAI211_X1 U15589 ( .C1(n6865), .C2(n13567), .A(n13515), .B(n13514), .ZN(
        P1_U3228) );
  XOR2_X1 U15590 ( .A(n13517), .B(n13516), .Z(n13522) );
  AOI22_X1 U15591 ( .A1(n13551), .A2(n13826), .B1(n13824), .B2(n14645), .ZN(
        n14041) );
  OAI22_X1 U15592 ( .A1(n14649), .A2(n14041), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13518), .ZN(n13519) );
  AOI21_X1 U15593 ( .B1(n14046), .B2(n13563), .A(n13519), .ZN(n13521) );
  NAND2_X1 U15594 ( .A1(n14200), .A2(n14657), .ZN(n13520) );
  OAI211_X1 U15595 ( .C1(n13522), .C2(n14651), .A(n13521), .B(n13520), .ZN(
        P1_U3229) );
  OAI211_X1 U15596 ( .C1(n13525), .C2(n13524), .A(n13523), .B(n14576), .ZN(
        n13531) );
  INV_X1 U15597 ( .A(n13526), .ZN(n14102) );
  AND2_X1 U15598 ( .A1(n13828), .A2(n14645), .ZN(n13527) );
  AOI21_X1 U15599 ( .B1(n13830), .B2(n13551), .A(n13527), .ZN(n14223) );
  INV_X1 U15600 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13528) );
  OAI22_X1 U15601 ( .A1(n14223), .A2(n14649), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13528), .ZN(n13529) );
  AOI21_X1 U15602 ( .B1(n14102), .B2(n13563), .A(n13529), .ZN(n13530) );
  OAI211_X1 U15603 ( .C1(n14225), .C2(n13567), .A(n13531), .B(n13530), .ZN(
        P1_U3233) );
  OAI21_X1 U15604 ( .B1(n13534), .B2(n13533), .A(n13532), .ZN(n13535) );
  NAND2_X1 U15605 ( .A1(n13535), .A2(n14576), .ZN(n13539) );
  AOI22_X1 U15606 ( .A1(n13551), .A2(n13828), .B1(n13826), .B2(n14645), .ZN(
        n14068) );
  OAI22_X1 U15607 ( .A1(n14649), .A2(n14068), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13536), .ZN(n13537) );
  AOI21_X1 U15608 ( .B1(n14077), .B2(n13563), .A(n13537), .ZN(n13538) );
  OAI211_X1 U15609 ( .C1(n13567), .C2(n14080), .A(n13539), .B(n13538), .ZN(
        P1_U3235) );
  XOR2_X1 U15610 ( .A(n13541), .B(n13540), .Z(n13548) );
  OAI22_X1 U15611 ( .A1(n13577), .A2(n13544), .B1(n13543), .B2(n13542), .ZN(
        n14132) );
  NAND2_X1 U15612 ( .A1(n14132), .A2(n14578), .ZN(n13545) );
  NAND2_X1 U15613 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13928)
         );
  OAI211_X1 U15614 ( .C1(n14659), .C2(n14135), .A(n13545), .B(n13928), .ZN(
        n13546) );
  AOI21_X1 U15615 ( .B1(n14238), .B2(n14657), .A(n13546), .ZN(n13547) );
  OAI21_X1 U15616 ( .B1(n13548), .B2(n14651), .A(n13547), .ZN(P1_U3238) );
  XOR2_X1 U15617 ( .A(n13550), .B(n13549), .Z(n13558) );
  NAND2_X1 U15618 ( .A1(n13824), .A2(n13551), .ZN(n13553) );
  NAND2_X1 U15619 ( .A1(n13822), .A2(n14645), .ZN(n13552) );
  AND2_X1 U15620 ( .A1(n13553), .A2(n13552), .ZN(n14185) );
  OAI22_X1 U15621 ( .A1(n14649), .A2(n14185), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13554), .ZN(n13555) );
  AOI21_X1 U15622 ( .B1(n14014), .B2(n13563), .A(n13555), .ZN(n13557) );
  NAND2_X1 U15623 ( .A1(n13717), .A2(n14657), .ZN(n13556) );
  OAI211_X1 U15624 ( .C1(n13558), .C2(n14651), .A(n13557), .B(n13556), .ZN(
        P1_U3240) );
  OAI211_X1 U15625 ( .C1(n13561), .C2(n13560), .A(n13559), .B(n14576), .ZN(
        n13566) );
  NAND2_X1 U15626 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14692)
         );
  OAI21_X1 U15627 ( .B1(n14649), .B2(n14592), .A(n14692), .ZN(n13562) );
  AOI21_X1 U15628 ( .B1(n13564), .B2(n13563), .A(n13562), .ZN(n13565) );
  OAI211_X1 U15629 ( .C1(n14594), .C2(n13567), .A(n13566), .B(n13565), .ZN(
        P1_U3241) );
  NAND2_X1 U15630 ( .A1(n9561), .A2(n13568), .ZN(n13570) );
  NAND2_X1 U15631 ( .A1(n13573), .A2(n13572), .ZN(n13736) );
  MUX2_X1 U15632 ( .A(n13717), .B(n13823), .S(n13607), .Z(n13719) );
  MUX2_X1 U15633 ( .A(n12046), .B(n13574), .S(n13607), .Z(n13710) );
  NOR2_X1 U15634 ( .A1(n13831), .A2(n13768), .ZN(n13684) );
  INV_X1 U15635 ( .A(n13684), .ZN(n13576) );
  NAND3_X1 U15636 ( .A1(n14138), .A2(n13768), .A3(n13831), .ZN(n13575) );
  OAI21_X1 U15637 ( .B1(n14138), .B2(n13576), .A(n13575), .ZN(n13689) );
  NOR2_X1 U15638 ( .A1(n13577), .A2(n13607), .ZN(n13579) );
  NOR2_X1 U15639 ( .A1(n13830), .A2(n13768), .ZN(n13578) );
  MUX2_X1 U15640 ( .A(n13579), .B(n13578), .S(n14233), .Z(n13688) );
  NAND2_X1 U15641 ( .A1(n13768), .A2(n14647), .ZN(n13583) );
  NAND2_X1 U15642 ( .A1(n13580), .A2(n13587), .ZN(n13582) );
  MUX2_X1 U15643 ( .A(n13583), .B(n13582), .S(n6453), .Z(n13595) );
  XNOR2_X1 U15644 ( .A(n14722), .B(n13768), .ZN(n13585) );
  MUX2_X1 U15645 ( .A(n6656), .B(n13846), .S(n13587), .Z(n13588) );
  AOI21_X1 U15646 ( .B1(n13591), .B2(n13589), .A(n13588), .ZN(n13593) );
  OAI21_X1 U15647 ( .B1(n13593), .B2(n13592), .A(n13777), .ZN(n13594) );
  NAND2_X1 U15648 ( .A1(n13768), .A2(n6457), .ZN(n13597) );
  NAND2_X1 U15649 ( .A1(n13607), .A2(n14760), .ZN(n13596) );
  MUX2_X1 U15650 ( .A(n13597), .B(n13596), .S(n13845), .Z(n13598) );
  NAND2_X1 U15651 ( .A1(n13599), .A2(n13598), .ZN(n13604) );
  INV_X1 U15652 ( .A(n14646), .ZN(n13600) );
  MUX2_X1 U15653 ( .A(n13600), .B(n14768), .S(n13607), .Z(n13603) );
  MUX2_X1 U15654 ( .A(n13601), .B(n14646), .S(n13607), .Z(n13602) );
  NAND2_X1 U15655 ( .A1(n13604), .A2(n13603), .ZN(n13605) );
  MUX2_X1 U15656 ( .A(n13608), .B(n13844), .S(n13607), .Z(n13612) );
  NAND2_X1 U15657 ( .A1(n13611), .A2(n13612), .ZN(n13610) );
  MUX2_X1 U15658 ( .A(n13844), .B(n13608), .S(n13607), .Z(n13609) );
  INV_X1 U15659 ( .A(n13611), .ZN(n13614) );
  INV_X1 U15660 ( .A(n13612), .ZN(n13613) );
  NAND2_X1 U15661 ( .A1(n13614), .A2(n13613), .ZN(n13615) );
  MUX2_X1 U15662 ( .A(n13843), .B(n13616), .S(n13607), .Z(n13618) );
  MUX2_X1 U15663 ( .A(n13616), .B(n13843), .S(n13607), .Z(n13617) );
  INV_X1 U15664 ( .A(n13618), .ZN(n13619) );
  MUX2_X1 U15665 ( .A(n13842), .B(n13620), .S(n13768), .Z(n13624) );
  NAND2_X1 U15666 ( .A1(n13623), .A2(n13624), .ZN(n13622) );
  MUX2_X1 U15667 ( .A(n13842), .B(n13620), .S(n13607), .Z(n13621) );
  NAND2_X1 U15668 ( .A1(n13622), .A2(n13621), .ZN(n13628) );
  INV_X1 U15669 ( .A(n13623), .ZN(n13626) );
  INV_X1 U15670 ( .A(n13624), .ZN(n13625) );
  NAND2_X1 U15671 ( .A1(n13626), .A2(n13625), .ZN(n13627) );
  MUX2_X1 U15672 ( .A(n13841), .B(n14787), .S(n13607), .Z(n13632) );
  NAND2_X1 U15673 ( .A1(n13631), .A2(n13632), .ZN(n13630) );
  MUX2_X1 U15674 ( .A(n13841), .B(n14787), .S(n13768), .Z(n13629) );
  NAND2_X1 U15675 ( .A1(n13630), .A2(n13629), .ZN(n13636) );
  INV_X1 U15676 ( .A(n13631), .ZN(n13634) );
  INV_X1 U15677 ( .A(n13632), .ZN(n13633) );
  NAND2_X1 U15678 ( .A1(n13634), .A2(n13633), .ZN(n13635) );
  MUX2_X1 U15679 ( .A(n13840), .B(n14698), .S(n13768), .Z(n13638) );
  MUX2_X1 U15680 ( .A(n13840), .B(n14698), .S(n13607), .Z(n13637) );
  INV_X1 U15681 ( .A(n13638), .ZN(n13639) );
  MUX2_X1 U15682 ( .A(n13839), .B(n13640), .S(n13607), .Z(n13644) );
  NAND2_X1 U15683 ( .A1(n13643), .A2(n13644), .ZN(n13642) );
  MUX2_X1 U15684 ( .A(n13839), .B(n13640), .S(n13768), .Z(n13641) );
  NAND2_X1 U15685 ( .A1(n13642), .A2(n13641), .ZN(n13648) );
  INV_X1 U15686 ( .A(n13643), .ZN(n13646) );
  INV_X1 U15687 ( .A(n13644), .ZN(n13645) );
  NAND2_X1 U15688 ( .A1(n13646), .A2(n13645), .ZN(n13647) );
  MUX2_X1 U15689 ( .A(n13838), .B(n13649), .S(n13768), .Z(n13651) );
  MUX2_X1 U15690 ( .A(n13838), .B(n13649), .S(n13607), .Z(n13650) );
  INV_X1 U15691 ( .A(n13651), .ZN(n13652) );
  MUX2_X1 U15692 ( .A(n13837), .B(n14564), .S(n13607), .Z(n13656) );
  NAND2_X1 U15693 ( .A1(n13655), .A2(n13656), .ZN(n13654) );
  MUX2_X1 U15694 ( .A(n14564), .B(n13837), .S(n13607), .Z(n13653) );
  NAND2_X1 U15695 ( .A1(n13654), .A2(n13653), .ZN(n13660) );
  INV_X1 U15696 ( .A(n13655), .ZN(n13658) );
  INV_X1 U15697 ( .A(n13656), .ZN(n13657) );
  NAND2_X1 U15698 ( .A1(n13658), .A2(n13657), .ZN(n13659) );
  MUX2_X1 U15699 ( .A(n13836), .B(n13661), .S(n13607), .Z(n13662) );
  MUX2_X1 U15700 ( .A(n13661), .B(n13836), .S(n13607), .Z(n13663) );
  NAND2_X1 U15701 ( .A1(n13672), .A2(n13664), .ZN(n13667) );
  NAND2_X1 U15702 ( .A1(n13671), .A2(n13665), .ZN(n13666) );
  MUX2_X1 U15703 ( .A(n13667), .B(n13666), .S(n13607), .Z(n13668) );
  AOI21_X1 U15704 ( .B1(n13670), .B2(n13669), .A(n13668), .ZN(n13676) );
  INV_X1 U15705 ( .A(n13671), .ZN(n13674) );
  INV_X1 U15706 ( .A(n13672), .ZN(n13673) );
  MUX2_X1 U15707 ( .A(n13674), .B(n13673), .S(n13607), .Z(n13675) );
  MUX2_X1 U15708 ( .A(n14585), .B(n13677), .S(n13607), .Z(n13679) );
  MUX2_X1 U15709 ( .A(n13833), .B(n14575), .S(n13607), .Z(n13678) );
  OAI21_X1 U15710 ( .B1(n13680), .B2(n13679), .A(n13678), .ZN(n13681) );
  MUX2_X1 U15711 ( .A(n13683), .B(n13682), .S(n13607), .Z(n13686) );
  MUX2_X1 U15712 ( .A(n13768), .B(n13831), .S(n14238), .Z(n13685) );
  MUX2_X1 U15713 ( .A(n14105), .B(n13829), .S(n13607), .Z(n13690) );
  MUX2_X1 U15714 ( .A(n13829), .B(n14105), .S(n13607), .Z(n13692) );
  INV_X1 U15715 ( .A(n13690), .ZN(n13691) );
  MUX2_X1 U15716 ( .A(n13693), .B(n14218), .S(n13607), .Z(n13695) );
  MUX2_X1 U15717 ( .A(n14090), .B(n13828), .S(n13607), .Z(n13694) );
  OAI21_X1 U15718 ( .B1(n6483), .B2(n13695), .A(n13694), .ZN(n13698) );
  AOI21_X1 U15719 ( .B1(n6483), .B2(n13695), .A(n13696), .ZN(n13697) );
  NAND2_X1 U15720 ( .A1(n13698), .A2(n13697), .ZN(n13702) );
  MUX2_X1 U15721 ( .A(n13700), .B(n13699), .S(n13607), .Z(n13701) );
  MUX2_X1 U15722 ( .A(n13826), .B(n14059), .S(n13607), .Z(n13704) );
  NAND2_X1 U15723 ( .A1(n13703), .A2(n13704), .ZN(n13708) );
  MUX2_X1 U15724 ( .A(n14059), .B(n13826), .S(n13607), .Z(n13707) );
  INV_X1 U15725 ( .A(n13703), .ZN(n13706) );
  INV_X1 U15726 ( .A(n13704), .ZN(n13705) );
  MUX2_X1 U15727 ( .A(n13825), .B(n14200), .S(n13607), .Z(n13709) );
  MUX2_X1 U15728 ( .A(n13824), .B(n6693), .S(n13607), .Z(n13715) );
  INV_X1 U15729 ( .A(n13824), .ZN(n13713) );
  MUX2_X1 U15730 ( .A(n14193), .B(n13713), .S(n13607), .Z(n13714) );
  MUX2_X1 U15731 ( .A(n13823), .B(n13717), .S(n13607), .Z(n13718) );
  MUX2_X1 U15732 ( .A(n13822), .B(n13998), .S(n13607), .Z(n13723) );
  MUX2_X1 U15733 ( .A(n13998), .B(n13822), .S(n13587), .Z(n13720) );
  NAND2_X1 U15734 ( .A1(n13721), .A2(n13720), .ZN(n13725) );
  MUX2_X1 U15735 ( .A(n14174), .B(n13821), .S(n13607), .Z(n13743) );
  MUX2_X1 U15736 ( .A(n13821), .B(n14174), .S(n13607), .Z(n13726) );
  NAND2_X1 U15737 ( .A1(n13728), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13729) );
  NAND2_X1 U15738 ( .A1(n11930), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U15739 ( .A1(n6456), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U15740 ( .A1(n13730), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n13731) );
  NAND3_X1 U15741 ( .A1(n13733), .A2(n13732), .A3(n13731), .ZN(n13968) );
  NAND2_X1 U15742 ( .A1(n13607), .A2(n13968), .ZN(n13735) );
  INV_X1 U15743 ( .A(n13819), .ZN(n13734) );
  AOI21_X1 U15744 ( .B1(n13736), .B2(n13735), .A(n13734), .ZN(n13737) );
  AOI21_X1 U15745 ( .B1(n13973), .B2(n13768), .A(n13737), .ZN(n13749) );
  OAI21_X1 U15746 ( .B1(n13968), .B2(n13738), .A(n13819), .ZN(n13739) );
  INV_X1 U15747 ( .A(n13739), .ZN(n13740) );
  MUX2_X1 U15748 ( .A(n13741), .B(n14169), .S(n13768), .Z(n13745) );
  INV_X1 U15749 ( .A(n13741), .ZN(n13820) );
  INV_X1 U15750 ( .A(n13744), .ZN(n13747) );
  INV_X1 U15751 ( .A(n13745), .ZN(n13746) );
  NAND2_X1 U15752 ( .A1(n13752), .A2(n13748), .ZN(n13754) );
  INV_X1 U15753 ( .A(n13750), .ZN(n13751) );
  OAI21_X1 U15754 ( .B1(n13752), .B2(n13748), .A(n13751), .ZN(n13753) );
  NAND2_X1 U15755 ( .A1(n13757), .A2(n13756), .ZN(n13760) );
  NAND2_X1 U15756 ( .A1(n13728), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n13759) );
  XNOR2_X1 U15757 ( .A(n13970), .B(n13968), .ZN(n13806) );
  NAND2_X1 U15758 ( .A1(n13762), .A2(n13761), .ZN(n13764) );
  AND2_X1 U15759 ( .A1(n13764), .A2(n13763), .ZN(n13772) );
  INV_X1 U15760 ( .A(n13772), .ZN(n13766) );
  NOR2_X1 U15761 ( .A1(n13768), .A2(n13968), .ZN(n13771) );
  INV_X1 U15762 ( .A(n13968), .ZN(n13769) );
  NOR3_X1 U15763 ( .A1(n13970), .A2(n13769), .A3(n13587), .ZN(n13770) );
  AOI21_X1 U15764 ( .B1(n13771), .B2(n13970), .A(n13770), .ZN(n13774) );
  NAND3_X1 U15765 ( .A1(n13773), .A2(n13772), .A3(n13774), .ZN(n13812) );
  INV_X1 U15766 ( .A(n13774), .ZN(n13775) );
  AOI21_X1 U15767 ( .B1(n13775), .B2(n7429), .A(n13817), .ZN(n13811) );
  INV_X1 U15768 ( .A(n13776), .ZN(n13778) );
  NAND4_X1 U15769 ( .A1(n13778), .A2(n14706), .A3(n13777), .A4(n10256), .ZN(
        n13781) );
  NOR3_X1 U15770 ( .A1(n13781), .A2(n13780), .A3(n13779), .ZN(n13784) );
  NAND4_X1 U15771 ( .A1(n13785), .A2(n13784), .A3(n13783), .A4(n13782), .ZN(
        n13786) );
  NOR2_X1 U15772 ( .A1(n13787), .A2(n13786), .ZN(n13790) );
  NAND4_X1 U15773 ( .A1(n13791), .A2(n13790), .A3(n13789), .A4(n13788), .ZN(
        n13792) );
  OR4_X1 U15774 ( .A1(n13794), .A2(n13793), .A3(n7217), .A4(n13792), .ZN(
        n13795) );
  NOR2_X1 U15775 ( .A1(n6680), .A2(n13795), .ZN(n13797) );
  NAND4_X1 U15776 ( .A1(n13798), .A2(n14128), .A3(n13797), .A4(n13796), .ZN(
        n13799) );
  NOR4_X1 U15777 ( .A1(n13696), .A2(n13800), .A3(n14085), .A4(n13799), .ZN(
        n13801) );
  NAND4_X1 U15778 ( .A1(n14025), .A2(n13801), .A3(n14038), .A4(n14056), .ZN(
        n13802) );
  NOR4_X1 U15779 ( .A1(n13983), .A2(n13995), .A3(n14008), .A4(n13802), .ZN(
        n13805) );
  XNOR2_X1 U15780 ( .A(n13973), .B(n13819), .ZN(n13803) );
  NAND4_X1 U15781 ( .A1(n13806), .A2(n13805), .A3(n13804), .A4(n13803), .ZN(
        n13807) );
  XNOR2_X1 U15782 ( .A(n13807), .B(n14155), .ZN(n13809) );
  NAND2_X1 U15783 ( .A1(n13809), .A2(n13808), .ZN(n13810) );
  NOR2_X1 U15784 ( .A1(n6455), .A2(P1_U3086), .ZN(n13814) );
  NAND3_X1 U15785 ( .A1(n13815), .A2(n13551), .A3(n13814), .ZN(n13816) );
  OAI211_X1 U15786 ( .C1(n9565), .C2(n13817), .A(n13816), .B(P1_B_REG_SCAN_IN), 
        .ZN(n13818) );
  MUX2_X1 U15787 ( .A(n13968), .B(P1_DATAO_REG_31__SCAN_IN), .S(n13847), .Z(
        P1_U3591) );
  MUX2_X1 U15788 ( .A(n13819), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13847), .Z(
        P1_U3590) );
  MUX2_X1 U15789 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13820), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15790 ( .A(n13821), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13847), .Z(
        P1_U3588) );
  MUX2_X1 U15791 ( .A(n13822), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13847), .Z(
        P1_U3587) );
  MUX2_X1 U15792 ( .A(n13823), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13847), .Z(
        P1_U3586) );
  MUX2_X1 U15793 ( .A(n13824), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13847), .Z(
        P1_U3585) );
  MUX2_X1 U15794 ( .A(n13825), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13847), .Z(
        P1_U3584) );
  MUX2_X1 U15795 ( .A(n13826), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13847), .Z(
        P1_U3583) );
  MUX2_X1 U15796 ( .A(n13827), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13847), .Z(
        P1_U3582) );
  MUX2_X1 U15797 ( .A(n13828), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13847), .Z(
        P1_U3581) );
  MUX2_X1 U15798 ( .A(n13829), .B(P1_DATAO_REG_20__SCAN_IN), .S(n13847), .Z(
        P1_U3580) );
  MUX2_X1 U15799 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13830), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15800 ( .A(n13831), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13847), .Z(
        P1_U3578) );
  MUX2_X1 U15801 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13832), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15802 ( .A(n13833), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13847), .Z(
        P1_U3576) );
  MUX2_X1 U15803 ( .A(n13834), .B(P1_DATAO_REG_15__SCAN_IN), .S(n13847), .Z(
        P1_U3575) );
  MUX2_X1 U15804 ( .A(n13835), .B(P1_DATAO_REG_14__SCAN_IN), .S(n13847), .Z(
        P1_U3574) );
  MUX2_X1 U15805 ( .A(n13836), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13847), .Z(
        P1_U3573) );
  MUX2_X1 U15806 ( .A(n13837), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13847), .Z(
        P1_U3572) );
  MUX2_X1 U15807 ( .A(n13838), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13847), .Z(
        P1_U3571) );
  MUX2_X1 U15808 ( .A(n13839), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13847), .Z(
        P1_U3570) );
  MUX2_X1 U15809 ( .A(n13840), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13847), .Z(
        P1_U3569) );
  MUX2_X1 U15810 ( .A(n13841), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13847), .Z(
        P1_U3568) );
  MUX2_X1 U15811 ( .A(n13842), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13847), .Z(
        P1_U3567) );
  MUX2_X1 U15812 ( .A(n13843), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13847), .Z(
        P1_U3566) );
  MUX2_X1 U15813 ( .A(n13844), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13847), .Z(
        P1_U3565) );
  MUX2_X1 U15814 ( .A(n14646), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13847), .Z(
        P1_U3564) );
  MUX2_X1 U15815 ( .A(n13845), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13847), .Z(
        P1_U3563) );
  MUX2_X1 U15816 ( .A(n14647), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13847), .Z(
        P1_U3562) );
  MUX2_X1 U15817 ( .A(n13846), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13847), .Z(
        P1_U3561) );
  MUX2_X1 U15818 ( .A(n13848), .B(P1_DATAO_REG_0__SCAN_IN), .S(n13847), .Z(
        P1_U3560) );
  OAI211_X1 U15819 ( .C1(n13858), .C2(n13849), .A(n14690), .B(n13865), .ZN(
        n13856) );
  OAI211_X1 U15820 ( .C1(n13851), .C2(n13850), .A(n14689), .B(n13870), .ZN(
        n13855) );
  NAND2_X1 U15821 ( .A1(n14686), .A2(n13852), .ZN(n13854) );
  AOI22_X1 U15822 ( .A1(n14673), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13853) );
  NAND4_X1 U15823 ( .A1(n13856), .A2(n13855), .A3(n13854), .A4(n13853), .ZN(
        P1_U3244) );
  MUX2_X1 U15824 ( .A(n13859), .B(n13858), .S(n13857), .Z(n13861) );
  NAND2_X1 U15825 ( .A1(n13861), .A2(n13860), .ZN(n13862) );
  OAI211_X1 U15826 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n13863), .A(n13862), .B(
        P1_U4016), .ZN(n14678) );
  AOI22_X1 U15827 ( .A1(n14673), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13878) );
  MUX2_X1 U15828 ( .A(n9448), .B(P1_REG2_REG_2__SCAN_IN), .S(n13868), .Z(
        n13866) );
  NAND3_X1 U15829 ( .A1(n13866), .A2(n13865), .A3(n13864), .ZN(n13867) );
  NAND3_X1 U15830 ( .A1(n14690), .A2(n13888), .A3(n13867), .ZN(n13874) );
  MUX2_X1 U15831 ( .A(n9407), .B(P1_REG1_REG_2__SCAN_IN), .S(n13868), .Z(
        n13871) );
  NAND3_X1 U15832 ( .A1(n13871), .A2(n13870), .A3(n13869), .ZN(n13872) );
  NAND3_X1 U15833 ( .A1(n14689), .A2(n13883), .A3(n13872), .ZN(n13873) );
  OAI211_X1 U15834 ( .C1(n13955), .C2(n13875), .A(n13874), .B(n13873), .ZN(
        n13876) );
  INV_X1 U15835 ( .A(n13876), .ZN(n13877) );
  NAND3_X1 U15836 ( .A1(n14678), .A2(n13878), .A3(n13877), .ZN(P1_U3245) );
  INV_X1 U15837 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n13879) );
  NAND2_X1 U15838 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14648) );
  OAI21_X1 U15839 ( .B1(n14694), .B2(n13879), .A(n14648), .ZN(n13880) );
  AOI21_X1 U15840 ( .B1(n13885), .B2(n14686), .A(n13880), .ZN(n13892) );
  MUX2_X1 U15841 ( .A(n9414), .B(P1_REG1_REG_3__SCAN_IN), .S(n13885), .Z(
        n13882) );
  NAND3_X1 U15842 ( .A1(n13883), .A2(n13882), .A3(n13881), .ZN(n13884) );
  NAND3_X1 U15843 ( .A1(n14689), .A2(n14668), .A3(n13884), .ZN(n13891) );
  MUX2_X1 U15844 ( .A(n9452), .B(P1_REG2_REG_3__SCAN_IN), .S(n13885), .Z(
        n13887) );
  NAND3_X1 U15845 ( .A1(n13888), .A2(n13887), .A3(n13886), .ZN(n13889) );
  NAND3_X1 U15846 ( .A1(n14690), .A2(n14662), .A3(n13889), .ZN(n13890) );
  NAND3_X1 U15847 ( .A1(n13892), .A2(n13891), .A3(n13890), .ZN(P1_U3246) );
  INV_X1 U15848 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n13894) );
  OAI21_X1 U15849 ( .B1(n14694), .B2(n13894), .A(n13893), .ZN(n13895) );
  AOI21_X1 U15850 ( .B1(n13897), .B2(n14686), .A(n13895), .ZN(n13910) );
  INV_X1 U15851 ( .A(n13896), .ZN(n13899) );
  MUX2_X1 U15852 ( .A(n14813), .B(P1_REG1_REG_7__SCAN_IN), .S(n13897), .Z(
        n13898) );
  NAND2_X1 U15853 ( .A1(n13899), .A2(n13898), .ZN(n13901) );
  OAI211_X1 U15854 ( .C1(n13902), .C2(n13901), .A(n14689), .B(n13900), .ZN(
        n13909) );
  NAND3_X1 U15855 ( .A1(n13905), .A2(n13904), .A3(n13903), .ZN(n13906) );
  NAND3_X1 U15856 ( .A1(n14690), .A2(n13907), .A3(n13906), .ZN(n13908) );
  NAND3_X1 U15857 ( .A1(n13910), .A2(n13909), .A3(n13908), .ZN(P1_U3250) );
  AOI21_X1 U15858 ( .B1(n13912), .B2(P1_REG1_REG_16__SCAN_IN), .A(n13911), 
        .ZN(n13915) );
  XNOR2_X1 U15859 ( .A(n13936), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n13914) );
  NOR2_X1 U15860 ( .A1(n13915), .A2(n13914), .ZN(n13935) );
  AOI211_X1 U15861 ( .C1(n13915), .C2(n13914), .A(n13935), .B(n13913), .ZN(
        n13916) );
  INV_X1 U15862 ( .A(n13916), .ZN(n13927) );
  INV_X1 U15863 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n13918) );
  OAI21_X1 U15864 ( .B1(n14694), .B2(n13918), .A(n13917), .ZN(n13919) );
  AOI21_X1 U15865 ( .B1(n13936), .B2(n14686), .A(n13919), .ZN(n13926) );
  XNOR2_X1 U15866 ( .A(n13932), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n13924) );
  OAI21_X1 U15867 ( .B1(n13922), .B2(n13921), .A(n13920), .ZN(n13923) );
  NAND2_X1 U15868 ( .A1(n13924), .A2(n13923), .ZN(n13931) );
  OAI211_X1 U15869 ( .C1(n13924), .C2(n13923), .A(n14690), .B(n13931), .ZN(
        n13925) );
  NAND3_X1 U15870 ( .A1(n13927), .A2(n13926), .A3(n13925), .ZN(P1_U3260) );
  INV_X1 U15871 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n13929) );
  OAI21_X1 U15872 ( .B1(n14694), .B2(n13929), .A(n13928), .ZN(n13930) );
  AOI21_X1 U15873 ( .B1(n13951), .B2(n14686), .A(n13930), .ZN(n13943) );
  INV_X1 U15874 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13933) );
  OAI21_X1 U15875 ( .B1(n13933), .B2(n13932), .A(n13931), .ZN(n13950) );
  XNOR2_X1 U15876 ( .A(n13944), .B(n13950), .ZN(n13934) );
  NAND2_X1 U15877 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13934), .ZN(n13953) );
  OAI211_X1 U15878 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13934), .A(n14690), 
        .B(n13953), .ZN(n13942) );
  AOI21_X1 U15879 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13936), .A(n13935), 
        .ZN(n13945) );
  XNOR2_X1 U15880 ( .A(n13944), .B(n13945), .ZN(n13937) );
  INV_X1 U15881 ( .A(n13937), .ZN(n13940) );
  NOR2_X1 U15882 ( .A1(n13938), .A2(n13937), .ZN(n13946) );
  INV_X1 U15883 ( .A(n13946), .ZN(n13939) );
  OAI211_X1 U15884 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13940), .A(n14689), 
        .B(n13939), .ZN(n13941) );
  NAND3_X1 U15885 ( .A1(n13943), .A2(n13942), .A3(n13941), .ZN(P1_U3261) );
  NOR2_X1 U15886 ( .A1(n13945), .A2(n13944), .ZN(n13947) );
  NOR2_X1 U15887 ( .A1(n13947), .A2(n13946), .ZN(n13949) );
  XOR2_X1 U15888 ( .A(n13949), .B(n13948), .Z(n13960) );
  INV_X1 U15889 ( .A(n13960), .ZN(n13958) );
  NAND2_X1 U15890 ( .A1(n13951), .A2(n13950), .ZN(n13952) );
  NAND2_X1 U15891 ( .A1(n13953), .A2(n13952), .ZN(n13954) );
  XOR2_X1 U15892 ( .A(n13954), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13959) );
  OAI21_X1 U15893 ( .B1(n13959), .B2(n13956), .A(n13955), .ZN(n13957) );
  AOI21_X1 U15894 ( .B1(n13958), .B2(n14689), .A(n13957), .ZN(n13962) );
  AOI22_X1 U15895 ( .A1(n13960), .A2(n14689), .B1(n14690), .B2(n13959), .ZN(
        n13961) );
  MUX2_X1 U15896 ( .A(n13962), .B(n13961), .S(n14155), .Z(n13965) );
  INV_X1 U15897 ( .A(n13963), .ZN(n13964) );
  OAI211_X1 U15898 ( .C1(n13966), .C2(n14694), .A(n13965), .B(n13964), .ZN(
        P1_U3262) );
  NAND2_X1 U15899 ( .A1(n13974), .A2(n14164), .ZN(n13967) );
  NAND2_X1 U15900 ( .A1(n13969), .A2(n13968), .ZN(n14162) );
  NOR2_X1 U15901 ( .A1(n14739), .A2(n14162), .ZN(n13977) );
  NOR2_X1 U15902 ( .A1(n6856), .A2(n14712), .ZN(n13971) );
  AOI211_X1 U15903 ( .C1(P1_REG2_REG_31__SCAN_IN), .C2(n14739), .A(n13977), 
        .B(n13971), .ZN(n13972) );
  OAI21_X1 U15904 ( .B1(n14161), .B2(n14732), .A(n13972), .ZN(P1_U3263) );
  XNOR2_X1 U15905 ( .A(n13973), .B(n13974), .ZN(n13975) );
  NAND2_X1 U15906 ( .A1(n13975), .A2(n14730), .ZN(n14163) );
  NOR2_X1 U15907 ( .A1(n14164), .A2(n14712), .ZN(n13976) );
  AOI211_X1 U15908 ( .C1(n14697), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13977), 
        .B(n13976), .ZN(n13978) );
  OAI21_X1 U15909 ( .B1(n14163), .B2(n14732), .A(n13978), .ZN(P1_U3264) );
  INV_X1 U15910 ( .A(n13983), .ZN(n13984) );
  INV_X1 U15911 ( .A(n14177), .ZN(n13993) );
  AOI21_X1 U15912 ( .B1(n14174), .B2(n13997), .A(n14789), .ZN(n13988) );
  NAND2_X1 U15913 ( .A1(n13988), .A2(n13987), .ZN(n14175) );
  AOI22_X1 U15914 ( .A1(n14739), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14728), 
        .B2(n13989), .ZN(n13991) );
  NAND2_X1 U15915 ( .A1(n14174), .A2(n14735), .ZN(n13990) );
  OAI211_X1 U15916 ( .C1(n14175), .C2(n14732), .A(n13991), .B(n13990), .ZN(
        n13992) );
  AOI21_X1 U15917 ( .B1(n13993), .B2(n14124), .A(n13992), .ZN(n13994) );
  OAI21_X1 U15918 ( .B1(n14739), .B2(n7436), .A(n13994), .ZN(P1_U3265) );
  XNOR2_X1 U15919 ( .A(n13996), .B(n13995), .ZN(n14184) );
  AOI211_X1 U15920 ( .C1(n13998), .C2(n14013), .A(n14789), .B(n13986), .ZN(
        n14181) );
  INV_X1 U15921 ( .A(n13998), .ZN(n14179) );
  INV_X1 U15922 ( .A(n13999), .ZN(n14000) );
  OAI22_X1 U15923 ( .A1(n14697), .A2(n14178), .B1(n14000), .B2(n14116), .ZN(
        n14001) );
  AOI21_X1 U15924 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(n14739), .A(n14001), 
        .ZN(n14002) );
  OAI21_X1 U15925 ( .B1(n14179), .B2(n14712), .A(n14002), .ZN(n14003) );
  AOI21_X1 U15926 ( .B1(n14181), .B2(n14717), .A(n14003), .ZN(n14007) );
  XNOR2_X1 U15927 ( .A(n14005), .B(n14004), .ZN(n14182) );
  NAND2_X1 U15928 ( .A1(n14182), .A2(n14093), .ZN(n14006) );
  OAI211_X1 U15929 ( .C1(n14184), .C2(n14160), .A(n14007), .B(n14006), .ZN(
        P1_U3266) );
  XNOR2_X1 U15930 ( .A(n14009), .B(n14008), .ZN(n14191) );
  OAI21_X1 U15931 ( .B1(n14012), .B2(n14011), .A(n14010), .ZN(n14189) );
  OAI211_X1 U15932 ( .C1(n14187), .C2(n6484), .A(n14730), .B(n14013), .ZN(
        n14186) );
  INV_X1 U15933 ( .A(n14014), .ZN(n14015) );
  OAI22_X1 U15934 ( .A1(n14697), .A2(n14185), .B1(n14015), .B2(n14116), .ZN(
        n14017) );
  NOR2_X1 U15935 ( .A1(n14187), .A2(n14712), .ZN(n14016) );
  AOI211_X1 U15936 ( .C1(n14739), .C2(P1_REG2_REG_26__SCAN_IN), .A(n14017), 
        .B(n14016), .ZN(n14018) );
  OAI21_X1 U15937 ( .B1(n14732), .B2(n14186), .A(n14018), .ZN(n14019) );
  AOI21_X1 U15938 ( .B1(n14189), .B2(n14093), .A(n14019), .ZN(n14020) );
  OAI21_X1 U15939 ( .B1(n14191), .B2(n14160), .A(n14020), .ZN(P1_U3267) );
  XNOR2_X1 U15940 ( .A(n14025), .B(n14021), .ZN(n14198) );
  INV_X1 U15941 ( .A(n14022), .ZN(n14023) );
  AOI21_X1 U15942 ( .B1(n14025), .B2(n14024), .A(n14023), .ZN(n14196) );
  AOI211_X1 U15943 ( .C1(n6693), .C2(n14044), .A(n14789), .B(n6484), .ZN(
        n14195) );
  INV_X1 U15944 ( .A(n14026), .ZN(n14027) );
  OAI21_X1 U15945 ( .B1(n14116), .B2(n14027), .A(n14192), .ZN(n14028) );
  AOI21_X1 U15946 ( .B1(n14195), .B2(n14155), .A(n14028), .ZN(n14031) );
  AOI22_X1 U15947 ( .A1(n6693), .A2(n14735), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n14697), .ZN(n14030) );
  OAI21_X1 U15948 ( .B1(n14031), .B2(n14697), .A(n14030), .ZN(n14032) );
  AOI21_X1 U15949 ( .B1(n14196), .B2(n14124), .A(n14032), .ZN(n14033) );
  OAI21_X1 U15950 ( .B1(n14126), .B2(n14198), .A(n14033), .ZN(P1_U3268) );
  NAND2_X1 U15951 ( .A1(n14034), .A2(n14035), .ZN(n14036) );
  AOI21_X2 U15952 ( .B1(n14038), .B2(n14036), .A(n6494), .ZN(n14203) );
  OAI211_X1 U15953 ( .C1(n14039), .C2(n14038), .A(n14037), .B(n14784), .ZN(
        n14040) );
  OAI211_X1 U15954 ( .C1(n14203), .C2(n14130), .A(n14041), .B(n14040), .ZN(
        n14042) );
  INV_X1 U15955 ( .A(n14042), .ZN(n14202) );
  INV_X1 U15956 ( .A(n14044), .ZN(n14045) );
  AOI211_X1 U15957 ( .C1(n14200), .C2(n14058), .A(n14789), .B(n14045), .ZN(
        n14199) );
  AOI22_X1 U15958 ( .A1(n14697), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14046), 
        .B2(n14728), .ZN(n14047) );
  OAI21_X1 U15959 ( .B1(n12046), .B2(n14712), .A(n14047), .ZN(n14049) );
  NOR2_X1 U15960 ( .A1(n14203), .A2(n14139), .ZN(n14048) );
  AOI211_X1 U15961 ( .C1(n14199), .C2(n14717), .A(n14049), .B(n14048), .ZN(
        n14050) );
  OAI21_X1 U15962 ( .B1(n14739), .B2(n14202), .A(n14050), .ZN(P1_U3269) );
  INV_X1 U15963 ( .A(n14051), .ZN(n14053) );
  INV_X1 U15964 ( .A(n14056), .ZN(n14052) );
  OAI21_X1 U15965 ( .B1(n14053), .B2(n14052), .A(n14034), .ZN(n14210) );
  INV_X1 U15966 ( .A(n14054), .ZN(n14055) );
  OAI21_X1 U15967 ( .B1(n14057), .B2(n14056), .A(n14055), .ZN(n14208) );
  INV_X1 U15968 ( .A(n14059), .ZN(n14205) );
  AOI211_X1 U15969 ( .C1(n14059), .C2(n14075), .A(n14789), .B(n14043), .ZN(
        n14207) );
  NAND2_X1 U15970 ( .A1(n14207), .A2(n14717), .ZN(n14064) );
  INV_X1 U15971 ( .A(n14060), .ZN(n14061) );
  OAI22_X1 U15972 ( .A1(n14739), .A2(n14204), .B1(n14061), .B2(n14116), .ZN(
        n14062) );
  AOI21_X1 U15973 ( .B1(P1_REG2_REG_23__SCAN_IN), .B2(n14697), .A(n14062), 
        .ZN(n14063) );
  OAI211_X1 U15974 ( .C1(n14205), .C2(n14712), .A(n14064), .B(n14063), .ZN(
        n14065) );
  AOI21_X1 U15975 ( .B1(n14208), .B2(n14093), .A(n14065), .ZN(n14066) );
  OAI21_X1 U15976 ( .B1(n14210), .B2(n14160), .A(n14066), .ZN(P1_U3270) );
  XNOR2_X1 U15977 ( .A(n14067), .B(n13696), .ZN(n14070) );
  INV_X1 U15978 ( .A(n14068), .ZN(n14069) );
  AOI21_X1 U15979 ( .B1(n14070), .B2(n14784), .A(n14069), .ZN(n14214) );
  INV_X1 U15980 ( .A(n14071), .ZN(n14072) );
  AOI21_X1 U15981 ( .B1(n14074), .B2(n14073), .A(n14072), .ZN(n14215) );
  INV_X1 U15982 ( .A(n14215), .ZN(n14082) );
  INV_X1 U15983 ( .A(n14075), .ZN(n14076) );
  AOI211_X1 U15984 ( .C1(n14212), .C2(n14086), .A(n14789), .B(n14076), .ZN(
        n14211) );
  NAND2_X1 U15985 ( .A1(n14211), .A2(n14717), .ZN(n14079) );
  AOI22_X1 U15986 ( .A1(n14739), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14077), 
        .B2(n14728), .ZN(n14078) );
  OAI211_X1 U15987 ( .C1(n14712), .C2(n14080), .A(n14079), .B(n14078), .ZN(
        n14081) );
  AOI21_X1 U15988 ( .B1(n14082), .B2(n14124), .A(n14081), .ZN(n14083) );
  OAI21_X1 U15989 ( .B1(n14739), .B2(n14214), .A(n14083), .ZN(P1_U3271) );
  XOR2_X1 U15990 ( .A(n14085), .B(n6471), .Z(n14222) );
  XOR2_X1 U15991 ( .A(n14085), .B(n14084), .Z(n14220) );
  OAI211_X1 U15992 ( .C1(n14099), .C2(n14218), .A(n14730), .B(n14086), .ZN(
        n14217) );
  AOI22_X1 U15993 ( .A1(n14697), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14087), 
        .B2(n14728), .ZN(n14088) );
  OAI21_X1 U15994 ( .B1(n14216), .B2(n14697), .A(n14088), .ZN(n14089) );
  AOI21_X1 U15995 ( .B1(n14090), .B2(n14735), .A(n14089), .ZN(n14091) );
  OAI21_X1 U15996 ( .B1(n14217), .B2(n14732), .A(n14091), .ZN(n14092) );
  AOI21_X1 U15997 ( .B1(n14220), .B2(n14093), .A(n14092), .ZN(n14094) );
  OAI21_X1 U15998 ( .B1(n14222), .B2(n14160), .A(n14094), .ZN(P1_U3272) );
  XNOR2_X1 U15999 ( .A(n14095), .B(n14098), .ZN(n14229) );
  AOI21_X1 U16000 ( .B1(n14098), .B2(n14097), .A(n14096), .ZN(n14227) );
  INV_X1 U16001 ( .A(n14099), .ZN(n14101) );
  AOI21_X1 U16002 ( .B1(n14115), .B2(n14105), .A(n14789), .ZN(n14100) );
  NAND2_X1 U16003 ( .A1(n14101), .A2(n14100), .ZN(n14224) );
  AOI22_X1 U16004 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n14697), .B1(n14102), 
        .B2(n14728), .ZN(n14103) );
  OAI21_X1 U16005 ( .B1(n14223), .B2(n14697), .A(n14103), .ZN(n14104) );
  AOI21_X1 U16006 ( .B1(n14105), .B2(n14735), .A(n14104), .ZN(n14106) );
  OAI21_X1 U16007 ( .B1(n14224), .B2(n14732), .A(n14106), .ZN(n14107) );
  AOI21_X1 U16008 ( .B1(n14227), .B2(n14124), .A(n14107), .ZN(n14108) );
  OAI21_X1 U16009 ( .B1(n14229), .B2(n14126), .A(n14108), .ZN(P1_U3273) );
  AOI21_X1 U16010 ( .B1(n14112), .B2(n14110), .A(n14109), .ZN(n14236) );
  OAI21_X1 U16011 ( .B1(n14113), .B2(n14112), .A(n6695), .ZN(n14230) );
  AOI21_X1 U16012 ( .B1(n14233), .B2(n14134), .A(n14789), .ZN(n14114) );
  AND2_X1 U16013 ( .A1(n14115), .A2(n14114), .ZN(n14231) );
  NAND2_X1 U16014 ( .A1(n14231), .A2(n14717), .ZN(n14122) );
  INV_X1 U16015 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14118) );
  OAI22_X1 U16016 ( .A1(n14120), .A2(n14118), .B1(n14117), .B2(n14116), .ZN(
        n14119) );
  AOI21_X1 U16017 ( .B1(n14120), .B2(n14232), .A(n14119), .ZN(n14121) );
  OAI211_X1 U16018 ( .C1(n6863), .C2(n14712), .A(n14122), .B(n14121), .ZN(
        n14123) );
  AOI21_X1 U16019 ( .B1(n14230), .B2(n14124), .A(n14123), .ZN(n14125) );
  OAI21_X1 U16020 ( .B1(n14236), .B2(n14126), .A(n14125), .ZN(P1_U3274) );
  XNOR2_X1 U16021 ( .A(n14127), .B(n14128), .ZN(n14133) );
  XNOR2_X1 U16022 ( .A(n14129), .B(n14128), .ZN(n14241) );
  NOR2_X1 U16023 ( .A1(n14241), .A2(n14130), .ZN(n14131) );
  AOI211_X1 U16024 ( .C1(n14784), .C2(n14133), .A(n14132), .B(n14131), .ZN(
        n14240) );
  AOI211_X1 U16025 ( .C1(n14238), .C2(n14151), .A(n14789), .B(n6864), .ZN(
        n14237) );
  INV_X1 U16026 ( .A(n14135), .ZN(n14136) );
  AOI22_X1 U16027 ( .A1(n14697), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14136), 
        .B2(n14728), .ZN(n14137) );
  OAI21_X1 U16028 ( .B1(n14138), .B2(n14712), .A(n14137), .ZN(n14141) );
  NOR2_X1 U16029 ( .A1(n14241), .A2(n14139), .ZN(n14140) );
  AOI211_X1 U16030 ( .C1(n14237), .C2(n14717), .A(n14141), .B(n14140), .ZN(
        n14142) );
  OAI21_X1 U16031 ( .B1(n14240), .B2(n14697), .A(n14142), .ZN(P1_U3275) );
  AOI21_X1 U16032 ( .B1(n14145), .B2(n14144), .A(n14143), .ZN(n14146) );
  INV_X1 U16033 ( .A(n14146), .ZN(n14246) );
  AOI22_X1 U16034 ( .A1(n14243), .A2(n14735), .B1(n14739), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n14159) );
  XNOR2_X1 U16035 ( .A(n14147), .B(n6680), .ZN(n14150) );
  INV_X1 U16036 ( .A(n14148), .ZN(n14149) );
  AOI21_X1 U16037 ( .B1(n14150), .B2(n14784), .A(n14149), .ZN(n14245) );
  INV_X1 U16038 ( .A(n14151), .ZN(n14152) );
  AOI211_X1 U16039 ( .C1(n14243), .C2(n14153), .A(n14789), .B(n14152), .ZN(
        n14242) );
  AOI22_X1 U16040 ( .A1(n14242), .A2(n14155), .B1(n14728), .B2(n14154), .ZN(
        n14156) );
  AOI21_X1 U16041 ( .B1(n14245), .B2(n14156), .A(n14739), .ZN(n14157) );
  INV_X1 U16042 ( .A(n14157), .ZN(n14158) );
  OAI211_X1 U16043 ( .C1(n14246), .C2(n14160), .A(n14159), .B(n14158), .ZN(
        P1_U3276) );
  OAI211_X1 U16044 ( .C1(n14164), .C2(n14799), .A(n14163), .B(n14162), .ZN(
        n14256) );
  MUX2_X1 U16045 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14256), .S(n14819), .Z(
        P1_U3558) );
  NAND2_X1 U16046 ( .A1(n14165), .A2(n14803), .ZN(n14173) );
  OAI211_X1 U16047 ( .C1(n14169), .C2(n14799), .A(n14168), .B(n14167), .ZN(
        n14170) );
  AOI21_X1 U16048 ( .B1(n14171), .B2(n14730), .A(n14170), .ZN(n14172) );
  NAND2_X1 U16049 ( .A1(n14174), .A2(n14786), .ZN(n14176) );
  MUX2_X1 U16050 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14258), .S(n14819), .Z(
        P1_U3556) );
  OAI21_X1 U16051 ( .B1(n14179), .B2(n14799), .A(n14178), .ZN(n14180) );
  OAI21_X1 U16052 ( .B1(n14184), .B2(n14769), .A(n14183), .ZN(n14259) );
  MUX2_X1 U16053 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14259), .S(n14819), .Z(
        P1_U3555) );
  OAI211_X1 U16054 ( .C1(n14187), .C2(n14799), .A(n14186), .B(n14185), .ZN(
        n14188) );
  AOI21_X1 U16055 ( .B1(n14189), .B2(n14784), .A(n14188), .ZN(n14190) );
  OAI21_X1 U16056 ( .B1(n14191), .B2(n14769), .A(n14190), .ZN(n14260) );
  MUX2_X1 U16057 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14260), .S(n14819), .Z(
        P1_U3554) );
  OAI21_X1 U16058 ( .B1(n14193), .B2(n14799), .A(n14192), .ZN(n14194) );
  AOI211_X1 U16059 ( .C1(n14196), .C2(n14803), .A(n14195), .B(n14194), .ZN(
        n14197) );
  OAI21_X1 U16060 ( .B1(n14795), .B2(n14198), .A(n14197), .ZN(n14261) );
  MUX2_X1 U16061 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14261), .S(n14819), .Z(
        P1_U3553) );
  AOI21_X1 U16062 ( .B1(n14786), .B2(n14200), .A(n14199), .ZN(n14201) );
  OAI211_X1 U16063 ( .C1(n14203), .C2(n14745), .A(n14202), .B(n14201), .ZN(
        n14262) );
  MUX2_X1 U16064 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14262), .S(n14819), .Z(
        P1_U3552) );
  OAI21_X1 U16065 ( .B1(n14205), .B2(n14799), .A(n14204), .ZN(n14206) );
  AOI211_X1 U16066 ( .C1(n14208), .C2(n14784), .A(n14207), .B(n14206), .ZN(
        n14209) );
  OAI21_X1 U16067 ( .B1(n14210), .B2(n14769), .A(n14209), .ZN(n14263) );
  MUX2_X1 U16068 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14263), .S(n14819), .Z(
        P1_U3551) );
  AOI21_X1 U16069 ( .B1(n14786), .B2(n14212), .A(n14211), .ZN(n14213) );
  OAI211_X1 U16070 ( .C1(n14215), .C2(n14769), .A(n14214), .B(n14213), .ZN(
        n14264) );
  MUX2_X1 U16071 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14264), .S(n14819), .Z(
        P1_U3550) );
  OAI211_X1 U16072 ( .C1(n14218), .C2(n14799), .A(n14217), .B(n14216), .ZN(
        n14219) );
  AOI21_X1 U16073 ( .B1(n14220), .B2(n14784), .A(n14219), .ZN(n14221) );
  OAI21_X1 U16074 ( .B1(n14222), .B2(n14769), .A(n14221), .ZN(n14265) );
  MUX2_X1 U16075 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14265), .S(n14819), .Z(
        P1_U3549) );
  OAI211_X1 U16076 ( .C1(n14225), .C2(n14799), .A(n14224), .B(n14223), .ZN(
        n14226) );
  AOI21_X1 U16077 ( .B1(n14227), .B2(n14803), .A(n14226), .ZN(n14228) );
  OAI21_X1 U16078 ( .B1(n14795), .B2(n14229), .A(n14228), .ZN(n14266) );
  MUX2_X1 U16079 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14266), .S(n14819), .Z(
        P1_U3548) );
  NAND2_X1 U16080 ( .A1(n14230), .A2(n14803), .ZN(n14235) );
  AOI211_X1 U16081 ( .C1(n14786), .C2(n14233), .A(n14232), .B(n14231), .ZN(
        n14234) );
  OAI211_X1 U16082 ( .C1(n14795), .C2(n14236), .A(n14235), .B(n14234), .ZN(
        n14267) );
  MUX2_X1 U16083 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14267), .S(n14819), .Z(
        P1_U3547) );
  AOI21_X1 U16084 ( .B1(n14786), .B2(n14238), .A(n14237), .ZN(n14239) );
  OAI211_X1 U16085 ( .C1(n14745), .C2(n14241), .A(n14240), .B(n14239), .ZN(
        n14268) );
  MUX2_X1 U16086 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14268), .S(n14819), .Z(
        P1_U3546) );
  AOI21_X1 U16087 ( .B1(n14786), .B2(n14243), .A(n14242), .ZN(n14244) );
  OAI211_X1 U16088 ( .C1(n14246), .C2(n14769), .A(n14245), .B(n14244), .ZN(
        n14269) );
  MUX2_X1 U16089 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14269), .S(n14819), .Z(
        P1_U3545) );
  NAND2_X1 U16090 ( .A1(n14247), .A2(n14730), .ZN(n14249) );
  OAI211_X1 U16091 ( .C1(n6857), .C2(n14799), .A(n14249), .B(n14248), .ZN(
        n14250) );
  AOI21_X1 U16092 ( .B1(n14251), .B2(n14803), .A(n14250), .ZN(n14252) );
  OAI21_X1 U16093 ( .B1(n14795), .B2(n14253), .A(n14252), .ZN(n14270) );
  MUX2_X1 U16094 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n14270), .S(n14819), .Z(
        P1_U3541) );
  MUX2_X1 U16095 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14254), .S(n14819), .Z(
        P1_U3528) );
  MUX2_X1 U16096 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14256), .S(n14807), .Z(
        P1_U3526) );
  MUX2_X1 U16097 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14258), .S(n14807), .Z(
        P1_U3524) );
  MUX2_X1 U16098 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14259), .S(n14807), .Z(
        P1_U3523) );
  MUX2_X1 U16099 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14260), .S(n14807), .Z(
        P1_U3522) );
  MUX2_X1 U16100 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14261), .S(n14807), .Z(
        P1_U3521) );
  MUX2_X1 U16101 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14262), .S(n14807), .Z(
        P1_U3520) );
  MUX2_X1 U16102 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14263), .S(n14807), .Z(
        P1_U3519) );
  MUX2_X1 U16103 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14264), .S(n14807), .Z(
        P1_U3518) );
  MUX2_X1 U16104 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14265), .S(n14807), .Z(
        P1_U3517) );
  MUX2_X1 U16105 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14266), .S(n14807), .Z(
        P1_U3516) );
  MUX2_X1 U16106 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14267), .S(n14807), .Z(
        P1_U3515) );
  MUX2_X1 U16107 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14268), .S(n14807), .Z(
        P1_U3513) );
  MUX2_X1 U16108 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14269), .S(n14807), .Z(
        P1_U3510) );
  MUX2_X1 U16109 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n14270), .S(n14807), .Z(
        P1_U3498) );
  NOR4_X1 U16110 ( .A1(n14273), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14272), .A4(
        P1_U3086), .ZN(n14274) );
  AOI21_X1 U16111 ( .B1(n14275), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14274), 
        .ZN(n14276) );
  OAI21_X1 U16112 ( .B1(n14277), .B2(n14286), .A(n14276), .ZN(P1_U3324) );
  OAI222_X1 U16113 ( .A1(P1_U3086), .A2(n14280), .B1(n14286), .B2(n14279), 
        .C1(n14278), .C2(n6454), .ZN(P1_U3329) );
  OAI222_X1 U16114 ( .A1(n6454), .A2(n14283), .B1(n14286), .B2(n14282), .C1(
        P1_U3086), .C2(n14281), .ZN(P1_U3330) );
  OAI222_X1 U16115 ( .A1(n6454), .A2(n14287), .B1(n14286), .B2(n14285), .C1(
        P1_U3086), .C2(n14284), .ZN(P1_U3331) );
  MUX2_X1 U16116 ( .A(n9565), .B(n14288), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16117 ( .A(n14289), .ZN(n14290) );
  MUX2_X1 U16118 ( .A(n14290), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16119 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14454) );
  INV_X1 U16120 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U16121 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P3_ADDR_REG_16__SCAN_IN), 
        .B1(n14291), .B2(n14320), .ZN(n14374) );
  INV_X1 U16122 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14695) );
  XNOR2_X1 U16123 ( .A(n14318), .B(n14695), .ZN(n14321) );
  INV_X1 U16124 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14316) );
  INV_X1 U16125 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14312) );
  XOR2_X1 U16126 ( .A(n14312), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14326) );
  INV_X1 U16127 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14310) );
  INV_X1 U16128 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14306) );
  XOR2_X1 U16129 ( .A(n14306), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14328) );
  INV_X1 U16130 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14304) );
  NAND2_X1 U16131 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n14331), .ZN(n14292) );
  INV_X1 U16132 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14293) );
  INV_X1 U16133 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14295) );
  NOR2_X1 U16134 ( .A1(n14296), .A2(n14295), .ZN(n14298) );
  NOR2_X1 U16135 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14347), .ZN(n14301) );
  INV_X1 U16136 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14300) );
  NOR2_X1 U16137 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14302), .ZN(n14303) );
  XOR2_X1 U16138 ( .A(n14302), .B(P3_ADDR_REG_7__SCAN_IN), .Z(n14351) );
  XOR2_X1 U16139 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n14355) );
  NAND2_X1 U16140 ( .A1(n14328), .A2(n14327), .ZN(n14305) );
  NOR2_X1 U16141 ( .A1(n6808), .A2(n14307), .ZN(n14308) );
  XNOR2_X1 U16142 ( .A(n14310), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n14363) );
  NAND2_X1 U16143 ( .A1(n14326), .A2(n14325), .ZN(n14311) );
  XOR2_X1 U16144 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14367) );
  XNOR2_X1 U16145 ( .A(n14316), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14323) );
  NAND2_X1 U16146 ( .A1(n14321), .A2(n14322), .ZN(n14317) );
  XNOR2_X1 U16147 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14376), .ZN(n14377) );
  XOR2_X1 U16148 ( .A(n14454), .B(n14377), .Z(n14444) );
  XOR2_X1 U16149 ( .A(n14322), .B(n14321), .Z(n14640) );
  XOR2_X1 U16150 ( .A(n14324), .B(n14323), .Z(n14372) );
  XOR2_X1 U16151 ( .A(n14328), .B(n14327), .Z(n14359) );
  INV_X1 U16152 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14853) );
  NOR2_X1 U16153 ( .A1(n14330), .A2(n14853), .ZN(n14341) );
  XNOR2_X1 U16154 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n14331), .ZN(n14332) );
  XNOR2_X1 U16155 ( .A(n14332), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n14401) );
  XOR2_X1 U16156 ( .A(n14335), .B(n14333), .Z(n14336) );
  NOR2_X1 U16157 ( .A1(n14336), .A2(n14334), .ZN(n14337) );
  OAI21_X1 U16158 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9511), .A(n14335), .ZN(
        n15140) );
  NAND2_X1 U16159 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15140), .ZN(n15150) );
  XOR2_X1 U16160 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n14336), .Z(n15149) );
  NOR2_X1 U16161 ( .A1(n15150), .A2(n15149), .ZN(n15148) );
  NAND2_X1 U16162 ( .A1(n14401), .A2(n14400), .ZN(n14338) );
  NOR2_X1 U16163 ( .A1(n14401), .A2(n14400), .ZN(n14399) );
  XOR2_X1 U16164 ( .A(n14339), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15145) );
  NOR2_X1 U16165 ( .A1(n15146), .A2(n15145), .ZN(n14340) );
  NAND2_X1 U16166 ( .A1(n15146), .A2(n15145), .ZN(n15144) );
  OAI21_X1 U16167 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14340), .A(n15144), .ZN(
        n15135) );
  NOR2_X1 U16168 ( .A1(n15136), .A2(n15135), .ZN(n15134) );
  NAND2_X1 U16169 ( .A1(n14343), .A2(n14344), .ZN(n14345) );
  INV_X1 U16170 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15138) );
  NOR2_X1 U16171 ( .A1(n14346), .A2(n6682), .ZN(n14350) );
  XOR2_X1 U16172 ( .A(n14347), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14349) );
  XNOR2_X1 U16173 ( .A(n14349), .B(n14348), .ZN(n14411) );
  NOR2_X1 U16174 ( .A1(n14412), .A2(n14411), .ZN(n14410) );
  INV_X1 U16175 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14881) );
  NOR2_X1 U16176 ( .A1(n14352), .A2(n14881), .ZN(n14353) );
  XNOR2_X1 U16177 ( .A(n14351), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15143) );
  XNOR2_X1 U16178 ( .A(n14355), .B(n14354), .ZN(n14357) );
  NAND2_X1 U16179 ( .A1(n14356), .A2(n14357), .ZN(n14358) );
  NAND2_X1 U16180 ( .A1(n14358), .A2(n14419), .ZN(n14360) );
  NOR2_X1 U16181 ( .A1(n14359), .A2(n14360), .ZN(n14361) );
  XNOR2_X1 U16182 ( .A(n14360), .B(n14359), .ZN(n14427) );
  NOR2_X1 U16183 ( .A1(n14428), .A2(n14427), .ZN(n14426) );
  INV_X1 U16184 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15105) );
  XOR2_X1 U16185 ( .A(n15105), .B(n14362), .Z(n14431) );
  XOR2_X1 U16186 ( .A(n14364), .B(n14363), .Z(n14365) );
  INV_X1 U16187 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14896) );
  NAND2_X1 U16188 ( .A1(n14366), .A2(n14365), .ZN(n14623) );
  XOR2_X1 U16189 ( .A(n14368), .B(n14367), .Z(n14369) );
  INV_X1 U16190 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14632) );
  NAND2_X1 U16191 ( .A1(n6480), .A2(n14369), .ZN(n14631) );
  NAND2_X1 U16192 ( .A1(n14632), .A2(n14631), .ZN(n14628) );
  INV_X1 U16193 ( .A(n14628), .ZN(n14370) );
  INV_X1 U16194 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14637) );
  NAND2_X1 U16195 ( .A1(n14372), .A2(n14371), .ZN(n14636) );
  XNOR2_X1 U16196 ( .A(n14374), .B(n14373), .ZN(n14642) );
  NAND2_X1 U16197 ( .A1(n14444), .A2(n14443), .ZN(n14375) );
  NOR2_X1 U16198 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14376), .ZN(n14379) );
  NOR2_X1 U16199 ( .A1(n14454), .A2(n14377), .ZN(n14378) );
  NOR2_X1 U16200 ( .A1(n14379), .A2(n14378), .ZN(n14382) );
  XOR2_X1 U16201 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14381) );
  XOR2_X1 U16202 ( .A(n14382), .B(n14381), .Z(n14390) );
  NOR2_X1 U16203 ( .A1(n14391), .A2(n14390), .ZN(n14380) );
  NAND2_X1 U16204 ( .A1(n14391), .A2(n14390), .ZN(n14389) );
  OAI21_X1 U16205 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n14380), .A(n14389), 
        .ZN(n14388) );
  NOR2_X1 U16206 ( .A1(n14382), .A2(n14381), .ZN(n14383) );
  AOI21_X1 U16207 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n13929), .A(n14383), 
        .ZN(n14386) );
  XNOR2_X1 U16208 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n14384) );
  XNOR2_X1 U16209 ( .A(n14384), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14385) );
  XNOR2_X1 U16210 ( .A(n14386), .B(n14385), .ZN(n14387) );
  XNOR2_X1 U16211 ( .A(n14388), .B(n14387), .ZN(SUB_1596_U4) );
  OAI21_X1 U16212 ( .B1(n14391), .B2(n14390), .A(n14389), .ZN(n14392) );
  XNOR2_X1 U16213 ( .A(n14392), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16214 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14393) );
  OAI21_X1 U16215 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14393), 
        .ZN(U28) );
  AOI21_X1 U16216 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14394) );
  OAI21_X1 U16217 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14394), 
        .ZN(U29) );
  INV_X1 U16218 ( .A(n14395), .ZN(n14396) );
  AOI22_X1 U16219 ( .A1(n14396), .A2(n14422), .B1(SI_17_), .B2(n14421), .ZN(
        n14397) );
  OAI21_X1 U16220 ( .B1(P3_U3151), .B2(n14398), .A(n14397), .ZN(P3_U3278) );
  AOI21_X1 U16221 ( .B1(n14401), .B2(n14400), .A(n14399), .ZN(n14402) );
  XOR2_X1 U16222 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n14402), .Z(SUB_1596_U61) );
  INV_X1 U16223 ( .A(n14403), .ZN(n14404) );
  AOI22_X1 U16224 ( .A1(n14404), .A2(n14422), .B1(SI_12_), .B2(n14421), .ZN(
        n14405) );
  OAI21_X1 U16225 ( .B1(P3_U3151), .B2(n14406), .A(n14405), .ZN(P3_U3283) );
  AOI22_X1 U16226 ( .A1(n14407), .A2(n14422), .B1(SI_13_), .B2(n14421), .ZN(
        n14408) );
  OAI21_X1 U16227 ( .B1(P3_U3151), .B2(n14409), .A(n14408), .ZN(P3_U3282) );
  AOI21_X1 U16228 ( .B1(n14412), .B2(n14411), .A(n14410), .ZN(SUB_1596_U57) );
  AOI22_X1 U16229 ( .A1(n14413), .A2(n14422), .B1(SI_15_), .B2(n14421), .ZN(
        n14414) );
  OAI21_X1 U16230 ( .B1(P3_U3151), .B2(n14415), .A(n14414), .ZN(P3_U3280) );
  AOI22_X1 U16231 ( .A1(n14416), .A2(n14422), .B1(SI_16_), .B2(n14421), .ZN(
        n14417) );
  OAI21_X1 U16232 ( .B1(P3_U3151), .B2(n14418), .A(n14417), .ZN(P3_U3279) );
  OAI21_X1 U16233 ( .B1(n14420), .B2(n9846), .A(n14419), .ZN(SUB_1596_U55) );
  AOI22_X1 U16234 ( .A1(n14423), .A2(n14422), .B1(SI_18_), .B2(n14421), .ZN(
        n14424) );
  OAI21_X1 U16235 ( .B1(P3_U3151), .B2(n14425), .A(n14424), .ZN(P3_U3277) );
  AOI21_X1 U16236 ( .B1(n14428), .B2(n14427), .A(n14426), .ZN(SUB_1596_U54) );
  OAI21_X1 U16237 ( .B1(n14431), .B2(n14430), .A(n14429), .ZN(n14432) );
  XNOR2_X1 U16238 ( .A(n14432), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  NOR2_X1 U16239 ( .A1(n14433), .A2(n14795), .ZN(n14438) );
  INV_X1 U16240 ( .A(n14564), .ZN(n14436) );
  OAI211_X1 U16241 ( .C1(n14436), .C2(n14799), .A(n14435), .B(n14434), .ZN(
        n14437) );
  AOI211_X1 U16242 ( .C1(n14439), .C2(n14803), .A(n14438), .B(n14437), .ZN(
        n14441) );
  INV_X1 U16243 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14440) );
  AOI22_X1 U16244 ( .A1(n14807), .A2(n14441), .B1(n14440), .B2(n14805), .ZN(
        P1_U3495) );
  AOI22_X1 U16245 ( .A1(n14819), .A2(n14441), .B1(n9684), .B2(n14816), .ZN(
        P1_U3540) );
  AOI21_X1 U16246 ( .B1(n14444), .B2(n14443), .A(n14442), .ZN(n14445) );
  XOR2_X1 U16247 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14445), .Z(SUB_1596_U63)
         );
  AOI21_X1 U16248 ( .B1(n14448), .B2(n14447), .A(n14446), .ZN(n14462) );
  OAI21_X1 U16249 ( .B1(n14450), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14449), 
        .ZN(n14460) );
  NAND2_X1 U16250 ( .A1(n15102), .A2(n14451), .ZN(n14453) );
  OAI211_X1 U16251 ( .C1(n14454), .C2(n15106), .A(n14453), .B(n14452), .ZN(
        n14459) );
  AOI211_X1 U16252 ( .C1(n14457), .C2(n14456), .A(n15096), .B(n14455), .ZN(
        n14458) );
  AOI211_X1 U16253 ( .C1(n15086), .C2(n14460), .A(n14459), .B(n14458), .ZN(
        n14461) );
  OAI21_X1 U16254 ( .B1(n14462), .B2(n15091), .A(n14461), .ZN(P3_U3199) );
  AOI22_X1 U16255 ( .A1(n14468), .A2(n14463), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15119), .ZN(n14464) );
  NAND2_X1 U16256 ( .A1(n14465), .A2(n14464), .ZN(P3_U3203) );
  AOI21_X1 U16257 ( .B1(n14468), .B2(n14467), .A(n14466), .ZN(n14477) );
  AOI22_X1 U16258 ( .A1(n15133), .A2(n14477), .B1(n14469), .B2(n15131), .ZN(
        P3_U3489) );
  NOR2_X1 U16259 ( .A1(n14471), .A2(n14470), .ZN(n14473) );
  AOI211_X1 U16260 ( .C1(n14475), .C2(n14474), .A(n14473), .B(n14472), .ZN(
        n14479) );
  AOI22_X1 U16261 ( .A1(n15133), .A2(n14479), .B1(n14476), .B2(n15131), .ZN(
        P3_U3471) );
  INV_X1 U16262 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14478) );
  AOI22_X1 U16263 ( .A1(n15127), .A2(n14478), .B1(n14477), .B2(n15129), .ZN(
        P3_U3457) );
  INV_X1 U16264 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14480) );
  AOI22_X1 U16265 ( .A1(n15127), .A2(n14480), .B1(n14479), .B2(n15129), .ZN(
        P3_U3426) );
  AOI22_X1 U16266 ( .A1(n14484), .A2(n14483), .B1(n14482), .B2(n14481), .ZN(
        n14497) );
  AOI21_X1 U16267 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(n14489) );
  OAI222_X1 U16268 ( .A1(n14491), .A2(n14497), .B1(n14490), .B2(n14489), .C1(
        n14488), .C2(n14523), .ZN(n14492) );
  INV_X1 U16269 ( .A(n14492), .ZN(n14494) );
  OAI211_X1 U16270 ( .C1(n14495), .C2(n14500), .A(n14494), .B(n14493), .ZN(
        P2_U3187) );
  XNOR2_X1 U16271 ( .A(n14496), .B(n14505), .ZN(n14499) );
  INV_X1 U16272 ( .A(n14497), .ZN(n14498) );
  AOI21_X1 U16273 ( .B1(n14499), .B2(n14535), .A(n14498), .ZN(n14522) );
  INV_X1 U16274 ( .A(n14500), .ZN(n14501) );
  AOI222_X1 U16275 ( .A1(n14503), .A2(n14502), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n14951), .C1(n14941), .C2(n14501), .ZN(n14512) );
  XOR2_X1 U16276 ( .A(n14504), .B(n14505), .Z(n14525) );
  INV_X1 U16277 ( .A(n14506), .ZN(n14507) );
  OAI211_X1 U16278 ( .C1(n14523), .C2(n6590), .A(n14507), .B(n6452), .ZN(
        n14521) );
  INV_X1 U16279 ( .A(n14521), .ZN(n14508) );
  AOI22_X1 U16280 ( .A1(n14525), .A2(n14510), .B1(n14509), .B2(n14508), .ZN(
        n14511) );
  OAI211_X1 U16281 ( .C1(n14951), .C2(n14522), .A(n14512), .B(n14511), .ZN(
        P2_U3251) );
  INV_X1 U16282 ( .A(n14513), .ZN(n14520) );
  OAI211_X1 U16283 ( .C1(n14516), .C2(n14986), .A(n14515), .B(n14514), .ZN(
        n14519) );
  INV_X1 U16284 ( .A(n14517), .ZN(n14518) );
  AOI211_X1 U16285 ( .C1(n14520), .C2(n14983), .A(n14519), .B(n14518), .ZN(
        n14545) );
  AOI22_X1 U16286 ( .A1(n15002), .A2(n14545), .B1(n14913), .B2(n14999), .ZN(
        P2_U3514) );
  OAI211_X1 U16287 ( .C1(n14523), .C2(n14986), .A(n14522), .B(n14521), .ZN(
        n14524) );
  AOI21_X1 U16288 ( .B1(n14983), .B2(n14525), .A(n14524), .ZN(n14547) );
  AOI22_X1 U16289 ( .A1(n15002), .A2(n14547), .B1(n14526), .B2(n14999), .ZN(
        P2_U3513) );
  OAI211_X1 U16290 ( .C1(n6877), .C2(n14986), .A(n14529), .B(n14528), .ZN(
        n14533) );
  NOR2_X1 U16291 ( .A1(n14531), .A2(n14530), .ZN(n14532) );
  AOI211_X1 U16292 ( .C1(n14535), .C2(n14534), .A(n14533), .B(n14532), .ZN(
        n14549) );
  AOI22_X1 U16293 ( .A1(n15002), .A2(n14549), .B1(n14536), .B2(n14999), .ZN(
        P2_U3512) );
  OAI21_X1 U16294 ( .B1(n14538), .B2(n14986), .A(n14537), .ZN(n14539) );
  AOI21_X1 U16295 ( .B1(n14540), .B2(n8957), .A(n14539), .ZN(n14541) );
  INV_X1 U16296 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14543) );
  AOI22_X1 U16297 ( .A1(n15002), .A2(n14551), .B1(n14543), .B2(n14999), .ZN(
        P2_U3511) );
  AOI22_X1 U16298 ( .A1(n10105), .A2(n14545), .B1(n14544), .B2(n14991), .ZN(
        P2_U3475) );
  INV_X1 U16299 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14546) );
  AOI22_X1 U16300 ( .A1(n10105), .A2(n14547), .B1(n14546), .B2(n14991), .ZN(
        P2_U3472) );
  INV_X1 U16301 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14548) );
  AOI22_X1 U16302 ( .A1(n10105), .A2(n14549), .B1(n14548), .B2(n14991), .ZN(
        P2_U3469) );
  INV_X1 U16303 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14550) );
  AOI22_X1 U16304 ( .A1(n10105), .A2(n14551), .B1(n14550), .B2(n14991), .ZN(
        P2_U3466) );
  INV_X1 U16305 ( .A(n14552), .ZN(n14555) );
  OAI21_X1 U16306 ( .B1(n14555), .B2(n14554), .A(n14553), .ZN(n14557) );
  NAND2_X1 U16307 ( .A1(n14557), .A2(n14556), .ZN(n14558) );
  AOI222_X1 U16308 ( .A1(n14599), .A2(n14578), .B1(n14558), .B2(n14576), .C1(
        n14600), .C2(n14657), .ZN(n14560) );
  OAI211_X1 U16309 ( .C1(n14659), .C2(n14561), .A(n14560), .B(n14559), .ZN(
        P1_U3215) );
  XNOR2_X1 U16310 ( .A(n14563), .B(n14562), .ZN(n14565) );
  AOI222_X1 U16311 ( .A1(n14566), .A2(n14578), .B1(n14576), .B2(n14565), .C1(
        n14564), .C2(n14657), .ZN(n14568) );
  OAI211_X1 U16312 ( .C1(n14659), .C2(n14569), .A(n14568), .B(n14567), .ZN(
        P1_U3224) );
  INV_X1 U16313 ( .A(n13559), .ZN(n14572) );
  OAI21_X1 U16314 ( .B1(n14572), .B2(n14571), .A(n14570), .ZN(n14574) );
  NAND2_X1 U16315 ( .A1(n14574), .A2(n14573), .ZN(n14577) );
  AOI222_X1 U16316 ( .A1(n14582), .A2(n14578), .B1(n14577), .B2(n14576), .C1(
        n14575), .C2(n14657), .ZN(n14580) );
  OAI211_X1 U16317 ( .C1(n14659), .C2(n14581), .A(n14580), .B(n14579), .ZN(
        P1_U3226) );
  INV_X1 U16318 ( .A(n14582), .ZN(n14583) );
  OAI211_X1 U16319 ( .C1(n14585), .C2(n14799), .A(n14584), .B(n14583), .ZN(
        n14588) );
  NOR2_X1 U16320 ( .A1(n14586), .A2(n14795), .ZN(n14587) );
  AOI211_X1 U16321 ( .C1(n14589), .C2(n14803), .A(n14588), .B(n14587), .ZN(
        n14614) );
  AOI22_X1 U16322 ( .A1(n14819), .A2(n14614), .B1(n14590), .B2(n14816), .ZN(
        P1_U3544) );
  NOR2_X1 U16323 ( .A1(n14591), .A2(n14795), .ZN(n14596) );
  OAI211_X1 U16324 ( .C1(n14594), .C2(n14799), .A(n14593), .B(n14592), .ZN(
        n14595) );
  AOI211_X1 U16325 ( .C1(n14597), .C2(n14803), .A(n14596), .B(n14595), .ZN(
        n14616) );
  AOI22_X1 U16326 ( .A1(n14819), .A2(n14616), .B1(n14684), .B2(n14816), .ZN(
        P1_U3543) );
  INV_X1 U16327 ( .A(n14598), .ZN(n14605) );
  AOI21_X1 U16328 ( .B1(n14600), .B2(n14786), .A(n14599), .ZN(n14602) );
  OAI211_X1 U16329 ( .C1(n14603), .C2(n14769), .A(n14602), .B(n14601), .ZN(
        n14604) );
  AOI21_X1 U16330 ( .B1(n14605), .B2(n14784), .A(n14604), .ZN(n14618) );
  AOI22_X1 U16331 ( .A1(n14819), .A2(n14618), .B1(n14606), .B2(n14816), .ZN(
        P1_U3542) );
  OAI22_X1 U16332 ( .A1(n14608), .A2(n14789), .B1(n14607), .B2(n14799), .ZN(
        n14609) );
  AOI211_X1 U16333 ( .C1(n14611), .C2(n14803), .A(n14610), .B(n14609), .ZN(
        n14620) );
  AOI22_X1 U16334 ( .A1(n14819), .A2(n14620), .B1(n14612), .B2(n14816), .ZN(
        P1_U3539) );
  INV_X1 U16335 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14613) );
  AOI22_X1 U16336 ( .A1(n14807), .A2(n14614), .B1(n14613), .B2(n14805), .ZN(
        P1_U3507) );
  INV_X1 U16337 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14615) );
  AOI22_X1 U16338 ( .A1(n14807), .A2(n14616), .B1(n14615), .B2(n14805), .ZN(
        P1_U3504) );
  INV_X1 U16339 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14617) );
  AOI22_X1 U16340 ( .A1(n14807), .A2(n14618), .B1(n14617), .B2(n14805), .ZN(
        P1_U3501) );
  INV_X1 U16341 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14619) );
  AOI22_X1 U16342 ( .A1(n14807), .A2(n14620), .B1(n14619), .B2(n14805), .ZN(
        P1_U3492) );
  OAI222_X1 U16343 ( .A1(n14896), .A2(n14623), .B1(n14896), .B2(n7326), .C1(
        n14622), .C2(n14621), .ZN(SUB_1596_U69) );
  OAI21_X1 U16344 ( .B1(n14626), .B2(n14625), .A(n14624), .ZN(n14627) );
  XNOR2_X1 U16345 ( .A(n14627), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  INV_X1 U16346 ( .A(n14629), .ZN(n14630) );
  OAI222_X1 U16347 ( .A1(n14632), .A2(n14631), .B1(n14632), .B2(n14630), .C1(
        n14629), .C2(n14628), .ZN(SUB_1596_U67) );
  OAI222_X1 U16348 ( .A1(n14637), .A2(n14636), .B1(n14637), .B2(n14635), .C1(
        n14634), .C2(n14633), .ZN(SUB_1596_U66) );
  AOI21_X1 U16349 ( .B1(n14640), .B2(n14639), .A(n14638), .ZN(n14641) );
  XOR2_X1 U16350 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14641), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16351 ( .B1(n14643), .B2(n14642), .A(n6565), .ZN(n14644) );
  XOR2_X1 U16352 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14644), .Z(SUB_1596_U64)
         );
  AOI22_X1 U16353 ( .A1(n13551), .A2(n14647), .B1(n14646), .B2(n14645), .ZN(
        n14707) );
  OAI21_X1 U16354 ( .B1(n14649), .B2(n14707), .A(n14648), .ZN(n14655) );
  AOI211_X1 U16355 ( .C1(n14653), .C2(n14652), .A(n14651), .B(n14650), .ZN(
        n14654) );
  AOI211_X1 U16356 ( .C1(n14657), .C2(n6457), .A(n14655), .B(n14654), .ZN(
        n14658) );
  OAI21_X1 U16357 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(n14659), .A(n14658), .ZN(
        P1_U3218) );
  MUX2_X1 U16358 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10485), .S(n14665), .Z(
        n14660) );
  NAND3_X1 U16359 ( .A1(n14662), .A2(n14661), .A3(n14660), .ZN(n14663) );
  NAND3_X1 U16360 ( .A1(n14690), .A2(n14664), .A3(n14663), .ZN(n14677) );
  MUX2_X1 U16361 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n14811), .S(n14665), .Z(
        n14666) );
  NAND3_X1 U16362 ( .A1(n14668), .A2(n14667), .A3(n14666), .ZN(n14669) );
  NAND3_X1 U16363 ( .A1(n14689), .A2(n14670), .A3(n14669), .ZN(n14676) );
  NAND2_X1 U16364 ( .A1(n14686), .A2(n14671), .ZN(n14675) );
  AOI21_X1 U16365 ( .B1(n14673), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14672), .ZN(
        n14674) );
  AND4_X1 U16366 ( .A1(n14677), .A2(n14676), .A3(n14675), .A4(n14674), .ZN(
        n14679) );
  NAND2_X1 U16367 ( .A1(n14679), .A2(n14678), .ZN(P1_U3247) );
  AOI21_X1 U16368 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14681), .A(n14680), 
        .ZN(n14682) );
  INV_X1 U16369 ( .A(n14682), .ZN(n14691) );
  OAI21_X1 U16370 ( .B1(n14685), .B2(n14684), .A(n14683), .ZN(n14688) );
  AOI222_X1 U16371 ( .A1(n14691), .A2(n14690), .B1(n14689), .B2(n14688), .C1(
        n14687), .C2(n14686), .ZN(n14693) );
  OAI211_X1 U16372 ( .C1(n14695), .C2(n14694), .A(n14693), .B(n14692), .ZN(
        P1_U3258) );
  AOI222_X1 U16373 ( .A1(n14698), .A2(n14735), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n14697), .C1(n14728), .C2(n14696), .ZN(n14702) );
  AOI22_X1 U16374 ( .A1(n14700), .A2(n14718), .B1(n14717), .B2(n14699), .ZN(
        n14701) );
  OAI211_X1 U16375 ( .C1(n14739), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        P1_U3284) );
  XNOR2_X1 U16376 ( .A(n14704), .B(n14706), .ZN(n14764) );
  XOR2_X1 U16377 ( .A(n14705), .B(n14706), .Z(n14708) );
  OAI21_X1 U16378 ( .B1(n14708), .B2(n14795), .A(n14707), .ZN(n14709) );
  AOI21_X1 U16379 ( .B1(n14723), .B2(n14764), .A(n14709), .ZN(n14761) );
  AOI22_X1 U16380 ( .A1(n14739), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n14728), 
        .B2(n14710), .ZN(n14711) );
  OAI21_X1 U16381 ( .B1(n14712), .B2(n14760), .A(n14711), .ZN(n14713) );
  INV_X1 U16382 ( .A(n14713), .ZN(n14720) );
  OAI211_X1 U16383 ( .C1(n14715), .C2(n14760), .A(n14714), .B(n14730), .ZN(
        n14759) );
  INV_X1 U16384 ( .A(n14759), .ZN(n14716) );
  AOI22_X1 U16385 ( .A1(n14764), .A2(n14718), .B1(n14717), .B2(n14716), .ZN(
        n14719) );
  OAI211_X1 U16386 ( .C1(n14739), .C2(n14761), .A(n14720), .B(n14719), .ZN(
        P1_U3290) );
  XNOR2_X1 U16387 ( .A(n10256), .B(n14721), .ZN(n14750) );
  XNOR2_X1 U16388 ( .A(n14722), .B(n10256), .ZN(n14726) );
  NAND2_X1 U16389 ( .A1(n14750), .A2(n14723), .ZN(n14725) );
  OAI211_X1 U16390 ( .C1(n14726), .C2(n14795), .A(n14725), .B(n14724), .ZN(
        n14748) );
  AOI21_X1 U16391 ( .B1(n14727), .B2(n14750), .A(n14748), .ZN(n14738) );
  AOI22_X1 U16392 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n14728), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n14739), .ZN(n14737) );
  OAI211_X1 U16393 ( .C1(n6664), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        n14747) );
  OAI22_X1 U16394 ( .A1(n14739), .A2(n14746), .B1(n14747), .B2(n14732), .ZN(
        n14733) );
  AOI21_X1 U16395 ( .B1(n14735), .B2(n6656), .A(n14733), .ZN(n14736) );
  OAI211_X1 U16396 ( .C1(n14739), .C2(n14738), .A(n14737), .B(n14736), .ZN(
        P1_U3292) );
  AND2_X1 U16397 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14744), .ZN(P1_U3294) );
  AND2_X1 U16398 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14744), .ZN(P1_U3295) );
  AND2_X1 U16399 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14744), .ZN(P1_U3296) );
  NOR2_X1 U16400 ( .A1(n14743), .A2(n14740), .ZN(P1_U3297) );
  AND2_X1 U16401 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14744), .ZN(P1_U3298) );
  AND2_X1 U16402 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14744), .ZN(P1_U3299) );
  AND2_X1 U16403 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14744), .ZN(P1_U3300) );
  NOR2_X1 U16404 ( .A1(n14743), .A2(n14741), .ZN(P1_U3301) );
  AND2_X1 U16405 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14744), .ZN(P1_U3302) );
  AND2_X1 U16406 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14744), .ZN(P1_U3303) );
  AND2_X1 U16407 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14744), .ZN(P1_U3304) );
  AND2_X1 U16408 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14744), .ZN(P1_U3305) );
  AND2_X1 U16409 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14744), .ZN(P1_U3306) );
  AND2_X1 U16410 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14744), .ZN(P1_U3307) );
  AND2_X1 U16411 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14744), .ZN(P1_U3308) );
  AND2_X1 U16412 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14744), .ZN(P1_U3309) );
  AND2_X1 U16413 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14744), .ZN(P1_U3310) );
  AND2_X1 U16414 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14744), .ZN(P1_U3311) );
  AND2_X1 U16415 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14744), .ZN(P1_U3312) );
  AND2_X1 U16416 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14744), .ZN(P1_U3313) );
  AND2_X1 U16417 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14744), .ZN(P1_U3314) );
  AND2_X1 U16418 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14744), .ZN(P1_U3315) );
  AND2_X1 U16419 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14744), .ZN(P1_U3316) );
  AND2_X1 U16420 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14744), .ZN(P1_U3317) );
  AND2_X1 U16421 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14744), .ZN(P1_U3318) );
  AND2_X1 U16422 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14744), .ZN(P1_U3319) );
  AND2_X1 U16423 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14744), .ZN(P1_U3320) );
  AND2_X1 U16424 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14744), .ZN(P1_U3321) );
  NOR2_X1 U16425 ( .A1(n14743), .A2(n14742), .ZN(P1_U3322) );
  AND2_X1 U16426 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14744), .ZN(P1_U3323) );
  INV_X1 U16427 ( .A(n14745), .ZN(n14781) );
  OAI211_X1 U16428 ( .C1(n6664), .C2(n14799), .A(n14747), .B(n14746), .ZN(
        n14749) );
  AOI211_X1 U16429 ( .C1(n14781), .C2(n14750), .A(n14749), .B(n14748), .ZN(
        n14808) );
  INV_X1 U16430 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14751) );
  AOI22_X1 U16431 ( .A1(n14807), .A2(n14808), .B1(n14751), .B2(n14805), .ZN(
        P1_U3462) );
  OAI21_X1 U16432 ( .B1(n14753), .B2(n14799), .A(n14752), .ZN(n14754) );
  AOI21_X1 U16433 ( .B1(n14755), .B2(n14781), .A(n14754), .ZN(n14756) );
  AND2_X1 U16434 ( .A1(n14757), .A2(n14756), .ZN(n14809) );
  INV_X1 U16435 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14758) );
  AOI22_X1 U16436 ( .A1(n14807), .A2(n14809), .B1(n14758), .B2(n14805), .ZN(
        P1_U3465) );
  OAI21_X1 U16437 ( .B1(n14760), .B2(n14799), .A(n14759), .ZN(n14763) );
  INV_X1 U16438 ( .A(n14761), .ZN(n14762) );
  AOI211_X1 U16439 ( .C1(n14781), .C2(n14764), .A(n14763), .B(n14762), .ZN(
        n14810) );
  INV_X1 U16440 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14765) );
  AOI22_X1 U16441 ( .A1(n14807), .A2(n14810), .B1(n14765), .B2(n14805), .ZN(
        P1_U3468) );
  OAI211_X1 U16442 ( .C1(n14768), .C2(n14799), .A(n14767), .B(n14766), .ZN(
        n14773) );
  NOR3_X1 U16443 ( .A1(n14771), .A2(n14770), .A3(n14769), .ZN(n14772) );
  AOI211_X1 U16444 ( .C1(n14784), .C2(n14774), .A(n14773), .B(n14772), .ZN(
        n14812) );
  INV_X1 U16445 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14775) );
  AOI22_X1 U16446 ( .A1(n14807), .A2(n14812), .B1(n14775), .B2(n14805), .ZN(
        P1_U3471) );
  OAI22_X1 U16447 ( .A1(n14777), .A2(n14789), .B1(n14776), .B2(n14799), .ZN(
        n14779) );
  AOI211_X1 U16448 ( .C1(n14781), .C2(n14780), .A(n14779), .B(n14778), .ZN(
        n14814) );
  INV_X1 U16449 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14782) );
  AOI22_X1 U16450 ( .A1(n14807), .A2(n14814), .B1(n14782), .B2(n14805), .ZN(
        P1_U3480) );
  AND3_X1 U16451 ( .A1(n11015), .A2(n14784), .A3(n14783), .ZN(n14792) );
  AOI21_X1 U16452 ( .B1(n14787), .B2(n14786), .A(n14785), .ZN(n14788) );
  OAI21_X1 U16453 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n14791) );
  AOI211_X1 U16454 ( .C1(n14793), .C2(n14803), .A(n14792), .B(n14791), .ZN(
        n14815) );
  INV_X1 U16455 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14794) );
  AOI22_X1 U16456 ( .A1(n14807), .A2(n14815), .B1(n14794), .B2(n14805), .ZN(
        P1_U3483) );
  NOR3_X1 U16457 ( .A1(n6479), .A2(n14796), .A3(n14795), .ZN(n14802) );
  OAI211_X1 U16458 ( .C1(n14800), .C2(n14799), .A(n14798), .B(n14797), .ZN(
        n14801) );
  AOI211_X1 U16459 ( .C1(n14804), .C2(n14803), .A(n14802), .B(n14801), .ZN(
        n14818) );
  INV_X1 U16460 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14806) );
  AOI22_X1 U16461 ( .A1(n14807), .A2(n14818), .B1(n14806), .B2(n14805), .ZN(
        P1_U3489) );
  AOI22_X1 U16462 ( .A1(n14819), .A2(n14808), .B1(n9409), .B2(n14816), .ZN(
        P1_U3529) );
  AOI22_X1 U16463 ( .A1(n14819), .A2(n14809), .B1(n9407), .B2(n14816), .ZN(
        P1_U3530) );
  AOI22_X1 U16464 ( .A1(n14819), .A2(n14810), .B1(n9414), .B2(n14816), .ZN(
        P1_U3531) );
  AOI22_X1 U16465 ( .A1(n14819), .A2(n14812), .B1(n14811), .B2(n14816), .ZN(
        P1_U3532) );
  AOI22_X1 U16466 ( .A1(n14819), .A2(n14814), .B1(n14813), .B2(n14816), .ZN(
        P1_U3535) );
  AOI22_X1 U16467 ( .A1(n14819), .A2(n14815), .B1(n9617), .B2(n14816), .ZN(
        P1_U3536) );
  AOI22_X1 U16468 ( .A1(n14819), .A2(n14818), .B1(n14817), .B2(n14816), .ZN(
        P1_U3538) );
  NOR2_X1 U16469 ( .A1(n14929), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16470 ( .A(n14820), .ZN(n14821) );
  AOI21_X1 U16471 ( .B1(n14900), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14821), .ZN(
        n14825) );
  AOI22_X1 U16472 ( .A1(n14929), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14824) );
  OAI22_X1 U16473 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14862), .B1(n14923), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n14822) );
  OAI21_X1 U16474 ( .B1(n14889), .B2(n14822), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14823) );
  OAI211_X1 U16475 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14825), .A(n14824), .B(
        n14823), .ZN(P2_U3214) );
  AOI22_X1 U16476 ( .A1(n14929), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14838) );
  OAI21_X1 U16477 ( .B1(n14829), .B2(n14828), .A(n14827), .ZN(n14830) );
  INV_X1 U16478 ( .A(n14830), .ZN(n14832) );
  AOI22_X1 U16479 ( .A1(n14900), .A2(n14832), .B1(n14831), .B2(n14889), .ZN(
        n14837) );
  OAI211_X1 U16480 ( .C1(n14835), .C2(n14834), .A(n14931), .B(n14833), .ZN(
        n14836) );
  NAND3_X1 U16481 ( .A1(n14838), .A2(n14837), .A3(n14836), .ZN(P2_U3216) );
  OAI211_X1 U16482 ( .C1(n14841), .C2(n14840), .A(n14900), .B(n14839), .ZN(
        n14846) );
  INV_X1 U16483 ( .A(n14842), .ZN(n14843) );
  AOI21_X1 U16484 ( .B1(n14889), .B2(n14844), .A(n14843), .ZN(n14845) );
  AND2_X1 U16485 ( .A1(n14846), .A2(n14845), .ZN(n14852) );
  AOI211_X1 U16486 ( .C1(n14849), .C2(n14848), .A(n14847), .B(n14862), .ZN(
        n14850) );
  INV_X1 U16487 ( .A(n14850), .ZN(n14851) );
  OAI211_X1 U16488 ( .C1(n14897), .C2(n14853), .A(n14852), .B(n14851), .ZN(
        P2_U3218) );
  OAI211_X1 U16489 ( .C1(n14856), .C2(n14855), .A(n14900), .B(n14854), .ZN(
        n14861) );
  OAI21_X1 U16490 ( .B1(n14937), .B2(n14858), .A(n14857), .ZN(n14859) );
  INV_X1 U16491 ( .A(n14859), .ZN(n14860) );
  AND2_X1 U16492 ( .A1(n14861), .A2(n14860), .ZN(n14868) );
  AOI211_X1 U16493 ( .C1(n14865), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14866) );
  INV_X1 U16494 ( .A(n14866), .ZN(n14867) );
  OAI211_X1 U16495 ( .C1(n14897), .C2(n15138), .A(n14868), .B(n14867), .ZN(
        P2_U3219) );
  OAI211_X1 U16496 ( .C1(n14871), .C2(n14870), .A(n14900), .B(n14869), .ZN(
        n14875) );
  AOI21_X1 U16497 ( .B1(n14889), .B2(n14873), .A(n14872), .ZN(n14874) );
  AND2_X1 U16498 ( .A1(n14875), .A2(n14874), .ZN(n14880) );
  OAI211_X1 U16499 ( .C1(n14878), .C2(n14877), .A(n14876), .B(n14931), .ZN(
        n14879) );
  OAI211_X1 U16500 ( .C1(n14897), .C2(n14881), .A(n14880), .B(n14879), .ZN(
        P2_U3221) );
  OAI211_X1 U16501 ( .C1(n14884), .C2(n14883), .A(n14882), .B(n14900), .ZN(
        n14885) );
  INV_X1 U16502 ( .A(n14885), .ZN(n14886) );
  AOI211_X1 U16503 ( .C1(n14889), .C2(n14888), .A(n14887), .B(n14886), .ZN(
        n14895) );
  OAI21_X1 U16504 ( .B1(n14892), .B2(n14891), .A(n14890), .ZN(n14893) );
  NAND2_X1 U16505 ( .A1(n14893), .A2(n14931), .ZN(n14894) );
  OAI211_X1 U16506 ( .C1(n14897), .C2(n14896), .A(n14895), .B(n14894), .ZN(
        P2_U3225) );
  NOR2_X1 U16507 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7688), .ZN(n14905) );
  NAND2_X1 U16508 ( .A1(n14899), .A2(n14898), .ZN(n14901) );
  NAND2_X1 U16509 ( .A1(n14901), .A2(n14900), .ZN(n14902) );
  NOR2_X1 U16510 ( .A1(n14903), .A2(n14902), .ZN(n14904) );
  AOI211_X1 U16511 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n14929), .A(n14905), 
        .B(n14904), .ZN(n14910) );
  OAI211_X1 U16512 ( .C1(n14908), .C2(n14907), .A(n14906), .B(n14931), .ZN(
        n14909) );
  OAI211_X1 U16513 ( .C1(n14937), .C2(n14911), .A(n14910), .B(n14909), .ZN(
        P2_U3227) );
  NOR2_X1 U16514 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7733), .ZN(n14916) );
  AOI211_X1 U16515 ( .C1(n14914), .C2(n14913), .A(n14912), .B(n14923), .ZN(
        n14915) );
  AOI211_X1 U16516 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n14929), .A(n14916), 
        .B(n14915), .ZN(n14920) );
  OAI211_X1 U16517 ( .C1(n14918), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14931), 
        .B(n14917), .ZN(n14919) );
  OAI211_X1 U16518 ( .C1(n14937), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        P2_U3229) );
  INV_X1 U16519 ( .A(n14922), .ZN(n14928) );
  AOI211_X1 U16520 ( .C1(n14926), .C2(n14925), .A(n14924), .B(n14923), .ZN(
        n14927) );
  AOI211_X1 U16521 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n14929), .A(n14928), 
        .B(n14927), .ZN(n14935) );
  OAI211_X1 U16522 ( .C1(n14933), .C2(n14932), .A(n14931), .B(n14930), .ZN(
        n14934) );
  OAI211_X1 U16523 ( .C1(n14937), .C2(n14936), .A(n14935), .B(n14934), .ZN(
        P2_U3230) );
  INV_X1 U16524 ( .A(n14938), .ZN(n14943) );
  AOI22_X1 U16525 ( .A1(n14941), .A2(n13050), .B1(n14940), .B2(n14939), .ZN(
        n14942) );
  OAI21_X1 U16526 ( .B1(n14943), .B2(n6463), .A(n14942), .ZN(n14944) );
  AOI211_X1 U16527 ( .C1(n14947), .C2(n14946), .A(n14945), .B(n14944), .ZN(
        n14949) );
  AOI22_X1 U16528 ( .A1(n14951), .A2(n14950), .B1(n14949), .B2(n14948), .ZN(
        P2_U3262) );
  NOR2_X1 U16529 ( .A1(n14961), .A2(n14952), .ZN(n14955) );
  AND2_X1 U16530 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14956), .ZN(P2_U3266) );
  AND2_X1 U16531 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14956), .ZN(P2_U3267) );
  AND2_X1 U16532 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14956), .ZN(P2_U3268) );
  AND2_X1 U16533 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14956), .ZN(P2_U3269) );
  AND2_X1 U16534 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14956), .ZN(P2_U3270) );
  NOR2_X1 U16535 ( .A1(n14955), .A2(n14953), .ZN(P2_U3271) );
  AND2_X1 U16536 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14956), .ZN(P2_U3272) );
  AND2_X1 U16537 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14956), .ZN(P2_U3273) );
  AND2_X1 U16538 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14956), .ZN(P2_U3274) );
  AND2_X1 U16539 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14956), .ZN(P2_U3275) );
  AND2_X1 U16540 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14956), .ZN(P2_U3276) );
  AND2_X1 U16541 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14956), .ZN(P2_U3277) );
  AND2_X1 U16542 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14956), .ZN(P2_U3278) );
  AND2_X1 U16543 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14956), .ZN(P2_U3279) );
  AND2_X1 U16544 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14956), .ZN(P2_U3280) );
  AND2_X1 U16545 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14956), .ZN(P2_U3281) );
  NOR2_X1 U16546 ( .A1(n14955), .A2(n14954), .ZN(P2_U3282) );
  AND2_X1 U16547 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14956), .ZN(P2_U3283) );
  AND2_X1 U16548 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14956), .ZN(P2_U3284) );
  AND2_X1 U16549 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14956), .ZN(P2_U3285) );
  AND2_X1 U16550 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14956), .ZN(P2_U3286) );
  AND2_X1 U16551 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14956), .ZN(P2_U3287) );
  AND2_X1 U16552 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14956), .ZN(P2_U3288) );
  AND2_X1 U16553 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14956), .ZN(P2_U3289) );
  AND2_X1 U16554 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14956), .ZN(P2_U3290) );
  AND2_X1 U16555 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14956), .ZN(P2_U3291) );
  AND2_X1 U16556 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14956), .ZN(P2_U3292) );
  AND2_X1 U16557 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14956), .ZN(P2_U3293) );
  AND2_X1 U16558 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14956), .ZN(P2_U3294) );
  AND2_X1 U16559 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14956), .ZN(P2_U3295) );
  AOI22_X1 U16560 ( .A1(n14959), .A2(n14958), .B1(n14957), .B2(n14961), .ZN(
        P2_U3416) );
  AOI21_X1 U16561 ( .B1(n14962), .B2(n14961), .A(n14960), .ZN(P2_U3417) );
  OAI211_X1 U16562 ( .C1(n14965), .C2(n14986), .A(n14964), .B(n14963), .ZN(
        n14966) );
  AOI21_X1 U16563 ( .B1(n14983), .B2(n14967), .A(n14966), .ZN(n14994) );
  INV_X1 U16564 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14968) );
  AOI22_X1 U16565 ( .A1(n10105), .A2(n14994), .B1(n14968), .B2(n14991), .ZN(
        P2_U3448) );
  OAI21_X1 U16566 ( .B1(n14970), .B2(n14986), .A(n14969), .ZN(n14971) );
  AOI21_X1 U16567 ( .B1(n14972), .B2(n8957), .A(n14971), .ZN(n14973) );
  INV_X1 U16568 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14975) );
  AOI22_X1 U16569 ( .A1(n10105), .A2(n14996), .B1(n14975), .B2(n14991), .ZN(
        P2_U3454) );
  OAI21_X1 U16570 ( .B1(n14977), .B2(n14986), .A(n14976), .ZN(n14978) );
  AOI21_X1 U16571 ( .B1(n14979), .B2(n8957), .A(n14978), .ZN(n14980) );
  AND2_X1 U16572 ( .A1(n14981), .A2(n14980), .ZN(n14998) );
  INV_X1 U16573 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14982) );
  AOI22_X1 U16574 ( .A1(n10105), .A2(n14998), .B1(n14982), .B2(n14991), .ZN(
        P2_U3460) );
  AND2_X1 U16575 ( .A1(n14984), .A2(n14983), .ZN(n14989) );
  OAI21_X1 U16576 ( .B1(n14987), .B2(n14986), .A(n14985), .ZN(n14988) );
  NOR3_X1 U16577 ( .A1(n14990), .A2(n14989), .A3(n14988), .ZN(n15001) );
  INV_X1 U16578 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U16579 ( .A1(n10105), .A2(n15001), .B1(n14992), .B2(n14991), .ZN(
        P2_U3463) );
  AOI22_X1 U16580 ( .A1(n15002), .A2(n14994), .B1(n14993), .B2(n14999), .ZN(
        P2_U3505) );
  AOI22_X1 U16581 ( .A1(n15002), .A2(n14996), .B1(n14995), .B2(n14999), .ZN(
        P2_U3507) );
  AOI22_X1 U16582 ( .A1(n15002), .A2(n14998), .B1(n14997), .B2(n14999), .ZN(
        P2_U3509) );
  AOI22_X1 U16583 ( .A1(n15002), .A2(n15001), .B1(n15000), .B2(n14999), .ZN(
        P2_U3510) );
  NOR2_X1 U16584 ( .A1(P3_U3897), .A2(n15075), .ZN(P3_U3150) );
  INV_X1 U16585 ( .A(n15003), .ZN(n15004) );
  AOI21_X1 U16586 ( .B1(n9998), .B2(n15005), .A(n15004), .ZN(n15021) );
  INV_X1 U16587 ( .A(n15006), .ZN(n15007) );
  OAI21_X1 U16588 ( .B1(n15106), .B2(n14293), .A(n15007), .ZN(n15015) );
  INV_X1 U16589 ( .A(n15008), .ZN(n15009) );
  NAND3_X1 U16590 ( .A1(n15011), .A2(n15010), .A3(n15009), .ZN(n15012) );
  AOI21_X1 U16591 ( .B1(n15013), .B2(n15012), .A(n15096), .ZN(n15014) );
  AOI211_X1 U16592 ( .C1(n15102), .C2(n15016), .A(n15015), .B(n15014), .ZN(
        n15020) );
  XNOR2_X1 U16593 ( .A(n15017), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n15018) );
  NAND2_X1 U16594 ( .A1(n15086), .A2(n15018), .ZN(n15019) );
  OAI211_X1 U16595 ( .C1(n15021), .C2(n15091), .A(n15020), .B(n15019), .ZN(
        P3_U3185) );
  OAI21_X1 U16596 ( .B1(n15024), .B2(n15023), .A(n15022), .ZN(n15025) );
  INV_X1 U16597 ( .A(n15025), .ZN(n15043) );
  NOR2_X1 U16598 ( .A1(n15027), .A2(n15026), .ZN(n15028) );
  OAI21_X1 U16599 ( .B1(n15029), .B2(n15028), .A(n15055), .ZN(n15032) );
  AOI21_X1 U16600 ( .B1(n15075), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n15030), .ZN(
        n15031) );
  OAI211_X1 U16601 ( .C1(n15070), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        n15034) );
  INV_X1 U16602 ( .A(n15034), .ZN(n15042) );
  INV_X1 U16603 ( .A(n15035), .ZN(n15036) );
  AOI21_X1 U16604 ( .B1(n15038), .B2(n15037), .A(n15036), .ZN(n15039) );
  OR2_X1 U16605 ( .A1(n15040), .A2(n15039), .ZN(n15041) );
  OAI211_X1 U16606 ( .C1(n15043), .C2(n15091), .A(n15042), .B(n15041), .ZN(
        P3_U3186) );
  AOI21_X1 U16607 ( .B1(n10474), .B2(n15045), .A(n15044), .ZN(n15062) );
  INV_X1 U16608 ( .A(n15046), .ZN(n15048) );
  NAND2_X1 U16609 ( .A1(n15048), .A2(n15047), .ZN(n15049) );
  XNOR2_X1 U16610 ( .A(n15050), .B(n15049), .ZN(n15056) );
  AOI21_X1 U16611 ( .B1(n15075), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n15051), .ZN(
        n15052) );
  OAI21_X1 U16612 ( .B1(n15070), .B2(n15053), .A(n15052), .ZN(n15054) );
  AOI21_X1 U16613 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(n15061) );
  XNOR2_X1 U16614 ( .A(n15058), .B(n15057), .ZN(n15059) );
  NAND2_X1 U16615 ( .A1(n15086), .A2(n15059), .ZN(n15060) );
  OAI211_X1 U16616 ( .C1(n15062), .C2(n15091), .A(n15061), .B(n15060), .ZN(
        P3_U3187) );
  AOI21_X1 U16617 ( .B1(n15065), .B2(n15064), .A(n15063), .ZN(n15081) );
  INV_X1 U16618 ( .A(n15094), .ZN(n15069) );
  OR2_X1 U16619 ( .A1(n15066), .A2(n15094), .ZN(n15067) );
  AOI22_X1 U16620 ( .A1(n15095), .A2(n15069), .B1(n15068), .B2(n15067), .ZN(
        n15072) );
  OAI22_X1 U16621 ( .A1(n15072), .A2(n15096), .B1(n15071), .B2(n15070), .ZN(
        n15073) );
  AOI211_X1 U16622 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15075), .A(n15074), .B(
        n15073), .ZN(n15080) );
  OAI21_X1 U16623 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15077), .A(n15076), .ZN(
        n15078) );
  NAND2_X1 U16624 ( .A1(n15078), .A2(n15086), .ZN(n15079) );
  OAI211_X1 U16625 ( .C1(n15081), .C2(n15091), .A(n15080), .B(n15079), .ZN(
        P3_U3191) );
  OAI21_X1 U16626 ( .B1(n15084), .B2(n15083), .A(n15082), .ZN(n15087) );
  AOI21_X1 U16627 ( .B1(n15087), .B2(n15086), .A(n15085), .ZN(n15104) );
  AOI21_X1 U16628 ( .B1(n15090), .B2(n15089), .A(n15088), .ZN(n15092) );
  NOR2_X1 U16629 ( .A1(n15092), .A2(n15091), .ZN(n15100) );
  OR3_X1 U16630 ( .A1(n15095), .A2(n15094), .A3(n15093), .ZN(n15097) );
  AOI21_X1 U16631 ( .B1(n15098), .B2(n15097), .A(n15096), .ZN(n15099) );
  AOI211_X1 U16632 ( .C1(n15102), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        n15103) );
  OAI211_X1 U16633 ( .C1(n15106), .C2(n15105), .A(n15104), .B(n15103), .ZN(
        P3_U3192) );
  INV_X1 U16634 ( .A(n15107), .ZN(n15108) );
  AOI21_X1 U16635 ( .B1(n15110), .B2(n15109), .A(n15108), .ZN(n15118) );
  INV_X1 U16636 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15112) );
  OAI22_X1 U16637 ( .A1(n15114), .A2(n15113), .B1(n15112), .B2(n15111), .ZN(
        n15115) );
  INV_X1 U16638 ( .A(n15115), .ZN(n15116) );
  OAI221_X1 U16639 ( .B1(n15119), .B2(n15118), .C1(n15117), .C2(n9744), .A(
        n15116), .ZN(P3_U3232) );
  AOI22_X1 U16640 ( .A1(n15127), .A2(n8139), .B1(n15120), .B2(n15129), .ZN(
        P3_U3393) );
  NAND2_X1 U16641 ( .A1(n15122), .A2(n15121), .ZN(n15124) );
  NAND2_X1 U16642 ( .A1(n15124), .A2(n15123), .ZN(n15125) );
  NOR2_X1 U16643 ( .A1(n15126), .A2(n15125), .ZN(n15132) );
  INV_X1 U16644 ( .A(n15132), .ZN(n15128) );
  OAI22_X1 U16645 ( .A1(n15129), .A2(P3_REG0_REG_2__SCAN_IN), .B1(n15128), 
        .B2(n15127), .ZN(n15130) );
  INV_X1 U16646 ( .A(n15130), .ZN(P3_U3396) );
  AOI22_X1 U16647 ( .A1(n15133), .A2(n15132), .B1(n9760), .B2(n15131), .ZN(
        P3_U3461) );
  AOI21_X1 U16648 ( .B1(n15136), .B2(n15135), .A(n15134), .ZN(SUB_1596_U59) );
  OAI21_X1 U16649 ( .B1(n15139), .B2(n15138), .A(n15137), .ZN(SUB_1596_U58) );
  XOR2_X1 U16650 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15140), .Z(SUB_1596_U53) );
  AOI21_X1 U16651 ( .B1(n15143), .B2(n15142), .A(n15141), .ZN(SUB_1596_U56) );
  OAI21_X1 U16652 ( .B1(n15146), .B2(n15145), .A(n15144), .ZN(n15147) );
  XNOR2_X1 U16653 ( .A(n15147), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U16654 ( .B1(n15150), .B2(n15149), .A(n15148), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7202 ( .A(n10229), .Z(n6451) );
  CLKBUF_X1 U7216 ( .A(n8557), .Z(n6449) );
  CLKBUF_X2 U7218 ( .A(n10235), .Z(n6456) );
  CLKBUF_X1 U7226 ( .A(n14111), .Z(n6695) );
  CLKBUF_X1 U7229 ( .A(n9561), .Z(n13569) );
  CLKBUF_X1 U7297 ( .A(n10014), .Z(n6450) );
  CLKBUF_X1 U7560 ( .A(n14029), .Z(n6693) );
  CLKBUF_X2 U8410 ( .A(n13581), .Z(n6453) );
endmodule

