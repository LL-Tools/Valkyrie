

module b15_C_SARLock_k_128_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3100, n3101, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018;

  INV_X2 U3549 ( .A(n4297), .ZN(n5808) );
  CLKBUF_X2 U3550 ( .A(n3433), .Z(n4128) );
  CLKBUF_X2 U3551 ( .A(n3350), .Z(n4142) );
  INV_X2 U3552 ( .A(n3402), .ZN(n3374) );
  NAND4_X2 U3553 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n3345), .ZN(n4281)
         );
  AND2_X1 U3554 ( .A1(n3266), .A2(n3265), .ZN(n3363) );
  AND2_X1 U3555 ( .A1(n3259), .A2(n4747), .ZN(n3356) );
  CLKBUF_X1 U3556 ( .A(n4199), .Z(n3100) );
  AND2_X1 U3557 ( .A1(n4583), .A2(n4747), .ZN(n3340) );
  CLKBUF_X2 U3558 ( .A(n3434), .Z(n4198) );
  AND2_X1 U3559 ( .A1(n4583), .A2(n4746), .ZN(n3452) );
  AND2_X1 U3560 ( .A1(n4746), .A2(n4582), .ZN(n3465) );
  INV_X1 U3561 ( .A(n4317), .ZN(n4564) );
  BUF_X1 U3562 ( .A(n3379), .Z(n3531) );
  NAND2_X1 U3564 ( .A1(n5514), .A2(n5569), .ZN(n4474) );
  NAND2_X2 U3565 ( .A1(n3296), .A2(n3138), .ZN(n4893) );
  NOR2_X2 U3566 ( .A1(n4474), .A2(n3228), .ZN(n4533) );
  INV_X1 U3567 ( .A(n6071), .ZN(n6104) );
  INV_X1 U3568 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3194) );
  BUF_X1 U3569 ( .A(n3402), .Z(n3120) );
  OR2_X2 U3570 ( .A1(n5121), .A2(n3233), .ZN(n3867) );
  NAND2_X2 U3571 ( .A1(n5120), .A2(n5122), .ZN(n5121) );
  NAND2_X2 U3572 ( .A1(n3287), .A2(n3286), .ZN(n3379) );
  XNOR2_X2 U3573 ( .A(n4249), .B(n5821), .ZN(n5677) );
  BUF_X8 U3574 ( .A(n4199), .Z(n3101) );
  AND2_X2 U3575 ( .A1(n4588), .A2(n4751), .ZN(n4199) );
  BUF_X1 U3576 ( .A(n5561), .Z(n3121) );
  CLKBUF_X1 U3577 ( .A(n5677), .Z(n3107) );
  CLKBUF_X1 U3578 ( .A(n5127), .Z(n3104) );
  NAND2_X1 U3579 ( .A1(n6181), .A2(n6180), .ZN(n6179) );
  INV_X1 U3580 ( .A(n3140), .ZN(n6164) );
  NAND2_X1 U3581 ( .A1(n4674), .A2(n4673), .ZN(n3744) );
  NAND2_X1 U3582 ( .A1(n3518), .A2(n5222), .ZN(n3582) );
  INV_X1 U3583 ( .A(n3517), .ZN(n3518) );
  NAND2_X1 U3584 ( .A1(n3527), .A2(n3526), .ZN(n3517) );
  OR2_X1 U3585 ( .A1(n3527), .A2(n3526), .ZN(n3528) );
  NAND2_X1 U3586 ( .A1(n3159), .A2(n3158), .ZN(n3526) );
  OAI21_X1 U3588 ( .B1(n3547), .B2(n3545), .A(n3546), .ZN(n3159) );
  CLKBUF_X2 U3589 ( .A(n4646), .Z(n6159) );
  OAI21_X1 U3590 ( .B1(n3536), .B2(n3730), .A(n3181), .ZN(n3183) );
  NAND2_X1 U3591 ( .A1(n6117), .A2(n4893), .ZN(n5592) );
  BUF_X1 U3592 ( .A(n3730), .Z(n3130) );
  NOR2_X1 U3593 ( .A1(n4868), .A2(n3408), .ZN(n4410) );
  NAND2_X1 U3594 ( .A1(n3365), .A2(n3364), .ZN(n4868) );
  NOR2_X1 U3595 ( .A1(n3671), .A2(n3119), .ZN(n4577) );
  CLKBUF_X1 U3596 ( .A(n3380), .Z(n4268) );
  NAND2_X2 U3597 ( .A1(n3374), .A2(n3408), .ZN(n3671) );
  INV_X2 U3598 ( .A(n3386), .ZN(n3399) );
  NAND2_X1 U3599 ( .A1(n3722), .A2(n4893), .ZN(n3407) );
  CLKBUF_X2 U3600 ( .A(n3375), .Z(n3119) );
  AND3_X1 U3601 ( .A1(n3381), .A2(STATE2_REG_0__SCAN_IN), .A3(n4281), .ZN(
        n3687) );
  NAND2_X2 U3602 ( .A1(n3307), .A2(n3249), .ZN(n3381) );
  NAND2_X1 U3603 ( .A1(n3276), .A2(n3275), .ZN(n3366) );
  BUF_X2 U3606 ( .A(n3314), .Z(n4123) );
  BUF_X2 U3607 ( .A(n3351), .Z(n4200) );
  BUF_X2 U3608 ( .A(n3356), .Z(n3117) );
  CLKBUF_X2 U3610 ( .A(n3301), .Z(n4753) );
  INV_X1 U3611 ( .A(n3124), .ZN(n3125) );
  AND2_X1 U3612 ( .A1(n4583), .A2(n4747), .ZN(n3134) );
  INV_X4 U3613 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4838) );
  AND2_X1 U3614 ( .A1(n4248), .A2(n4247), .ZN(n3226) );
  OR2_X1 U3615 ( .A1(n5729), .A2(n6172), .ZN(n4407) );
  AND2_X1 U3616 ( .A1(n4185), .A2(n4184), .ZN(n5434) );
  XNOR2_X1 U3617 ( .A(n3246), .B(n4223), .ZN(n5595) );
  NAND2_X1 U3618 ( .A1(n3186), .A2(n3187), .ZN(n5546) );
  CLKBUF_X1 U3619 ( .A(n5530), .Z(n5531) );
  CLKBUF_X1 U3620 ( .A(n5452), .Z(n5453) );
  NAND2_X1 U3621 ( .A1(n3173), .A2(n3155), .ZN(n4251) );
  NAND2_X1 U3622 ( .A1(n3219), .A2(n3174), .ZN(n3173) );
  OR2_X1 U3623 ( .A1(n3867), .A2(n3868), .ZN(n3882) );
  OAI21_X1 U3624 ( .B1(n3216), .B2(n3142), .A(n3651), .ZN(n3177) );
  INV_X1 U3625 ( .A(n3217), .ZN(n3216) );
  NAND2_X1 U3626 ( .A1(n6179), .A2(n3581), .ZN(n5114) );
  OR2_X1 U3627 ( .A1(n4512), .A2(n4511), .ZN(n5731) );
  NOR3_X1 U3628 ( .A1(n5495), .A2(n3212), .A3(n3210), .ZN(n4448) );
  INV_X2 U3629 ( .A(n3140), .ZN(n5643) );
  AND2_X1 U3630 ( .A1(n3560), .A2(n3559), .ZN(n4828) );
  AND2_X1 U3631 ( .A1(n3516), .A2(n3515), .ZN(n4883) );
  CLKBUF_X1 U3632 ( .A(n5436), .Z(n6129) );
  XNOR2_X1 U3633 ( .A(n3160), .B(n3443), .ZN(n3527) );
  NAND2_X1 U3634 ( .A1(n3161), .A2(n3441), .ZN(n3160) );
  NAND2_X1 U3635 ( .A1(n6134), .A2(n4694), .ZN(n6135) );
  NAND2_X1 U3636 ( .A1(n3183), .A2(n3640), .ZN(n3546) );
  INV_X1 U3637 ( .A(n3444), .ZN(n3447) );
  NOR2_X1 U3638 ( .A1(n4805), .A2(n4806), .ZN(n4881) );
  NAND2_X1 U3639 ( .A1(n3391), .A2(n3390), .ZN(n3421) );
  AOI21_X1 U3640 ( .B1(n6091), .B2(n4564), .A(n4302), .ZN(n4738) );
  NAND2_X1 U3641 ( .A1(n3136), .A2(n3400), .ZN(n4374) );
  NAND2_X1 U3642 ( .A1(n4438), .A2(n4297), .ZN(n4597) );
  INV_X1 U3643 ( .A(n4304), .ZN(n4438) );
  AND2_X1 U3644 ( .A1(n3376), .A2(n4578), .ZN(n3414) );
  AND2_X1 U3645 ( .A1(n4577), .A2(n3368), .ZN(n4280) );
  AND2_X1 U3646 ( .A1(n3405), .A2(n4893), .ZN(n3327) );
  NAND2_X1 U3647 ( .A1(n4564), .A2(n4297), .ZN(n4430) );
  AND3_X1 U3648 ( .A1(n4504), .A2(n3379), .A3(n4893), .ZN(n3385) );
  NAND2_X1 U3649 ( .A1(n3367), .A2(n4893), .ZN(n5435) );
  INV_X1 U3650 ( .A(n3363), .ZN(n3375) );
  INV_X2 U3651 ( .A(n4281), .ZN(n3408) );
  OR2_X1 U3652 ( .A1(n3471), .A2(n3470), .ZN(n3642) );
  OR2_X1 U3653 ( .A1(n3489), .A2(n3488), .ZN(n3540) );
  CLKBUF_X1 U3654 ( .A(n3366), .Z(n3367) );
  NAND2_X1 U3655 ( .A1(n3362), .A2(n3361), .ZN(n3402) );
  AND4_X1 U3656 ( .A1(n3285), .A2(n3284), .A3(n3283), .A4(n3282), .ZN(n3286)
         );
  AND4_X1 U3657 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3287)
         );
  AND4_X1 U3658 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3307)
         );
  AND4_X1 U3659 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3348)
         );
  AND3_X1 U3660 ( .A1(n3250), .A2(n3291), .A3(n3290), .ZN(n3296) );
  AND4_X1 U3661 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3361)
         );
  AND4_X1 U3662 ( .A1(n3258), .A2(n3257), .A3(n3256), .A4(n3255), .ZN(n3266)
         );
  AND4_X1 U3663 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3276)
         );
  AND4_X1 U3664 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3275)
         );
  AND4_X1 U3666 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3362)
         );
  AND4_X1 U3667 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3345)
         );
  AND4_X1 U3668 ( .A1(n3339), .A2(n3338), .A3(n3337), .A4(n3336), .ZN(n3346)
         );
  AND4_X1 U3669 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3347)
         );
  AND4_X1 U3670 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3265)
         );
  AND2_X1 U3671 ( .A1(n3172), .A2(n3171), .ZN(n3300) );
  BUF_X2 U3672 ( .A(n4201), .Z(n4062) );
  BUF_X2 U3673 ( .A(n3315), .Z(n4029) );
  INV_X2 U3674 ( .A(n5696), .ZN(n3103) );
  BUF_X2 U3675 ( .A(n3465), .Z(n3483) );
  AND2_X2 U3676 ( .A1(n4583), .A2(n3260), .ZN(n3302) );
  AND2_X4 U3677 ( .A1(n4588), .A2(n4747), .ZN(n4129) );
  AND2_X2 U3678 ( .A1(n3194), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4751)
         );
  AND2_X2 U3679 ( .A1(n4747), .A2(n4582), .ZN(n3316) );
  AND2_X2 U3680 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4747) );
  NOR2_X2 U3681 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4746) );
  AND2_X2 U3682 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4582) );
  NOR2_X2 U3683 ( .A1(n5021), .A2(n5072), .ZN(n5120) );
  NOR2_X2 U3684 ( .A1(n4803), .A2(n4811), .ZN(n4812) );
  NAND2_X1 U3685 ( .A1(n3418), .A2(n3417), .ZN(n3477) );
  INV_X1 U3686 ( .A(n3558), .ZN(n3105) );
  INV_X1 U3687 ( .A(n3668), .ZN(n3106) );
  NAND2_X1 U3688 ( .A1(n5129), .A2(n5128), .ZN(n5127) );
  NAND2_X1 U3689 ( .A1(n3375), .A2(n3402), .ZN(n3520) );
  NAND2_X1 U3690 ( .A1(n3104), .A2(n3639), .ZN(n3108) );
  CLKBUF_X1 U3691 ( .A(n4827), .Z(n3109) );
  NAND2_X1 U3692 ( .A1(n3460), .A2(n3459), .ZN(n3110) );
  NAND2_X1 U3693 ( .A1(n3460), .A2(n3459), .ZN(n3111) );
  AND2_X1 U3694 ( .A1(n5643), .A2(n6723), .ZN(n3112) );
  NOR2_X1 U3695 ( .A1(n3112), .A2(n5660), .ZN(n5655) );
  NAND2_X1 U3696 ( .A1(n5127), .A2(n3639), .ZN(n5309) );
  NAND2_X1 U3697 ( .A1(n3460), .A2(n3459), .ZN(n3547) );
  NAND2_X2 U3698 ( .A1(n4575), .A2(n6952), .ZN(n3460) );
  XNOR2_X1 U3699 ( .A(n4774), .B(n5187), .ZN(n4742) );
  NAND2_X1 U3700 ( .A1(n3498), .A2(n3497), .ZN(n4774) );
  NAND2_X1 U3701 ( .A1(n3525), .A2(n3524), .ZN(n3561) );
  NAND2_X1 U3702 ( .A1(n3363), .A2(n3366), .ZN(n4504) );
  AND2_X2 U3703 ( .A1(n3254), .A2(n4838), .ZN(n4583) );
  BUF_X8 U3704 ( .A(n4129), .Z(n3113) );
  INV_X1 U3705 ( .A(n3125), .ZN(n3114) );
  INV_X1 U3706 ( .A(n3125), .ZN(n3115) );
  OAI21_X2 U3707 ( .B1(n5136), .B2(n3106), .A(n3542), .ZN(n4638) );
  INV_X2 U3708 ( .A(n3381), .ZN(n3382) );
  AND2_X2 U3709 ( .A1(n3254), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4588)
         );
  AND4_X1 U3710 ( .A1(n3414), .A2(n3413), .A3(n3412), .A4(n4762), .ZN(n3415)
         );
  XNOR2_X1 U3711 ( .A(n3548), .B(n3111), .ZN(n3723) );
  AND2_X4 U3712 ( .A1(n4281), .A2(n3374), .ZN(n3406) );
  NOR2_X2 U3713 ( .A1(n5515), .A2(n4009), .ZN(n5514) );
  AND2_X2 U3714 ( .A1(n3519), .A2(n3582), .ZN(n4914) );
  OAI21_X1 U3715 ( .B1(n5385), .B2(n3225), .A(n5386), .ZN(n5922) );
  AND2_X1 U3716 ( .A1(n4838), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3259)
         );
  XNOR2_X1 U3717 ( .A(n3561), .B(n6273), .ZN(n3215) );
  NOR2_X2 U3718 ( .A1(n3404), .A2(n3386), .ZN(n3718) );
  NAND2_X2 U3719 ( .A1(n3528), .A2(n3517), .ZN(n4782) );
  OAI21_X2 U3720 ( .B1(n3179), .B2(n3142), .A(n3176), .ZN(n5385) );
  AND2_X2 U3721 ( .A1(n4533), .A2(n3192), .ZN(n4234) );
  AND2_X1 U3722 ( .A1(n4583), .A2(n3260), .ZN(n3122) );
  AND2_X2 U3723 ( .A1(n4583), .A2(n3260), .ZN(n3123) );
  AND2_X1 U3724 ( .A1(n4583), .A2(n4746), .ZN(n3124) );
  INV_X1 U3725 ( .A(n3723), .ZN(n3127) );
  INV_X1 U3726 ( .A(n3127), .ZN(n3128) );
  INV_X1 U3727 ( .A(n3127), .ZN(n3129) );
  XNOR2_X1 U3728 ( .A(n3478), .B(n3477), .ZN(n3730) );
  AND2_X1 U3729 ( .A1(n4747), .A2(n4582), .ZN(n3131) );
  AND2_X2 U3730 ( .A1(n4747), .A2(n4582), .ZN(n3132) );
  AND2_X1 U3731 ( .A1(n4583), .A2(n4747), .ZN(n3133) );
  AND2_X2 U3732 ( .A1(n3195), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3260)
         );
  NOR2_X1 U3733 ( .A1(n4267), .A2(n6952), .ZN(n4214) );
  NOR2_X1 U3734 ( .A1(n3492), .A2(n6952), .ZN(n3495) );
  NAND2_X1 U3735 ( .A1(n3642), .A2(n3382), .ZN(n3492) );
  NAND2_X1 U3736 ( .A1(n3236), .A2(n3234), .ZN(n3233) );
  NOR2_X1 U3737 ( .A1(n3237), .A2(n3235), .ZN(n3234) );
  INV_X1 U3738 ( .A(n5623), .ZN(n3227) );
  NAND2_X1 U3739 ( .A1(n5519), .A2(n3204), .ZN(n3203) );
  INV_X1 U3740 ( .A(n5533), .ZN(n3204) );
  INV_X1 U3741 ( .A(n3618), .ZN(n3616) );
  INV_X1 U3742 ( .A(n3619), .ZN(n3617) );
  NOR2_X1 U3743 ( .A1(n3657), .A2(n3175), .ZN(n3174) );
  INV_X1 U3744 ( .A(n3655), .ZN(n3175) );
  INV_X1 U3745 ( .A(n5358), .ZN(n3178) );
  OAI21_X1 U3746 ( .B1(n3647), .B2(n3218), .A(n5316), .ZN(n3217) );
  INV_X1 U3747 ( .A(n3495), .ZN(n3640) );
  OR2_X1 U3748 ( .A1(n3407), .A2(n3719), .ZN(n4267) );
  AOI22_X1 U3749 ( .A1(n3314), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3264) );
  AND2_X1 U3750 ( .A1(n3389), .A2(n3349), .ZN(n4273) );
  AND2_X1 U3751 ( .A1(n6084), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5262) );
  NOR2_X1 U3752 ( .A1(n4576), .A2(n4378), .ZN(n4745) );
  OR2_X1 U3753 ( .A1(n4611), .A2(n4549), .ZN(n4594) );
  INV_X2 U3754 ( .A(n4076), .ZN(n4221) );
  OR2_X1 U3755 ( .A1(n3230), .A2(n3229), .ZN(n3228) );
  NAND2_X1 U3756 ( .A1(n4225), .A2(n4224), .ZN(n5615) );
  NAND2_X1 U3757 ( .A1(n5635), .A2(n5634), .ZN(n5633) );
  NAND2_X1 U3758 ( .A1(n3716), .A2(n3715), .ZN(n4589) );
  NAND2_X1 U3759 ( .A1(n4257), .A2(n3714), .ZN(n3715) );
  AOI22_X1 U3760 ( .A1(n3302), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3291) );
  INV_X1 U3761 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6952) );
  INV_X1 U3762 ( .A(n6582), .ZN(n4865) );
  AND2_X1 U3763 ( .A1(n6084), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6094) );
  NOR2_X1 U3764 ( .A1(n4454), .A2(n6981), .ZN(n4416) );
  AND2_X1 U3765 ( .A1(n4454), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4455) );
  AND2_X1 U3766 ( .A1(n3699), .A2(n3698), .ZN(n3701) );
  INV_X1 U3767 ( .A(n5366), .ZN(n3235) );
  AND2_X1 U3768 ( .A1(n5222), .A2(n3231), .ZN(n3180) );
  AND2_X1 U3769 ( .A1(n3605), .A2(n3583), .ZN(n3231) );
  NAND2_X1 U3770 ( .A1(n3375), .A2(n3722), .ZN(n3380) );
  OAI22_X1 U3771 ( .A1(n4187), .A2(n5182), .B1(n3717), .B2(n6358), .ZN(n3392)
         );
  NOR2_X1 U3772 ( .A1(n3245), .A2(n4183), .ZN(n3244) );
  INV_X1 U3773 ( .A(n4236), .ZN(n3245) );
  NOR2_X1 U3774 ( .A1(n5481), .A2(n3193), .ZN(n3192) );
  INV_X1 U3775 ( .A(n5493), .ZN(n3193) );
  INV_X1 U3776 ( .A(n4214), .ZN(n4180) );
  NOR2_X1 U3777 ( .A1(n3188), .A2(n5585), .ZN(n3187) );
  INV_X1 U3778 ( .A(n5547), .ZN(n3188) );
  NAND2_X1 U3779 ( .A1(n3832), .A2(n3239), .ZN(n3238) );
  INV_X1 U3780 ( .A(n5301), .ZN(n3832) );
  AND2_X1 U3781 ( .A1(n3724), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3752) );
  INV_X1 U3782 ( .A(n3200), .ZN(n3199) );
  NAND2_X1 U3783 ( .A1(n4914), .A2(n3668), .ZN(n3525) );
  NAND2_X1 U3784 ( .A1(n3399), .A2(n4281), .ZN(n3400) );
  NAND2_X1 U3785 ( .A1(n3408), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3503) );
  NOR2_X1 U3786 ( .A1(n3129), .A2(n6703), .ZN(n6360) );
  AOI22_X1 U3787 ( .A1(n4201), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3311) );
  OR2_X1 U3788 ( .A1(n6673), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4187) );
  INV_X1 U3789 ( .A(n4355), .ZN(n3205) );
  AND2_X1 U3790 ( .A1(n4456), .A2(n4158), .ZN(n4218) );
  NAND2_X1 U3791 ( .A1(n4094), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4096)
         );
  AND2_X1 U3792 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n4025), .ZN(n4026)
         );
  INV_X1 U3793 ( .A(n5517), .ZN(n4009) );
  NOR2_X1 U3794 ( .A1(n3989), .A2(n5680), .ZN(n3990) );
  NAND2_X1 U3795 ( .A1(n3990), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4024)
         );
  INV_X1 U3796 ( .A(n5367), .ZN(n3191) );
  NAND2_X1 U3797 ( .A1(n3847), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3862)
         );
  INV_X1 U3798 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5405) );
  OR2_X1 U3799 ( .A1(n3799), .A2(n5291), .ZN(n3800) );
  NOR2_X1 U3800 ( .A1(n6782), .A2(n3800), .ZN(n3818) );
  OR2_X1 U3801 ( .A1(n4589), .A2(n6582), .ZN(n4611) );
  AND2_X1 U3802 ( .A1(n3227), .A2(n3157), .ZN(n3164) );
  OR2_X1 U3803 ( .A1(n5496), .A2(n3211), .ZN(n3210) );
  OR2_X1 U3804 ( .A1(n4484), .A2(n4444), .ZN(n3211) );
  NOR2_X1 U3805 ( .A1(n5495), .A2(n5496), .ZN(n5494) );
  AND2_X1 U3806 ( .A1(n4290), .A2(n4289), .ZN(n5533) );
  NOR2_X1 U3807 ( .A1(n3640), .A2(n3106), .ZN(n3641) );
  INV_X1 U3808 ( .A(n3252), .ZN(n3225) );
  NAND2_X1 U3809 ( .A1(n3108), .A2(n5308), .ZN(n5307) );
  NAND2_X1 U3810 ( .A1(n4278), .A2(n4865), .ZN(n4385) );
  AOI21_X1 U3811 ( .B1(n3491), .B2(STATE2_REG_0__SCAN_IN), .A(n3182), .ZN(
        n3181) );
  INV_X1 U3812 ( .A(n3537), .ZN(n3182) );
  AND2_X1 U3813 ( .A1(n3129), .A2(n5136), .ZN(n6430) );
  OR2_X1 U3814 ( .A1(n3129), .A2(n5181), .ZN(n6368) );
  OR2_X1 U3815 ( .A1(n3129), .A2(n5136), .ZN(n6403) );
  AND2_X1 U3816 ( .A1(n4761), .A2(n4575), .ZN(n6439) );
  INV_X1 U3817 ( .A(n5184), .ZN(n5079) );
  OR2_X1 U3818 ( .A1(n4279), .A2(n3721), .ZN(n4859) );
  AND3_X1 U3819 ( .A1(n3399), .A2(n3363), .A3(n3379), .ZN(n3364) );
  INV_X1 U3820 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6695) );
  AND2_X1 U3821 ( .A1(n6090), .A2(EBX_REG_30__SCAN_IN), .ZN(n3207) );
  AND2_X1 U3822 ( .A1(n5262), .A2(n4419), .ZN(n6090) );
  OR2_X1 U3823 ( .A1(n6685), .A2(n4415), .ZN(n6084) );
  NAND2_X1 U3824 ( .A1(n4509), .A2(n4508), .ZN(n6117) );
  OR2_X1 U3825 ( .A1(n4689), .A2(n4676), .ZN(n4508) );
  INV_X1 U3826 ( .A(n6134), .ZN(n6128) );
  INV_X1 U3827 ( .A(n6195), .ZN(n6168) );
  OR2_X1 U3828 ( .A1(n4611), .A2(n4859), .ZN(n6172) );
  AND2_X1 U3829 ( .A1(n4242), .A2(n4243), .ZN(n5748) );
  INV_X1 U3830 ( .A(n3238), .ZN(n3236) );
  NAND2_X1 U3831 ( .A1(n3574), .A2(n3573), .ZN(n3583) );
  OR2_X1 U3832 ( .A1(n3593), .A2(n3592), .ZN(n3621) );
  NAND2_X1 U3833 ( .A1(n3687), .A2(n3668), .ZN(n3705) );
  AND2_X1 U3834 ( .A1(n3401), .A2(n3378), .ZN(n3387) );
  AOI22_X1 U3835 ( .A1(n4129), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U3836 ( .A1(n3100), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U3837 ( .A1(n3315), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U3838 ( .A1(n3122), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U3839 ( .A1(n3315), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3267) );
  AND2_X1 U3840 ( .A1(n3113), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U3841 ( .A1(n3433), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3280) );
  INV_X1 U3842 ( .A(n5484), .ZN(n3213) );
  OR2_X1 U3843 ( .A1(n5504), .A2(n4475), .ZN(n3230) );
  OR2_X1 U3844 ( .A1(n5532), .A2(n3185), .ZN(n3184) );
  INV_X1 U3845 ( .A(n3187), .ZN(n3185) );
  NAND2_X1 U3846 ( .A1(n3242), .A2(n3241), .ZN(n3240) );
  INV_X1 U3847 ( .A(n5580), .ZN(n3242) );
  INV_X1 U3848 ( .A(n5918), .ZN(n3241) );
  INV_X1 U3849 ( .A(n5345), .ZN(n3237) );
  INV_X1 U3850 ( .A(n3603), .ZN(n3224) );
  OR2_X1 U3851 ( .A1(n3213), .A2(n5469), .ZN(n3212) );
  NOR2_X1 U3852 ( .A1(n5073), .A2(n3201), .ZN(n3200) );
  INV_X1 U3853 ( .A(n5124), .ZN(n3201) );
  NAND2_X1 U3854 ( .A1(n4299), .A2(n3214), .ZN(n4301) );
  NAND2_X1 U3855 ( .A1(n3383), .A2(n3382), .ZN(n3384) );
  OR2_X1 U3856 ( .A1(n3458), .A2(n3457), .ZN(n3549) );
  NOR2_X1 U3857 ( .A1(n3381), .A2(n6952), .ZN(n4503) );
  OR2_X1 U3858 ( .A1(n3514), .A2(n3513), .ZN(n3575) );
  NAND2_X1 U3859 ( .A1(n3504), .A2(n3503), .ZN(n3714) );
  INV_X1 U3860 ( .A(n4503), .ZN(n3504) );
  INV_X1 U3861 ( .A(n3705), .ZN(n3711) );
  AOI221_X1 U3862 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3710), .C1(
        n5964), .C2(n3710), .A(n3709), .ZN(n4257) );
  AND2_X1 U3863 ( .A1(n3323), .A2(n4504), .ZN(n3324) );
  INV_X1 U3864 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6279) );
  AOI22_X1 U3865 ( .A1(n3315), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3352) );
  NAND2_X1 U3866 ( .A1(n4201), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3172) );
  NAND2_X1 U3867 ( .A1(n3433), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U3868 ( .A1(n3433), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3290) );
  INV_X1 U3869 ( .A(n4888), .ZN(n4940) );
  INV_X1 U3870 ( .A(n4410), .ZN(n4549) );
  OR2_X1 U3871 ( .A1(n3392), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3372)
         );
  AND2_X1 U3872 ( .A1(n5262), .A2(n4422), .ZN(n6063) );
  AOI22_X1 U3873 ( .A1(n4160), .A2(n4159), .B1(n4158), .B2(n5472), .ZN(n4236)
         );
  XNOR2_X1 U3874 ( .A(n4228), .B(n4227), .ZN(n4454) );
  AND2_X1 U3875 ( .A1(n4398), .A2(n3244), .ZN(n3243) );
  OR2_X1 U3876 ( .A1(n4164), .A2(n4163), .ZN(n4226) );
  OR2_X1 U3877 ( .A1(n4121), .A2(n5486), .ZN(n4161) );
  AND2_X1 U3878 ( .A1(n4118), .A2(n4117), .ZN(n5493) );
  NAND2_X1 U3879 ( .A1(n4071), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4093)
         );
  AND2_X1 U3880 ( .A1(n4028), .A2(n4027), .ZN(n5569) );
  AND2_X1 U3881 ( .A1(n4008), .A2(n4007), .ZN(n5517) );
  AND2_X1 U3882 ( .A1(n3992), .A2(n3991), .ZN(n5671) );
  NOR2_X1 U3883 ( .A1(n3956), .A2(n5998), .ZN(n3957) );
  NAND2_X1 U3884 ( .A1(n3926), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3956)
         );
  AND2_X1 U3885 ( .A1(n3913), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3926)
         );
  INV_X1 U3886 ( .A(n5452), .ZN(n3186) );
  NOR2_X1 U3887 ( .A1(n6020), .A2(n3897), .ZN(n3913) );
  NOR2_X1 U3888 ( .A1(n3862), .A2(n5405), .ZN(n3863) );
  NAND2_X1 U3889 ( .A1(n3863), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3897)
         );
  NAND2_X1 U3890 ( .A1(n3190), .A2(n3189), .ZN(n5428) );
  INV_X1 U3891 ( .A(n5430), .ZN(n3189) );
  NAND2_X1 U3892 ( .A1(n3861), .A2(n3860), .ZN(n5366) );
  NOR2_X1 U3893 ( .A1(n3833), .A2(n5360), .ZN(n3847) );
  NAND2_X1 U3894 ( .A1(n3818), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3833)
         );
  AND2_X1 U3895 ( .A1(n3831), .A2(n3830), .ZN(n5301) );
  OR2_X1 U3896 ( .A1(n3803), .A2(n3802), .ZN(n5122) );
  NOR2_X1 U3897 ( .A1(n3776), .A2(n5276), .ZN(n3777) );
  AOI21_X1 U3898 ( .B1(n3782), .B2(n3894), .A(n3781), .ZN(n5024) );
  CLKBUF_X1 U3899 ( .A(n5021), .Z(n5022) );
  CLKBUF_X1 U3900 ( .A(n4816), .Z(n4817) );
  AND3_X1 U3901 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .A3(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n3767) );
  INV_X1 U3902 ( .A(n3759), .ZN(n3760) );
  NAND2_X1 U3903 ( .A1(n4914), .A2(n3894), .ZN(n3761) );
  AND2_X1 U3904 ( .A1(n3164), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3163)
         );
  INV_X1 U3905 ( .A(n5615), .ZN(n3169) );
  NOR2_X1 U3906 ( .A1(n5743), .A2(n3168), .ZN(n3167) );
  NAND2_X1 U3907 ( .A1(n5707), .A2(n6776), .ZN(n3168) );
  INV_X1 U3908 ( .A(n5616), .ZN(n4238) );
  NAND2_X1 U3909 ( .A1(n3139), .A2(n3227), .ZN(n5616) );
  AND2_X1 U3910 ( .A1(n4436), .A2(n4435), .ZN(n5496) );
  OAI22_X1 U3911 ( .A1(n4249), .A2(n3162), .B1(n3156), .B2(n3140), .ZN(n5635)
         );
  NOR2_X1 U3912 ( .A1(n6164), .A2(n3663), .ZN(n3162) );
  AND2_X1 U3913 ( .A1(n4427), .A2(n4426), .ZN(n5506) );
  NOR2_X2 U3914 ( .A1(n5927), .A2(n3202), .ZN(n5573) );
  OR3_X1 U3915 ( .A1(n3205), .A2(n3203), .A3(n5571), .ZN(n3202) );
  OAI22_X1 U3916 ( .A1(n5670), .A2(n5669), .B1(n5643), .B2(n6935), .ZN(n5661)
         );
  AOI22_X1 U3917 ( .A1(n5677), .A2(n3140), .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n4249), .ZN(n5670) );
  NOR2_X1 U3918 ( .A1(n5927), .A2(n5533), .ZN(n5809) );
  NOR2_X1 U3919 ( .A1(n3144), .A2(n3221), .ZN(n3220) );
  INV_X1 U3920 ( .A(n3653), .ZN(n3221) );
  OR2_X1 U3921 ( .A1(n4385), .A2(n4377), .ZN(n5416) );
  INV_X1 U3922 ( .A(n3177), .ZN(n3176) );
  NOR2_X1 U3923 ( .A1(n3148), .A2(n3198), .ZN(n3197) );
  INV_X1 U3924 ( .A(n5303), .ZN(n3198) );
  NOR2_X1 U3925 ( .A1(n4525), .A2(n3148), .ZN(n6050) );
  NAND2_X1 U3926 ( .A1(n3196), .A2(n3200), .ZN(n6051) );
  NOR2_X1 U3927 ( .A1(n4525), .A2(n5073), .ZN(n5123) );
  NAND2_X1 U3928 ( .A1(n4827), .A2(n3562), .ZN(n6181) );
  NAND2_X1 U3929 ( .A1(n3215), .A2(n4828), .ZN(n4827) );
  AOI21_X1 U3930 ( .B1(n4680), .B2(n4679), .A(n3556), .ZN(n4792) );
  NAND2_X1 U3931 ( .A1(n3110), .A2(n3545), .ZN(n3158) );
  NAND2_X1 U3932 ( .A1(n6952), .A2(n4889), .ZN(n5184) );
  OR2_X1 U3933 ( .A1(n4573), .A2(n4572), .ZN(n4842) );
  OR2_X1 U3934 ( .A1(n4782), .A2(n5222), .ZN(n6432) );
  AND2_X1 U3935 ( .A1(n4914), .A2(n4782), .ZN(n6516) );
  AND2_X1 U3936 ( .A1(n4761), .A2(n5852), .ZN(n6362) );
  INV_X1 U3937 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6398) );
  OR2_X1 U3938 ( .A1(n4782), .A2(n4883), .ZN(n4888) );
  NOR2_X1 U3939 ( .A1(n3313), .A2(n3312), .ZN(n3321) );
  AND2_X1 U3940 ( .A1(n4890), .A2(n4889), .ZN(n4908) );
  NAND2_X1 U3941 ( .A1(n3130), .A2(n6952), .ZN(n3535) );
  AND2_X1 U3942 ( .A1(n6981), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3717) );
  INV_X1 U3943 ( .A(n6090), .ZN(n6080) );
  INV_X1 U3944 ( .A(n6063), .ZN(n6083) );
  INV_X1 U3945 ( .A(n6027), .ZN(n6053) );
  AND2_X1 U3946 ( .A1(n5260), .A2(n5873), .ZN(n6064) );
  NOR3_X1 U3947 ( .A1(n5927), .A2(n3205), .A3(n5533), .ZN(n5520) );
  INV_X1 U3948 ( .A(n6117), .ZN(n5588) );
  INV_X1 U3949 ( .A(n6135), .ZN(n6126) );
  INV_X1 U3950 ( .A(n6133), .ZN(n5613) );
  NAND2_X1 U3951 ( .A1(n4693), .A2(n4692), .ZN(n6134) );
  OR3_X1 U3952 ( .A1(n4611), .A2(n4610), .A3(n6689), .ZN(n4636) );
  INV_X1 U3953 ( .A(n4692), .ZN(n6146) );
  INV_X1 U3954 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5680) );
  INV_X1 U3955 ( .A(n6046), .ZN(n6169) );
  INV_X1 U3956 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5360) );
  INV_X1 U3957 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5276) );
  AND2_X1 U3958 ( .A1(n6172), .A2(n4188), .ZN(n6188) );
  INV_X1 U3959 ( .A(n6188), .ZN(n5686) );
  XNOR2_X1 U3960 ( .A(n3165), .B(n6991), .ZN(n5704) );
  NAND2_X1 U3961 ( .A1(n3170), .A2(n3166), .ZN(n3165) );
  NAND2_X1 U3962 ( .A1(n3169), .A2(n3167), .ZN(n3166) );
  NAND2_X1 U3963 ( .A1(n3139), .A2(n3163), .ZN(n3170) );
  XNOR2_X1 U3964 ( .A(n4406), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5729)
         );
  NAND2_X1 U3965 ( .A1(n4405), .A2(n3141), .ZN(n4406) );
  NAND2_X1 U3966 ( .A1(n5645), .A2(n5778), .ZN(n5646) );
  AND2_X1 U3967 ( .A1(n5790), .A2(n5798), .ZN(n5787) );
  NOR2_X1 U3968 ( .A1(n5394), .A2(n5420), .ZN(n5937) );
  NAND2_X1 U3969 ( .A1(n3654), .A2(n3653), .ZN(n5412) );
  NAND2_X1 U3970 ( .A1(n5357), .A2(n5358), .ZN(n6163) );
  NAND2_X1 U3971 ( .A1(n5307), .A2(n3647), .ZN(n5318) );
  NAND2_X1 U3972 ( .A1(n5112), .A2(n3603), .ZN(n4524) );
  OR2_X1 U3973 ( .A1(n4385), .A2(n4286), .ZN(n6255) );
  INV_X1 U3974 ( .A(n6223), .ZN(n6269) );
  XNOR2_X1 U3975 ( .A(n3546), .B(n3545), .ZN(n3548) );
  NOR2_X2 U3976 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6409) );
  AND2_X1 U3977 ( .A1(n3129), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6515) );
  CLKBUF_X1 U3978 ( .A(n4760), .Z(n4761) );
  INV_X1 U3979 ( .A(n6409), .ZN(n6527) );
  OR2_X1 U3980 ( .A1(n4589), .A2(n6665), .ZN(n5862) );
  NAND2_X1 U3981 ( .A1(n6981), .A2(n6665), .ZN(n6673) );
  OAI21_X1 U3982 ( .B1(n6284), .B2(n6299), .A(n6283), .ZN(n6302) );
  OAI21_X1 U3983 ( .B1(n6493), .B2(n6492), .A(n6491), .ZN(n6511) );
  INV_X1 U3984 ( .A(n5258), .ZN(n4937) );
  INV_X1 U3985 ( .A(n5144), .ZN(n5173) );
  INV_X1 U3986 ( .A(n6534), .ZN(n6437) );
  INV_X1 U3987 ( .A(n6309), .ZN(n6522) );
  INV_X1 U3988 ( .A(n6540), .ZN(n6450) );
  INV_X1 U3989 ( .A(n6322), .ZN(n6535) );
  INV_X1 U3990 ( .A(n6546), .ZN(n6454) );
  INV_X1 U3991 ( .A(n6552), .ZN(n6458) );
  INV_X1 U3992 ( .A(n6330), .ZN(n6547) );
  INV_X1 U3993 ( .A(n6558), .ZN(n6462) );
  INV_X1 U3994 ( .A(n6334), .ZN(n6553) );
  INV_X1 U3995 ( .A(n6564), .ZN(n6466) );
  INV_X1 U3996 ( .A(n6338), .ZN(n6559) );
  INV_X1 U3997 ( .A(n6570), .ZN(n6470) );
  INV_X1 U3998 ( .A(n6342), .ZN(n6565) );
  INV_X1 U3999 ( .A(n6580), .ZN(n6476) );
  NOR2_X2 U4000 ( .A1(n4888), .A2(n6368), .ZN(n5217) );
  OAI211_X1 U4001 ( .C1(n5082), .C2(n6665), .A(n5081), .B(n5080), .ZN(n5104)
         );
  INV_X1 U4002 ( .A(n5076), .ZN(n5108) );
  INV_X1 U4003 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6981) );
  NAND2_X1 U4004 ( .A1(n3717), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6582) );
  INV_X1 U4005 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6703) );
  INV_X1 U4006 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6665) );
  OR2_X1 U4007 ( .A1(n4870), .A2(n4869), .ZN(n6664) );
  AOI21_X1 U4008 ( .B1(n3208), .B2(n6092), .A(n3206), .ZN(n4471) );
  AOI21_X1 U4009 ( .B1(n4514), .B2(n6113), .A(n4513), .ZN(n4515) );
  NOR2_X1 U4010 ( .A1(n6117), .A2(n6916), .ZN(n4513) );
  OAI21_X1 U4011 ( .B1(n5748), .B2(n6172), .A(n3226), .ZN(U2958) );
  INV_X1 U4012 ( .A(n4480), .ZN(n4481) );
  OAI21_X1 U4013 ( .B1(n5874), .B2(n5696), .A(n4479), .ZN(n4480) );
  AND2_X2 U4014 ( .A1(n3631), .A2(n3641), .ZN(n3140) );
  AND2_X2 U4015 ( .A1(n3260), .A2(n4582), .ZN(n3301) );
  AND2_X2 U4016 ( .A1(n4588), .A2(n3260), .ZN(n3315) );
  NAND2_X1 U4017 ( .A1(n3173), .A2(n3656), .ZN(n5683) );
  NAND2_X1 U4018 ( .A1(n4533), .A2(n5493), .ZN(n5480) );
  NOR2_X1 U4019 ( .A1(n5121), .A2(n3238), .ZN(n5300) );
  OR2_X1 U4020 ( .A1(n4474), .A2(n4475), .ZN(n4473) );
  AND2_X1 U4021 ( .A1(n3398), .A2(n3397), .ZN(n3136) );
  NAND2_X1 U4022 ( .A1(n5366), .A2(n3882), .ZN(n3137) );
  NAND2_X1 U4023 ( .A1(n3722), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3911) );
  INV_X1 U4024 ( .A(n3911), .ZN(n3894) );
  INV_X1 U4025 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3195) );
  AND4_X1 U4026 ( .A1(n3295), .A2(n3294), .A3(n3293), .A4(n3292), .ZN(n3138)
         );
  AND2_X1 U4027 ( .A1(n5633), .A2(n3664), .ZN(n3139) );
  AND2_X1 U4028 ( .A1(n4588), .A2(n4746), .ZN(n3350) );
  NOR2_X1 U4029 ( .A1(n4474), .A2(n3230), .ZN(n4531) );
  NOR2_X1 U4030 ( .A1(n5452), .A2(n5585), .ZN(n5545) );
  NAND2_X1 U4031 ( .A1(n5530), .A2(n5671), .ZN(n5515) );
  NAND2_X1 U4032 ( .A1(n3139), .A2(n3164), .ZN(n3141) );
  OR2_X1 U4033 ( .A1(n3652), .A2(n3178), .ZN(n3142) );
  OR2_X1 U4034 ( .A1(n5546), .A2(n3240), .ZN(n5529) );
  OR3_X1 U4035 ( .A1(n5495), .A2(n5496), .A3(n3213), .ZN(n3143) );
  NAND2_X1 U4036 ( .A1(n3380), .A2(n3379), .ZN(n3405) );
  INV_X1 U4037 ( .A(n3209), .ZN(n5471) );
  NOR3_X1 U4038 ( .A1(n5495), .A2(n3212), .A3(n5496), .ZN(n3209) );
  OR2_X1 U4039 ( .A1(n5546), .A2(n5918), .ZN(n5579) );
  INV_X1 U4040 ( .A(n3208), .ZN(n5722) );
  OR2_X1 U4041 ( .A1(n4450), .A2(n4449), .ZN(n3208) );
  INV_X1 U4042 ( .A(n5315), .ZN(n3218) );
  NOR2_X1 U4043 ( .A1(n3520), .A2(n3381), .ZN(n3396) );
  AND2_X1 U4044 ( .A1(n5643), .A2(n5421), .ZN(n3144) );
  NAND2_X1 U4045 ( .A1(n3627), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3145)
         );
  AND2_X1 U4046 ( .A1(n5308), .A2(n5315), .ZN(n3146) );
  NOR2_X1 U4047 ( .A1(n5929), .A2(n5928), .ZN(n4348) );
  OR2_X1 U4048 ( .A1(n5121), .A2(n5268), .ZN(n3147) );
  OR2_X1 U4049 ( .A1(n3199), .A2(n6052), .ZN(n3148) );
  INV_X1 U4050 ( .A(n3366), .ZN(n3722) );
  NAND2_X1 U4051 ( .A1(n3179), .A2(n3216), .ZN(n5357) );
  NAND2_X1 U4052 ( .A1(n5573), .A2(n4365), .ZN(n4431) );
  OR3_X1 U4053 ( .A1(n5927), .A2(n3205), .A3(n3203), .ZN(n3149) );
  INV_X1 U4054 ( .A(n3190), .ZN(n5429) );
  OR2_X1 U4055 ( .A1(n3238), .A2(n3237), .ZN(n3150) );
  OR2_X1 U4056 ( .A1(n3184), .A2(n3240), .ZN(n3151) );
  NAND2_X1 U4057 ( .A1(n5643), .A2(n3658), .ZN(n3152) );
  NAND2_X1 U4058 ( .A1(n3219), .A2(n3655), .ZN(n5692) );
  AND2_X1 U4059 ( .A1(n4236), .A2(n3192), .ZN(n3153) );
  NOR2_X1 U4060 ( .A1(n4458), .A2(n3207), .ZN(n3154) );
  AND2_X1 U4061 ( .A1(n3152), .A2(n3656), .ZN(n3155) );
  INV_X1 U4062 ( .A(n5871), .ZN(n6092) );
  INV_X1 U4063 ( .A(n3739), .ZN(n4216) );
  NOR2_X1 U4064 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3739) );
  NOR2_X1 U4065 ( .A1(n6041), .A2(n6042), .ZN(n5368) );
  INV_X1 U4066 ( .A(n4532), .ZN(n3229) );
  AOI21_X1 U4067 ( .B1(n3788), .B2(n3894), .A(n3787), .ZN(n5072) );
  NOR2_X1 U4068 ( .A1(n5586), .A2(n5587), .ZN(n5548) );
  INV_X1 U4069 ( .A(n6172), .ZN(n6191) );
  AND3_X1 U4070 ( .A1(n3817), .A2(n3816), .A3(n3815), .ZN(n5268) );
  INV_X1 U4071 ( .A(n5268), .ZN(n3239) );
  AND3_X1 U4072 ( .A1(n5813), .A2(n5705), .A3(n4384), .ZN(n3156) );
  AND2_X1 U4073 ( .A1(n5706), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3157)
         );
  NAND2_X1 U4074 ( .A1(n4760), .A2(n6952), .ZN(n3161) );
  AND2_X2 U4075 ( .A1(n4583), .A2(n4751), .ZN(n3433) );
  AND2_X2 U4076 ( .A1(n3260), .A2(n3259), .ZN(n4201) );
  NAND2_X1 U4077 ( .A1(n3146), .A2(n5309), .ZN(n3179) );
  NAND2_X1 U4078 ( .A1(n3518), .A2(n3180), .ZN(n3619) );
  INV_X1 U4079 ( .A(n3582), .ZN(n3232) );
  NAND3_X1 U4080 ( .A1(n3631), .A2(n3668), .A3(n3782), .ZN(n3625) );
  NOR2_X2 U4081 ( .A1(n5452), .A2(n3151), .ZN(n5530) );
  OAI21_X2 U4082 ( .B1(n3137), .B2(n3191), .A(n3870), .ZN(n3190) );
  NOR2_X2 U4083 ( .A1(n5121), .A2(n3150), .ZN(n5367) );
  NAND2_X1 U4084 ( .A1(n4533), .A2(n3153), .ZN(n4235) );
  INV_X1 U4085 ( .A(n4525), .ZN(n3196) );
  NAND2_X1 U4086 ( .A1(n3196), .A2(n3197), .ZN(n6041) );
  NAND3_X1 U4087 ( .A1(n4457), .A2(n4470), .A3(n3154), .ZN(n3206) );
  XNOR2_X1 U4088 ( .A(n4300), .B(n4301), .ZN(n6091) );
  NAND3_X1 U4089 ( .A1(n5808), .A2(n6877), .A3(n4564), .ZN(n3214) );
  AND2_X2 U4090 ( .A1(n5808), .A2(n4564), .ZN(n4441) );
  OAI21_X1 U4091 ( .B1(n4828), .B2(n3215), .A(n3109), .ZN(n6267) );
  NAND3_X1 U4092 ( .A1(n3389), .A2(n3349), .A3(n3374), .ZN(n4282) );
  NAND2_X1 U4093 ( .A1(n3654), .A2(n3220), .ZN(n3219) );
  NAND3_X1 U4094 ( .A1(n3223), .A2(n3145), .A3(n3222), .ZN(n5129) );
  NAND3_X1 U4095 ( .A1(n5114), .A2(n5113), .A3(n4523), .ZN(n3222) );
  NAND2_X1 U4096 ( .A1(n5114), .A2(n5113), .ZN(n5112) );
  NAND2_X1 U4097 ( .A1(n4523), .A2(n3224), .ZN(n3223) );
  NAND2_X1 U4098 ( .A1(n4524), .A2(n4523), .ZN(n4522) );
  NAND2_X1 U4099 ( .A1(n3232), .A2(n3583), .ZN(n3604) );
  AND2_X1 U4100 ( .A1(n4234), .A2(n3244), .ZN(n4399) );
  NAND2_X1 U4101 ( .A1(n4234), .A2(n3243), .ZN(n3246) );
  NAND2_X1 U4102 ( .A1(n4237), .A2(n3103), .ZN(n4248) );
  NAND2_X1 U4103 ( .A1(n5434), .A2(n3103), .ZN(n4195) );
  NOR3_X2 U4104 ( .A1(n3139), .A2(n5743), .A3(n5624), .ZN(n4404) );
  XNOR2_X1 U4105 ( .A(n3631), .B(n3630), .ZN(n3788) );
  NAND2_X1 U4106 ( .A1(n3617), .A2(n3616), .ZN(n3631) );
  OR2_X1 U4107 ( .A1(n5787), .A2(n5778), .ZN(n3247) );
  AND2_X1 U4108 ( .A1(n4232), .A2(n4231), .ZN(n3248) );
  NAND2_X1 U4109 ( .A1(n3321), .A2(n3251), .ZN(n3386) );
  AND4_X1 U4110 ( .A1(n3306), .A2(n3305), .A3(n3304), .A4(n3303), .ZN(n3249)
         );
  INV_X1 U4111 ( .A(n3731), .ZN(n4076) );
  NOR2_X1 U4112 ( .A1(n4893), .A2(n6695), .ZN(n3731) );
  INV_X1 U4113 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5964) );
  AND2_X1 U4114 ( .A1(n3289), .A2(n3288), .ZN(n3250) );
  INV_X1 U4115 ( .A(n4717), .ZN(n6140) );
  AND4_X1 U4116 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3251)
         );
  OR2_X1 U4117 ( .A1(n5643), .A2(n4380), .ZN(n3252) );
  INV_X1 U4118 ( .A(n6142), .ZN(n6687) );
  AND2_X1 U4119 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3253) );
  NAND2_X1 U4120 ( .A1(n3120), .A2(n4281), .ZN(n4317) );
  NAND2_X1 U4121 ( .A1(n6117), .A2(n5593), .ZN(n5591) );
  INV_X1 U4122 ( .A(n3520), .ZN(n3668) );
  NAND2_X1 U4123 ( .A1(n6695), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4072) );
  INV_X1 U4124 ( .A(n4280), .ZN(n3369) );
  INV_X1 U4125 ( .A(n4072), .ZN(n3747) );
  NAND2_X1 U4126 ( .A1(n4503), .A2(n3521), .ZN(n3441) );
  OR2_X1 U4127 ( .A1(n3683), .A2(n3682), .ZN(n3685) );
  AND2_X1 U4128 ( .A1(n3671), .A2(n3672), .ZN(n3688) );
  OAI211_X1 U4129 ( .C1(n3475), .C2(n3503), .A(n3474), .B(n3473), .ZN(n3545)
         );
  NAND2_X1 U4130 ( .A1(n3882), .A2(n3869), .ZN(n3870) );
  OR2_X1 U4131 ( .A1(n3572), .A2(n3571), .ZN(n3596) );
  OR2_X1 U4132 ( .A1(n3440), .A2(n3439), .ZN(n3521) );
  INV_X1 U4133 ( .A(n3308), .ZN(n3313) );
  AOI21_X1 U4134 ( .B1(n3340), .B2(INSTQUEUE_REG_12__3__SCAN_IN), .A(n3281), 
        .ZN(n3282) );
  AOI22_X1 U4135 ( .A1(n3100), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U4136 ( .A1(n3761), .A2(n3760), .ZN(n4801) );
  OR2_X1 U4137 ( .A1(n4068), .A2(n4067), .ZN(n4112) );
  INV_X1 U4138 ( .A(n5024), .ZN(n3783) );
  OR2_X1 U4139 ( .A1(n3615), .A2(n3614), .ZN(n3633) );
  AOI21_X1 U4140 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6359), .A(n3701), 
        .ZN(n3710) );
  AOI22_X1 U4141 ( .A1(n3315), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3295) );
  NAND2_X1 U4142 ( .A1(n4287), .A2(n3399), .ZN(n3410) );
  INV_X1 U4143 ( .A(n4070), .ZN(n4071) );
  INV_X1 U4144 ( .A(n4801), .ZN(n4802) );
  INV_X1 U4145 ( .A(n3445), .ZN(n3446) );
  NAND2_X1 U4146 ( .A1(n3502), .A2(n3501), .ZN(n5187) );
  OR2_X1 U4147 ( .A1(n4226), .A2(n6803), .ZN(n4228) );
  OR2_X1 U4148 ( .A1(n4096), .A2(n4095), .ZN(n4119) );
  NAND2_X1 U4149 ( .A1(n4240), .A2(n4239), .ZN(n4241) );
  INV_X1 U4150 ( .A(n5644), .ZN(n5645) );
  NOR2_X1 U4151 ( .A1(n5926), .A2(n4381), .ZN(n5822) );
  INV_X1 U4152 ( .A(n3130), .ZN(n6484) );
  INV_X1 U4153 ( .A(n4977), .ZN(n5229) );
  INV_X1 U4154 ( .A(n3540), .ZN(n3550) );
  AND2_X1 U4155 ( .A1(n6063), .A2(n4460), .ZN(n5870) );
  INV_X1 U4156 ( .A(n4024), .ZN(n4025) );
  INV_X1 U4157 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6020) );
  INV_X1 U4158 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5291) );
  OR2_X1 U4159 ( .A1(n4871), .A2(n4414), .ZN(n4415) );
  INV_X1 U4160 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5998) );
  INV_X1 U4161 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U4162 ( .A1(n4404), .A2(n6776), .ZN(n4405) );
  OR2_X1 U4163 ( .A1(n5779), .A2(n5713), .ZN(n5773) );
  OR2_X1 U4164 ( .A1(n5795), .A2(n4384), .ZN(n5790) );
  OR2_X1 U4165 ( .A1(n5937), .A2(n4386), .ZN(n5926) );
  INV_X1 U4166 ( .A(n5838), .ZN(n6209) );
  AND2_X1 U4167 ( .A1(n5711), .A2(n5416), .ZN(n5413) );
  OR2_X1 U4168 ( .A1(n4385), .A2(n4554), .ZN(n5711) );
  OR2_X1 U4169 ( .A1(n4385), .A2(n4839), .ZN(n5952) );
  OAI21_X1 U4170 ( .B1(n5966), .B2(n4786), .A(n5862), .ZN(n4889) );
  INV_X1 U4171 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6358) );
  AND2_X1 U4172 ( .A1(n6400), .A2(n6399), .ZN(n6404) );
  INV_X1 U4173 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U4174 ( .A1(n3129), .A2(n5181), .ZN(n6305) );
  AOI21_X1 U4175 ( .B1(n6398), .B2(STATE2_REG_3__SCAN_IN), .A(n5184), .ZN(
        n6406) );
  NOR2_X1 U4176 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5966) );
  AND2_X1 U4177 ( .A1(n4497), .A2(REIP_REG_31__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U4178 ( .A1(n5262), .A2(n4453), .ZN(n5871) );
  NAND2_X1 U4179 ( .A1(n4026), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4070)
         );
  INV_X1 U4180 ( .A(n5873), .ZN(n6056) );
  AND2_X1 U4181 ( .A1(n6084), .A2(n4455), .ZN(n6071) );
  AOI21_X1 U4182 ( .B1(n4220), .B2(n4219), .A(n4218), .ZN(n4398) );
  INV_X1 U4183 ( .A(n5591), .ZN(n6113) );
  AOI21_X1 U4184 ( .B1(n4691), .B2(n4865), .A(n4690), .ZN(n4693) );
  NOR2_X1 U4185 ( .A1(n4636), .A2(n3408), .ZN(n4729) );
  AND2_X1 U4186 ( .A1(n4839), .A2(n4609), .ZN(n4610) );
  INV_X1 U4187 ( .A(n4636), .ZN(n6139) );
  OAI21_X1 U4188 ( .B1(n3374), .B2(n6690), .A(n4595), .ZN(n4646) );
  OR2_X1 U4189 ( .A1(n4594), .A2(n4593), .ZN(n4692) );
  NAND2_X1 U4190 ( .A1(n3957), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3989)
         );
  AND2_X1 U4191 ( .A1(n5428), .A2(n5431), .ZN(n6108) );
  NAND2_X1 U4192 ( .A1(n3777), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3799)
         );
  NAND2_X1 U4193 ( .A1(n3767), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3776)
         );
  AND2_X1 U4194 ( .A1(n6252), .A2(n4388), .ZN(n5420) );
  OR2_X1 U4195 ( .A1(n6673), .A2(n4191), .ZN(n6253) );
  NAND2_X1 U4196 ( .A1(n5413), .A2(n5952), .ZN(n5838) );
  INV_X1 U4197 ( .A(n5711), .ZN(n6252) );
  INV_X1 U4198 ( .A(n6255), .ZN(n6266) );
  INV_X1 U4199 ( .A(n3118), .ZN(n6354) );
  AND2_X1 U4200 ( .A1(n4985), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6355) );
  INV_X1 U4201 ( .A(n6406), .ZN(n6525) );
  NOR2_X2 U4202 ( .A1(n5033), .A2(n6403), .ZN(n6301) );
  NOR2_X1 U4203 ( .A1(n4914), .A2(n4978), .ZN(n6307) );
  NOR2_X2 U4204 ( .A1(n6432), .A2(n6403), .ZN(n6477) );
  INV_X1 U4205 ( .A(n6481), .ZN(n6510) );
  NOR2_X2 U4206 ( .A1(n6432), .A2(n6305), .ZN(n6509) );
  INV_X1 U4207 ( .A(n6368), .ZN(n4983) );
  INV_X1 U4208 ( .A(n5139), .ZN(n5177) );
  OAI21_X1 U4209 ( .B1(n6530), .B2(n6529), .A(n6528), .ZN(n6577) );
  AND2_X1 U4210 ( .A1(n6516), .A2(n6430), .ZN(n6574) );
  NOR2_X1 U4211 ( .A1(n5855), .A2(n6305), .ZN(n6575) );
  INV_X1 U4212 ( .A(n6326), .ZN(n6541) );
  INV_X1 U4213 ( .A(n6347), .ZN(n6572) );
  INV_X1 U4214 ( .A(n6383), .ZN(n6554) );
  AND2_X1 U4215 ( .A1(n3103), .A2(DATAI_24_), .ZN(n6531) );
  AND2_X1 U4216 ( .A1(n3103), .A2(DATAI_27_), .ZN(n6549) );
  NOR2_X1 U4217 ( .A1(n6981), .A2(n6695), .ZN(n4786) );
  INV_X1 U4218 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6602) );
  INV_X1 U4219 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U4220 ( .A1(n4594), .A2(n5867), .ZN(n6685) );
  INV_X1 U4221 ( .A(n6094), .ZN(n6019) );
  NAND2_X1 U4222 ( .A1(n6084), .A2(n4416), .ZN(n5873) );
  NAND2_X1 U4223 ( .A1(n6134), .A2(n4695), .ZN(n6133) );
  INV_X1 U4224 ( .A(n4729), .ZN(n4708) );
  OR2_X1 U4225 ( .A1(n6139), .A2(n6687), .ZN(n4717) );
  INV_X1 U4226 ( .A(n4193), .ZN(n4194) );
  OR2_X1 U4227 ( .A1(n6188), .A2(n4710), .ZN(n6195) );
  NAND2_X1 U4228 ( .A1(n4186), .A2(n6409), .ZN(n5696) );
  AND2_X1 U4229 ( .A1(n4395), .A2(n3247), .ZN(n4396) );
  OR2_X1 U4230 ( .A1(n4385), .A2(n4284), .ZN(n6223) );
  INV_X1 U4231 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U4232 ( .A1(n6307), .A2(n6430), .ZN(n6348) );
  NAND2_X1 U4233 ( .A1(n6307), .A2(n6306), .ZN(n6395) );
  AOI22_X1 U4234 ( .A1(n6405), .A2(n6402), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6408), .ZN(n6429) );
  OR2_X1 U4235 ( .A1(n6432), .A2(n6431), .ZN(n6481) );
  AOI22_X1 U4236 ( .A1(n6489), .A2(n6492), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6487), .ZN(n6514) );
  NAND2_X1 U4237 ( .A1(n6516), .A2(n4983), .ZN(n5258) );
  NAND2_X1 U4238 ( .A1(n6516), .A2(n4915), .ZN(n5139) );
  AOI22_X1 U4239 ( .A1(n5141), .A2(n6517), .B1(n6363), .B2(n5138), .ZN(n5180)
         );
  AOI22_X1 U4240 ( .A1(n6524), .A2(n6529), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6520), .ZN(n6581) );
  INV_X1 U4241 ( .A(n6575), .ZN(n5220) );
  OR2_X1 U4242 ( .A1(n4888), .A2(n6403), .ZN(n5076) );
  INV_X1 U4243 ( .A(n6543), .ZN(n6457) );
  INV_X1 U4244 ( .A(n6561), .ZN(n6469) );
  NAND2_X1 U4245 ( .A1(n4943), .A2(n5136), .ZN(n5111) );
  INV_X1 U4246 ( .A(n6661), .ZN(n6592) );
  INV_X1 U4247 ( .A(READY_N), .ZN(n6690) );
  AND2_X1 U4248 ( .A1(n6602), .A2(STATE_REG_1__SCAN_IN), .ZN(n6684) );
  INV_X1 U4249 ( .A(n6650), .ZN(n6655) );
  NAND2_X1 U4250 ( .A1(n4516), .A2(n4515), .ZN(U2830) );
  OAI211_X1 U4251 ( .C1(n5738), .C2(n6172), .A(n4195), .B(n4194), .ZN(U2957)
         );
  NAND2_X1 U4252 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5742) );
  INV_X1 U4253 ( .A(n5742), .ZN(n5706) );
  INV_X1 U4254 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3254) );
  AND2_X2 U4255 ( .A1(n3259), .A2(n4746), .ZN(n3434) );
  AOI22_X1 U4256 ( .A1(n4201), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4257 ( .A1(n3356), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3256) );
  AND2_X2 U4258 ( .A1(n4751), .A2(n3259), .ZN(n3314) );
  AND2_X2 U4259 ( .A1(n4751), .A2(n4582), .ZN(n3351) );
  AOI22_X1 U4260 ( .A1(n3351), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3124), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4261 ( .A1(n3113), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4262 ( .A1(n3100), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4263 ( .A1(n3301), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3124), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4264 ( .A1(n4201), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4265 ( .A1(n3314), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4266 ( .A1(n3433), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4267 ( .A1(n3351), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4268 ( .A1(n3101), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4269 ( .A1(n3302), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4270 ( .A1(n4201), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4271 ( .A1(n3314), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4272 ( .A1(n3351), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4273 ( .A1(n3315), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4274 ( .A1(n3351), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4275 ( .A1(n3314), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4276 ( .A1(n4201), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4277 ( .A1(n3113), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4278 ( .A1(n3101), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4279 ( .A1(n3356), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4280 ( .A1(n3113), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4281 ( .A1(n3302), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4282 ( .A1(n3314), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4283 ( .A1(n3351), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4284 ( .A1(n3315), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3303) );
  NAND3_X1 U4285 ( .A1(n3407), .A2(n4504), .A3(n3382), .ZN(n3322) );
  AOI22_X1 U4286 ( .A1(n3356), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4287 ( .A1(n3113), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4288 ( .A1(n3100), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3309) );
  NAND3_X1 U4289 ( .A1(n3311), .A2(n3310), .A3(n3309), .ZN(n3312) );
  AOI22_X1 U4290 ( .A1(n3351), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4291 ( .A1(n3314), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4292 ( .A1(n3302), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4293 ( .A1(n3315), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4294 ( .A1(n3322), .A2(n3386), .ZN(n3326) );
  NAND2_X1 U4295 ( .A1(n3722), .A2(n3381), .ZN(n3323) );
  NAND2_X1 U4296 ( .A1(n3399), .A2(n3324), .ZN(n3325) );
  AND3_X2 U4297 ( .A1(n3327), .A2(n3326), .A3(n3325), .ZN(n3389) );
  NAND2_X1 U4298 ( .A1(n3314), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3331)
         );
  NAND2_X1 U4299 ( .A1(n3315), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4300 ( .A1(n3113), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3329)
         );
  NAND2_X1 U4301 ( .A1(n3433), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4302 ( .A1(n3351), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3335)
         );
  NAND2_X1 U4303 ( .A1(n3302), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4304 ( .A1(n3301), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4305 ( .A1(n3452), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4306 ( .A1(n3101), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4307 ( .A1(n3350), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U4308 ( .A1(n3434), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U4309 ( .A1(n3316), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3336)
         );
  NAND2_X1 U4310 ( .A1(n4201), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4311 ( .A1(n3356), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3343)
         );
  NAND2_X1 U4312 ( .A1(n3340), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3342)
         );
  NAND2_X1 U4313 ( .A1(n3465), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3341) );
  AND3_X1 U4314 ( .A1(n3382), .A2(n3408), .A3(n3119), .ZN(n3349) );
  AOI22_X1 U4315 ( .A1(n3123), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4316 ( .A1(n3314), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4317 ( .A1(n3351), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4318 ( .A1(n4201), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4319 ( .A1(n3100), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4320 ( .A1(n3356), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4321 ( .A1(n4129), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3357) );
  NAND3_X1 U4322 ( .A1(n4504), .A2(n3382), .A3(n4893), .ZN(n4271) );
  INV_X1 U4323 ( .A(n4271), .ZN(n3365) );
  XNOR2_X1 U4324 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4253) );
  NAND2_X1 U4325 ( .A1(n3374), .A2(n4253), .ZN(n3377) );
  NAND2_X1 U4326 ( .A1(n4410), .A2(n3377), .ZN(n3370) );
  INV_X1 U4327 ( .A(n3379), .ZN(n4287) );
  NOR2_X1 U4328 ( .A1(n3410), .A2(n5435), .ZN(n3368) );
  NAND3_X1 U4329 ( .A1(n4282), .A2(n3370), .A3(n3369), .ZN(n3371) );
  NAND2_X1 U4330 ( .A1(n3371), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3393) );
  INV_X1 U4331 ( .A(n3393), .ZN(n3373) );
  NAND2_X1 U4332 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4843) );
  OAI21_X1 U4333 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n4843), .ZN(n5182) );
  NAND2_X1 U4334 ( .A1(n3373), .A2(n3372), .ZN(n3395) );
  NAND2_X1 U4335 ( .A1(n3406), .A2(n4271), .ZN(n3376) );
  NAND2_X1 U4336 ( .A1(n3396), .A2(n3531), .ZN(n4578) );
  NAND2_X1 U4337 ( .A1(n4268), .A2(n3381), .ZN(n3401) );
  NAND2_X1 U4338 ( .A1(n3377), .A2(n3363), .ZN(n3378) );
  INV_X1 U4339 ( .A(n3380), .ZN(n3383) );
  NAND2_X1 U4340 ( .A1(n3385), .A2(n3384), .ZN(n3404) );
  NAND3_X1 U4341 ( .A1(n3414), .A2(n3387), .A3(n3718), .ZN(n3388) );
  NAND2_X1 U4342 ( .A1(n3388), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4343 ( .A1(n3389), .A2(n3374), .ZN(n3398) );
  INV_X1 U4344 ( .A(n3503), .ZN(n3442) );
  NAND2_X1 U4345 ( .A1(n3398), .A2(n3442), .ZN(n3390) );
  AOI21_X1 U4346 ( .B1(n3421), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3392), 
        .ZN(n3394) );
  NAND2_X1 U4347 ( .A1(n3394), .A2(n3393), .ZN(n3419) );
  AND2_X2 U4348 ( .A1(n3395), .A2(n3419), .ZN(n3444) );
  INV_X1 U4349 ( .A(n3396), .ZN(n3397) );
  INV_X1 U4350 ( .A(n3401), .ZN(n3403) );
  OAI21_X1 U4351 ( .B1(n3404), .B2(n3403), .A(n3120), .ZN(n3413) );
  OR2_X1 U4352 ( .A1(n6673), .A2(n6952), .ZN(n6583) );
  AOI21_X1 U4353 ( .B1(n3405), .B2(n3406), .A(n6583), .ZN(n3412) );
  NAND2_X1 U4354 ( .A1(n3408), .A2(n3381), .ZN(n3409) );
  NOR2_X1 U4355 ( .A1(n3407), .A2(n3409), .ZN(n3411) );
  INV_X1 U4356 ( .A(n3410), .ZN(n4506) );
  NAND2_X1 U4357 ( .A1(n3411), .A2(n4506), .ZN(n4762) );
  NAND2_X1 U4358 ( .A1(n4374), .A2(n3415), .ZN(n3476) );
  NAND2_X1 U4359 ( .A1(n3421), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3418) );
  INV_X1 U4360 ( .A(n3717), .ZN(n3424) );
  INV_X1 U4361 ( .A(n4187), .ZN(n3425) );
  MUX2_X1 U4362 ( .A(n3424), .B(n3425), .S(n6398), .Z(n3416) );
  INV_X1 U4363 ( .A(n3416), .ZN(n3417) );
  NAND2_X1 U4364 ( .A1(n3476), .A2(n3477), .ZN(n3445) );
  NAND2_X1 U4365 ( .A1(n3444), .A2(n3445), .ZN(n3420) );
  NAND2_X1 U4366 ( .A1(n3420), .A2(n3419), .ZN(n3496) );
  NAND2_X1 U4367 ( .A1(n3421), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3427) );
  INV_X1 U4368 ( .A(n4843), .ZN(n3422) );
  NAND2_X1 U4369 ( .A1(n3422), .A2(n6279), .ZN(n6308) );
  NAND2_X1 U4370 ( .A1(n4843), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3423) );
  NAND2_X1 U4371 ( .A1(n6308), .A2(n3423), .ZN(n4985) );
  AOI22_X1 U4372 ( .A1(n3425), .A2(n4985), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3424), .ZN(n3426) );
  NAND2_X1 U4373 ( .A1(n3427), .A2(n3426), .ZN(n3497) );
  XNOR2_X1 U4374 ( .A(n3496), .B(n3497), .ZN(n4760) );
  AOI22_X1 U4375 ( .A1(n3302), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4376 ( .A1(n3314), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4377 ( .A1(n4200), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3430) );
  INV_X1 U4378 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4379 ( .A1(n3315), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3429) );
  NAND4_X1 U4380 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3440)
         );
  AOI22_X1 U4381 ( .A1(n4062), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4382 ( .A1(n3101), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U4383 ( .A1(n3117), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4384 ( .A1(n3113), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3435) );
  NAND4_X1 U4385 ( .A1(n3438), .A2(n3437), .A3(n3436), .A4(n3435), .ZN(n3439)
         );
  AOI22_X1 U4386 ( .A1(n3442), .A2(n3521), .B1(n3687), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3443) );
  XNOR2_X2 U4387 ( .A(n3447), .B(n3446), .ZN(n4575) );
  AOI22_X1 U4388 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n3101), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4389 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4128), .B1(n3113), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4390 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n3117), .B1(n4198), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4391 ( .A1(n4200), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4392 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3458)
         );
  AOI22_X1 U4393 ( .A1(n3315), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4394 ( .A1(n4753), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4395 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n4123), .B1(n3135), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4396 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n4062), .B1(n3483), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3453) );
  NAND4_X1 U4397 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3457)
         );
  NAND2_X1 U4398 ( .A1(n4503), .A2(n3549), .ZN(n3459) );
  INV_X1 U4399 ( .A(n3549), .ZN(n3475) );
  AOI22_X1 U4400 ( .A1(n3302), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4401 ( .A1(n4123), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4402 ( .A1(n4200), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3462) );
  INV_X1 U4403 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6818) );
  AOI22_X1 U4404 ( .A1(n4029), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3461) );
  NAND4_X1 U4405 ( .A1(n3464), .A2(n3463), .A3(n3462), .A4(n3461), .ZN(n3471)
         );
  AOI22_X1 U4406 ( .A1(n4062), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4407 ( .A1(n3101), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4408 ( .A1(n3116), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4409 ( .A1(n3113), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4410 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3470)
         );
  INV_X1 U4411 ( .A(n3642), .ZN(n3472) );
  AND2_X1 U4412 ( .A1(n4503), .A2(n3472), .ZN(n3490) );
  INV_X1 U4413 ( .A(n3490), .ZN(n3474) );
  NAND2_X1 U4414 ( .A1(n3687), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3473) );
  INV_X1 U4415 ( .A(n3476), .ZN(n3478) );
  AOI22_X1 U4416 ( .A1(n3302), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4417 ( .A1(n4062), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4418 ( .A1(n4128), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4419 ( .A1(n4753), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3479) );
  NAND4_X1 U4420 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3489)
         );
  AOI22_X1 U4421 ( .A1(n4029), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4422 ( .A1(n3101), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4423 ( .A1(n4200), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4424 ( .A1(n3134), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3484) );
  NAND4_X1 U4425 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3488)
         );
  MUX2_X1 U4426 ( .A(n3490), .B(n3495), .S(n3550), .Z(n3536) );
  INV_X1 U4427 ( .A(n3536), .ZN(n3491) );
  NAND2_X1 U4428 ( .A1(n3687), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3494) );
  AOI21_X1 U4429 ( .B1(n3408), .B2(n3540), .A(n6952), .ZN(n3493) );
  NAND3_X1 U4430 ( .A1(n3494), .A2(n3493), .A3(n3492), .ZN(n3537) );
  INV_X1 U4431 ( .A(n3496), .ZN(n3498) );
  NAND2_X1 U4432 ( .A1(n3421), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3502) );
  NAND3_X1 U4433 ( .A1(n6359), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6490) );
  INV_X1 U4434 ( .A(n6490), .ZN(n6487) );
  NAND2_X1 U4435 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6487), .ZN(n6488) );
  NAND2_X1 U4436 ( .A1(n6359), .A2(n6488), .ZN(n3499) );
  NAND3_X1 U4437 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5075) );
  INV_X1 U4438 ( .A(n5075), .ZN(n4948) );
  NAND2_X1 U4439 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4948), .ZN(n4972) );
  NAND2_X1 U4440 ( .A1(n3499), .A2(n4972), .ZN(n4980) );
  OAI22_X1 U4441 ( .A1(n4187), .A2(n4980), .B1(n3717), .B2(n6359), .ZN(n3500)
         );
  INV_X1 U4442 ( .A(n3500), .ZN(n3501) );
  NAND2_X1 U4443 ( .A1(n4742), .A2(n6952), .ZN(n3516) );
  AOI22_X1 U4444 ( .A1(n3314), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4445 ( .A1(n4128), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4446 ( .A1(n4753), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3506) );
  AOI22_X1 U4447 ( .A1(n4062), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3505) );
  NAND4_X1 U4448 ( .A1(n3508), .A2(n3507), .A3(n3506), .A4(n3505), .ZN(n3514)
         );
  AOI22_X1 U4449 ( .A1(n4200), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4450 ( .A1(n3113), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4451 ( .A1(n4029), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4452 ( .A1(n3101), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3509) );
  NAND4_X1 U4453 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3513)
         );
  AOI22_X1 U4454 ( .A1(n3714), .A2(n3575), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3687), .ZN(n3515) );
  NAND2_X1 U4455 ( .A1(n3517), .A2(n4883), .ZN(n3519) );
  INV_X1 U4456 ( .A(n4883), .ZN(n5222) );
  NAND2_X1 U4457 ( .A1(n3540), .A2(n3549), .ZN(n3530) );
  INV_X1 U4458 ( .A(n3521), .ZN(n3529) );
  NAND2_X1 U4459 ( .A1(n3530), .A2(n3529), .ZN(n3576) );
  INV_X1 U4460 ( .A(n3575), .ZN(n3522) );
  XNOR2_X1 U4461 ( .A(n3576), .B(n3522), .ZN(n3523) );
  NAND2_X1 U4462 ( .A1(n3523), .A2(n3406), .ZN(n3524) );
  INV_X1 U4463 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6273) );
  OR2_X1 U4464 ( .A1(n4782), .A2(n3106), .ZN(n3534) );
  XNOR2_X1 U4465 ( .A(n3530), .B(n3529), .ZN(n3532) );
  AND2_X1 U4466 ( .A1(n3408), .A2(n3531), .ZN(n3539) );
  AOI21_X1 U4467 ( .B1(n3532), .B2(n3406), .A(n3539), .ZN(n3533) );
  NAND2_X1 U4468 ( .A1(n3534), .A2(n3533), .ZN(n4790) );
  NAND2_X1 U4469 ( .A1(n4790), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3557)
         );
  NAND2_X1 U4470 ( .A1(n3535), .A2(n3537), .ZN(n3538) );
  MUX2_X2 U4471 ( .A(n3538), .B(n3537), .S(n3536), .Z(n5136) );
  INV_X1 U4472 ( .A(n3406), .ZN(n4867) );
  INV_X1 U4473 ( .A(n3539), .ZN(n4375) );
  OAI21_X1 U4474 ( .B1(n4867), .B2(n3540), .A(n4375), .ZN(n3541) );
  INV_X1 U4475 ( .A(n3541), .ZN(n3542) );
  NAND2_X1 U4476 ( .A1(n4638), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3543)
         );
  INV_X1 U4477 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U4478 ( .A1(n3543), .A2(n6795), .ZN(n3544) );
  AND2_X1 U4479 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4794) );
  NAND2_X1 U4480 ( .A1(n4638), .A2(n4794), .ZN(n3555) );
  AND2_X1 U4481 ( .A1(n3544), .A2(n3555), .ZN(n4680) );
  NAND2_X1 U4482 ( .A1(n3129), .A2(n3668), .ZN(n3554) );
  XNOR2_X1 U4483 ( .A(n3550), .B(n3549), .ZN(n3552) );
  NAND3_X1 U4484 ( .A1(n3399), .A2(n3119), .A3(n3531), .ZN(n3551) );
  AOI21_X1 U4485 ( .B1(n3552), .B2(n3406), .A(n3551), .ZN(n3553) );
  NAND2_X1 U4486 ( .A1(n3554), .A2(n3553), .ZN(n4679) );
  INV_X1 U4487 ( .A(n3555), .ZN(n3556) );
  NAND2_X1 U4488 ( .A1(n3557), .A2(n4792), .ZN(n3560) );
  INV_X1 U4489 ( .A(n4790), .ZN(n3558) );
  INV_X1 U4490 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4305) );
  NAND2_X1 U4491 ( .A1(n3558), .A2(n4305), .ZN(n3559) );
  NAND2_X1 U4492 ( .A1(n3561), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3562)
         );
  AOI22_X1 U4493 ( .A1(n3302), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4494 ( .A1(n4123), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4495 ( .A1(n4200), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4496 ( .A1(n4029), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4497 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3572)
         );
  AOI22_X1 U4498 ( .A1(n4062), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4499 ( .A1(n3101), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4500 ( .A1(n3117), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4501 ( .A1(n3113), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4502 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3571)
         );
  NAND2_X1 U4503 ( .A1(n3714), .A2(n3596), .ZN(n3574) );
  NAND2_X1 U4504 ( .A1(n3687), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3573) );
  XNOR2_X1 U4505 ( .A(n3582), .B(n3583), .ZN(n3771) );
  NAND2_X1 U4506 ( .A1(n3771), .A2(n3668), .ZN(n3579) );
  NAND2_X1 U4507 ( .A1(n3576), .A2(n3575), .ZN(n3598) );
  XNOR2_X1 U4508 ( .A(n3598), .B(n3596), .ZN(n3577) );
  NAND2_X1 U4509 ( .A1(n3577), .A2(n3406), .ZN(n3578) );
  NAND2_X1 U4510 ( .A1(n3579), .A2(n3578), .ZN(n3580) );
  INV_X1 U4511 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6263) );
  XNOR2_X1 U4512 ( .A(n3580), .B(n6263), .ZN(n6180) );
  NAND2_X1 U4513 ( .A1(n3580), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3581)
         );
  AOI22_X1 U4514 ( .A1(n4200), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4515 ( .A1(n4029), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4516 ( .A1(n3113), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4517 ( .A1(n3302), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3584) );
  NAND4_X1 U4518 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(n3593)
         );
  AOI22_X1 U4519 ( .A1(n4128), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4520 ( .A1(n4142), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4521 ( .A1(n3101), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4522 ( .A1(n4062), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3588) );
  NAND4_X1 U4523 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3592)
         );
  NAND2_X1 U4524 ( .A1(n3714), .A2(n3621), .ZN(n3595) );
  NAND2_X1 U4525 ( .A1(n3687), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4526 ( .A1(n3595), .A2(n3594), .ZN(n3605) );
  XNOR2_X1 U4527 ( .A(n3604), .B(n3605), .ZN(n3772) );
  NAND2_X1 U4528 ( .A1(n3772), .A2(n3668), .ZN(n3601) );
  INV_X1 U4529 ( .A(n3596), .ZN(n3597) );
  OR2_X1 U4530 ( .A1(n3598), .A2(n3597), .ZN(n3620) );
  XNOR2_X1 U4531 ( .A(n3620), .B(n3621), .ZN(n3599) );
  NAND2_X1 U4532 ( .A1(n3599), .A2(n3406), .ZN(n3600) );
  NAND2_X1 U4533 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  INV_X1 U4534 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6718) );
  XNOR2_X1 U4535 ( .A(n3602), .B(n6718), .ZN(n5113) );
  NAND2_X1 U4536 ( .A1(n3602), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3603)
         );
  AOI22_X1 U4537 ( .A1(n3123), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4538 ( .A1(n4123), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4539 ( .A1(n4200), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3607) );
  INV_X1 U4540 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6785) );
  AOI22_X1 U4541 ( .A1(n4029), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3606) );
  NAND4_X1 U4542 ( .A1(n3609), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(n3615)
         );
  AOI22_X1 U4543 ( .A1(n4062), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4544 ( .A1(n3101), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4545 ( .A1(n3117), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4546 ( .A1(n3113), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3610) );
  NAND4_X1 U4547 ( .A1(n3613), .A2(n3612), .A3(n3611), .A4(n3610), .ZN(n3614)
         );
  AOI22_X1 U4548 ( .A1(n3714), .A2(n3633), .B1(n3687), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3618) );
  NAND2_X1 U4549 ( .A1(n3619), .A2(n3618), .ZN(n3782) );
  INV_X1 U4550 ( .A(n3620), .ZN(n3622) );
  NAND2_X1 U4551 ( .A1(n3622), .A2(n3621), .ZN(n3632) );
  XNOR2_X1 U4552 ( .A(n3632), .B(n3633), .ZN(n3623) );
  NAND2_X1 U4553 ( .A1(n3623), .A2(n3406), .ZN(n3624) );
  NAND2_X1 U4554 ( .A1(n3625), .A2(n3624), .ZN(n3627) );
  INV_X1 U4555 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3626) );
  XNOR2_X1 U4556 ( .A(n3627), .B(n3626), .ZN(n4523) );
  NAND2_X1 U4557 ( .A1(n3714), .A2(n3642), .ZN(n3629) );
  NAND2_X1 U4558 ( .A1(n3687), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3628) );
  NAND2_X1 U4559 ( .A1(n3629), .A2(n3628), .ZN(n3630) );
  NAND2_X1 U4560 ( .A1(n3788), .A2(n3668), .ZN(n3637) );
  INV_X1 U4561 ( .A(n3632), .ZN(n3634) );
  NAND2_X1 U4562 ( .A1(n3634), .A2(n3633), .ZN(n3644) );
  XNOR2_X1 U4563 ( .A(n3644), .B(n3642), .ZN(n3635) );
  NAND2_X1 U4564 ( .A1(n3635), .A2(n3406), .ZN(n3636) );
  NAND2_X1 U4565 ( .A1(n3637), .A2(n3636), .ZN(n3638) );
  INV_X1 U4566 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6913) );
  XNOR2_X1 U4567 ( .A(n3638), .B(n6913), .ZN(n5128) );
  NAND2_X1 U4568 ( .A1(n3638), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3639)
         );
  NAND2_X1 U4569 ( .A1(n3406), .A2(n3642), .ZN(n3643) );
  OR2_X1 U4570 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  NAND2_X1 U4571 ( .A1(n5643), .A2(n3645), .ZN(n3646) );
  INV_X1 U4572 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6229) );
  XNOR2_X1 U4573 ( .A(n3646), .B(n6229), .ZN(n5308) );
  NAND2_X1 U4574 ( .A1(n3646), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3647)
         );
  INV_X1 U4575 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U4576 ( .A1(n5643), .A2(n6967), .ZN(n5315) );
  NAND2_X1 U4577 ( .A1(n3140), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5316)
         );
  INV_X1 U4578 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3648) );
  NAND2_X1 U4579 ( .A1(n5643), .A2(n3648), .ZN(n5358) );
  INV_X1 U4580 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3649) );
  AND2_X1 U4581 ( .A1(n5643), .A2(n3649), .ZN(n3652) );
  NAND2_X1 U4582 ( .A1(n3140), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U4583 ( .A1(n3140), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3650) );
  AND2_X1 U4584 ( .A1(n6162), .A2(n3650), .ZN(n3651) );
  INV_X1 U4585 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U4586 ( .A1(n5643), .A2(n4380), .ZN(n5386) );
  XNOR2_X1 U4587 ( .A(n6164), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5921)
         );
  NAND2_X1 U4588 ( .A1(n5922), .A2(n5921), .ZN(n3654) );
  INV_X1 U4589 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6721) );
  NAND2_X1 U4590 ( .A1(n5643), .A2(n6721), .ZN(n3653) );
  NAND2_X1 U4591 ( .A1(n3140), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3655) );
  INV_X1 U4592 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5942) );
  NOR2_X1 U4593 ( .A1(n6164), .A2(n5942), .ZN(n3657) );
  NAND2_X1 U4594 ( .A1(n5643), .A2(n5942), .ZN(n3656) );
  AND2_X1 U4595 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4392) );
  NAND2_X1 U4596 ( .A1(n4392), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3658) );
  INV_X1 U4597 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5840) );
  INV_X1 U4598 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5930) );
  INV_X1 U4599 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5832) );
  NAND3_X1 U4600 ( .A1(n5840), .A2(n5930), .A3(n5832), .ZN(n3659) );
  NAND2_X1 U4601 ( .A1(n3140), .A2(n3659), .ZN(n3660) );
  NAND2_X2 U4602 ( .A1(n4251), .A2(n3660), .ZN(n4249) );
  AND2_X1 U4603 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5813) );
  AND2_X1 U4604 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5705) );
  AND2_X1 U4605 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4384) );
  INV_X1 U4606 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5777) );
  INV_X1 U4607 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6723) );
  INV_X1 U4608 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5778) );
  INV_X1 U4609 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3661) );
  NAND4_X1 U4610 ( .A1(n5777), .A2(n6723), .A3(n5778), .A4(n3661), .ZN(n3662)
         );
  INV_X1 U4611 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5821) );
  INV_X1 U4612 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U4613 ( .A1(n5821), .A2(n6935), .ZN(n5814) );
  NOR2_X1 U4614 ( .A1(n3662), .A2(n5814), .ZN(n3663) );
  XNOR2_X1 U4615 ( .A(n6164), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5634)
         );
  INV_X1 U4616 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U4617 ( .A1(n5643), .A2(n5761), .ZN(n3664) );
  NAND2_X1 U4618 ( .A1(n5643), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5623) );
  INV_X1 U4619 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5752) );
  INV_X1 U4620 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U4621 ( .A1(n5752), .A2(n6983), .ZN(n5743) );
  NOR2_X1 U4622 ( .A1(n6164), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4224)
         );
  INV_X1 U4623 ( .A(n4224), .ZN(n5624) );
  AOI21_X1 U4624 ( .B1(n5706), .B2(n4238), .A(n4404), .ZN(n3665) );
  INV_X1 U4625 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6776) );
  XNOR2_X1 U4626 ( .A(n3665), .B(n6776), .ZN(n5738) );
  NAND2_X1 U4627 ( .A1(n6358), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3684) );
  NAND2_X1 U4628 ( .A1(n3254), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U4629 ( .A1(n3684), .A2(n3666), .ZN(n3683) );
  NAND2_X1 U4630 ( .A1(n6398), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3682) );
  INV_X1 U4631 ( .A(n3682), .ZN(n3667) );
  XNOR2_X1 U4632 ( .A(n3683), .B(n3667), .ZN(n4255) );
  NAND2_X1 U4633 ( .A1(n3714), .A2(n3120), .ZN(n3669) );
  NAND2_X1 U4634 ( .A1(n3669), .A2(n3119), .ZN(n3679) );
  NAND2_X1 U4635 ( .A1(n4838), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3670) );
  NAND2_X1 U4636 ( .A1(n3682), .A2(n3670), .ZN(n3674) );
  AOI21_X1 U4637 ( .B1(n4503), .B2(n3119), .A(n3674), .ZN(n3673) );
  NAND2_X1 U4638 ( .A1(n3374), .A2(n3119), .ZN(n3672) );
  OAI21_X1 U4639 ( .B1(n3673), .B2(n3408), .A(n3688), .ZN(n3678) );
  INV_X1 U4640 ( .A(n3674), .ZN(n3675) );
  NAND2_X1 U4641 ( .A1(n3714), .A2(n3675), .ZN(n3676) );
  NAND2_X1 U4642 ( .A1(n3676), .A2(n3705), .ZN(n3677) );
  OAI211_X1 U4643 ( .C1(n3679), .C2(n4255), .A(n3678), .B(n3677), .ZN(n3681)
         );
  NAND3_X1 U4644 ( .A1(n3679), .A2(n4255), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3680) );
  OAI211_X1 U4645 ( .C1(n4255), .C2(n3705), .A(n3681), .B(n3680), .ZN(n3692)
         );
  NAND2_X1 U4646 ( .A1(n3685), .A2(n3684), .ZN(n3695) );
  NAND2_X1 U4647 ( .A1(n6279), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3696) );
  NAND2_X1 U4648 ( .A1(n3194), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3686) );
  NAND2_X1 U4649 ( .A1(n3696), .A2(n3686), .ZN(n3693) );
  XNOR2_X1 U4650 ( .A(n3695), .B(n3693), .ZN(n4256) );
  INV_X1 U4651 ( .A(n3687), .ZN(n3704) );
  NAND2_X1 U4652 ( .A1(n3714), .A2(n4256), .ZN(n3689) );
  OAI211_X1 U4653 ( .C1(n4256), .C2(n3704), .A(n3689), .B(n3688), .ZN(n3691)
         );
  NOR2_X1 U4654 ( .A1(n3689), .A2(n3688), .ZN(n3690) );
  AOI21_X1 U4655 ( .B1(n3692), .B2(n3691), .A(n3690), .ZN(n3708) );
  INV_X1 U4656 ( .A(n3693), .ZN(n3694) );
  NAND2_X1 U4657 ( .A1(n3695), .A2(n3694), .ZN(n3697) );
  NAND2_X1 U4658 ( .A1(n3697), .A2(n3696), .ZN(n3699) );
  XNOR2_X1 U4659 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3698) );
  NAND3_X1 U4660 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3710), .A3(n5964), .ZN(n3703) );
  NOR2_X1 U4661 ( .A1(n3699), .A2(n3698), .ZN(n3700) );
  NOR2_X1 U4662 ( .A1(n3701), .A2(n3700), .ZN(n3702) );
  NAND2_X1 U4663 ( .A1(n3703), .A2(n3702), .ZN(n4260) );
  AND2_X1 U4664 ( .A1(n4260), .A2(n3704), .ZN(n3707) );
  AOI22_X1 U4665 ( .A1(n4260), .A2(n3711), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6952), .ZN(n3706) );
  OAI21_X1 U4666 ( .B1(n3708), .B2(n3707), .A(n3706), .ZN(n3713) );
  NOR2_X1 U4667 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6276), .ZN(n3709)
         );
  NAND2_X1 U4668 ( .A1(n4257), .A2(n3711), .ZN(n3712) );
  NAND2_X1 U4669 ( .A1(n3713), .A2(n3712), .ZN(n3716) );
  NAND2_X1 U4670 ( .A1(n3381), .A2(n3119), .ZN(n3719) );
  NAND2_X1 U4671 ( .A1(n4267), .A2(n3408), .ZN(n3720) );
  NAND2_X1 U4672 ( .A1(n3718), .A2(n3720), .ZN(n4279) );
  NAND2_X1 U4673 ( .A1(n3382), .A2(n3119), .ZN(n3721) );
  NAND2_X1 U4674 ( .A1(n3128), .A2(n3894), .ZN(n3728) );
  AOI22_X1 U4675 ( .A1(n3731), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6695), .ZN(n3726) );
  INV_X1 U4676 ( .A(n5435), .ZN(n3724) );
  NAND2_X1 U4677 ( .A1(n3752), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3725) );
  AND2_X1 U4678 ( .A1(n3726), .A2(n3725), .ZN(n3727) );
  NAND2_X1 U4679 ( .A1(n3728), .A2(n3727), .ZN(n4674) );
  INV_X1 U4680 ( .A(n3407), .ZN(n3729) );
  NAND2_X1 U4681 ( .A1(n5136), .A2(n3729), .ZN(n4600) );
  NAND2_X1 U4682 ( .A1(n3130), .A2(n3894), .ZN(n3735) );
  AOI22_X1 U4683 ( .A1(n3731), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6695), .ZN(n3733) );
  NAND2_X1 U4684 ( .A1(n3752), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3732) );
  AND2_X1 U4685 ( .A1(n3733), .A2(n3732), .ZN(n3734) );
  NAND2_X1 U4686 ( .A1(n3735), .A2(n3734), .ZN(n4602) );
  AND2_X1 U4687 ( .A1(n4602), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3736) );
  NAND2_X1 U4688 ( .A1(n4600), .A2(n3736), .ZN(n4601) );
  INV_X1 U4689 ( .A(n4602), .ZN(n3737) );
  NAND2_X1 U4690 ( .A1(n3737), .A2(n3739), .ZN(n3738) );
  NAND2_X1 U4691 ( .A1(n4601), .A2(n3738), .ZN(n4673) );
  NAND2_X1 U4692 ( .A1(n3752), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3743) );
  INV_X1 U4693 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6726) );
  NAND2_X1 U4694 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3753) );
  OAI21_X1 U4695 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3753), .ZN(n6196) );
  NAND2_X1 U4696 ( .A1(n3739), .A2(n6196), .ZN(n3740) );
  OAI21_X1 U4697 ( .B1(n6726), .B2(n4072), .A(n3740), .ZN(n3741) );
  AOI21_X1 U4698 ( .B1(n4221), .B2(EAX_REG_2__SCAN_IN), .A(n3741), .ZN(n3742)
         );
  AND2_X1 U4699 ( .A1(n3743), .A2(n3742), .ZN(n4733) );
  NAND2_X1 U4700 ( .A1(n3744), .A2(n4733), .ZN(n3751) );
  INV_X1 U4701 ( .A(n3744), .ZN(n3746) );
  INV_X1 U4702 ( .A(n4733), .ZN(n3745) );
  NAND2_X1 U4703 ( .A1(n3746), .A2(n3745), .ZN(n3749) );
  OAI21_X1 U4704 ( .B1(n4782), .B2(n3911), .A(n4072), .ZN(n3748) );
  INV_X1 U4705 ( .A(n3748), .ZN(n4732) );
  NAND2_X1 U4706 ( .A1(n3749), .A2(n4732), .ZN(n3750) );
  NAND2_X1 U4707 ( .A1(n3751), .A2(n3750), .ZN(n4731) );
  INV_X1 U4708 ( .A(n4731), .ZN(n3762) );
  INV_X1 U4709 ( .A(n3752), .ZN(n3765) );
  INV_X1 U4710 ( .A(n3753), .ZN(n3754) );
  NOR2_X1 U4711 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3754), .ZN(n3755)
         );
  NOR2_X1 U4712 ( .A1(n3767), .A2(n3755), .ZN(n6072) );
  INV_X1 U4713 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3756) );
  OAI22_X1 U4714 ( .A1(n6072), .A2(n4216), .B1(n4072), .B2(n3756), .ZN(n3757)
         );
  AOI21_X1 U4715 ( .B1(n4221), .B2(EAX_REG_3__SCAN_IN), .A(n3757), .ZN(n3758)
         );
  OAI21_X1 U4716 ( .B1(n3195), .B2(n3765), .A(n3758), .ZN(n3759) );
  NAND2_X1 U4717 ( .A1(n3762), .A2(n4801), .ZN(n4803) );
  NAND2_X1 U4718 ( .A1(n6695), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3764)
         );
  NAND2_X1 U4719 ( .A1(n4221), .A2(EAX_REG_4__SCAN_IN), .ZN(n3763) );
  OAI211_X1 U4720 ( .C1(n3765), .C2(n5964), .A(n3764), .B(n3763), .ZN(n3766)
         );
  NAND2_X1 U4721 ( .A1(n3766), .A2(n4216), .ZN(n3769) );
  OAI21_X1 U4722 ( .B1(n3767), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3776), 
        .ZN(n6187) );
  NAND2_X1 U4723 ( .A1(n6187), .A2(n3739), .ZN(n3768) );
  NAND2_X1 U4724 ( .A1(n3769), .A2(n3768), .ZN(n3770) );
  AOI21_X1 U4725 ( .B1(n3771), .B2(n3894), .A(n3770), .ZN(n4811) );
  NAND2_X1 U4726 ( .A1(n3772), .A2(n3894), .ZN(n3775) );
  XNOR2_X1 U4727 ( .A(n3776), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5273) );
  OAI22_X1 U4728 ( .A1(n5273), .A2(n4216), .B1(n4072), .B2(n5276), .ZN(n3773)
         );
  AOI21_X1 U4729 ( .B1(n4221), .B2(EAX_REG_5__SCAN_IN), .A(n3773), .ZN(n3774)
         );
  NAND2_X1 U4730 ( .A1(n3775), .A2(n3774), .ZN(n4818) );
  NAND2_X1 U4731 ( .A1(n4812), .A2(n4818), .ZN(n4816) );
  INV_X1 U4732 ( .A(n4816), .ZN(n3784) );
  OR2_X1 U4733 ( .A1(n3777), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3778) );
  NAND2_X1 U4734 ( .A1(n3799), .A2(n3778), .ZN(n6178) );
  INV_X1 U4735 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5025) );
  INV_X1 U4736 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3779) );
  OAI22_X1 U4737 ( .A1(n4076), .A2(n5025), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3779), .ZN(n3780) );
  MUX2_X1 U4738 ( .A(n6178), .B(n3780), .S(n4216), .Z(n3781) );
  NAND2_X1 U4739 ( .A1(n3784), .A2(n3783), .ZN(n5021) );
  INV_X1 U4740 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5118) );
  XNOR2_X1 U4741 ( .A(n3799), .B(n5291), .ZN(n5290) );
  NAND2_X1 U4742 ( .A1(n5290), .A2(n4158), .ZN(n3786) );
  NAND2_X1 U4743 ( .A1(n3747), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3785)
         );
  OAI211_X1 U4744 ( .C1(n4076), .C2(n5118), .A(n3786), .B(n3785), .ZN(n3787)
         );
  AOI22_X1 U4745 ( .A1(n4200), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4746 ( .A1(n4029), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4747 ( .A1(n4062), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4748 ( .A1(n4128), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4749 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3798)
         );
  AOI22_X1 U4750 ( .A1(n4123), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4751 ( .A1(n3101), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4752 ( .A1(n3115), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4753 ( .A1(n3135), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3793) );
  NAND4_X1 U4754 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n3797)
         );
  NOR2_X1 U4755 ( .A1(n3798), .A2(n3797), .ZN(n3801) );
  AOI21_X1 U4756 ( .B1(n3800), .B2(n6782), .A(n3818), .ZN(n5313) );
  OAI22_X1 U4757 ( .A1(n3911), .A2(n3801), .B1(n5313), .B2(n4216), .ZN(n3803)
         );
  INV_X1 U4758 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5135) );
  OAI22_X1 U4759 ( .A1(n4076), .A2(n5135), .B1(n4072), .B2(n6782), .ZN(n3802)
         );
  AOI22_X1 U4760 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n4029), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4761 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n3113), .B1(n3117), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4762 ( .A1(n4753), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4763 ( .A1(n3101), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4764 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3813)
         );
  AOI22_X1 U4765 ( .A1(n3302), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4766 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n4128), .B1(n4198), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4767 ( .A1(n3351), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4768 ( .A1(n4062), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4769 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812)
         );
  OAI21_X1 U4770 ( .B1(n3813), .B2(n3812), .A(n3894), .ZN(n3817) );
  INV_X1 U4771 ( .A(n4216), .ZN(n4158) );
  XOR2_X1 U4772 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3818), .Z(n6055) );
  INV_X1 U4773 ( .A(n6055), .ZN(n3814) );
  AOI22_X1 U4774 ( .A1(n3747), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n4158), 
        .B2(n3814), .ZN(n3816) );
  NAND2_X1 U4775 ( .A1(n4221), .A2(EAX_REG_9__SCAN_IN), .ZN(n3815) );
  XNOR2_X1 U4776 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3833), .ZN(n5362)
         );
  OAI22_X1 U4777 ( .A1(n4216), .A2(n5362), .B1(n4072), .B2(n5360), .ZN(n3819)
         );
  AOI21_X1 U4778 ( .B1(n4221), .B2(EAX_REG_10__SCAN_IN), .A(n3819), .ZN(n3831)
         );
  AOI22_X1 U4779 ( .A1(n4200), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4780 ( .A1(n4029), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4781 ( .A1(n4062), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4782 ( .A1(n4142), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4783 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4784 ( .A1(n3101), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4785 ( .A1(n4198), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4786 ( .A1(n3115), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4787 ( .A1(n4128), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4788 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  OAI21_X1 U4789 ( .B1(n3829), .B2(n3828), .A(n3894), .ZN(n3830) );
  XOR2_X1 U4790 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3847), .Z(n6167) );
  AOI22_X1 U4791 ( .A1(n4029), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4792 ( .A1(n4062), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4793 ( .A1(n4123), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4794 ( .A1(n3113), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4795 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3843)
         );
  AOI22_X1 U4796 ( .A1(n3101), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4797 ( .A1(n4753), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4798 ( .A1(n3117), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4799 ( .A1(n3302), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4800 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3842)
         );
  OR2_X1 U4801 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  AOI22_X1 U4802 ( .A1(n3894), .A2(n3844), .B1(n3747), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3846) );
  NAND2_X1 U4803 ( .A1(n4221), .A2(EAX_REG_11__SCAN_IN), .ZN(n3845) );
  OAI211_X1 U4804 ( .C1(n6167), .C2(n4216), .A(n3846), .B(n3845), .ZN(n5345)
         );
  XNOR2_X1 U4805 ( .A(n3862), .B(n5405), .ZN(n5403) );
  NAND2_X1 U4806 ( .A1(n5403), .A2(n4158), .ZN(n3861) );
  INV_X1 U4807 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5383) );
  OAI22_X1 U4808 ( .A1(n4076), .A2(n5383), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5405), .ZN(n3859) );
  AOI22_X1 U4809 ( .A1(n3123), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4810 ( .A1(n4029), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4811 ( .A1(n4128), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4812 ( .A1(n3117), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3848) );
  NAND4_X1 U4813 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3857)
         );
  AOI22_X1 U4814 ( .A1(n4123), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4815 ( .A1(n4200), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4816 ( .A1(n4062), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4817 ( .A1(n4142), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3852) );
  NAND4_X1 U4818 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3856)
         );
  OR2_X1 U4819 ( .A1(n3857), .A2(n3856), .ZN(n3858) );
  AOI22_X1 U4820 ( .A1(n3859), .A2(n4216), .B1(n3894), .B2(n3858), .ZN(n3860)
         );
  INV_X1 U4821 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3865) );
  OAI21_X1 U4822 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3863), .A(n3897), 
        .ZN(n6040) );
  NAND2_X1 U4823 ( .A1(n6040), .A2(n4158), .ZN(n3864) );
  OAI21_X1 U4824 ( .B1(n3865), .B2(n4072), .A(n3864), .ZN(n3866) );
  AOI21_X1 U4825 ( .B1(n4221), .B2(EAX_REG_13__SCAN_IN), .A(n3866), .ZN(n3868)
         );
  INV_X1 U4826 ( .A(n3868), .ZN(n3869) );
  AOI22_X1 U4827 ( .A1(n4029), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4828 ( .A1(n3101), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4829 ( .A1(n4062), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4830 ( .A1(n3113), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3871) );
  NAND4_X1 U4831 ( .A1(n3874), .A2(n3873), .A3(n3872), .A4(n3871), .ZN(n3880)
         );
  AOI22_X1 U4832 ( .A1(n4123), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4833 ( .A1(n4128), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4834 ( .A1(n3351), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4835 ( .A1(n3123), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3875) );
  NAND4_X1 U4836 ( .A1(n3878), .A2(n3877), .A3(n3876), .A4(n3875), .ZN(n3879)
         );
  OR2_X1 U4837 ( .A1(n3880), .A2(n3879), .ZN(n3881) );
  NAND2_X1 U4838 ( .A1(n3894), .A2(n3881), .ZN(n5430) );
  NAND2_X1 U4839 ( .A1(n5428), .A2(n3882), .ZN(n5451) );
  XOR2_X1 U4840 ( .A(n6020), .B(n3897), .Z(n6022) );
  AOI22_X1 U4841 ( .A1(n4029), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4842 ( .A1(n4062), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4843 ( .A1(n4200), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4844 ( .A1(n4753), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3883) );
  NAND4_X1 U4845 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3892)
         );
  AOI22_X1 U4846 ( .A1(n3302), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4847 ( .A1(n4128), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4848 ( .A1(n4123), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4849 ( .A1(n3113), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4850 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3891)
         );
  OR2_X1 U4851 ( .A1(n3892), .A2(n3891), .ZN(n3893) );
  AOI22_X1 U4852 ( .A1(n3894), .A2(n3893), .B1(n3747), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3896) );
  NAND2_X1 U4853 ( .A1(n4221), .A2(EAX_REG_14__SCAN_IN), .ZN(n3895) );
  OAI211_X1 U4854 ( .C1(n6022), .C2(n4216), .A(n3896), .B(n3895), .ZN(n5454)
         );
  NAND2_X1 U4855 ( .A1(n5451), .A2(n5454), .ZN(n5452) );
  XNOR2_X1 U4856 ( .A(n3913), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6006)
         );
  AOI22_X1 U4857 ( .A1(n4200), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4858 ( .A1(n3101), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4859 ( .A1(n4062), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4860 ( .A1(n4142), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3898) );
  NAND4_X1 U4861 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3907)
         );
  AOI22_X1 U4862 ( .A1(n4029), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4863 ( .A1(n4753), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4864 ( .A1(n4128), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4865 ( .A1(n3113), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4866 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3906)
         );
  NOR2_X1 U4867 ( .A1(n3907), .A2(n3906), .ZN(n3910) );
  NAND2_X1 U4868 ( .A1(n4221), .A2(EAX_REG_15__SCAN_IN), .ZN(n3909) );
  NAND2_X1 U4869 ( .A1(n3747), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3908)
         );
  OAI211_X1 U4870 ( .C1(n3911), .C2(n3910), .A(n3909), .B(n3908), .ZN(n3912)
         );
  AOI21_X1 U4871 ( .B1(n6006), .B2(n4158), .A(n3912), .ZN(n5585) );
  XOR2_X1 U4872 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3926), .Z(n5689) );
  AOI22_X1 U4873 ( .A1(n4221), .A2(EAX_REG_16__SCAN_IN), .B1(n3747), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4874 ( .A1(n4128), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4875 ( .A1(n3123), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4876 ( .A1(n3113), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4877 ( .A1(n4029), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4878 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3923)
         );
  AOI22_X1 U4879 ( .A1(n4200), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4880 ( .A1(n4123), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4881 ( .A1(n3101), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4882 ( .A1(n4062), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3918) );
  NAND4_X1 U4883 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n3922)
         );
  OAI21_X1 U4884 ( .B1(n3923), .B2(n3922), .A(n4214), .ZN(n3924) );
  OAI211_X1 U4885 ( .C1(n5689), .C2(n4216), .A(n3925), .B(n3924), .ZN(n5547)
         );
  XNOR2_X1 U4886 ( .A(n3956), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6000)
         );
  NAND2_X1 U4887 ( .A1(n6000), .A2(n4158), .ZN(n3941) );
  AOI22_X1 U4888 ( .A1(n3302), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4889 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n4142), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4890 ( .A1(n4200), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4891 ( .A1(n4029), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3927) );
  NAND4_X1 U4892 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3936)
         );
  AOI22_X1 U4893 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n4128), .B1(n4062), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4894 ( .A1(n3101), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4895 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n3117), .B1(n3135), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4896 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n3113), .B1(n3483), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3931) );
  NAND4_X1 U4897 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3935)
         );
  NOR2_X1 U4898 ( .A1(n3936), .A2(n3935), .ZN(n3939) );
  AOI21_X1 U4899 ( .B1(n5998), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3937) );
  AOI21_X1 U4900 ( .B1(n4221), .B2(EAX_REG_17__SCAN_IN), .A(n3937), .ZN(n3938)
         );
  OAI21_X1 U4901 ( .B1(n4180), .B2(n3939), .A(n3938), .ZN(n3940) );
  NAND2_X1 U4902 ( .A1(n3941), .A2(n3940), .ZN(n5918) );
  AOI22_X1 U4903 ( .A1(n4029), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4904 ( .A1(n4142), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4905 ( .A1(n4128), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4906 ( .A1(n4062), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4907 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3951)
         );
  AOI22_X1 U4908 ( .A1(n3101), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4909 ( .A1(n3113), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4910 ( .A1(n4753), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4911 ( .A1(n3123), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3946) );
  NAND4_X1 U4912 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3950)
         );
  NOR2_X1 U4913 ( .A1(n3951), .A2(n3950), .ZN(n3955) );
  OAI21_X1 U4914 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6703), .A(n6695), 
        .ZN(n3952) );
  INV_X1 U4915 ( .A(n3952), .ZN(n3953) );
  AOI21_X1 U4916 ( .B1(n4221), .B2(EAX_REG_18__SCAN_IN), .A(n3953), .ZN(n3954)
         );
  OAI21_X1 U4917 ( .B1(n4180), .B2(n3955), .A(n3954), .ZN(n3959) );
  OAI21_X1 U4918 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3957), .A(n3989), 
        .ZN(n5996) );
  OR2_X1 U4919 ( .A1(n4216), .A2(n5996), .ZN(n3958) );
  NAND2_X1 U4920 ( .A1(n3959), .A2(n3958), .ZN(n5580) );
  AOI22_X1 U4921 ( .A1(n3123), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4922 ( .A1(n4123), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4923 ( .A1(n3351), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4924 ( .A1(n4029), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U4925 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3969)
         );
  AOI22_X1 U4926 ( .A1(n4062), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4927 ( .A1(n3101), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4928 ( .A1(n3117), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4929 ( .A1(n3113), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3964) );
  NAND4_X1 U4930 ( .A1(n3967), .A2(n3966), .A3(n3965), .A4(n3964), .ZN(n3968)
         );
  NOR2_X1 U4931 ( .A1(n3969), .A2(n3968), .ZN(n3972) );
  AOI21_X1 U4932 ( .B1(n5680), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3970) );
  AOI21_X1 U4933 ( .B1(n4221), .B2(EAX_REG_19__SCAN_IN), .A(n3970), .ZN(n3971)
         );
  OAI21_X1 U4934 ( .B1(n4180), .B2(n3972), .A(n3971), .ZN(n3974) );
  XNOR2_X1 U4935 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3989), .ZN(n5678)
         );
  NAND2_X1 U4936 ( .A1(n4158), .A2(n5678), .ZN(n3973) );
  NAND2_X1 U4937 ( .A1(n3974), .A2(n3973), .ZN(n5532) );
  AOI22_X1 U4938 ( .A1(n3302), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4939 ( .A1(n4128), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4940 ( .A1(n4200), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4941 ( .A1(n3135), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4942 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3984)
         );
  AOI22_X1 U4943 ( .A1(n4029), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4944 ( .A1(n3101), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4945 ( .A1(n4198), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4946 ( .A1(n4062), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U4947 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3983)
         );
  NOR2_X1 U4948 ( .A1(n3984), .A2(n3983), .ZN(n3988) );
  OAI21_X1 U4949 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6703), .A(n6695), 
        .ZN(n3985) );
  INV_X1 U4950 ( .A(n3985), .ZN(n3986) );
  AOI21_X1 U4951 ( .B1(n4221), .B2(EAX_REG_20__SCAN_IN), .A(n3986), .ZN(n3987)
         );
  OAI21_X1 U4952 ( .B1(n4180), .B2(n3988), .A(n3987), .ZN(n3992) );
  OAI21_X1 U4953 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n3990), .A(n4024), 
        .ZN(n5896) );
  OR2_X1 U4954 ( .A1(n4216), .A2(n5896), .ZN(n3991) );
  AOI22_X1 U4955 ( .A1(n4029), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4956 ( .A1(n3101), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4957 ( .A1(n3351), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4958 ( .A1(n3113), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4959 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4002)
         );
  AOI22_X1 U4960 ( .A1(n4062), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4961 ( .A1(n4142), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4962 ( .A1(n4753), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4963 ( .A1(n3116), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U4964 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4001)
         );
  NOR2_X1 U4965 ( .A1(n4002), .A2(n4001), .ZN(n4006) );
  NAND2_X1 U4966 ( .A1(n6695), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4003)
         );
  NAND2_X1 U4967 ( .A1(n4216), .A2(n4003), .ZN(n4004) );
  AOI21_X1 U4968 ( .B1(n4221), .B2(EAX_REG_21__SCAN_IN), .A(n4004), .ZN(n4005)
         );
  OAI21_X1 U4969 ( .B1(n4180), .B2(n4006), .A(n4005), .ZN(n4008) );
  XNOR2_X1 U4970 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4024), .ZN(n5667)
         );
  NAND2_X1 U4971 ( .A1(n4158), .A2(n5667), .ZN(n4007) );
  AOI22_X1 U4972 ( .A1(n3302), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4973 ( .A1(n4142), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4974 ( .A1(n4200), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4975 ( .A1(n3315), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4976 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4019)
         );
  AOI22_X1 U4977 ( .A1(n3101), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4978 ( .A1(n4128), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4979 ( .A1(n4198), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4980 ( .A1(n4201), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U4981 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4018)
         );
  NOR2_X1 U4982 ( .A1(n4019), .A2(n4018), .ZN(n4023) );
  NAND2_X1 U4983 ( .A1(n6695), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4020)
         );
  NAND2_X1 U4984 ( .A1(n4216), .A2(n4020), .ZN(n4021) );
  AOI21_X1 U4985 ( .B1(n4221), .B2(EAX_REG_22__SCAN_IN), .A(n4021), .ZN(n4022)
         );
  OAI21_X1 U4986 ( .B1(n4180), .B2(n4023), .A(n4022), .ZN(n4028) );
  OAI21_X1 U4987 ( .B1(n4026), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n4070), 
        .ZN(n5888) );
  OR2_X1 U4988 ( .A1(n5888), .A2(n4216), .ZN(n4027) );
  AOI22_X1 U4989 ( .A1(n3123), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4990 ( .A1(n3314), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4991 ( .A1(n4200), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4992 ( .A1(n4029), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U4993 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4039)
         );
  AOI22_X1 U4994 ( .A1(n4062), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4995 ( .A1(n3101), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4996 ( .A1(n3117), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4997 ( .A1(n3113), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4034) );
  NAND4_X1 U4998 ( .A1(n4037), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(n4038)
         );
  NOR2_X1 U4999 ( .A1(n4039), .A2(n4038), .ZN(n4057) );
  AOI22_X1 U5000 ( .A1(n3101), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5001 ( .A1(n4128), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5002 ( .A1(n4753), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5003 ( .A1(n4062), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4040) );
  NAND4_X1 U5004 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4049)
         );
  AOI22_X1 U5005 ( .A1(n4029), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5006 ( .A1(n4142), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5007 ( .A1(n4200), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5008 ( .A1(n3113), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4044) );
  NAND4_X1 U5009 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4048)
         );
  NOR2_X1 U5010 ( .A1(n4049), .A2(n4048), .ZN(n4056) );
  XOR2_X1 U5011 ( .A(n4057), .B(n4056), .Z(n4050) );
  NAND2_X1 U5012 ( .A1(n4050), .A2(n4214), .ZN(n4053) );
  INV_X1 U5013 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5880) );
  AOI21_X1 U5014 ( .B1(n5880), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4051) );
  AOI21_X1 U5015 ( .B1(n4221), .B2(EAX_REG_23__SCAN_IN), .A(n4051), .ZN(n4052)
         );
  NAND2_X1 U5016 ( .A1(n4053), .A2(n4052), .ZN(n4055) );
  XNOR2_X1 U5017 ( .A(n4070), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5869)
         );
  NAND2_X1 U5018 ( .A1(n5869), .A2(n4158), .ZN(n4054) );
  NAND2_X1 U5019 ( .A1(n4055), .A2(n4054), .ZN(n4475) );
  NOR2_X1 U5020 ( .A1(n4057), .A2(n4056), .ZN(n4113) );
  AOI22_X1 U5021 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n4753), .B1(n3302), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5022 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4142), .B1(n4123), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5023 ( .A1(n3351), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5024 ( .A1(n4029), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U5025 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4068)
         );
  AOI22_X1 U5026 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n4062), .B1(n4128), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5027 ( .A1(n3101), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5028 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n3117), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5029 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n3113), .B1(n3483), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U5030 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4067)
         );
  INV_X1 U5031 ( .A(n4112), .ZN(n4069) );
  XNOR2_X1 U5032 ( .A(n4113), .B(n4069), .ZN(n4078) );
  INV_X1 U5033 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4075) );
  INV_X1 U5034 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5505) );
  XNOR2_X1 U5035 ( .A(n4093), .B(n5505), .ZN(n5650) );
  NOR2_X1 U5036 ( .A1(n4072), .A2(n5505), .ZN(n4073) );
  AOI21_X1 U5037 ( .B1(n5650), .B2(n4158), .A(n4073), .ZN(n4074) );
  OAI21_X1 U5038 ( .B1(n4076), .B2(n4075), .A(n4074), .ZN(n4077) );
  AOI21_X1 U5039 ( .B1(n4078), .B2(n4214), .A(n4077), .ZN(n5504) );
  AOI22_X1 U5040 ( .A1(n3122), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5041 ( .A1(n4123), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5042 ( .A1(n4200), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5043 ( .A1(n4029), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4079) );
  NAND4_X1 U5044 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4088)
         );
  AOI22_X1 U5045 ( .A1(n4062), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5046 ( .A1(n3101), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5047 ( .A1(n3117), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5048 ( .A1(n3113), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4083) );
  NAND4_X1 U5049 ( .A1(n4086), .A2(n4085), .A3(n4084), .A4(n4083), .ZN(n4087)
         );
  OR2_X1 U5050 ( .A1(n4088), .A2(n4087), .ZN(n4111) );
  NAND2_X1 U5051 ( .A1(n4112), .A2(n4113), .ZN(n4089) );
  XNOR2_X1 U5052 ( .A(n4111), .B(n4089), .ZN(n4090) );
  NAND2_X1 U5053 ( .A1(n4214), .A2(n4090), .ZN(n4100) );
  NAND2_X1 U5054 ( .A1(n6695), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4091)
         );
  NAND2_X1 U5055 ( .A1(n4216), .A2(n4091), .ZN(n4092) );
  AOI21_X1 U5056 ( .B1(n4221), .B2(EAX_REG_25__SCAN_IN), .A(n4092), .ZN(n4099)
         );
  INV_X1 U5057 ( .A(n4093), .ZN(n4094) );
  INV_X1 U5058 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4095) );
  NAND2_X1 U5059 ( .A1(n4096), .A2(n4095), .ZN(n4097) );
  NAND2_X1 U5060 ( .A1(n4119), .A2(n4097), .ZN(n5639) );
  NOR2_X1 U5061 ( .A1(n5639), .A2(n4216), .ZN(n4098) );
  AOI21_X1 U5062 ( .B1(n4100), .B2(n4099), .A(n4098), .ZN(n4532) );
  AOI22_X1 U5063 ( .A1(n3122), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5064 ( .A1(n4753), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5065 ( .A1(n3101), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5066 ( .A1(n4029), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U5067 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4110)
         );
  AOI22_X1 U5068 ( .A1(n4128), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5069 ( .A1(n4062), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5070 ( .A1(n3113), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5071 ( .A1(n4200), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4105) );
  NAND4_X1 U5072 ( .A1(n4108), .A2(n4107), .A3(n4106), .A4(n4105), .ZN(n4109)
         );
  NOR2_X1 U5073 ( .A1(n4110), .A2(n4109), .ZN(n4136) );
  NAND3_X1 U5074 ( .A1(n4113), .A2(n4112), .A3(n4111), .ZN(n4137) );
  XNOR2_X1 U5075 ( .A(n4136), .B(n4137), .ZN(n4116) );
  INV_X1 U5076 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6910) );
  OAI21_X1 U5077 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6910), .A(n4216), .ZN(
        n4114) );
  AOI21_X1 U5078 ( .B1(n4221), .B2(EAX_REG_26__SCAN_IN), .A(n4114), .ZN(n4115)
         );
  OAI21_X1 U5079 ( .B1(n4180), .B2(n4116), .A(n4115), .ZN(n4118) );
  XNOR2_X1 U5080 ( .A(n4119), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5627)
         );
  NAND2_X1 U5081 ( .A1(n5627), .A2(n4158), .ZN(n4117) );
  INV_X1 U5082 ( .A(n4119), .ZN(n4120) );
  NAND2_X1 U5083 ( .A1(n4120), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4121)
         );
  INV_X1 U5084 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U5085 ( .A1(n4121), .A2(n5486), .ZN(n4122) );
  NAND2_X1 U5086 ( .A1(n4161), .A2(n4122), .ZN(n5619) );
  AOI22_X1 U5087 ( .A1(n3123), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5088 ( .A1(n4029), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5089 ( .A1(n4200), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5090 ( .A1(n4062), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4124) );
  NAND4_X1 U5091 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4135)
         );
  AOI22_X1 U5092 ( .A1(n3101), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5093 ( .A1(n4128), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5094 ( .A1(n4142), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5095 ( .A1(n3113), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4130) );
  NAND4_X1 U5096 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4134)
         );
  NOR2_X1 U5097 ( .A1(n4135), .A2(n4134), .ZN(n4154) );
  OR2_X1 U5098 ( .A1(n4137), .A2(n4136), .ZN(n4153) );
  XNOR2_X1 U5099 ( .A(n4154), .B(n4153), .ZN(n4140) );
  AOI21_X1 U5100 ( .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6695), .A(n4158), 
        .ZN(n4139) );
  NAND2_X1 U5101 ( .A1(n4221), .A2(EAX_REG_27__SCAN_IN), .ZN(n4138) );
  OAI211_X1 U5102 ( .C1(n4140), .C2(n4180), .A(n4139), .B(n4138), .ZN(n4141)
         );
  OAI21_X1 U5103 ( .B1(n4216), .B2(n5619), .A(n4141), .ZN(n5481) );
  AOI22_X1 U5104 ( .A1(n3122), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5105 ( .A1(n4123), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5106 ( .A1(n4200), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5107 ( .A1(n4029), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4143) );
  NAND4_X1 U5108 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4152)
         );
  AOI22_X1 U5109 ( .A1(n4062), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5110 ( .A1(n3101), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5111 ( .A1(n3117), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5112 ( .A1(n3113), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U5113 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4151)
         );
  OR2_X1 U5114 ( .A1(n4152), .A2(n4151), .ZN(n4176) );
  NOR2_X1 U5115 ( .A1(n4154), .A2(n4153), .ZN(n4177) );
  XOR2_X1 U5116 ( .A(n4176), .B(n4177), .Z(n4155) );
  NAND2_X1 U5117 ( .A1(n4155), .A2(n4214), .ZN(n4160) );
  INV_X1 U5118 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4156) );
  NOR2_X1 U5119 ( .A1(n4156), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4157) );
  AOI211_X1 U5120 ( .C1(n4221), .C2(EAX_REG_28__SCAN_IN), .A(n4158), .B(n4157), 
        .ZN(n4159) );
  XNOR2_X1 U5121 ( .A(n4161), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5472)
         );
  INV_X1 U5122 ( .A(n4161), .ZN(n4162) );
  NAND2_X1 U5123 ( .A1(n4162), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4164)
         );
  INV_X1 U5124 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U5125 ( .A1(n4164), .A2(n4163), .ZN(n4165) );
  NAND2_X1 U5126 ( .A1(n4226), .A2(n4165), .ZN(n5439) );
  AOI22_X1 U5127 ( .A1(n4200), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5128 ( .A1(n4198), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5129 ( .A1(n4029), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U5130 ( .A1(n4062), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4166) );
  NAND4_X1 U5131 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4175)
         );
  AOI22_X1 U5132 ( .A1(n4123), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5133 ( .A1(n4128), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5134 ( .A1(n4753), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5135 ( .A1(n3101), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4170) );
  NAND4_X1 U5136 ( .A1(n4173), .A2(n4172), .A3(n4171), .A4(n4170), .ZN(n4174)
         );
  NOR2_X1 U5137 ( .A1(n4175), .A2(n4174), .ZN(n4197) );
  NAND2_X1 U5138 ( .A1(n4177), .A2(n4176), .ZN(n4196) );
  XNOR2_X1 U5139 ( .A(n4197), .B(n4196), .ZN(n4181) );
  AOI21_X1 U5140 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6695), .A(n4158), 
        .ZN(n4179) );
  NAND2_X1 U5141 ( .A1(n4221), .A2(EAX_REG_29__SCAN_IN), .ZN(n4178) );
  OAI211_X1 U5142 ( .C1(n4181), .C2(n4180), .A(n4179), .B(n4178), .ZN(n4182)
         );
  OAI21_X1 U5143 ( .B1(n4216), .B2(n5439), .A(n4182), .ZN(n4183) );
  NAND2_X1 U5144 ( .A1(n4235), .A2(n4183), .ZN(n4185) );
  INV_X1 U5145 ( .A(n4399), .ZN(n4184) );
  AND3_X1 U5146 ( .A1(n6952), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n4186) );
  NAND2_X1 U5147 ( .A1(n6527), .A2(n4187), .ZN(n6686) );
  NAND2_X1 U5148 ( .A1(n6686), .A2(n6952), .ZN(n4188) );
  NAND2_X1 U5149 ( .A1(n6952), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4190) );
  NAND2_X1 U5150 ( .A1(n6703), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4189) );
  AND2_X1 U5151 ( .A1(n4190), .A2(n4189), .ZN(n4710) );
  NOR2_X1 U5152 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6591) );
  INV_X1 U5153 ( .A(n6591), .ZN(n4191) );
  INV_X1 U5154 ( .A(REIP_REG_29__SCAN_IN), .ZN(n4494) );
  NOR2_X1 U5155 ( .A1(n6253), .A2(n4494), .ZN(n5732) );
  AOI21_X1 U5156 ( .B1(n6188), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5732), 
        .ZN(n4192) );
  OAI21_X1 U5157 ( .B1(n6195), .B2(n5439), .A(n4192), .ZN(n4193) );
  NOR2_X1 U5158 ( .A1(n4197), .A2(n4196), .ZN(n4213) );
  AOI22_X1 U5159 ( .A1(n3315), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5160 ( .A1(n3101), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U5161 ( .A1(n4200), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U5162 ( .A1(n4201), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4202) );
  NAND4_X1 U5163 ( .A1(n4205), .A2(n4204), .A3(n4203), .A4(n4202), .ZN(n4211)
         );
  AOI22_X1 U5164 ( .A1(n3302), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U5165 ( .A1(n3433), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U5166 ( .A1(n4753), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U5167 ( .A1(n3113), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4206) );
  NAND4_X1 U5168 ( .A1(n4209), .A2(n4208), .A3(n4207), .A4(n4206), .ZN(n4210)
         );
  NOR2_X1 U5169 ( .A1(n4211), .A2(n4210), .ZN(n4212) );
  XNOR2_X1 U5170 ( .A(n4213), .B(n4212), .ZN(n4215) );
  NAND2_X1 U5171 ( .A1(n4215), .A2(n4214), .ZN(n4220) );
  INV_X1 U5172 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6803) );
  OAI21_X1 U5173 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6803), .A(n4216), .ZN(
        n4217) );
  AOI21_X1 U5174 ( .B1(n4221), .B2(EAX_REG_30__SCAN_IN), .A(n4217), .ZN(n4219)
         );
  XNOR2_X1 U5175 ( .A(n4226), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4456)
         );
  AOI22_X1 U5176 ( .A1(n4221), .A2(EAX_REG_31__SCAN_IN), .B1(n3747), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4222) );
  INV_X1 U5177 ( .A(n4222), .ZN(n4223) );
  NAND2_X1 U5178 ( .A1(n5595), .A2(n3103), .ZN(n4233) );
  INV_X1 U5179 ( .A(n5633), .ZN(n4225) );
  NAND2_X1 U5180 ( .A1(n5704), .A2(n6191), .ZN(n4232) );
  INV_X1 U5181 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4227) );
  INV_X1 U5182 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6764) );
  NOR2_X1 U5183 ( .A1(n6253), .A2(n6764), .ZN(n5709) );
  AOI21_X1 U5184 ( .B1(n6188), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5709), 
        .ZN(n4229) );
  OAI21_X1 U5185 ( .B1(n6195), .B2(n4454), .A(n4229), .ZN(n4230) );
  INV_X1 U5186 ( .A(n4230), .ZN(n4231) );
  NAND2_X1 U5187 ( .A1(n4233), .A2(n3248), .ZN(U2955) );
  OAI21_X1 U5188 ( .B1(n4234), .B2(n4236), .A(n4235), .ZN(n5561) );
  INV_X1 U5189 ( .A(n3121), .ZN(n4237) );
  NAND3_X1 U5190 ( .A1(n4238), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n6983), .ZN(n4243) );
  NAND3_X1 U5191 ( .A1(n5615), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n5752), .ZN(n4240) );
  INV_X1 U5192 ( .A(n4404), .ZN(n4239) );
  AOI21_X1 U5193 ( .B1(n5616), .B2(n5706), .A(n4241), .ZN(n4242) );
  INV_X1 U5194 ( .A(n5472), .ZN(n4245) );
  INV_X1 U5195 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6649) );
  NOR2_X1 U5196 ( .A1(n6253), .A2(n6649), .ZN(n5740) );
  AOI21_X1 U5197 ( .B1(n6188), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5740), 
        .ZN(n4244) );
  OAI21_X1 U5198 ( .B1(n6195), .B2(n4245), .A(n4244), .ZN(n4246) );
  INV_X1 U5199 ( .A(n4246), .ZN(n4247) );
  AND2_X1 U5200 ( .A1(n5813), .A2(n4384), .ZN(n4382) );
  NAND2_X1 U5201 ( .A1(n5643), .A2(n4382), .ZN(n4250) );
  XNOR2_X1 U5202 ( .A(n6164), .B(n6935), .ZN(n5669) );
  XNOR2_X1 U5203 ( .A(n6164), .B(n6723), .ZN(n5662) );
  NOR2_X2 U5204 ( .A1(n5661), .A2(n5662), .ZN(n5660) );
  NOR2_X1 U5205 ( .A1(n6164), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5654)
         );
  NAND2_X1 U5206 ( .A1(n5660), .A2(n5654), .ZN(n5644) );
  OAI21_X1 U5207 ( .B1(n4251), .B2(n4250), .A(n5644), .ZN(n4252) );
  XNOR2_X1 U5208 ( .A(n4252), .B(n5778), .ZN(n4472) );
  INV_X1 U5209 ( .A(n4253), .ZN(n4254) );
  NAND2_X1 U5210 ( .A1(n4254), .A2(n6602), .ZN(n6689) );
  NAND2_X1 U5211 ( .A1(n3120), .A2(n6689), .ZN(n4261) );
  NAND2_X1 U5212 ( .A1(n4256), .A2(n4255), .ZN(n4259) );
  INV_X1 U5213 ( .A(n4257), .ZN(n4258) );
  OAI21_X1 U5214 ( .B1(n4260), .B2(n4259), .A(n4258), .ZN(n4551) );
  NOR2_X1 U5215 ( .A1(READY_N), .A2(n4551), .ZN(n4561) );
  NAND2_X1 U5216 ( .A1(n4261), .A2(n4561), .ZN(n4266) );
  NAND2_X1 U5217 ( .A1(n3374), .A2(n6689), .ZN(n4421) );
  NAND2_X1 U5218 ( .A1(n4421), .A2(n6690), .ZN(n4262) );
  OAI211_X1 U5219 ( .C1(n4868), .C2(n4262), .A(n4281), .B(n5435), .ZN(n4263)
         );
  INV_X1 U5220 ( .A(n4263), .ZN(n4264) );
  OR2_X1 U5221 ( .A1(n4589), .A2(n4264), .ZN(n4265) );
  MUX2_X1 U5222 ( .A(n4266), .B(n4265), .S(n3399), .Z(n4277) );
  INV_X1 U5223 ( .A(n4267), .ZN(n4835) );
  NAND2_X1 U5224 ( .A1(n4835), .A2(n3120), .ZN(n4378) );
  INV_X1 U5225 ( .A(n4378), .ZN(n4275) );
  NAND2_X1 U5226 ( .A1(n4268), .A2(n4281), .ZN(n4269) );
  NAND2_X1 U5227 ( .A1(n4867), .A2(n4269), .ZN(n4270) );
  OAI21_X1 U5228 ( .B1(n4271), .B2(n3383), .A(n4270), .ZN(n4369) );
  INV_X1 U5229 ( .A(n4369), .ZN(n4272) );
  NOR2_X1 U5230 ( .A1(n4279), .A2(n4272), .ZN(n4274) );
  NOR2_X1 U5231 ( .A1(n4274), .A2(n4273), .ZN(n4567) );
  AOI21_X1 U5232 ( .B1(n4589), .B2(n4275), .A(n4567), .ZN(n4276) );
  NAND2_X1 U5233 ( .A1(n4277), .A2(n4276), .ZN(n4278) );
  OR2_X1 U5234 ( .A1(n4279), .A2(n3671), .ZN(n4743) );
  AND2_X1 U5235 ( .A1(n4859), .A2(n4743), .ZN(n4550) );
  INV_X1 U5236 ( .A(n4868), .ZN(n4563) );
  AOI22_X1 U5237 ( .A1(n4280), .A2(n3381), .B1(n4563), .B2(n4564), .ZN(n4283)
         );
  AND3_X1 U5238 ( .A1(n4550), .A2(n4283), .A3(n4282), .ZN(n4284) );
  NAND2_X1 U5239 ( .A1(n4472), .A2(n6269), .ZN(n4397) );
  NAND2_X1 U5240 ( .A1(n4563), .A2(n3406), .ZN(n4609) );
  NAND2_X1 U5241 ( .A1(n4280), .A2(n3382), .ZN(n4285) );
  AND2_X1 U5242 ( .A1(n4609), .A2(n4285), .ZN(n4286) );
  NAND2_X1 U5243 ( .A1(n4287), .A2(n4281), .ZN(n4303) );
  AOI22_X1 U5244 ( .A1(n4304), .A2(EBX_REG_19__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n4676), .ZN(n4290) );
  NAND2_X2 U5245 ( .A1(n3531), .A2(n3120), .ZN(n4297) );
  INV_X1 U5246 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4288) );
  NAND2_X1 U5247 ( .A1(n4441), .A2(n4288), .ZN(n4289) );
  NAND2_X1 U5248 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4291) );
  OAI211_X1 U5249 ( .C1(n4676), .C2(EBX_REG_13__SCAN_IN), .A(n4438), .B(n4291), 
        .ZN(n4292) );
  OAI21_X1 U5250 ( .B1(n4430), .B2(EBX_REG_13__SCAN_IN), .A(n4292), .ZN(n5949)
         );
  INV_X1 U5251 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U5252 ( .A1(n4564), .A2(n6732), .ZN(n4293) );
  OAI211_X1 U5253 ( .C1(n5808), .C2(n6967), .A(n4438), .B(n4293), .ZN(n4294)
         );
  OAI21_X1 U5254 ( .B1(n4430), .B2(EBX_REG_9__SCAN_IN), .A(n4294), .ZN(n6052)
         );
  NAND2_X1 U5255 ( .A1(n4303), .A2(EBX_REG_0__SCAN_IN), .ZN(n4296) );
  INV_X1 U5256 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U5257 ( .A1(n4297), .A2(n6929), .ZN(n4295) );
  AND2_X1 U5258 ( .A1(n4296), .A2(n4295), .ZN(n4599) );
  INV_X1 U5259 ( .A(n4599), .ZN(n4300) );
  INV_X1 U5260 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U5261 ( .A1(n4303), .A2(n6795), .ZN(n4298) );
  OAI211_X1 U5262 ( .C1(n4317), .C2(EBX_REG_1__SCAN_IN), .A(n4298), .B(n4297), 
        .ZN(n4299) );
  INV_X1 U5263 ( .A(n4301), .ZN(n4302) );
  INV_X1 U5264 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U5265 ( .A1(n4441), .A2(n6081), .ZN(n4308) );
  INV_X1 U5266 ( .A(n4303), .ZN(n4304) );
  NAND2_X1 U5267 ( .A1(n4438), .A2(n4305), .ZN(n4306) );
  OAI211_X1 U5268 ( .C1(n4676), .C2(EBX_REG_2__SCAN_IN), .A(n4306), .B(n4297), 
        .ZN(n4307) );
  NAND2_X1 U5269 ( .A1(n4308), .A2(n4307), .ZN(n4737) );
  NAND2_X1 U5270 ( .A1(n4738), .A2(n4737), .ZN(n4805) );
  OR2_X1 U5271 ( .A1(n4597), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4312)
         );
  NAND2_X1 U5272 ( .A1(n5808), .A2(EBX_REG_3__SCAN_IN), .ZN(n4311) );
  INV_X1 U5273 ( .A(n4430), .ZN(n4483) );
  INV_X1 U5274 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4309) );
  NAND2_X1 U5275 ( .A1(n4483), .A2(n4309), .ZN(n4310) );
  NAND3_X1 U5276 ( .A1(n4312), .A2(n4311), .A3(n4310), .ZN(n4806) );
  OR2_X1 U5277 ( .A1(n4564), .A2(n4438), .ZN(n4345) );
  INV_X1 U5278 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U5279 ( .A1(n4441), .A2(n4313), .ZN(n4316) );
  OR2_X1 U5280 ( .A1(n4438), .A2(n4313), .ZN(n4315) );
  NAND2_X1 U5281 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n4676), .ZN(n4314)
         );
  NAND4_X1 U5282 ( .A1(n4345), .A2(n4316), .A3(n4315), .A4(n4314), .ZN(n4882)
         );
  NAND2_X1 U5283 ( .A1(n4881), .A2(n4882), .ZN(n4880) );
  NAND2_X1 U5284 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4318)
         );
  OAI211_X1 U5285 ( .C1(n4676), .C2(EBX_REG_5__SCAN_IN), .A(n4438), .B(n4318), 
        .ZN(n4319) );
  OAI21_X1 U5286 ( .B1(n4430), .B2(EBX_REG_5__SCAN_IN), .A(n4319), .ZN(n4820)
         );
  NOR2_X2 U5287 ( .A1(n4880), .A2(n4820), .ZN(n4819) );
  INV_X1 U5288 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U5289 ( .A1(n4441), .A2(n5071), .ZN(n4322) );
  OR2_X1 U5290 ( .A1(n4438), .A2(n5071), .ZN(n4321) );
  NAND2_X1 U5291 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4676), .ZN(n4320)
         );
  NAND4_X1 U5292 ( .A1(n4345), .A2(n4322), .A3(n4321), .A4(n4320), .ZN(n4526)
         );
  NAND2_X1 U5293 ( .A1(n4819), .A2(n4526), .ZN(n4525) );
  INV_X1 U5294 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6932) );
  NAND2_X1 U5295 ( .A1(n4564), .A2(n6932), .ZN(n4323) );
  OAI211_X1 U5296 ( .C1(n5808), .C2(n6913), .A(n4438), .B(n4323), .ZN(n4324)
         );
  OAI21_X1 U5297 ( .B1(n4430), .B2(EBX_REG_7__SCAN_IN), .A(n4324), .ZN(n5073)
         );
  INV_X1 U5298 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4325) );
  NAND2_X1 U5299 ( .A1(n4441), .A2(n4325), .ZN(n4328) );
  NAND2_X1 U5300 ( .A1(n4438), .A2(n6229), .ZN(n4326) );
  OAI211_X1 U5301 ( .C1(n4676), .C2(EBX_REG_8__SCAN_IN), .A(n4326), .B(n4297), 
        .ZN(n4327) );
  NAND2_X1 U5302 ( .A1(n4328), .A2(n4327), .ZN(n5124) );
  INV_X1 U5303 ( .A(n4441), .ZN(n4364) );
  INV_X1 U5304 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U5305 ( .A1(n4564), .A2(n6797), .ZN(n4329) );
  OAI211_X1 U5306 ( .C1(n4304), .C2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n4329), .B(n4297), .ZN(n4330) );
  OAI21_X1 U5307 ( .B1(n4364), .B2(EBX_REG_10__SCAN_IN), .A(n4330), .ZN(n5303)
         );
  NAND2_X1 U5308 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4331) );
  OAI211_X1 U5309 ( .C1(n4676), .C2(EBX_REG_11__SCAN_IN), .A(n4438), .B(n4331), 
        .ZN(n4332) );
  OAI21_X1 U5310 ( .B1(n4430), .B2(EBX_REG_11__SCAN_IN), .A(n4332), .ZN(n6042)
         );
  INV_X1 U5311 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U5312 ( .A1(n4441), .A2(n5376), .ZN(n4335) );
  NAND2_X1 U5313 ( .A1(n4438), .A2(n4380), .ZN(n4333) );
  OAI211_X1 U5314 ( .C1(n4676), .C2(EBX_REG_12__SCAN_IN), .A(n4333), .B(n4297), 
        .ZN(n4334) );
  NAND2_X1 U5315 ( .A1(n4335), .A2(n4334), .ZN(n5369) );
  NAND2_X1 U5316 ( .A1(n5368), .A2(n5369), .ZN(n5948) );
  NOR2_X2 U5317 ( .A1(n5949), .A2(n5948), .ZN(n5947) );
  INV_X1 U5318 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U5319 ( .A1(n4441), .A2(n5590), .ZN(n4338) );
  OR2_X1 U5320 ( .A1(n4438), .A2(n5590), .ZN(n4337) );
  NAND2_X1 U5321 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4676), .ZN(n4336) );
  NAND4_X1 U5322 ( .A1(n4345), .A2(n4338), .A3(n4337), .A4(n4336), .ZN(n5423)
         );
  NAND2_X1 U5323 ( .A1(n5947), .A2(n5423), .ZN(n5586) );
  NOR2_X1 U5324 ( .A1(n4430), .A2(EBX_REG_15__SCAN_IN), .ZN(n4339) );
  AOI21_X1 U5325 ( .B1(n5808), .B2(EBX_REG_15__SCAN_IN), .A(n4339), .ZN(n4340)
         );
  OAI21_X1 U5326 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4597), .A(n4340), 
        .ZN(n5587) );
  INV_X1 U5327 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4341) );
  NAND2_X1 U5328 ( .A1(n4441), .A2(n4341), .ZN(n4344) );
  OR2_X1 U5329 ( .A1(n4438), .A2(n4341), .ZN(n4343) );
  NAND2_X1 U5330 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4676), .ZN(n4342) );
  NAND4_X1 U5331 ( .A1(n4345), .A2(n4344), .A3(n4343), .A4(n4342), .ZN(n5549)
         );
  NAND2_X1 U5332 ( .A1(n5548), .A2(n5549), .ZN(n5929) );
  NAND2_X1 U5333 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4346) );
  OAI211_X1 U5334 ( .C1(n4676), .C2(EBX_REG_17__SCAN_IN), .A(n4438), .B(n4346), 
        .ZN(n4347) );
  OAI21_X1 U5335 ( .B1(n4430), .B2(EBX_REG_17__SCAN_IN), .A(n4347), .ZN(n5928)
         );
  INV_X1 U5336 ( .A(n4348), .ZN(n5927) );
  NAND2_X1 U5337 ( .A1(n4597), .A2(EBX_REG_20__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U5338 ( .A1(n4676), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4349) );
  NAND2_X1 U5339 ( .A1(n4350), .A2(n4349), .ZN(n5810) );
  NOR2_X1 U5340 ( .A1(n5810), .A2(n4297), .ZN(n4354) );
  AND2_X1 U5341 ( .A1(n5810), .A2(n4297), .ZN(n4353) );
  NAND2_X1 U5342 ( .A1(n4597), .A2(EBX_REG_18__SCAN_IN), .ZN(n4352) );
  NAND2_X1 U5343 ( .A1(n4676), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U5344 ( .A1(n4352), .A2(n4351), .ZN(n5805) );
  MUX2_X1 U5345 ( .A(n4354), .B(n4353), .S(n5805), .Z(n4355) );
  INV_X1 U5346 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U5347 ( .A1(n4441), .A2(n6800), .ZN(n4359) );
  NAND2_X1 U5348 ( .A1(n4438), .A2(n6723), .ZN(n4357) );
  NAND2_X1 U5349 ( .A1(n4564), .A2(n6800), .ZN(n4356) );
  NAND3_X1 U5350 ( .A1(n4357), .A2(n4297), .A3(n4356), .ZN(n4358) );
  NAND2_X1 U5351 ( .A1(n4359), .A2(n4358), .ZN(n5519) );
  OR2_X1 U5352 ( .A1(n4597), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4361)
         );
  NAND2_X1 U5353 ( .A1(n5808), .A2(EBX_REG_22__SCAN_IN), .ZN(n4360) );
  OAI211_X1 U5354 ( .C1(n4430), .C2(EBX_REG_22__SCAN_IN), .A(n4361), .B(n4360), 
        .ZN(n5571) );
  NAND2_X1 U5355 ( .A1(n4676), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U5356 ( .A1(n4304), .A2(EBX_REG_23__SCAN_IN), .ZN(n4362) );
  OAI211_X1 U5357 ( .C1(n4364), .C2(EBX_REG_23__SCAN_IN), .A(n4363), .B(n4362), 
        .ZN(n4365) );
  OR2_X1 U5358 ( .A1(n5573), .A2(n4365), .ZN(n4366) );
  AND2_X1 U5359 ( .A1(n4431), .A2(n4366), .ZN(n5568) );
  INV_X1 U5360 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4367) );
  NOR2_X1 U5361 ( .A1(n6253), .A2(n4367), .ZN(n4478) );
  NAND2_X1 U5362 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U5363 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U5364 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4368) );
  NOR3_X1 U5365 ( .A1(n4517), .A2(n6260), .A3(n4368), .ZN(n5389) );
  NAND2_X1 U5366 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6226) );
  INV_X1 U5367 ( .A(n6226), .ZN(n6208) );
  NAND3_X1 U5368 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6208), .ZN(n4379) );
  INV_X1 U5369 ( .A(n4379), .ZN(n5393) );
  NAND2_X1 U5370 ( .A1(n5389), .A2(n5393), .ZN(n5944) );
  INV_X1 U5371 ( .A(n4597), .ZN(n4371) );
  AND2_X1 U5372 ( .A1(n3408), .A2(n3120), .ZN(n6688) );
  AOI22_X1 U5373 ( .A1(n4506), .A2(n6688), .B1(n3386), .B2(n5435), .ZN(n4370)
         );
  OAI211_X1 U5374 ( .C1(n3718), .C2(n4371), .A(n4370), .B(n4369), .ZN(n4372)
         );
  INV_X1 U5375 ( .A(n4372), .ZN(n4373) );
  NAND2_X1 U5376 ( .A1(n4374), .A2(n4373), .ZN(n4576) );
  OAI21_X1 U5377 ( .B1(n3106), .B2(n4375), .A(n4762), .ZN(n4376) );
  NOR2_X1 U5378 ( .A1(n4576), .A2(n4376), .ZN(n4377) );
  NAND2_X1 U5379 ( .A1(n4273), .A2(n3120), .ZN(n4839) );
  NAND2_X1 U5380 ( .A1(n5416), .A2(n5952), .ZN(n5388) );
  INV_X1 U5381 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U5382 ( .A1(n5417), .A2(n5952), .ZN(n4681) );
  NAND2_X1 U5383 ( .A1(n5388), .A2(n4681), .ZN(n5712) );
  NOR2_X1 U5384 ( .A1(n5944), .A2(n5712), .ZN(n5394) );
  INV_X1 U5385 ( .A(n4745), .ZN(n4554) );
  AOI21_X1 U5386 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6259) );
  NOR2_X1 U5387 ( .A1(n6259), .A2(n6260), .ZN(n6239) );
  NAND3_X1 U5388 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6239), .ZN(n6204) );
  NOR2_X1 U5389 ( .A1(n4379), .A2(n6204), .ZN(n4388) );
  NOR2_X1 U5390 ( .A1(n3649), .A2(n4380), .ZN(n5414) );
  INV_X1 U5391 ( .A(n5414), .ZN(n5418) );
  NOR2_X1 U5392 ( .A1(n6721), .A2(n5418), .ZN(n5422) );
  NAND2_X1 U5393 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5422), .ZN(n5936) );
  NAND2_X1 U5394 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5841) );
  NOR2_X1 U5395 ( .A1(n5936), .A2(n5841), .ZN(n4387) );
  INV_X1 U5396 ( .A(n4387), .ZN(n4386) );
  INV_X1 U5397 ( .A(n4392), .ZN(n4381) );
  NAND2_X1 U5398 ( .A1(n5822), .A2(n4382), .ZN(n5779) );
  NOR2_X1 U5399 ( .A1(n5779), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4383)
         );
  AOI211_X1 U5400 ( .C1(n6266), .C2(n5568), .A(n4478), .B(n4383), .ZN(n4395)
         );
  NAND2_X1 U5401 ( .A1(n5822), .A2(n5813), .ZN(n5795) );
  NAND2_X1 U5402 ( .A1(n6253), .A2(n4385), .ZN(n4682) );
  OAI21_X1 U5403 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5416), .A(n4682), 
        .ZN(n5391) );
  AOI221_X1 U5404 ( .B1(n5944), .B2(n5388), .C1(n4386), .C2(n5388), .A(n5391), 
        .ZN(n4391) );
  NAND2_X1 U5405 ( .A1(n4388), .A2(n4387), .ZN(n4389) );
  NAND2_X1 U5406 ( .A1(n6252), .A2(n4389), .ZN(n4390) );
  NAND2_X1 U5407 ( .A1(n4391), .A2(n4390), .ZN(n5925) );
  NAND2_X1 U5408 ( .A1(n5813), .A2(n4392), .ZN(n4393) );
  AND2_X1 U5409 ( .A1(n5838), .A2(n4393), .ZN(n4394) );
  NOR2_X1 U5410 ( .A1(n5925), .A2(n4394), .ZN(n5798) );
  NAND2_X1 U5411 ( .A1(n4397), .A2(n4396), .ZN(U2995) );
  XNOR2_X2 U5412 ( .A(n4399), .B(n4398), .ZN(n5450) );
  INV_X1 U5413 ( .A(n5450), .ZN(n4400) );
  NAND2_X1 U5414 ( .A1(n4400), .A2(n3103), .ZN(n4409) );
  INV_X1 U5415 ( .A(n4456), .ZN(n4402) );
  INV_X1 U5416 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6656) );
  NOR2_X1 U5417 ( .A1(n6253), .A2(n6656), .ZN(n5724) );
  AOI21_X1 U5418 ( .B1(n6188), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5724), 
        .ZN(n4401) );
  OAI21_X1 U5419 ( .B1(n6195), .B2(n4402), .A(n4401), .ZN(n4403) );
  INV_X1 U5420 ( .A(n4403), .ZN(n4408) );
  NAND3_X1 U5421 ( .A1(n4409), .A2(n4408), .A3(n4407), .ZN(U2956) );
  INV_X1 U5422 ( .A(n4273), .ZN(n4411) );
  NOR2_X1 U5423 ( .A1(n4551), .A2(n4411), .ZN(n4545) );
  NAND2_X1 U5424 ( .A1(n4545), .A2(n4865), .ZN(n5867) );
  INV_X1 U5425 ( .A(n5966), .ZN(n6589) );
  NOR3_X1 U5426 ( .A1(n6665), .A2(n6952), .A3(n6589), .ZN(n4871) );
  NAND2_X1 U5427 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6952), .ZN(n6694) );
  INV_X1 U5428 ( .A(n6694), .ZN(n4412) );
  AND2_X1 U5429 ( .A1(n4158), .A2(n4412), .ZN(n6585) );
  INV_X1 U5430 ( .A(n6585), .ZN(n4413) );
  NAND2_X1 U5431 ( .A1(n4413), .A2(n6253), .ZN(n4414) );
  NAND2_X1 U5432 ( .A1(n6690), .A2(n6703), .ZN(n4451) );
  OR2_X1 U5433 ( .A1(n6689), .A2(n4451), .ZN(n4866) );
  AND2_X1 U5434 ( .A1(n3406), .A2(n4866), .ZN(n4491) );
  INV_X1 U5435 ( .A(n4491), .ZN(n4418) );
  INV_X1 U5436 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5467) );
  NAND3_X1 U5437 ( .A1(n4281), .A2(n4451), .A3(n5467), .ZN(n4417) );
  NAND2_X1 U5438 ( .A1(n4418), .A2(n4417), .ZN(n4419) );
  INV_X1 U5439 ( .A(n4451), .ZN(n4420) );
  AND3_X1 U5440 ( .A1(n4421), .A2(n4281), .A3(n4420), .ZN(n4422) );
  INV_X1 U5441 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6739) );
  INV_X1 U5442 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6628) );
  INV_X1 U5443 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6626) );
  INV_X1 U5444 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6619) );
  INV_X1 U5445 ( .A(REIP_REG_7__SCAN_IN), .ZN(n5337) );
  INV_X1 U5446 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6615) );
  INV_X1 U5447 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6613) );
  NAND3_X1 U5448 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5351) );
  NOR3_X1 U5449 ( .A1(n6615), .A2(n6613), .A3(n5351), .ZN(n5328) );
  NAND2_X1 U5450 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5328), .ZN(n5336) );
  NOR3_X1 U5451 ( .A1(n6619), .A2(n5337), .A3(n5336), .ZN(n5281) );
  NAND4_X1 U5452 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5281), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n5375) );
  NOR2_X1 U5453 ( .A1(n6626), .A2(n5375), .ZN(n6029) );
  NAND2_X1 U5454 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6029), .ZN(n6018) );
  NOR2_X1 U5455 ( .A1(n6628), .A2(n6018), .ZN(n5552) );
  NAND4_X1 U5456 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(n5552), .ZN(n5538) );
  INV_X1 U5457 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6635) );
  INV_X1 U5458 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6633) );
  NOR2_X1 U5459 ( .A1(n6635), .A2(n6633), .ZN(n5889) );
  INV_X1 U5460 ( .A(n5889), .ZN(n5539) );
  NOR3_X1 U5461 ( .A1(n6739), .A2(n5538), .A3(n5539), .ZN(n4460) );
  NAND3_X1 U5462 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4459) );
  INV_X1 U5463 ( .A(n4459), .ZN(n4423) );
  NAND2_X1 U5464 ( .A1(n5870), .A2(n4423), .ZN(n5511) );
  NAND3_X1 U5465 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4464) );
  NOR2_X1 U5466 ( .A1(n5511), .A2(n4464), .ZN(n5483) );
  AND2_X1 U5467 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n4466) );
  NAND2_X1 U5468 ( .A1(n5483), .A2(n4466), .ZN(n4495) );
  NOR3_X1 U5469 ( .A1(n4495), .A2(REIP_REG_30__SCAN_IN), .A3(n4494), .ZN(n4458) );
  INV_X1 U5470 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U5471 ( .A1(n4441), .A2(n6809), .ZN(n4427) );
  NAND2_X1 U5472 ( .A1(n4438), .A2(n5777), .ZN(n4425) );
  NAND2_X1 U5473 ( .A1(n4564), .A2(n6809), .ZN(n4424) );
  NAND3_X1 U5474 ( .A1(n4425), .A2(n4297), .A3(n4424), .ZN(n4426) );
  NAND2_X1 U5475 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4428) );
  OAI211_X1 U5476 ( .C1(n4676), .C2(EBX_REG_25__SCAN_IN), .A(n4438), .B(n4428), 
        .ZN(n4429) );
  OAI21_X1 U5477 ( .B1(n4430), .B2(EBX_REG_25__SCAN_IN), .A(n4429), .ZN(n4536)
         );
  OR3_X2 U5478 ( .A1(n4431), .A2(n5506), .A3(n4536), .ZN(n5495) );
  INV_X1 U5479 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4432) );
  NAND2_X1 U5480 ( .A1(n4441), .A2(n4432), .ZN(n4436) );
  INV_X1 U5481 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U5482 ( .A1(n4438), .A2(n5762), .ZN(n4434) );
  NAND2_X1 U5483 ( .A1(n4564), .A2(n4432), .ZN(n4433) );
  NAND3_X1 U5484 ( .A1(n4434), .A2(n4297), .A3(n4433), .ZN(n4435) );
  INV_X1 U5485 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U5486 ( .A1(n4483), .A2(n5563), .ZN(n4440) );
  NAND2_X1 U5487 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4437) );
  OAI211_X1 U5488 ( .C1(n4676), .C2(EBX_REG_27__SCAN_IN), .A(n4438), .B(n4437), 
        .ZN(n4439) );
  AND2_X1 U5489 ( .A1(n4440), .A2(n4439), .ZN(n5484) );
  AOI22_X1 U5490 ( .A1(n4304), .A2(EBX_REG_28__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n4676), .ZN(n4443) );
  INV_X1 U5491 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U5492 ( .A1(n4441), .A2(n5562), .ZN(n4442) );
  AND2_X1 U5493 ( .A1(n4443), .A2(n4442), .ZN(n5469) );
  NOR2_X1 U5494 ( .A1(n4597), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4484)
         );
  INV_X1 U5495 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6916) );
  AND2_X1 U5496 ( .A1(n4564), .A2(n6916), .ZN(n4444) );
  INV_X1 U5497 ( .A(n4448), .ZN(n4447) );
  AND2_X1 U5498 ( .A1(n4676), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4445)
         );
  AOI21_X1 U5499 ( .B1(n4597), .B2(EBX_REG_30__SCAN_IN), .A(n4445), .ZN(n4488)
         );
  INV_X1 U5500 ( .A(n4488), .ZN(n4446) );
  NOR2_X1 U5501 ( .A1(n4448), .A2(n5808), .ZN(n4487) );
  AOI211_X1 U5502 ( .C1(n3209), .C2(n4447), .A(n4446), .B(n4487), .ZN(n4450)
         );
  AOI211_X1 U5503 ( .C1(n5808), .C2(n5471), .A(n4488), .B(n4448), .ZN(n4449)
         );
  NAND2_X1 U5504 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4451), .ZN(n4452) );
  NOR2_X1 U5505 ( .A1(n4676), .A2(n4452), .ZN(n4453) );
  AOI22_X1 U5506 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6094), .B1(n6071), 
        .B2(n4456), .ZN(n4457) );
  NOR2_X1 U5507 ( .A1(n4495), .A2(REIP_REG_29__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U5508 ( .A1(n6083), .A2(n6084), .ZN(n6086) );
  NAND2_X1 U5509 ( .A1(n6086), .A2(n4459), .ZN(n4463) );
  INV_X1 U5510 ( .A(n4460), .ZN(n4461) );
  NAND2_X1 U5511 ( .A1(n6063), .A2(n4461), .ZN(n4462) );
  AND2_X1 U5512 ( .A1(n4462), .A2(n6084), .ZN(n5890) );
  NAND2_X1 U5513 ( .A1(n4463), .A2(n5890), .ZN(n5877) );
  AND2_X1 U5514 ( .A1(n6086), .A2(n4464), .ZN(n4465) );
  NOR2_X1 U5515 ( .A1(n5877), .A2(n4465), .ZN(n5482) );
  INV_X1 U5516 ( .A(n4466), .ZN(n4467) );
  NAND2_X1 U5517 ( .A1(n6063), .A2(n4467), .ZN(n4468) );
  NAND2_X1 U5518 ( .A1(n5482), .A2(n4468), .ZN(n5474) );
  NOR2_X1 U5519 ( .A1(n5444), .A2(n5474), .ZN(n4496) );
  INV_X1 U5520 ( .A(n4496), .ZN(n4469) );
  NAND2_X1 U5521 ( .A1(n4469), .A2(REIP_REG_30__SCAN_IN), .ZN(n4470) );
  OAI21_X1 U5522 ( .B1(n5450), .B2(n5873), .A(n4471), .ZN(U2797) );
  NAND2_X1 U5523 ( .A1(n4472), .A2(n6191), .ZN(n4482) );
  NAND2_X1 U5524 ( .A1(n4474), .A2(n4475), .ZN(n4476) );
  NAND2_X1 U5525 ( .A1(n4473), .A2(n4476), .ZN(n5874) );
  NOR2_X1 U5526 ( .A1(n5686), .A2(n5880), .ZN(n4477) );
  AOI211_X1 U5527 ( .C1(n6168), .C2(n5869), .A(n4478), .B(n4477), .ZN(n4479)
         );
  NAND2_X1 U5528 ( .A1(n4482), .A2(n4481), .ZN(U2963) );
  NAND2_X1 U5529 ( .A1(n5595), .A2(n6056), .ZN(n4502) );
  AOI22_X1 U5530 ( .A1(n4483), .A2(n6916), .B1(n5808), .B2(EBX_REG_29__SCAN_IN), .ZN(n4486) );
  INV_X1 U5531 ( .A(n4484), .ZN(n4485) );
  NAND2_X1 U5532 ( .A1(n4486), .A2(n4485), .ZN(n4510) );
  NOR2_X1 U5533 ( .A1(n5471), .A2(n4510), .ZN(n4511) );
  AOI21_X1 U5534 ( .B1(n4488), .B2(n4511), .A(n4487), .ZN(n4490) );
  AOI22_X1 U5535 ( .A1(n4597), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4676), .ZN(n4489) );
  XNOR2_X1 U5536 ( .A(n4490), .B(n4489), .ZN(n5710) );
  INV_X1 U5537 ( .A(n5710), .ZN(n5468) );
  NAND3_X1 U5538 ( .A1(n5262), .A2(EBX_REG_31__SCAN_IN), .A3(n4491), .ZN(n4493) );
  NAND2_X1 U5539 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4492)
         );
  OAI211_X1 U5540 ( .C1(n5468), .C2(n5871), .A(n4493), .B(n4492), .ZN(n4500)
         );
  NOR4_X1 U5541 ( .A1(n4495), .A2(REIP_REG_31__SCAN_IN), .A3(n6656), .A4(n4494), .ZN(n4499) );
  OAI21_X1 U5542 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6083), .A(n4496), .ZN(n4497) );
  NOR3_X1 U5543 ( .A1(n4500), .A2(n4499), .A3(n4498), .ZN(n4501) );
  NAND2_X1 U5544 ( .A1(n4502), .A2(n4501), .ZN(U2796) );
  NAND3_X1 U5545 ( .A1(n4745), .A2(n4865), .A3(n4589), .ZN(n4509) );
  AND2_X1 U5546 ( .A1(n4503), .A2(n6981), .ZN(n4507) );
  INV_X1 U5547 ( .A(n4504), .ZN(n4505) );
  NAND4_X1 U5548 ( .A1(n4507), .A2(n4506), .A3(n4505), .A4(n4221), .ZN(n4689)
         );
  NAND2_X1 U5549 ( .A1(n5434), .A2(n6114), .ZN(n4516) );
  AND2_X1 U5550 ( .A1(n5471), .A2(n4510), .ZN(n4512) );
  INV_X1 U5551 ( .A(n5731), .ZN(n4514) );
  INV_X1 U5552 ( .A(n4893), .ZN(n5593) );
  NOR2_X1 U5553 ( .A1(n4517), .A2(n5712), .ZN(n6244) );
  NOR2_X1 U5554 ( .A1(n6252), .A2(n6244), .ZN(n6258) );
  NAND2_X1 U5555 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6239), .ZN(n4519)
         );
  NOR2_X1 U5556 ( .A1(n6258), .A2(n4519), .ZN(n4521) );
  AOI21_X1 U5557 ( .B1(n5388), .B2(n4517), .A(n5391), .ZN(n4518) );
  INV_X1 U5558 ( .A(n4518), .ZN(n6251) );
  AOI21_X1 U5559 ( .B1(n5838), .B2(n4519), .A(n6251), .ZN(n6250) );
  INV_X1 U5560 ( .A(n6250), .ZN(n4520) );
  MUX2_X1 U5561 ( .A(n4521), .B(n4520), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4530) );
  OAI21_X1 U5562 ( .B1(n4524), .B2(n4523), .A(n4522), .ZN(n6173) );
  NOR2_X1 U5563 ( .A1(n6173), .A2(n6223), .ZN(n4529) );
  OAI21_X1 U5564 ( .B1(n4526), .B2(n4819), .A(n4525), .ZN(n5330) );
  INV_X1 U5565 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4527) );
  OAI22_X1 U5566 ( .A1(n6255), .A2(n5330), .B1(n6253), .B2(n4527), .ZN(n4528)
         );
  OR3_X1 U5567 ( .A1(n4530), .A2(n4529), .A3(n4528), .ZN(U3012) );
  INV_X1 U5568 ( .A(n4531), .ZN(n4534) );
  AOI21_X1 U5569 ( .B1(n4534), .B2(n3229), .A(n4533), .ZN(n5641) );
  INV_X1 U5570 ( .A(n5641), .ZN(n5607) );
  NOR2_X1 U5571 ( .A1(n5607), .A2(n5873), .ZN(n4544) );
  AND2_X1 U5572 ( .A1(n5877), .A2(REIP_REG_25__SCAN_IN), .ZN(n4543) );
  XNOR2_X1 U5573 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n4535) );
  NOR2_X1 U5574 ( .A1(n5511), .A2(n4535), .ZN(n4542) );
  OAI21_X1 U5575 ( .B1(n4431), .B2(n5506), .A(n4536), .ZN(n4537) );
  NAND2_X1 U5576 ( .A1(n4537), .A2(n5495), .ZN(n5769) );
  INV_X1 U5577 ( .A(n5639), .ZN(n4538) );
  AOI22_X1 U5578 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6094), .B1(n6071), 
        .B2(n4538), .ZN(n4540) );
  NAND2_X1 U5579 ( .A1(n6090), .A2(EBX_REG_25__SCAN_IN), .ZN(n4539) );
  OAI211_X1 U5580 ( .C1(n5769), .C2(n5871), .A(n4540), .B(n4539), .ZN(n4541)
         );
  OR4_X1 U5581 ( .A1(n4544), .A2(n4543), .A3(n4542), .A4(n4541), .ZN(U2802) );
  NAND2_X1 U5582 ( .A1(n4589), .A2(n3671), .ZN(n4547) );
  OR2_X1 U5583 ( .A1(n4545), .A2(n4410), .ZN(n4546) );
  NAND2_X1 U5584 ( .A1(n4547), .A2(n4546), .ZN(n5967) );
  OR2_X1 U5585 ( .A1(n3406), .A2(n6688), .ZN(n4559) );
  AOI21_X1 U5586 ( .B1(n4559), .B2(n6689), .A(READY_N), .ZN(n4548) );
  NOR2_X1 U5587 ( .A1(n5967), .A2(n4548), .ZN(n4857) );
  NOR2_X1 U5588 ( .A1(n4857), .A2(n6582), .ZN(n5974) );
  INV_X1 U5589 ( .A(MORE_REG_SCAN_IN), .ZN(n4556) );
  NAND2_X1 U5590 ( .A1(n4550), .A2(n4549), .ZN(n4552) );
  AOI22_X1 U5591 ( .A1(n4589), .A2(n4552), .B1(n4551), .B2(n4273), .ZN(n4553)
         );
  OAI21_X1 U5592 ( .B1(n4554), .B2(n4589), .A(n4553), .ZN(n4856) );
  NAND2_X1 U5593 ( .A1(n5974), .A2(n4856), .ZN(n4555) );
  OAI21_X1 U5594 ( .B1(n5974), .B2(n4556), .A(n4555), .ZN(U3471) );
  AND2_X1 U5595 ( .A1(n6409), .A2(n6981), .ZN(n5272) );
  INV_X1 U5596 ( .A(n5272), .ZN(n4557) );
  NAND2_X1 U5597 ( .A1(n4594), .A2(n4557), .ZN(n5866) );
  NOR2_X1 U5598 ( .A1(n5866), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4558) );
  AND2_X1 U5599 ( .A1(n4558), .A2(n5867), .ZN(n4560) );
  OAI22_X1 U5600 ( .A1(n4560), .A2(n4559), .B1(n4558), .B2(n6685), .ZN(U3474)
         );
  INV_X1 U5601 ( .A(n4561), .ZN(n4562) );
  OAI22_X1 U5602 ( .A1(n4589), .A2(n4743), .B1(n4562), .B2(n4282), .ZN(n4691)
         );
  INV_X1 U5603 ( .A(n6689), .ZN(n6692) );
  OAI21_X1 U5604 ( .B1(n6692), .B2(n4564), .A(n4563), .ZN(n4565) );
  OAI21_X1 U5605 ( .B1(n4839), .B2(n6689), .A(n4565), .ZN(n4566) );
  NAND2_X1 U5606 ( .A1(n4566), .A2(n6690), .ZN(n4570) );
  INV_X1 U5607 ( .A(n4567), .ZN(n4569) );
  NAND2_X1 U5608 ( .A1(n6688), .A2(n3399), .ZN(n4568) );
  OAI211_X1 U5609 ( .C1(n4589), .C2(n4570), .A(n4569), .B(n4568), .ZN(n4571)
         );
  OR2_X1 U5610 ( .A1(n4691), .A2(n4571), .ZN(n4573) );
  AND2_X1 U5611 ( .A1(n4745), .A2(n4589), .ZN(n4572) );
  NAND2_X1 U5612 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4786), .ZN(n6662) );
  INV_X1 U5613 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5973) );
  NOR2_X1 U5614 ( .A1(n6662), .A2(n5973), .ZN(n4574) );
  AOI21_X1 U5615 ( .B1(n4842), .B2(n4865), .A(n4574), .ZN(n5961) );
  NAND2_X1 U5616 ( .A1(n6952), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U5617 ( .A1(n5961), .A2(n6663), .ZN(n6669) );
  INV_X1 U5618 ( .A(n6669), .ZN(n5465) );
  INV_X1 U5619 ( .A(n4576), .ZN(n4581) );
  INV_X1 U5620 ( .A(n4577), .ZN(n4579) );
  AND4_X1 U5621 ( .A1(n4282), .A2(n4868), .A3(n4579), .A4(n4578), .ZN(n4580)
         );
  NAND2_X1 U5622 ( .A1(n4581), .A2(n4580), .ZN(n4834) );
  NAND2_X1 U5623 ( .A1(n4575), .A2(n4834), .ZN(n4587) );
  INV_X1 U5624 ( .A(n4582), .ZN(n5456) );
  INV_X1 U5625 ( .A(n4583), .ZN(n4780) );
  NAND3_X1 U5626 ( .A1(n4835), .A2(n5456), .A3(n4780), .ZN(n4584) );
  OAI21_X1 U5627 ( .B1(n4839), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4584), 
        .ZN(n4585) );
  INV_X1 U5628 ( .A(n4585), .ZN(n4586) );
  NAND2_X1 U5629 ( .A1(n4587), .A2(n4586), .ZN(n4841) );
  INV_X1 U5630 ( .A(n6673), .ZN(n6667) );
  INV_X1 U5631 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6991) );
  AOI22_X1 U5632 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6991), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6795), .ZN(n5460) );
  NOR2_X1 U5633 ( .A1(n6981), .A2(n5417), .ZN(n5457) );
  INV_X1 U5634 ( .A(n5862), .ZN(n5458) );
  AOI222_X1 U5635 ( .A1(n4841), .A2(n6667), .B1(n5460), .B2(n5457), .C1(n4588), 
        .C2(n5458), .ZN(n4592) );
  NAND2_X1 U5636 ( .A1(n5458), .A2(n4838), .ZN(n6666) );
  INV_X1 U5637 ( .A(n6666), .ZN(n4590) );
  OAI21_X1 U5638 ( .B1(n5465), .B2(n4590), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4591) );
  OAI21_X1 U5639 ( .B1(n5465), .B2(n4592), .A(n4591), .ZN(U3460) );
  INV_X1 U5640 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6894) );
  OR2_X1 U5641 ( .A1(n4594), .A2(n3120), .ZN(n4671) );
  NAND2_X1 U5642 ( .A1(n3120), .A2(n6690), .ZN(n4593) );
  NAND2_X1 U5643 ( .A1(n6146), .A2(DATAI_10_), .ZN(n6152) );
  INV_X1 U5644 ( .A(n4594), .ZN(n4595) );
  NAND2_X1 U5645 ( .A1(n4646), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4596) );
  OAI211_X1 U5646 ( .C1(n6894), .C2(n4671), .A(n6152), .B(n4596), .ZN(U2934)
         );
  NOR2_X1 U5647 ( .A1(n4597), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4598)
         );
  OR2_X1 U5648 ( .A1(n4599), .A2(n4598), .ZN(n4639) );
  AND2_X1 U5649 ( .A1(n4600), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4603) );
  OAI21_X1 U5650 ( .B1(n4603), .B2(n4602), .A(n4601), .ZN(n6136) );
  OAI222_X1 U5651 ( .A1(n4639), .A2(n5591), .B1(n6929), .B2(n6117), .C1(n6136), 
        .C2(n5592), .ZN(U2859) );
  INV_X2 U5652 ( .A(n4671), .ZN(n6158) );
  AOI22_X1 U5653 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n4646), .B1(n6158), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n4604) );
  INV_X1 U5654 ( .A(DATAI_3_), .ZN(n4809) );
  OR2_X1 U5655 ( .A1(n4692), .A2(n4809), .ZN(n4647) );
  NAND2_X1 U5656 ( .A1(n4604), .A2(n4647), .ZN(U2927) );
  AOI22_X1 U5657 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n4646), .B1(n6158), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n4605) );
  INV_X1 U5658 ( .A(DATAI_0_), .ZN(n6132) );
  OR2_X1 U5659 ( .A1(n4692), .A2(n6132), .ZN(n4649) );
  NAND2_X1 U5660 ( .A1(n4605), .A2(n4649), .ZN(U2924) );
  AOI22_X1 U5661 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n4646), .B1(n6158), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U5662 ( .A1(n6146), .A2(DATAI_2_), .ZN(n4653) );
  NAND2_X1 U5663 ( .A1(n4606), .A2(n4653), .ZN(U2926) );
  AOI22_X1 U5664 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n4646), .B1(n6158), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n4607) );
  NAND2_X1 U5665 ( .A1(n6146), .A2(DATAI_1_), .ZN(n4662) );
  NAND2_X1 U5666 ( .A1(n4607), .A2(n4662), .ZN(U2925) );
  AOI22_X1 U5667 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n4646), .B1(n6158), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n4608) );
  INV_X1 U5668 ( .A(DATAI_4_), .ZN(n4815) );
  OR2_X1 U5669 ( .A1(n4692), .A2(n4815), .ZN(n4658) );
  NAND2_X1 U5670 ( .A1(n4608), .A2(n4658), .ZN(U2928) );
  INV_X1 U5671 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4614) );
  NAND2_X1 U5672 ( .A1(n4786), .A2(n6952), .ZN(n6142) );
  INV_X1 U5673 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4613) );
  INV_X1 U5674 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4612) );
  OAI222_X1 U5675 ( .A1(n4614), .A2(n4717), .B1(n4708), .B2(n4613), .C1(n4612), 
        .C2(n6142), .ZN(U2906) );
  INV_X1 U5676 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4616) );
  INV_X1 U5677 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6705) );
  INV_X1 U5678 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n4615) );
  OAI222_X1 U5679 ( .A1(n4616), .A2(n4717), .B1(n4636), .B2(n6705), .C1(n4615), 
        .C2(n6142), .ZN(U2909) );
  INV_X1 U5680 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4619) );
  INV_X1 U5681 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4618) );
  INV_X1 U5682 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4617) );
  OAI222_X1 U5683 ( .A1(n4619), .A2(n4717), .B1(n4708), .B2(n4618), .C1(n4617), 
        .C2(n6142), .ZN(U2901) );
  INV_X1 U5684 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4622) );
  INV_X1 U5685 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4621) );
  INV_X1 U5686 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4620) );
  OAI222_X1 U5687 ( .A1(n4622), .A2(n4717), .B1(n4708), .B2(n4621), .C1(n4620), 
        .C2(n6142), .ZN(U2902) );
  INV_X1 U5688 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4625) );
  INV_X1 U5689 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4624) );
  INV_X1 U5690 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4623) );
  OAI222_X1 U5691 ( .A1(n4625), .A2(n4717), .B1(n4708), .B2(n4624), .C1(n4623), 
        .C2(n6142), .ZN(U2900) );
  INV_X1 U5692 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n4628) );
  INV_X1 U5693 ( .A(EAX_REG_13__SCAN_IN), .ZN(n4627) );
  INV_X1 U5694 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4626) );
  OAI222_X1 U5695 ( .A1(n4628), .A2(n6142), .B1(n4636), .B2(n4627), .C1(n4717), 
        .C2(n4626), .ZN(U2910) );
  INV_X1 U5696 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n4631) );
  INV_X1 U5697 ( .A(EAX_REG_11__SCAN_IN), .ZN(n4630) );
  INV_X1 U5698 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4629) );
  OAI222_X1 U5699 ( .A1(n4631), .A2(n6142), .B1(n4636), .B2(n4630), .C1(n4717), 
        .C2(n4629), .ZN(U2912) );
  INV_X1 U5700 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n4634) );
  INV_X1 U5701 ( .A(EAX_REG_9__SCAN_IN), .ZN(n4633) );
  INV_X1 U5702 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4632) );
  OAI222_X1 U5703 ( .A1(n4634), .A2(n6142), .B1(n4636), .B2(n4633), .C1(n4717), 
        .C2(n4632), .ZN(U2914) );
  INV_X1 U5704 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n4637) );
  INV_X1 U5705 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4635) );
  OAI222_X1 U5706 ( .A1(n4637), .A2(n6142), .B1(n4636), .B2(n5383), .C1(n4717), 
        .C2(n4635), .ZN(U2911) );
  XOR2_X1 U5707 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .B(n4638), .Z(n4709) );
  INV_X1 U5708 ( .A(n4709), .ZN(n4645) );
  INV_X1 U5709 ( .A(n4639), .ZN(n5261) );
  INV_X1 U5710 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6680) );
  INV_X1 U5711 ( .A(n5413), .ZN(n4640) );
  NAND2_X1 U5712 ( .A1(n5417), .A2(n4640), .ZN(n4641) );
  OAI21_X1 U5713 ( .B1(n6253), .B2(n6680), .A(n4641), .ZN(n4643) );
  AOI21_X1 U5714 ( .B1(n5952), .B2(n4682), .A(n5417), .ZN(n4642) );
  AOI211_X1 U5715 ( .C1(n6266), .C2(n5261), .A(n4643), .B(n4642), .ZN(n4644)
         );
  OAI21_X1 U5716 ( .B1(n4645), .B2(n6223), .A(n4644), .ZN(U3018) );
  AOI22_X1 U5717 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U5718 ( .A1(n4648), .A2(n4647), .ZN(U2942) );
  AOI22_X1 U5719 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n4650) );
  NAND2_X1 U5720 ( .A1(n4650), .A2(n4649), .ZN(U2939) );
  AOI22_X1 U5721 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n4651) );
  INV_X1 U5722 ( .A(DATAI_6_), .ZN(n6744) );
  OR2_X1 U5723 ( .A1(n4692), .A2(n6744), .ZN(n4656) );
  NAND2_X1 U5724 ( .A1(n4651), .A2(n4656), .ZN(U2930) );
  AOI22_X1 U5725 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n4652) );
  INV_X1 U5726 ( .A(DATAI_5_), .ZN(n4913) );
  OR2_X1 U5727 ( .A1(n4692), .A2(n4913), .ZN(n4660) );
  NAND2_X1 U5728 ( .A1(n4652), .A2(n4660), .ZN(U2929) );
  AOI22_X1 U5729 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U5730 ( .A1(n4654), .A2(n4653), .ZN(U2941) );
  AOI22_X1 U5731 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n4655) );
  OR2_X1 U5732 ( .A1(n4692), .A2(n5119), .ZN(n4664) );
  NAND2_X1 U5733 ( .A1(n4655), .A2(n4664), .ZN(U2931) );
  AOI22_X1 U5734 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U5735 ( .A1(n4657), .A2(n4656), .ZN(U2945) );
  AOI22_X1 U5736 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4659) );
  NAND2_X1 U5737 ( .A1(n4659), .A2(n4658), .ZN(U2943) );
  AOI22_X1 U5738 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4661) );
  NAND2_X1 U5739 ( .A1(n4661), .A2(n4660), .ZN(U2944) );
  AOI22_X1 U5740 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4663) );
  NAND2_X1 U5741 ( .A1(n4663), .A2(n4662), .ZN(U2940) );
  AOI22_X1 U5742 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U5743 ( .A1(n4665), .A2(n4664), .ZN(U2946) );
  INV_X1 U5744 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6812) );
  NAND2_X1 U5745 ( .A1(n6146), .A2(DATAI_13_), .ZN(n6160) );
  NAND2_X1 U5746 ( .A1(n6159), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4666) );
  OAI211_X1 U5747 ( .C1(n6812), .C2(n4671), .A(n6160), .B(n4666), .ZN(U2937)
         );
  NAND2_X1 U5748 ( .A1(n6146), .A2(DATAI_14_), .ZN(n4669) );
  NAND2_X1 U5749 ( .A1(n6159), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4667) );
  OAI211_X1 U5750 ( .C1(n6705), .C2(n4671), .A(n4669), .B(n4667), .ZN(U2953)
         );
  INV_X1 U5751 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U5752 ( .A1(n6159), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4668) );
  OAI211_X1 U5753 ( .C1(n6887), .C2(n4671), .A(n4669), .B(n4668), .ZN(U2938)
         );
  INV_X1 U5754 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4672) );
  AOI22_X1 U5755 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6159), .B1(n6146), .B2(
        DATAI_15_), .ZN(n4670) );
  OAI21_X1 U5756 ( .B1(n4672), .B2(n4671), .A(n4670), .ZN(U2954) );
  OR2_X1 U5757 ( .A1(n4674), .A2(n4673), .ZN(n4675) );
  AND2_X1 U5758 ( .A1(n3744), .A2(n4675), .ZN(n6102) );
  INV_X1 U5759 ( .A(n6102), .ZN(n4696) );
  XNOR2_X1 U5760 ( .A(n6091), .B(n4676), .ZN(n4686) );
  INV_X1 U5761 ( .A(n4686), .ZN(n4677) );
  AOI22_X1 U5762 ( .A1(n6113), .A2(n4677), .B1(n5588), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4678) );
  OAI21_X1 U5763 ( .B1(n4696), .B2(n5592), .A(n4678), .ZN(U2858) );
  XOR2_X1 U5764 ( .A(n4680), .B(n4679), .Z(n4822) );
  NAND3_X1 U5765 ( .A1(n5838), .A2(n4681), .A3(n6795), .ZN(n4685) );
  INV_X2 U5766 ( .A(n6253), .ZN(n6197) );
  OAI21_X1 U5767 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5413), .A(n4682), 
        .ZN(n4683) );
  AOI22_X1 U5768 ( .A1(n6197), .A2(REIP_REG_1__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n4683), .ZN(n4684) );
  OAI211_X1 U5769 ( .C1(n6255), .C2(n4686), .A(n4685), .B(n4684), .ZN(n4687)
         );
  AOI21_X1 U5770 ( .B1(n4822), .B2(n6269), .A(n4687), .ZN(n4688) );
  INV_X1 U5771 ( .A(n4688), .ZN(U3017) );
  NOR2_X1 U5772 ( .A1(n4689), .A2(n3671), .ZN(n4690) );
  NAND2_X1 U5773 ( .A1(n4268), .A2(n4893), .ZN(n4694) );
  INV_X1 U5774 ( .A(n4694), .ZN(n4695) );
  INV_X1 U5775 ( .A(DATAI_1_), .ZN(n6738) );
  INV_X1 U5776 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6903) );
  OAI222_X1 U5777 ( .A1(n4696), .A2(n6135), .B1(n6133), .B2(n6738), .C1(n6134), 
        .C2(n6903), .ZN(U2890) );
  INV_X1 U5778 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U5779 ( .A1(n6140), .A2(DATAO_REG_27__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U5780 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6687), .ZN(n4697) );
  OAI211_X1 U5781 ( .C1(n4708), .C2(n4699), .A(n4698), .B(n4697), .ZN(U2896)
         );
  INV_X1 U5782 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4702) );
  NAND2_X1 U5783 ( .A1(n6140), .A2(DATAO_REG_25__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U5784 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6687), .ZN(n4700) );
  OAI211_X1 U5785 ( .C1(n4708), .C2(n4702), .A(n4701), .B(n4700), .ZN(U2898)
         );
  NAND2_X1 U5786 ( .A1(n6140), .A2(DATAO_REG_24__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U5787 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n6687), .ZN(n4703) );
  OAI211_X1 U5788 ( .C1(n4708), .C2(n4075), .A(n4704), .B(n4703), .ZN(U2899)
         );
  INV_X1 U5789 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U5790 ( .A1(n6140), .A2(DATAO_REG_28__SCAN_IN), .ZN(n4706) );
  NAND2_X1 U5791 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6687), .ZN(n4705) );
  OAI211_X1 U5792 ( .C1(n4708), .C2(n4707), .A(n4706), .B(n4705), .ZN(U2895)
         );
  NAND2_X1 U5793 ( .A1(n4709), .A2(n6191), .ZN(n4713) );
  NAND2_X1 U5794 ( .A1(n5686), .A2(n4710), .ZN(n4711) );
  AOI22_X1 U5795 ( .A1(n4711), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6197), 
        .B2(REIP_REG_0__SCAN_IN), .ZN(n4712) );
  OAI211_X1 U5796 ( .C1(n5696), .C2(n6136), .A(n4713), .B(n4712), .ZN(U2986)
         );
  AOI222_X1 U5797 ( .A1(n6140), .A2(DATAO_REG_20__SCAN_IN), .B1(n4729), .B2(
        EAX_REG_20__SCAN_IN), .C1(UWORD_REG_4__SCAN_IN), .C2(n6687), .ZN(n4714) );
  INV_X1 U5798 ( .A(n4714), .ZN(U2903) );
  AOI222_X1 U5799 ( .A1(n6140), .A2(DATAO_REG_18__SCAN_IN), .B1(n4729), .B2(
        EAX_REG_18__SCAN_IN), .C1(UWORD_REG_2__SCAN_IN), .C2(n6687), .ZN(n4715) );
  INV_X1 U5800 ( .A(n4715), .ZN(U2905) );
  AOI222_X1 U5801 ( .A1(EAX_REG_30__SCAN_IN), .A2(n4729), .B1(
        DATAO_REG_30__SCAN_IN), .B2(n6140), .C1(UWORD_REG_14__SCAN_IN), .C2(
        n6687), .ZN(n4716) );
  INV_X1 U5802 ( .A(n4716), .ZN(U2893) );
  AOI222_X1 U5803 ( .A1(EAX_REG_0__SCAN_IN), .A2(n6139), .B1(n6140), .B2(
        DATAO_REG_0__SCAN_IN), .C1(LWORD_REG_0__SCAN_IN), .C2(n6687), .ZN(
        n4718) );
  INV_X1 U5804 ( .A(n4718), .ZN(U2923) );
  AOI222_X1 U5805 ( .A1(EAX_REG_1__SCAN_IN), .A2(n6139), .B1(n6140), .B2(
        DATAO_REG_1__SCAN_IN), .C1(n6687), .C2(LWORD_REG_1__SCAN_IN), .ZN(
        n4719) );
  INV_X1 U5806 ( .A(n4719), .ZN(U2922) );
  AOI222_X1 U5807 ( .A1(EAX_REG_2__SCAN_IN), .A2(n6139), .B1(n6140), .B2(
        DATAO_REG_2__SCAN_IN), .C1(n6687), .C2(LWORD_REG_2__SCAN_IN), .ZN(
        n4720) );
  INV_X1 U5808 ( .A(n4720), .ZN(U2921) );
  AOI222_X1 U5809 ( .A1(EAX_REG_3__SCAN_IN), .A2(n6139), .B1(n6140), .B2(
        DATAO_REG_3__SCAN_IN), .C1(n6687), .C2(LWORD_REG_3__SCAN_IN), .ZN(
        n4721) );
  INV_X1 U5810 ( .A(n4721), .ZN(U2920) );
  AOI222_X1 U5811 ( .A1(EAX_REG_4__SCAN_IN), .A2(n6139), .B1(n6140), .B2(
        DATAO_REG_4__SCAN_IN), .C1(n6687), .C2(LWORD_REG_4__SCAN_IN), .ZN(
        n4722) );
  INV_X1 U5812 ( .A(n4722), .ZN(U2919) );
  AOI222_X1 U5813 ( .A1(EAX_REG_5__SCAN_IN), .A2(n6139), .B1(n6140), .B2(
        DATAO_REG_5__SCAN_IN), .C1(n6687), .C2(LWORD_REG_5__SCAN_IN), .ZN(
        n4723) );
  INV_X1 U5814 ( .A(n4723), .ZN(U2918) );
  AOI222_X1 U5815 ( .A1(EAX_REG_7__SCAN_IN), .A2(n6139), .B1(n6140), .B2(
        DATAO_REG_7__SCAN_IN), .C1(LWORD_REG_7__SCAN_IN), .C2(n6687), .ZN(
        n4724) );
  INV_X1 U5816 ( .A(n4724), .ZN(U2916) );
  AOI222_X1 U5817 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6139), .B1(n6140), .B2(
        DATAO_REG_15__SCAN_IN), .C1(n6687), .C2(LWORD_REG_15__SCAN_IN), .ZN(
        n4725) );
  INV_X1 U5818 ( .A(n4725), .ZN(U2908) );
  AOI222_X1 U5819 ( .A1(EAX_REG_16__SCAN_IN), .A2(n4729), .B1(n6140), .B2(
        DATAO_REG_16__SCAN_IN), .C1(UWORD_REG_0__SCAN_IN), .C2(n6687), .ZN(
        n4726) );
  INV_X1 U5820 ( .A(n4726), .ZN(U2907) );
  AOI222_X1 U5821 ( .A1(EAX_REG_19__SCAN_IN), .A2(n4729), .B1(n6140), .B2(
        DATAO_REG_19__SCAN_IN), .C1(UWORD_REG_3__SCAN_IN), .C2(n6687), .ZN(
        n4727) );
  INV_X1 U5822 ( .A(n4727), .ZN(U2904) );
  AOI222_X1 U5823 ( .A1(EAX_REG_26__SCAN_IN), .A2(n4729), .B1(n6140), .B2(
        DATAO_REG_26__SCAN_IN), .C1(UWORD_REG_10__SCAN_IN), .C2(n6687), .ZN(
        n4728) );
  INV_X1 U5824 ( .A(n4728), .ZN(U2897) );
  AOI222_X1 U5825 ( .A1(EAX_REG_29__SCAN_IN), .A2(n4729), .B1(n6140), .B2(
        DATAO_REG_29__SCAN_IN), .C1(UWORD_REG_13__SCAN_IN), .C2(n6687), .ZN(
        n4730) );
  INV_X1 U5826 ( .A(n4730), .ZN(U2894) );
  NAND3_X1 U5827 ( .A1(n4732), .A2(n4733), .A3(n3744), .ZN(n4734) );
  AND2_X1 U5828 ( .A1(n4731), .A2(n4734), .ZN(n6190) );
  INV_X1 U5829 ( .A(n6190), .ZN(n4736) );
  INV_X1 U5830 ( .A(DATAI_2_), .ZN(n6810) );
  INV_X1 U5831 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4735) );
  OAI222_X1 U5832 ( .A1(n4736), .A2(n6135), .B1(n6133), .B2(n6810), .C1(n6134), 
        .C2(n4735), .ZN(U2889) );
  INV_X1 U5833 ( .A(n5592), .ZN(n6114) );
  OR2_X1 U5834 ( .A1(n4738), .A2(n4737), .ZN(n4739) );
  NAND2_X1 U5835 ( .A1(n4739), .A2(n4805), .ZN(n6076) );
  OAI22_X1 U5836 ( .A1(n6076), .A2(n5591), .B1(n6081), .B2(n6117), .ZN(n4740)
         );
  AOI21_X1 U5837 ( .B1(n6190), .B2(n6114), .A(n4740), .ZN(n4741) );
  INV_X1 U5838 ( .A(n4741), .ZN(U2857) );
  NAND2_X1 U5839 ( .A1(n3118), .A2(n4834), .ZN(n4759) );
  INV_X1 U5840 ( .A(n4743), .ZN(n4744) );
  OR2_X1 U5841 ( .A1(n4745), .A2(n4744), .ZN(n4766) );
  MUX2_X1 U5842 ( .A(n4746), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4582), 
        .Z(n4748) );
  NOR2_X1 U5843 ( .A1(n4748), .A2(n4747), .ZN(n4757) );
  AND2_X1 U5844 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4749) );
  INV_X1 U5845 ( .A(n4749), .ZN(n4750) );
  MUX2_X1 U5846 ( .A(n4750), .B(n4749), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4755) );
  INV_X1 U5847 ( .A(n4751), .ZN(n4752) );
  OAI21_X1 U5848 ( .B1(n4582), .B2(n3195), .A(n4752), .ZN(n4754) );
  NOR2_X1 U5849 ( .A1(n4754), .A2(n4753), .ZN(n5863) );
  OAI22_X1 U5850 ( .A1(n4839), .A2(n4755), .B1(n5863), .B2(n4762), .ZN(n4756)
         );
  AOI21_X1 U5851 ( .B1(n4766), .B2(n4757), .A(n4756), .ZN(n4758) );
  NAND2_X1 U5852 ( .A1(n4759), .A2(n4758), .ZN(n5861) );
  MUX2_X1 U5853 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5861), .S(n4842), 
        .Z(n4851) );
  INV_X1 U5854 ( .A(n4851), .ZN(n4854) );
  NAND2_X1 U5855 ( .A1(n4761), .A2(n4834), .ZN(n4768) );
  XNOR2_X1 U5856 ( .A(n4582), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4765)
         );
  XNOR2_X1 U5857 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4763) );
  OAI22_X1 U5858 ( .A1(n4839), .A2(n4763), .B1(n4762), .B2(n4765), .ZN(n4764)
         );
  AOI21_X1 U5859 ( .B1(n4766), .B2(n4765), .A(n4764), .ZN(n4767) );
  NAND2_X1 U5860 ( .A1(n4768), .A2(n4767), .ZN(n5463) );
  NAND2_X1 U5861 ( .A1(n5463), .A2(n4842), .ZN(n4771) );
  INV_X1 U5862 ( .A(n4842), .ZN(n4769) );
  NAND2_X1 U5863 ( .A1(n4769), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4770) );
  NAND2_X1 U5864 ( .A1(n4771), .A2(n4770), .ZN(n4848) );
  NAND2_X1 U5865 ( .A1(n4848), .A2(n6981), .ZN(n4773) );
  NAND2_X1 U5866 ( .A1(n5973), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4776) );
  INV_X1 U5867 ( .A(n4747), .ZN(n4772) );
  OAI22_X1 U5868 ( .A1(n4854), .A2(n4773), .B1(n4776), .B2(n4772), .ZN(n4862)
         );
  INV_X1 U5869 ( .A(n5187), .ZN(n6438) );
  NOR2_X1 U5870 ( .A1(n4774), .A2(n6438), .ZN(n4775) );
  XNOR2_X1 U5871 ( .A(n4775), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5962)
         );
  OAI22_X1 U5872 ( .A1(n5962), .A2(n4282), .B1(n5964), .B2(n4842), .ZN(n4778)
         );
  INV_X1 U5873 ( .A(n4776), .ZN(n4777) );
  AOI22_X1 U5874 ( .A1(n4778), .A2(n6981), .B1(n4777), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4861) );
  INV_X1 U5875 ( .A(n4861), .ZN(n4779) );
  AOI21_X1 U5876 ( .B1(n4780), .B2(n4862), .A(n4779), .ZN(n4873) );
  AND2_X1 U5877 ( .A1(n4873), .A2(n5973), .ZN(n4781) );
  OAI21_X1 U5878 ( .B1(n4781), .B2(n6662), .A(n5184), .ZN(n6275) );
  INV_X1 U5879 ( .A(n6275), .ZN(n4789) );
  XNOR2_X1 U5880 ( .A(n4782), .B(n6515), .ZN(n4783) );
  NAND2_X1 U5881 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6665), .ZN(n5850) );
  AOI22_X1 U5882 ( .A1(n4783), .A2(n6409), .B1(n5850), .B2(n4761), .ZN(n4785)
         );
  NAND2_X1 U5883 ( .A1(n4789), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4784) );
  OAI21_X1 U5884 ( .B1(n4789), .B2(n4785), .A(n4784), .ZN(U3463) );
  INV_X1 U5885 ( .A(n5136), .ZN(n5181) );
  AOI222_X1 U5886 ( .A1(n4873), .A2(n4786), .B1(n3130), .B2(n5850), .C1(n5181), 
        .C2(n6409), .ZN(n4788) );
  NAND2_X1 U5887 ( .A1(n4789), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4787) );
  OAI21_X1 U5888 ( .B1(n4789), .B2(n4788), .A(n4787), .ZN(U3465) );
  XNOR2_X1 U5889 ( .A(n3105), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4791)
         );
  XNOR2_X1 U5890 ( .A(n4792), .B(n4791), .ZN(n6189) );
  INV_X1 U5891 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4793) );
  OAI22_X1 U5892 ( .A1(n6076), .A2(n6255), .B1(n6253), .B2(n4793), .ZN(n4799)
         );
  NOR2_X1 U5893 ( .A1(n6795), .A2(n5712), .ZN(n4797) );
  AOI21_X1 U5894 ( .B1(n6252), .B2(n4794), .A(n6251), .ZN(n4795) );
  INV_X1 U5895 ( .A(n4795), .ZN(n4796) );
  MUX2_X1 U5896 ( .A(n4797), .B(n4796), .S(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .Z(n4798) );
  AOI211_X1 U5897 ( .C1(n6252), .C2(n6259), .A(n4799), .B(n4798), .ZN(n4800)
         );
  OAI21_X1 U5898 ( .B1(n6223), .B2(n6189), .A(n4800), .ZN(U3016) );
  INV_X1 U5899 ( .A(n4803), .ZN(n4804) );
  AOI21_X1 U5900 ( .B1(n4802), .B2(n4731), .A(n4804), .ZN(n6065) );
  INV_X1 U5901 ( .A(n6065), .ZN(n4810) );
  AOI21_X1 U5902 ( .B1(n4806), .B2(n4805), .A(n4881), .ZN(n6265) );
  AOI22_X1 U5903 ( .A1(n6113), .A2(n6265), .B1(n5588), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4807) );
  OAI21_X1 U5904 ( .B1(n4810), .B2(n5592), .A(n4807), .ZN(U2856) );
  INV_X1 U5905 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4808) );
  OAI222_X1 U5906 ( .A1(n4810), .A2(n6135), .B1(n6133), .B2(n4809), .C1(n6134), 
        .C2(n4808), .ZN(U2888) );
  AND2_X1 U5907 ( .A1(n4803), .A2(n4811), .ZN(n4813) );
  OR2_X1 U5908 ( .A1(n4813), .A2(n4812), .ZN(n6183) );
  INV_X1 U5909 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4814) );
  OAI222_X1 U5910 ( .A1(n6183), .A2(n6135), .B1(n6133), .B2(n4815), .C1(n6134), 
        .C2(n4814), .ZN(U2887) );
  OAI21_X1 U5911 ( .B1(n4812), .B2(n4818), .A(n4817), .ZN(n5280) );
  AOI21_X1 U5912 ( .B1(n4820), .B2(n4880), .A(n4819), .ZN(n6242) );
  AOI22_X1 U5913 ( .A1(n6113), .A2(n6242), .B1(n5588), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4821) );
  OAI21_X1 U5914 ( .B1(n5280), .B2(n5592), .A(n4821), .ZN(U2854) );
  INV_X1 U5915 ( .A(n4822), .ZN(n4826) );
  AOI22_X1 U5916 ( .A1(n6188), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6197), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4823) );
  OAI21_X1 U5917 ( .B1(n6195), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4823), 
        .ZN(n4824) );
  AOI21_X1 U5918 ( .B1(n6102), .B2(n3103), .A(n4824), .ZN(n4825) );
  OAI21_X1 U5919 ( .B1(n4826), .B2(n6172), .A(n4825), .ZN(U2985) );
  INV_X1 U5920 ( .A(n6072), .ZN(n4831) );
  INV_X1 U5921 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4829) );
  NOR2_X1 U5922 ( .A1(n6253), .A2(n4829), .ZN(n6264) );
  AOI21_X1 U5923 ( .B1(n6188), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6264), 
        .ZN(n4830) );
  OAI21_X1 U5924 ( .B1(n6195), .B2(n4831), .A(n4830), .ZN(n4832) );
  AOI21_X1 U5925 ( .B1(n6065), .B2(n3103), .A(n4832), .ZN(n4833) );
  OAI21_X1 U5926 ( .B1(n6172), .B2(n6267), .A(n4833), .ZN(U2983) );
  AOI21_X1 U5927 ( .B1(n5966), .B2(n5458), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n4878) );
  NAND2_X1 U5928 ( .A1(n4848), .A2(n6279), .ZN(n4847) );
  NAND2_X1 U5929 ( .A1(n3130), .A2(n4834), .ZN(n4837) );
  NAND2_X1 U5930 ( .A1(n4835), .A2(n4838), .ZN(n4836) );
  NAND2_X1 U5931 ( .A1(n4837), .A2(n4836), .ZN(n6668) );
  OR2_X1 U5932 ( .A1(n4839), .A2(n4838), .ZN(n6674) );
  INV_X1 U5933 ( .A(n6674), .ZN(n4840) );
  OR2_X1 U5934 ( .A1(n6668), .A2(n4840), .ZN(n4844) );
  OAI211_X1 U5935 ( .C1(n4844), .C2(n4843), .A(n4842), .B(n4841), .ZN(n4846)
         );
  OAI21_X1 U5936 ( .B1(n4844), .B2(n6398), .A(n6358), .ZN(n4845) );
  NAND3_X1 U5937 ( .A1(n4847), .A2(n4846), .A3(n4845), .ZN(n4850) );
  OR2_X1 U5938 ( .A1(n4848), .A2(n6279), .ZN(n4849) );
  AND2_X1 U5939 ( .A1(n4850), .A2(n4849), .ZN(n4852) );
  INV_X1 U5940 ( .A(n4852), .ZN(n4855) );
  OAI21_X1 U5941 ( .B1(n4852), .B2(n4851), .A(n6359), .ZN(n4853) );
  OAI21_X1 U5942 ( .B1(n4855), .B2(n4854), .A(n4853), .ZN(n4864) );
  INV_X1 U5943 ( .A(n4856), .ZN(n4860) );
  OAI21_X1 U5944 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n4857), 
        .ZN(n4858) );
  NAND4_X1 U5945 ( .A1(n4861), .A2(n4860), .A3(n4859), .A4(n4858), .ZN(n4863)
         );
  AOI211_X1 U5946 ( .C1(n6276), .C2(n4864), .A(n4863), .B(n4862), .ZN(n4875)
         );
  AOI22_X1 U5947 ( .A1(n4875), .A2(n4865), .B1(READY_N), .B2(n6687), .ZN(n4870) );
  NOR3_X1 U5948 ( .A1(n4868), .A2(n4867), .A3(n4866), .ZN(n4869) );
  INV_X1 U5949 ( .A(n6662), .ZN(n4872) );
  AOI21_X1 U5950 ( .B1(n4873), .B2(n4872), .A(n4871), .ZN(n4874) );
  OAI21_X1 U5951 ( .B1(n4875), .B2(n6582), .A(n4874), .ZN(n4877) );
  NAND2_X1 U5952 ( .A1(READY_N), .A2(n6695), .ZN(n6588) );
  AOI21_X1 U5953 ( .B1(n6588), .B2(n6664), .A(n6952), .ZN(n4876) );
  AOI211_X1 U5954 ( .C1(n4878), .C2(n6664), .A(n4877), .B(n4876), .ZN(n4879)
         );
  INV_X1 U5955 ( .A(n4879), .ZN(U3148) );
  OAI21_X1 U5956 ( .B1(n4882), .B2(n4881), .A(n4880), .ZN(n6254) );
  OAI222_X1 U5957 ( .A1(n6254), .A2(n5591), .B1(n6117), .B2(n4313), .C1(n5592), 
        .C2(n6183), .ZN(U2855) );
  AND2_X1 U5958 ( .A1(n3103), .A2(DATAI_19_), .ZN(n6548) );
  INV_X1 U5959 ( .A(n6548), .ZN(n6461) );
  NOR3_X1 U5960 ( .A1(n6279), .A2(n6359), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5185) );
  NOR2_X1 U5961 ( .A1(n6354), .A2(n6484), .ZN(n4942) );
  INV_X1 U5962 ( .A(n4575), .ZN(n5852) );
  INV_X1 U5963 ( .A(n5185), .ZN(n4885) );
  NOR2_X1 U5964 ( .A1(n6398), .A2(n4885), .ZN(n4909) );
  AOI21_X1 U5965 ( .B1(n4942), .B2(n6362), .A(n4909), .ZN(n4887) );
  NAND2_X1 U5966 ( .A1(n4940), .A2(n6360), .ZN(n5854) );
  NAND3_X1 U5967 ( .A1(n6409), .A2(n4887), .A3(n5854), .ZN(n4884) );
  OAI211_X1 U5968 ( .C1(n6409), .C2(n5185), .A(n6406), .B(n4884), .ZN(n4907)
         );
  NAND2_X1 U5969 ( .A1(DATAI_3_), .A2(n5079), .ZN(n6552) );
  NAND2_X1 U5970 ( .A1(n6409), .A2(n5854), .ZN(n4886) );
  OAI22_X1 U5971 ( .A1(n4887), .A2(n4886), .B1(n6695), .B2(n4885), .ZN(n4906)
         );
  AOI22_X1 U5972 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4907), .B1(n6458), 
        .B2(n4906), .ZN(n4892) );
  INV_X1 U5973 ( .A(n6663), .ZN(n4890) );
  NAND2_X1 U5974 ( .A1(n4908), .A2(n3531), .ZN(n6330) );
  AOI22_X1 U5975 ( .A1(n5217), .A2(n6549), .B1(n6547), .B2(n4909), .ZN(n4891)
         );
  OAI211_X1 U5976 ( .C1(n6461), .C2(n5076), .A(n4892), .B(n4891), .ZN(U3127)
         );
  AND2_X1 U5977 ( .A1(n3103), .A2(DATAI_23_), .ZN(n6576) );
  INV_X1 U5978 ( .A(n6576), .ZN(n6482) );
  NAND2_X1 U5979 ( .A1(DATAI_7_), .A2(n5079), .ZN(n6580) );
  AOI22_X1 U5980 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4907), .B1(n6476), 
        .B2(n4906), .ZN(n4895) );
  AND2_X1 U5981 ( .A1(n3103), .A2(DATAI_31_), .ZN(n6573) );
  NAND2_X1 U5982 ( .A1(n4908), .A2(n4893), .ZN(n6347) );
  AOI22_X1 U5983 ( .A1(n5217), .A2(n6573), .B1(n6572), .B2(n4909), .ZN(n4894)
         );
  OAI211_X1 U5984 ( .C1(n6482), .C2(n5076), .A(n4895), .B(n4894), .ZN(U3131)
         );
  AND2_X1 U5985 ( .A1(n3103), .A2(DATAI_21_), .ZN(n6561) );
  NAND2_X1 U5986 ( .A1(DATAI_5_), .A2(n5079), .ZN(n6564) );
  AOI22_X1 U5987 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4907), .B1(n6466), 
        .B2(n4906), .ZN(n4897) );
  AND2_X1 U5988 ( .A1(n3103), .A2(DATAI_29_), .ZN(n6560) );
  NAND2_X1 U5989 ( .A1(n4908), .A2(n3119), .ZN(n6338) );
  AOI22_X1 U5990 ( .A1(n5217), .A2(n6560), .B1(n6559), .B2(n4909), .ZN(n4896)
         );
  OAI211_X1 U5991 ( .C1(n6469), .C2(n5076), .A(n4897), .B(n4896), .ZN(U3129)
         );
  AND2_X1 U5992 ( .A1(n3103), .A2(DATAI_20_), .ZN(n6555) );
  INV_X1 U5993 ( .A(n6555), .ZN(n6465) );
  NAND2_X1 U5994 ( .A1(DATAI_4_), .A2(n5079), .ZN(n6558) );
  AOI22_X1 U5995 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4907), .B1(n6462), 
        .B2(n4906), .ZN(n4899) );
  NAND2_X1 U5996 ( .A1(n3103), .A2(DATAI_28_), .ZN(n6383) );
  NAND2_X1 U5997 ( .A1(n4908), .A2(n3381), .ZN(n6334) );
  AOI22_X1 U5998 ( .A1(n5217), .A2(n6554), .B1(n6553), .B2(n4909), .ZN(n4898)
         );
  OAI211_X1 U5999 ( .C1(n6465), .C2(n5076), .A(n4899), .B(n4898), .ZN(U3128)
         );
  AND2_X1 U6000 ( .A1(n3103), .A2(DATAI_22_), .ZN(n6566) );
  INV_X1 U6001 ( .A(n6566), .ZN(n6473) );
  NAND2_X1 U6002 ( .A1(DATAI_6_), .A2(n5079), .ZN(n6570) );
  AOI22_X1 U6003 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4907), .B1(n6470), 
        .B2(n4906), .ZN(n4901) );
  AND2_X1 U6004 ( .A1(n3103), .A2(DATAI_30_), .ZN(n6567) );
  NAND2_X1 U6005 ( .A1(n4908), .A2(n3367), .ZN(n6342) );
  AOI22_X1 U6006 ( .A1(n5217), .A2(n6567), .B1(n6565), .B2(n4909), .ZN(n4900)
         );
  OAI211_X1 U6007 ( .C1(n6473), .C2(n5076), .A(n4901), .B(n4900), .ZN(U3130)
         );
  AND2_X1 U6008 ( .A1(n3103), .A2(DATAI_18_), .ZN(n6543) );
  NAND2_X1 U6009 ( .A1(DATAI_2_), .A2(n5079), .ZN(n6546) );
  AOI22_X1 U6010 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4907), .B1(n6454), 
        .B2(n4906), .ZN(n4903) );
  AND2_X1 U6011 ( .A1(n3103), .A2(DATAI_26_), .ZN(n6542) );
  NAND2_X1 U6012 ( .A1(n4908), .A2(n3386), .ZN(n6326) );
  AOI22_X1 U6013 ( .A1(n5217), .A2(n6542), .B1(n6541), .B2(n4909), .ZN(n4902)
         );
  OAI211_X1 U6014 ( .C1(n6457), .C2(n5076), .A(n4903), .B(n4902), .ZN(U3126)
         );
  NAND2_X1 U6015 ( .A1(n3103), .A2(DATAI_17_), .ZN(n6453) );
  NAND2_X1 U6016 ( .A1(DATAI_1_), .A2(n5079), .ZN(n6540) );
  AOI22_X1 U6017 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4907), .B1(n6450), 
        .B2(n4906), .ZN(n4905) );
  AND2_X1 U6018 ( .A1(n3103), .A2(DATAI_25_), .ZN(n6537) );
  NAND2_X1 U6019 ( .A1(n4908), .A2(n3120), .ZN(n6322) );
  AOI22_X1 U6020 ( .A1(n5217), .A2(n6537), .B1(n6535), .B2(n4909), .ZN(n4904)
         );
  OAI211_X1 U6021 ( .C1(n6453), .C2(n5076), .A(n4905), .B(n4904), .ZN(U3125)
         );
  NAND2_X1 U6022 ( .A1(n3103), .A2(DATAI_16_), .ZN(n6449) );
  NAND2_X1 U6023 ( .A1(DATAI_0_), .A2(n5079), .ZN(n6534) );
  AOI22_X1 U6024 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4907), .B1(n6437), 
        .B2(n4906), .ZN(n4911) );
  NAND2_X1 U6025 ( .A1(n4908), .A2(n4281), .ZN(n6309) );
  AOI22_X1 U6026 ( .A1(n5217), .A2(n6531), .B1(n6522), .B2(n4909), .ZN(n4910)
         );
  OAI211_X1 U6027 ( .C1(n6449), .C2(n5076), .A(n4911), .B(n4910), .ZN(U3124)
         );
  INV_X1 U6028 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4912) );
  OAI222_X1 U6029 ( .A1(n5280), .A2(n6135), .B1(n6133), .B2(n4913), .C1(n6134), 
        .C2(n4912), .ZN(U2886) );
  INV_X1 U6030 ( .A(n6403), .ZN(n4915) );
  OR2_X1 U6031 ( .A1(n4761), .A2(n4575), .ZN(n4977) );
  NAND3_X1 U6032 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6279), .A3(n6358), .ZN(n5221) );
  NOR2_X1 U6033 ( .A1(n6398), .A2(n5221), .ZN(n4936) );
  AOI21_X1 U6034 ( .B1(n4942), .B2(n5229), .A(n4936), .ZN(n4919) );
  AOI21_X1 U6035 ( .B1(n6516), .B2(n6360), .A(n6527), .ZN(n4917) );
  AOI22_X1 U6036 ( .A1(n4919), .A2(n4917), .B1(n6527), .B2(n5221), .ZN(n4916)
         );
  NAND2_X1 U6037 ( .A1(n6406), .A2(n4916), .ZN(n4935) );
  INV_X1 U6038 ( .A(n4917), .ZN(n4918) );
  OAI22_X1 U6039 ( .A1(n4919), .A2(n4918), .B1(n6695), .B2(n5221), .ZN(n4934)
         );
  AOI22_X1 U6040 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4935), .B1(n6476), 
        .B2(n4934), .ZN(n4921) );
  AOI22_X1 U6041 ( .A1(n4937), .A2(n6573), .B1(n6572), .B2(n4936), .ZN(n4920)
         );
  OAI211_X1 U6042 ( .C1(n6482), .C2(n5139), .A(n4921), .B(n4920), .ZN(U3099)
         );
  AOI22_X1 U6043 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4935), .B1(n6470), 
        .B2(n4934), .ZN(n4923) );
  AOI22_X1 U6044 ( .A1(n4937), .A2(n6567), .B1(n6565), .B2(n4936), .ZN(n4922)
         );
  OAI211_X1 U6045 ( .C1(n6473), .C2(n5139), .A(n4923), .B(n4922), .ZN(U3098)
         );
  AOI22_X1 U6046 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4935), .B1(n6462), 
        .B2(n4934), .ZN(n4925) );
  AOI22_X1 U6047 ( .A1(n4937), .A2(n6554), .B1(n6553), .B2(n4936), .ZN(n4924)
         );
  OAI211_X1 U6048 ( .C1(n6465), .C2(n5139), .A(n4925), .B(n4924), .ZN(U3096)
         );
  AOI22_X1 U6049 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4935), .B1(n6458), 
        .B2(n4934), .ZN(n4927) );
  AOI22_X1 U6050 ( .A1(n4937), .A2(n6549), .B1(n6547), .B2(n4936), .ZN(n4926)
         );
  OAI211_X1 U6051 ( .C1(n6461), .C2(n5139), .A(n4927), .B(n4926), .ZN(U3095)
         );
  AOI22_X1 U6052 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4935), .B1(n6466), 
        .B2(n4934), .ZN(n4929) );
  AOI22_X1 U6053 ( .A1(n4937), .A2(n6560), .B1(n6559), .B2(n4936), .ZN(n4928)
         );
  OAI211_X1 U6054 ( .C1(n6469), .C2(n5139), .A(n4929), .B(n4928), .ZN(U3097)
         );
  AOI22_X1 U6055 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4935), .B1(n6450), 
        .B2(n4934), .ZN(n4931) );
  AOI22_X1 U6056 ( .A1(n4937), .A2(n6537), .B1(n6535), .B2(n4936), .ZN(n4930)
         );
  OAI211_X1 U6057 ( .C1(n6453), .C2(n5139), .A(n4931), .B(n4930), .ZN(U3093)
         );
  AOI22_X1 U6058 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4935), .B1(n6437), 
        .B2(n4934), .ZN(n4933) );
  AOI22_X1 U6059 ( .A1(n4937), .A2(n6531), .B1(n6522), .B2(n4936), .ZN(n4932)
         );
  OAI211_X1 U6060 ( .C1(n6449), .C2(n5139), .A(n4933), .B(n4932), .ZN(U3092)
         );
  AOI22_X1 U6061 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4935), .B1(n6454), 
        .B2(n4934), .ZN(n4939) );
  AOI22_X1 U6062 ( .A1(n4937), .A2(n6542), .B1(n6541), .B2(n4936), .ZN(n4938)
         );
  OAI211_X1 U6063 ( .C1(n6457), .C2(n5139), .A(n4939), .B(n4938), .ZN(U3094)
         );
  NAND2_X1 U6064 ( .A1(n4940), .A2(n3129), .ZN(n4946) );
  INV_X1 U6065 ( .A(n4946), .ZN(n4943) );
  INV_X1 U6066 ( .A(n6549), .ZN(n6380) );
  INV_X1 U6067 ( .A(n4972), .ZN(n4941) );
  AOI21_X1 U6068 ( .B1(n4942), .B2(n6439), .A(n4941), .ZN(n4947) );
  NAND2_X1 U6069 ( .A1(n6409), .A2(n6703), .ZN(n6280) );
  OAI21_X1 U6070 ( .B1(n4943), .B2(n5696), .A(n6280), .ZN(n4944) );
  AOI22_X1 U6071 ( .A1(n4947), .A2(n4944), .B1(n5075), .B2(n6527), .ZN(n4945)
         );
  NAND2_X1 U6072 ( .A1(n6406), .A2(n4945), .ZN(n4971) );
  NAND2_X1 U6073 ( .A1(n4971), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4952)
         );
  NOR2_X2 U6074 ( .A1(n4946), .A2(n5136), .ZN(n5017) );
  INV_X1 U6075 ( .A(n4947), .ZN(n4949) );
  AOI22_X1 U6076 ( .A1(n4949), .A2(n6409), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4948), .ZN(n4973) );
  OAI22_X1 U6077 ( .A1(n6552), .A2(n4973), .B1(n4972), .B2(n6330), .ZN(n4950)
         );
  AOI21_X1 U6078 ( .B1(n6548), .B2(n5017), .A(n4950), .ZN(n4951) );
  OAI211_X1 U6079 ( .C1(n5111), .C2(n6380), .A(n4952), .B(n4951), .ZN(U3143)
         );
  NAND2_X1 U6080 ( .A1(n4971), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4955)
         );
  OAI22_X1 U6081 ( .A1(n6558), .A2(n4973), .B1(n4972), .B2(n6334), .ZN(n4953)
         );
  AOI21_X1 U6082 ( .B1(n6555), .B2(n5017), .A(n4953), .ZN(n4954) );
  OAI211_X1 U6083 ( .C1(n5111), .C2(n6383), .A(n4955), .B(n4954), .ZN(U3144)
         );
  INV_X1 U6084 ( .A(n6560), .ZN(n6386) );
  NAND2_X1 U6085 ( .A1(n4971), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4958)
         );
  OAI22_X1 U6086 ( .A1(n6564), .A2(n4973), .B1(n4972), .B2(n6338), .ZN(n4956)
         );
  AOI21_X1 U6087 ( .B1(n6561), .B2(n5017), .A(n4956), .ZN(n4957) );
  OAI211_X1 U6088 ( .C1(n5111), .C2(n6386), .A(n4958), .B(n4957), .ZN(U3145)
         );
  INV_X1 U6089 ( .A(n6567), .ZN(n6389) );
  NAND2_X1 U6090 ( .A1(n4971), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4961)
         );
  OAI22_X1 U6091 ( .A1(n6570), .A2(n4973), .B1(n4972), .B2(n6342), .ZN(n4959)
         );
  AOI21_X1 U6092 ( .B1(n6566), .B2(n5017), .A(n4959), .ZN(n4960) );
  OAI211_X1 U6093 ( .C1(n5111), .C2(n6389), .A(n4961), .B(n4960), .ZN(U3146)
         );
  INV_X1 U6094 ( .A(n6542), .ZN(n6377) );
  NAND2_X1 U6095 ( .A1(n4971), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4964)
         );
  OAI22_X1 U6096 ( .A1(n6546), .A2(n4973), .B1(n4972), .B2(n6326), .ZN(n4962)
         );
  AOI21_X1 U6097 ( .B1(n6543), .B2(n5017), .A(n4962), .ZN(n4963) );
  OAI211_X1 U6098 ( .C1(n5111), .C2(n6377), .A(n4964), .B(n4963), .ZN(U3142)
         );
  INV_X1 U6099 ( .A(n6537), .ZN(n6374) );
  NAND2_X1 U6100 ( .A1(n4971), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4967)
         );
  INV_X1 U6101 ( .A(n6453), .ZN(n6536) );
  OAI22_X1 U6102 ( .A1(n6540), .A2(n4973), .B1(n4972), .B2(n6322), .ZN(n4965)
         );
  AOI21_X1 U6103 ( .B1(n6536), .B2(n5017), .A(n4965), .ZN(n4966) );
  OAI211_X1 U6104 ( .C1(n5111), .C2(n6374), .A(n4967), .B(n4966), .ZN(U3141)
         );
  INV_X1 U6105 ( .A(n6531), .ZN(n6371) );
  NAND2_X1 U6106 ( .A1(n4971), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4970)
         );
  INV_X1 U6107 ( .A(n6449), .ZN(n6523) );
  OAI22_X1 U6108 ( .A1(n6534), .A2(n4973), .B1(n4972), .B2(n6309), .ZN(n4968)
         );
  AOI21_X1 U6109 ( .B1(n6523), .B2(n5017), .A(n4968), .ZN(n4969) );
  OAI211_X1 U6110 ( .C1(n6371), .C2(n5111), .A(n4970), .B(n4969), .ZN(U3140)
         );
  INV_X1 U6111 ( .A(n6573), .ZN(n6396) );
  NAND2_X1 U6112 ( .A1(n4971), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4976)
         );
  OAI22_X1 U6113 ( .A1(n6580), .A2(n4973), .B1(n4972), .B2(n6347), .ZN(n4974)
         );
  AOI21_X1 U6114 ( .B1(n6576), .B2(n5017), .A(n4974), .ZN(n4975) );
  OAI211_X1 U6115 ( .C1(n5111), .C2(n6396), .A(n4976), .B(n4975), .ZN(U3147)
         );
  NOR2_X1 U6116 ( .A1(n3118), .A2(n4977), .ZN(n4984) );
  INV_X1 U6117 ( .A(n4782), .ZN(n4978) );
  NAND2_X1 U6118 ( .A1(n6307), .A2(n6360), .ZN(n4979) );
  NAND2_X1 U6119 ( .A1(n4979), .A2(n6409), .ZN(n5032) );
  AOI211_X1 U6120 ( .C1(n5017), .C2(n6280), .A(n4984), .B(n5032), .ZN(n4982)
         );
  INV_X1 U6121 ( .A(n4980), .ZN(n5183) );
  INV_X1 U6122 ( .A(n5182), .ZN(n6278) );
  NOR2_X1 U6123 ( .A1(n5183), .A2(n6278), .ZN(n4986) );
  OAI21_X1 U6124 ( .B1(n4986), .B2(n6695), .A(n5079), .ZN(n6364) );
  NAND3_X1 U6125 ( .A1(n6359), .A2(n6279), .A3(n6358), .ZN(n5030) );
  NOR2_X1 U6126 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5030), .ZN(n5013)
         );
  NOR2_X1 U6127 ( .A1(n6665), .A2(n5013), .ZN(n4981) );
  NOR4_X2 U6128 ( .A1(n4982), .A2(n6355), .A3(n6364), .A4(n4981), .ZN(n5020)
         );
  INV_X1 U6129 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U6130 ( .A1(n6307), .A2(n4983), .ZN(n5064) );
  INV_X1 U6131 ( .A(n4984), .ZN(n5027) );
  NOR2_X1 U6132 ( .A1(n4985), .A2(n6695), .ZN(n6363) );
  INV_X1 U6133 ( .A(n6363), .ZN(n6444) );
  INV_X1 U6134 ( .A(n4986), .ZN(n6356) );
  OAI22_X1 U6135 ( .A1(n5027), .A2(n6527), .B1(n6444), .B2(n6356), .ZN(n5014)
         );
  AOI22_X1 U6136 ( .A1(n6462), .A2(n5014), .B1(n6553), .B2(n5013), .ZN(n4987)
         );
  OAI21_X1 U6137 ( .B1(n5064), .B2(n6465), .A(n4987), .ZN(n4988) );
  AOI21_X1 U6138 ( .B1(n6554), .B2(n5017), .A(n4988), .ZN(n4989) );
  OAI21_X1 U6139 ( .B1(n5020), .B2(n4990), .A(n4989), .ZN(U3024) );
  AOI22_X1 U6140 ( .A1(n6476), .A2(n5014), .B1(n6572), .B2(n5013), .ZN(n4991)
         );
  OAI21_X1 U6141 ( .B1(n5064), .B2(n6482), .A(n4991), .ZN(n4992) );
  AOI21_X1 U6142 ( .B1(n6573), .B2(n5017), .A(n4992), .ZN(n4993) );
  OAI21_X1 U6143 ( .B1(n5020), .B2(n6818), .A(n4993), .ZN(U3027) );
  INV_X1 U6144 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4997) );
  AOI22_X1 U6145 ( .A1(n6450), .A2(n5014), .B1(n6535), .B2(n5013), .ZN(n4994)
         );
  OAI21_X1 U6146 ( .B1(n5064), .B2(n6453), .A(n4994), .ZN(n4995) );
  AOI21_X1 U6147 ( .B1(n6537), .B2(n5017), .A(n4995), .ZN(n4996) );
  OAI21_X1 U6148 ( .B1(n5020), .B2(n4997), .A(n4996), .ZN(U3021) );
  AOI22_X1 U6149 ( .A1(n6454), .A2(n5014), .B1(n6541), .B2(n5013), .ZN(n4998)
         );
  OAI21_X1 U6150 ( .B1(n5064), .B2(n6457), .A(n4998), .ZN(n4999) );
  AOI21_X1 U6151 ( .B1(n6542), .B2(n5017), .A(n4999), .ZN(n5000) );
  OAI21_X1 U6152 ( .B1(n5020), .B2(n3428), .A(n5000), .ZN(U3022) );
  INV_X1 U6153 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5004) );
  AOI22_X1 U6154 ( .A1(n6458), .A2(n5014), .B1(n6547), .B2(n5013), .ZN(n5001)
         );
  OAI21_X1 U6155 ( .B1(n5064), .B2(n6461), .A(n5001), .ZN(n5002) );
  AOI21_X1 U6156 ( .B1(n6549), .B2(n5017), .A(n5002), .ZN(n5003) );
  OAI21_X1 U6157 ( .B1(n5020), .B2(n5004), .A(n5003), .ZN(U3023) );
  INV_X1 U6158 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5008) );
  AOI22_X1 U6159 ( .A1(n6470), .A2(n5014), .B1(n6565), .B2(n5013), .ZN(n5005)
         );
  OAI21_X1 U6160 ( .B1(n5064), .B2(n6473), .A(n5005), .ZN(n5006) );
  AOI21_X1 U6161 ( .B1(n6567), .B2(n5017), .A(n5006), .ZN(n5007) );
  OAI21_X1 U6162 ( .B1(n5020), .B2(n5008), .A(n5007), .ZN(U3026) );
  INV_X1 U6163 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5012) );
  AOI22_X1 U6164 ( .A1(n6466), .A2(n5014), .B1(n6559), .B2(n5013), .ZN(n5009)
         );
  OAI21_X1 U6165 ( .B1(n5064), .B2(n6469), .A(n5009), .ZN(n5010) );
  AOI21_X1 U6166 ( .B1(n6560), .B2(n5017), .A(n5010), .ZN(n5011) );
  OAI21_X1 U6167 ( .B1(n5020), .B2(n5012), .A(n5011), .ZN(U3025) );
  INV_X1 U6168 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5019) );
  AOI22_X1 U6169 ( .A1(n6437), .A2(n5014), .B1(n6522), .B2(n5013), .ZN(n5015)
         );
  OAI21_X1 U6170 ( .B1(n5064), .B2(n6449), .A(n5015), .ZN(n5016) );
  AOI21_X1 U6171 ( .B1(n6531), .B2(n5017), .A(n5016), .ZN(n5018) );
  OAI21_X1 U6172 ( .B1(n5020), .B2(n5019), .A(n5018), .ZN(U3020) );
  INV_X1 U6173 ( .A(n5022), .ZN(n5023) );
  AOI21_X1 U6174 ( .B1(n5024), .B2(n4817), .A(n5023), .ZN(n6174) );
  INV_X1 U6175 ( .A(n6174), .ZN(n5070) );
  OAI222_X1 U6176 ( .A1(n5070), .A2(n6135), .B1(n6134), .B2(n5025), .C1(n6133), 
        .C2(n6744), .ZN(U2885) );
  NOR2_X1 U6177 ( .A1(n6398), .A2(n5030), .ZN(n5062) );
  INV_X1 U6178 ( .A(n5062), .ZN(n5026) );
  OAI21_X1 U6179 ( .B1(n5027), .B2(n6484), .A(n5026), .ZN(n5029) );
  NOR2_X1 U6180 ( .A1(n5032), .A2(n5029), .ZN(n5028) );
  AOI211_X2 U6181 ( .C1(n5030), .C2(n6527), .A(n6525), .B(n5028), .ZN(n5069)
         );
  INV_X1 U6182 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5037) );
  INV_X1 U6183 ( .A(n5029), .ZN(n5031) );
  OAI22_X1 U6184 ( .A1(n5032), .A2(n5031), .B1(n5030), .B2(n6695), .ZN(n5066)
         );
  INV_X1 U6185 ( .A(n6307), .ZN(n5033) );
  AOI22_X1 U6186 ( .A1(n6301), .A2(n6566), .B1(n6565), .B2(n5062), .ZN(n5034)
         );
  OAI21_X1 U6187 ( .B1(n6389), .B2(n5064), .A(n5034), .ZN(n5035) );
  AOI21_X1 U6188 ( .B1(n6470), .B2(n5066), .A(n5035), .ZN(n5036) );
  OAI21_X1 U6189 ( .B1(n5069), .B2(n5037), .A(n5036), .ZN(U3034) );
  INV_X1 U6190 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5041) );
  AOI22_X1 U6191 ( .A1(n6301), .A2(n6561), .B1(n6559), .B2(n5062), .ZN(n5038)
         );
  OAI21_X1 U6192 ( .B1(n6386), .B2(n5064), .A(n5038), .ZN(n5039) );
  AOI21_X1 U6193 ( .B1(n6466), .B2(n5066), .A(n5039), .ZN(n5040) );
  OAI21_X1 U6194 ( .B1(n5069), .B2(n5041), .A(n5040), .ZN(U3033) );
  INV_X1 U6195 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5045) );
  AOI22_X1 U6196 ( .A1(n6301), .A2(n6548), .B1(n6547), .B2(n5062), .ZN(n5042)
         );
  OAI21_X1 U6197 ( .B1(n6380), .B2(n5064), .A(n5042), .ZN(n5043) );
  AOI21_X1 U6198 ( .B1(n6458), .B2(n5066), .A(n5043), .ZN(n5044) );
  OAI21_X1 U6199 ( .B1(n5069), .B2(n5045), .A(n5044), .ZN(U3031) );
  INV_X1 U6200 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5049) );
  AOI22_X1 U6201 ( .A1(n6301), .A2(n6555), .B1(n6553), .B2(n5062), .ZN(n5046)
         );
  OAI21_X1 U6202 ( .B1(n6383), .B2(n5064), .A(n5046), .ZN(n5047) );
  AOI21_X1 U6203 ( .B1(n6462), .B2(n5066), .A(n5047), .ZN(n5048) );
  OAI21_X1 U6204 ( .B1(n5069), .B2(n5049), .A(n5048), .ZN(U3032) );
  INV_X1 U6205 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5053) );
  AOI22_X1 U6206 ( .A1(n6301), .A2(n6543), .B1(n6541), .B2(n5062), .ZN(n5050)
         );
  OAI21_X1 U6207 ( .B1(n6377), .B2(n5064), .A(n5050), .ZN(n5051) );
  AOI21_X1 U6208 ( .B1(n6454), .B2(n5066), .A(n5051), .ZN(n5052) );
  OAI21_X1 U6209 ( .B1(n5069), .B2(n5053), .A(n5052), .ZN(U3030) );
  INV_X1 U6210 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5057) );
  AOI22_X1 U6211 ( .A1(n6301), .A2(n6536), .B1(n6535), .B2(n5062), .ZN(n5054)
         );
  OAI21_X1 U6212 ( .B1(n6374), .B2(n5064), .A(n5054), .ZN(n5055) );
  AOI21_X1 U6213 ( .B1(n6450), .B2(n5066), .A(n5055), .ZN(n5056) );
  OAI21_X1 U6214 ( .B1(n5069), .B2(n5057), .A(n5056), .ZN(U3029) );
  INV_X1 U6215 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5061) );
  AOI22_X1 U6216 ( .A1(n6301), .A2(n6576), .B1(n6572), .B2(n5062), .ZN(n5058)
         );
  OAI21_X1 U6217 ( .B1(n6396), .B2(n5064), .A(n5058), .ZN(n5059) );
  AOI21_X1 U6218 ( .B1(n6476), .B2(n5066), .A(n5059), .ZN(n5060) );
  OAI21_X1 U6219 ( .B1(n5069), .B2(n5061), .A(n5060), .ZN(U3035) );
  INV_X1 U6220 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5068) );
  AOI22_X1 U6221 ( .A1(n6301), .A2(n6523), .B1(n6522), .B2(n5062), .ZN(n5063)
         );
  OAI21_X1 U6222 ( .B1(n6371), .B2(n5064), .A(n5063), .ZN(n5065) );
  AOI21_X1 U6223 ( .B1(n6437), .B2(n5066), .A(n5065), .ZN(n5067) );
  OAI21_X1 U6224 ( .B1(n5069), .B2(n5068), .A(n5067), .ZN(U3028) );
  OAI222_X1 U6225 ( .A1(n5330), .A2(n5591), .B1(n5071), .B2(n6117), .C1(n5592), 
        .C2(n5070), .ZN(U2853) );
  XOR2_X1 U6226 ( .A(n5072), .B(n5022), .Z(n5132) );
  INV_X1 U6227 ( .A(n5132), .ZN(n5299) );
  AOI21_X1 U6228 ( .B1(n5073), .B2(n4525), .A(n5123), .ZN(n6232) );
  AOI22_X1 U6229 ( .A1(n6113), .A2(n6232), .B1(n5588), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5074) );
  OAI21_X1 U6230 ( .B1(n5299), .B2(n5592), .A(n5074), .ZN(U2852) );
  NOR2_X1 U6231 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5075), .ZN(n5082)
         );
  INV_X1 U6232 ( .A(n5111), .ZN(n5077) );
  NOR3_X1 U6233 ( .A1(n5077), .A2(n5108), .A3(n6527), .ZN(n5078) );
  INV_X1 U6234 ( .A(n6280), .ZN(n6440) );
  INV_X1 U6235 ( .A(n6439), .ZN(n6435) );
  OAI21_X1 U6236 ( .B1(n5078), .B2(n6440), .A(n6435), .ZN(n5081) );
  OAI21_X1 U6237 ( .B1(n6278), .B2(n6695), .A(n5079), .ZN(n6442) );
  NOR3_X1 U6238 ( .A1(n6442), .A2(n6359), .A3(n6363), .ZN(n5080) );
  NAND2_X1 U6239 ( .A1(n5104), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5085)
         );
  NOR2_X1 U6240 ( .A1(n6354), .A2(n6527), .ZN(n5230) );
  NOR2_X1 U6241 ( .A1(n5182), .A2(n6359), .ZN(n5138) );
  AOI22_X1 U6242 ( .A1(n5230), .A2(n6439), .B1(n6355), .B2(n5138), .ZN(n5106)
         );
  INV_X1 U6243 ( .A(n5082), .ZN(n5105) );
  OAI22_X1 U6244 ( .A1(n6564), .A2(n5106), .B1(n6338), .B2(n5105), .ZN(n5083)
         );
  AOI21_X1 U6245 ( .B1(n6560), .B2(n5108), .A(n5083), .ZN(n5084) );
  OAI211_X1 U6246 ( .C1(n5111), .C2(n6469), .A(n5085), .B(n5084), .ZN(U3137)
         );
  NAND2_X1 U6247 ( .A1(n5104), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5088)
         );
  OAI22_X1 U6248 ( .A1(n6558), .A2(n5106), .B1(n6334), .B2(n5105), .ZN(n5086)
         );
  AOI21_X1 U6249 ( .B1(n6554), .B2(n5108), .A(n5086), .ZN(n5087) );
  OAI211_X1 U6250 ( .C1(n5111), .C2(n6465), .A(n5088), .B(n5087), .ZN(U3136)
         );
  NAND2_X1 U6251 ( .A1(n5104), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5091)
         );
  OAI22_X1 U6252 ( .A1(n6540), .A2(n5106), .B1(n6322), .B2(n5105), .ZN(n5089)
         );
  AOI21_X1 U6253 ( .B1(n6537), .B2(n5108), .A(n5089), .ZN(n5090) );
  OAI211_X1 U6254 ( .C1(n5111), .C2(n6453), .A(n5091), .B(n5090), .ZN(U3133)
         );
  NAND2_X1 U6255 ( .A1(n5104), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5094)
         );
  OAI22_X1 U6256 ( .A1(n6580), .A2(n5106), .B1(n6347), .B2(n5105), .ZN(n5092)
         );
  AOI21_X1 U6257 ( .B1(n6573), .B2(n5108), .A(n5092), .ZN(n5093) );
  OAI211_X1 U6258 ( .C1(n5111), .C2(n6482), .A(n5094), .B(n5093), .ZN(U3139)
         );
  NAND2_X1 U6259 ( .A1(n5104), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5097)
         );
  OAI22_X1 U6260 ( .A1(n6534), .A2(n5106), .B1(n6309), .B2(n5105), .ZN(n5095)
         );
  AOI21_X1 U6261 ( .B1(n6531), .B2(n5108), .A(n5095), .ZN(n5096) );
  OAI211_X1 U6262 ( .C1(n5111), .C2(n6449), .A(n5097), .B(n5096), .ZN(U3132)
         );
  NAND2_X1 U6263 ( .A1(n5104), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5100)
         );
  OAI22_X1 U6264 ( .A1(n6570), .A2(n5106), .B1(n6342), .B2(n5105), .ZN(n5098)
         );
  AOI21_X1 U6265 ( .B1(n6567), .B2(n5108), .A(n5098), .ZN(n5099) );
  OAI211_X1 U6266 ( .C1(n5111), .C2(n6473), .A(n5100), .B(n5099), .ZN(U3138)
         );
  NAND2_X1 U6267 ( .A1(n5104), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5103)
         );
  OAI22_X1 U6268 ( .A1(n6552), .A2(n5106), .B1(n6330), .B2(n5105), .ZN(n5101)
         );
  AOI21_X1 U6269 ( .B1(n6549), .B2(n5108), .A(n5101), .ZN(n5102) );
  OAI211_X1 U6270 ( .C1(n5111), .C2(n6461), .A(n5103), .B(n5102), .ZN(U3135)
         );
  NAND2_X1 U6271 ( .A1(n5104), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5110)
         );
  OAI22_X1 U6272 ( .A1(n6546), .A2(n5106), .B1(n6326), .B2(n5105), .ZN(n5107)
         );
  AOI21_X1 U6273 ( .B1(n6542), .B2(n5108), .A(n5107), .ZN(n5109) );
  OAI211_X1 U6274 ( .C1(n5111), .C2(n6457), .A(n5110), .B(n5109), .ZN(U3134)
         );
  OAI21_X1 U6275 ( .B1(n5114), .B2(n5113), .A(n5112), .ZN(n6243) );
  NAND2_X1 U6276 ( .A1(n6197), .A2(REIP_REG_5__SCAN_IN), .ZN(n6240) );
  OAI21_X1 U6277 ( .B1(n5686), .B2(n5276), .A(n6240), .ZN(n5116) );
  NOR2_X1 U6278 ( .A1(n5280), .A2(n5696), .ZN(n5115) );
  AOI211_X1 U6279 ( .C1(n6168), .C2(n5273), .A(n5116), .B(n5115), .ZN(n5117)
         );
  OAI21_X1 U6280 ( .B1(n6172), .B2(n6243), .A(n5117), .ZN(U2981) );
  INV_X1 U6281 ( .A(DATAI_7_), .ZN(n5119) );
  OAI222_X1 U6282 ( .A1(n6133), .A2(n5119), .B1(n6135), .B2(n5299), .C1(n5118), 
        .C2(n6134), .ZN(U2884) );
  OAI21_X1 U6283 ( .B1(n5120), .B2(n5122), .A(n5121), .ZN(n5310) );
  OR2_X1 U6284 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  NAND2_X1 U6285 ( .A1(n5125), .A2(n6051), .ZN(n6224) );
  INV_X1 U6286 ( .A(n6224), .ZN(n5282) );
  AOI22_X1 U6287 ( .A1(n6113), .A2(n5282), .B1(n5588), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5126) );
  OAI21_X1 U6288 ( .B1(n5310), .B2(n5592), .A(n5126), .ZN(U2851) );
  OAI21_X1 U6289 ( .B1(n5129), .B2(n5128), .A(n3104), .ZN(n6233) );
  NAND2_X1 U6290 ( .A1(n6197), .A2(REIP_REG_7__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U6291 ( .A1(n6188), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5130)
         );
  OAI211_X1 U6292 ( .C1(n6195), .C2(n5290), .A(n6230), .B(n5130), .ZN(n5131)
         );
  AOI21_X1 U6293 ( .B1(n5132), .B2(n3103), .A(n5131), .ZN(n5133) );
  OAI21_X1 U6294 ( .B1(n6233), .B2(n6172), .A(n5133), .ZN(U2979) );
  INV_X1 U6295 ( .A(DATAI_8_), .ZN(n5134) );
  OAI222_X1 U6296 ( .A1(n5310), .A2(n6135), .B1(n6134), .B2(n5135), .C1(n6133), 
        .C2(n5134), .ZN(U2883) );
  NAND2_X1 U6297 ( .A1(n5139), .A2(n6409), .ZN(n5137) );
  OAI21_X1 U6298 ( .B1(n5137), .B2(n6574), .A(n6280), .ZN(n5141) );
  NOR2_X1 U6299 ( .A1(n4761), .A2(n5852), .ZN(n6277) );
  AND2_X1 U6300 ( .A1(n6277), .A2(n3118), .ZN(n6517) );
  NAND3_X1 U6301 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6279), .ZN(n6526) );
  NOR2_X1 U6302 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6526), .ZN(n5143)
         );
  INV_X1 U6303 ( .A(n5143), .ZN(n5175) );
  INV_X1 U6304 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5145) );
  NOR2_X1 U6305 ( .A1(n6355), .A2(n6442), .ZN(n6283) );
  INV_X1 U6306 ( .A(n6517), .ZN(n5140) );
  AOI22_X1 U6307 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6359), .B1(n5141), .B2(
        n5140), .ZN(n5142) );
  OAI211_X1 U6308 ( .C1(n5143), .C2(n6665), .A(n6283), .B(n5142), .ZN(n5144)
         );
  OAI22_X1 U6309 ( .A1(n6334), .A2(n5175), .B1(n5145), .B2(n5173), .ZN(n5146)
         );
  AOI21_X1 U6310 ( .B1(n5177), .B2(n6554), .A(n5146), .ZN(n5148) );
  NAND2_X1 U6311 ( .A1(n6574), .A2(n6555), .ZN(n5147) );
  OAI211_X1 U6312 ( .C1(n5180), .C2(n6558), .A(n5148), .B(n5147), .ZN(U3104)
         );
  INV_X1 U6313 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5149) );
  OAI22_X1 U6314 ( .A1(n6326), .A2(n5175), .B1(n5149), .B2(n5173), .ZN(n5150)
         );
  AOI21_X1 U6315 ( .B1(n5177), .B2(n6542), .A(n5150), .ZN(n5152) );
  NAND2_X1 U6316 ( .A1(n6574), .A2(n6543), .ZN(n5151) );
  OAI211_X1 U6317 ( .C1(n5180), .C2(n6546), .A(n5152), .B(n5151), .ZN(U3102)
         );
  INV_X1 U6318 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5153) );
  OAI22_X1 U6319 ( .A1(n6338), .A2(n5175), .B1(n5153), .B2(n5173), .ZN(n5154)
         );
  AOI21_X1 U6320 ( .B1(n5177), .B2(n6560), .A(n5154), .ZN(n5156) );
  NAND2_X1 U6321 ( .A1(n6574), .A2(n6561), .ZN(n5155) );
  OAI211_X1 U6322 ( .C1(n5180), .C2(n6564), .A(n5156), .B(n5155), .ZN(U3105)
         );
  INV_X1 U6323 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5157) );
  OAI22_X1 U6324 ( .A1(n6342), .A2(n5175), .B1(n5157), .B2(n5173), .ZN(n5158)
         );
  AOI21_X1 U6325 ( .B1(n5177), .B2(n6567), .A(n5158), .ZN(n5160) );
  NAND2_X1 U6326 ( .A1(n6574), .A2(n6566), .ZN(n5159) );
  OAI211_X1 U6327 ( .C1(n5180), .C2(n6570), .A(n5160), .B(n5159), .ZN(U3106)
         );
  INV_X1 U6328 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5161) );
  OAI22_X1 U6329 ( .A1(n6322), .A2(n5175), .B1(n5161), .B2(n5173), .ZN(n5162)
         );
  AOI21_X1 U6330 ( .B1(n5177), .B2(n6537), .A(n5162), .ZN(n5164) );
  NAND2_X1 U6331 ( .A1(n6574), .A2(n6536), .ZN(n5163) );
  OAI211_X1 U6332 ( .C1(n5180), .C2(n6540), .A(n5164), .B(n5163), .ZN(U3101)
         );
  INV_X1 U6333 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5165) );
  OAI22_X1 U6334 ( .A1(n6330), .A2(n5175), .B1(n5165), .B2(n5173), .ZN(n5166)
         );
  AOI21_X1 U6335 ( .B1(n5177), .B2(n6549), .A(n5166), .ZN(n5168) );
  NAND2_X1 U6336 ( .A1(n6574), .A2(n6548), .ZN(n5167) );
  OAI211_X1 U6337 ( .C1(n5180), .C2(n6552), .A(n5168), .B(n5167), .ZN(U3103)
         );
  INV_X1 U6338 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5169) );
  OAI22_X1 U6339 ( .A1(n6347), .A2(n5175), .B1(n5169), .B2(n5173), .ZN(n5170)
         );
  AOI21_X1 U6340 ( .B1(n5177), .B2(n6573), .A(n5170), .ZN(n5172) );
  NAND2_X1 U6341 ( .A1(n6574), .A2(n6576), .ZN(n5171) );
  OAI211_X1 U6342 ( .C1(n5180), .C2(n6580), .A(n5172), .B(n5171), .ZN(U3107)
         );
  INV_X1 U6343 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5174) );
  OAI22_X1 U6344 ( .A1(n6309), .A2(n5175), .B1(n5174), .B2(n5173), .ZN(n5176)
         );
  AOI21_X1 U6345 ( .B1(n5177), .B2(n6531), .A(n5176), .ZN(n5179) );
  NAND2_X1 U6346 ( .A1(n6574), .A2(n6523), .ZN(n5178) );
  OAI211_X1 U6347 ( .C1(n5180), .C2(n6534), .A(n5179), .B(n5178), .ZN(U3100)
         );
  INV_X1 U6348 ( .A(n6516), .ZN(n5855) );
  NAND2_X1 U6349 ( .A1(n5183), .A2(n5182), .ZN(n5191) );
  AOI21_X1 U6350 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5191), .A(n5184), .ZN(
        n5227) );
  NAND2_X1 U6351 ( .A1(n6398), .A2(n5185), .ZN(n5214) );
  INV_X1 U6352 ( .A(n5217), .ZN(n5186) );
  NAND3_X1 U6353 ( .A1(n5220), .A2(n6409), .A3(n5186), .ZN(n5188) );
  AOI22_X1 U6354 ( .A1(n5188), .A2(n6280), .B1(n6362), .B2(n5187), .ZN(n5189)
         );
  AOI211_X1 U6355 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5214), .A(n6363), .B(
        n5189), .ZN(n5190) );
  NAND2_X1 U6356 ( .A1(n5227), .A2(n5190), .ZN(n5213) );
  NAND2_X1 U6357 ( .A1(n5213), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5194)
         );
  INV_X1 U6358 ( .A(n5191), .ZN(n5228) );
  AOI22_X1 U6359 ( .A1(n5230), .A2(n6362), .B1(n5228), .B2(n6355), .ZN(n5215)
         );
  OAI22_X1 U6360 ( .A1(n6534), .A2(n5215), .B1(n6309), .B2(n5214), .ZN(n5192)
         );
  AOI21_X1 U6361 ( .B1(n6523), .B2(n5217), .A(n5192), .ZN(n5193) );
  OAI211_X1 U6362 ( .C1(n6371), .C2(n5220), .A(n5194), .B(n5193), .ZN(U3116)
         );
  NAND2_X1 U6363 ( .A1(n5213), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5197)
         );
  OAI22_X1 U6364 ( .A1(n6540), .A2(n5215), .B1(n6322), .B2(n5214), .ZN(n5195)
         );
  AOI21_X1 U6365 ( .B1(n6536), .B2(n5217), .A(n5195), .ZN(n5196) );
  OAI211_X1 U6366 ( .C1(n5220), .C2(n6374), .A(n5197), .B(n5196), .ZN(U3117)
         );
  NAND2_X1 U6367 ( .A1(n5213), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5200)
         );
  OAI22_X1 U6368 ( .A1(n6546), .A2(n5215), .B1(n6326), .B2(n5214), .ZN(n5198)
         );
  AOI21_X1 U6369 ( .B1(n6543), .B2(n5217), .A(n5198), .ZN(n5199) );
  OAI211_X1 U6370 ( .C1(n5220), .C2(n6377), .A(n5200), .B(n5199), .ZN(U3118)
         );
  NAND2_X1 U6371 ( .A1(n5213), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5203)
         );
  OAI22_X1 U6372 ( .A1(n6580), .A2(n5215), .B1(n6347), .B2(n5214), .ZN(n5201)
         );
  AOI21_X1 U6373 ( .B1(n6576), .B2(n5217), .A(n5201), .ZN(n5202) );
  OAI211_X1 U6374 ( .C1(n5220), .C2(n6396), .A(n5203), .B(n5202), .ZN(U3123)
         );
  NAND2_X1 U6375 ( .A1(n5213), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5206)
         );
  OAI22_X1 U6376 ( .A1(n6570), .A2(n5215), .B1(n6342), .B2(n5214), .ZN(n5204)
         );
  AOI21_X1 U6377 ( .B1(n6566), .B2(n5217), .A(n5204), .ZN(n5205) );
  OAI211_X1 U6378 ( .C1(n5220), .C2(n6389), .A(n5206), .B(n5205), .ZN(U3122)
         );
  NAND2_X1 U6379 ( .A1(n5213), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5209)
         );
  OAI22_X1 U6380 ( .A1(n6564), .A2(n5215), .B1(n6338), .B2(n5214), .ZN(n5207)
         );
  AOI21_X1 U6381 ( .B1(n6561), .B2(n5217), .A(n5207), .ZN(n5208) );
  OAI211_X1 U6382 ( .C1(n5220), .C2(n6386), .A(n5209), .B(n5208), .ZN(U3121)
         );
  NAND2_X1 U6383 ( .A1(n5213), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5212)
         );
  OAI22_X1 U6384 ( .A1(n6552), .A2(n5215), .B1(n6330), .B2(n5214), .ZN(n5210)
         );
  AOI21_X1 U6385 ( .B1(n6548), .B2(n5217), .A(n5210), .ZN(n5211) );
  OAI211_X1 U6386 ( .C1(n5220), .C2(n6380), .A(n5212), .B(n5211), .ZN(U3119)
         );
  NAND2_X1 U6387 ( .A1(n5213), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5219)
         );
  OAI22_X1 U6388 ( .A1(n6558), .A2(n5215), .B1(n6334), .B2(n5214), .ZN(n5216)
         );
  AOI21_X1 U6389 ( .B1(n6555), .B2(n5217), .A(n5216), .ZN(n5218) );
  OAI211_X1 U6390 ( .C1(n5220), .C2(n6383), .A(n5219), .B(n5218), .ZN(U3120)
         );
  OR2_X1 U6391 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5221), .ZN(n5253)
         );
  INV_X1 U6392 ( .A(n6509), .ZN(n5223) );
  AOI21_X1 U6393 ( .B1(n5223), .B2(n5258), .A(n6703), .ZN(n5224) );
  AOI211_X1 U6394 ( .C1(n5229), .C2(n3118), .A(n6527), .B(n5224), .ZN(n5225)
         );
  AOI211_X1 U6395 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5253), .A(n6355), .B(
        n5225), .ZN(n5226) );
  NAND2_X1 U6396 ( .A1(n5227), .A2(n5226), .ZN(n5252) );
  NAND2_X1 U6397 ( .A1(n5252), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5233) );
  AOI22_X1 U6398 ( .A1(n5230), .A2(n5229), .B1(n6363), .B2(n5228), .ZN(n5254)
         );
  OAI22_X1 U6399 ( .A1(n6552), .A2(n5254), .B1(n5253), .B2(n6330), .ZN(n5231)
         );
  AOI21_X1 U6400 ( .B1(n6509), .B2(n6549), .A(n5231), .ZN(n5232) );
  OAI211_X1 U6401 ( .C1(n5258), .C2(n6461), .A(n5233), .B(n5232), .ZN(U3087)
         );
  NAND2_X1 U6402 ( .A1(n5252), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5236) );
  OAI22_X1 U6403 ( .A1(n6558), .A2(n5254), .B1(n5253), .B2(n6334), .ZN(n5234)
         );
  AOI21_X1 U6404 ( .B1(n6509), .B2(n6554), .A(n5234), .ZN(n5235) );
  OAI211_X1 U6405 ( .C1(n5258), .C2(n6465), .A(n5236), .B(n5235), .ZN(U3088)
         );
  NAND2_X1 U6406 ( .A1(n5252), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5239) );
  OAI22_X1 U6407 ( .A1(n6570), .A2(n5254), .B1(n5253), .B2(n6342), .ZN(n5237)
         );
  AOI21_X1 U6408 ( .B1(n6509), .B2(n6567), .A(n5237), .ZN(n5238) );
  OAI211_X1 U6409 ( .C1(n5258), .C2(n6473), .A(n5239), .B(n5238), .ZN(U3090)
         );
  NAND2_X1 U6410 ( .A1(n5252), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5242) );
  OAI22_X1 U6411 ( .A1(n6580), .A2(n5254), .B1(n5253), .B2(n6347), .ZN(n5240)
         );
  AOI21_X1 U6412 ( .B1(n6509), .B2(n6573), .A(n5240), .ZN(n5241) );
  OAI211_X1 U6413 ( .C1(n5258), .C2(n6482), .A(n5242), .B(n5241), .ZN(U3091)
         );
  NAND2_X1 U6414 ( .A1(n5252), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5245) );
  OAI22_X1 U6415 ( .A1(n6546), .A2(n5254), .B1(n5253), .B2(n6326), .ZN(n5243)
         );
  AOI21_X1 U6416 ( .B1(n6509), .B2(n6542), .A(n5243), .ZN(n5244) );
  OAI211_X1 U6417 ( .C1(n5258), .C2(n6457), .A(n5245), .B(n5244), .ZN(U3086)
         );
  NAND2_X1 U6418 ( .A1(n5252), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5248) );
  OAI22_X1 U6419 ( .A1(n6564), .A2(n5254), .B1(n5253), .B2(n6338), .ZN(n5246)
         );
  AOI21_X1 U6420 ( .B1(n6509), .B2(n6560), .A(n5246), .ZN(n5247) );
  OAI211_X1 U6421 ( .C1(n5258), .C2(n6469), .A(n5248), .B(n5247), .ZN(U3089)
         );
  NAND2_X1 U6422 ( .A1(n5252), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5251) );
  OAI22_X1 U6423 ( .A1(n6540), .A2(n5254), .B1(n5253), .B2(n6322), .ZN(n5249)
         );
  AOI21_X1 U6424 ( .B1(n6509), .B2(n6537), .A(n5249), .ZN(n5250) );
  OAI211_X1 U6425 ( .C1(n5258), .C2(n6453), .A(n5251), .B(n5250), .ZN(U3085)
         );
  NAND2_X1 U6426 ( .A1(n5252), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5257) );
  OAI22_X1 U6427 ( .A1(n6534), .A2(n5254), .B1(n6309), .B2(n5253), .ZN(n5255)
         );
  AOI21_X1 U6428 ( .B1(n6531), .B2(n6509), .A(n5255), .ZN(n5256) );
  OAI211_X1 U6429 ( .C1(n6449), .C2(n5258), .A(n5257), .B(n5256), .ZN(U3084)
         );
  INV_X1 U6430 ( .A(n3671), .ZN(n5259) );
  NAND2_X1 U6431 ( .A1(n5262), .A2(n5259), .ZN(n5260) );
  NAND2_X1 U6432 ( .A1(n6086), .A2(REIP_REG_0__SCAN_IN), .ZN(n5266) );
  AOI22_X1 U6433 ( .A1(n6092), .A2(n5261), .B1(n6090), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5265) );
  AND2_X1 U6434 ( .A1(n5262), .A2(n6688), .ZN(n6095) );
  NAND2_X1 U6435 ( .A1(n6095), .A2(n3130), .ZN(n5264) );
  OAI21_X1 U6436 ( .B1(n6094), .B2(n6071), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5263) );
  AND4_X1 U6437 ( .A1(n5266), .A2(n5265), .A3(n5264), .A4(n5263), .ZN(n5267)
         );
  OAI21_X1 U6438 ( .B1(n6064), .B2(n6136), .A(n5267), .ZN(U2827) );
  INV_X1 U6439 ( .A(n5121), .ZN(n5269) );
  OAI21_X1 U6440 ( .B1(n5269), .B2(n3239), .A(n3147), .ZN(n6054) );
  AOI22_X1 U6441 ( .A1(n5613), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6128), .ZN(n5270) );
  OAI21_X1 U6442 ( .B1(n6054), .B2(n6135), .A(n5270), .ZN(U2882) );
  INV_X1 U6443 ( .A(n5351), .ZN(n5271) );
  NAND2_X1 U6444 ( .A1(n6063), .A2(n5271), .ZN(n5352) );
  OAI21_X1 U6445 ( .B1(n6613), .B2(n5352), .A(n6615), .ZN(n5278) );
  OAI21_X1 U6446 ( .B1(n6083), .B2(n5328), .A(n6084), .ZN(n5324) );
  AOI22_X1 U6447 ( .A1(n6092), .A2(n6242), .B1(n6090), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n5275) );
  NAND2_X1 U6448 ( .A1(n6084), .A2(n5272), .ZN(n6027) );
  AOI21_X1 U6449 ( .B1(n6071), .B2(n5273), .A(n6053), .ZN(n5274) );
  OAI211_X1 U6450 ( .C1(n5276), .C2(n6019), .A(n5275), .B(n5274), .ZN(n5277)
         );
  AOI21_X1 U6451 ( .B1(n5278), .B2(n5324), .A(n5277), .ZN(n5279) );
  OAI21_X1 U6452 ( .B1(n6064), .B2(n5280), .A(n5279), .ZN(U2822) );
  OR2_X1 U6453 ( .A1(n6083), .A2(n5281), .ZN(n5286) );
  NAND2_X1 U6454 ( .A1(n5286), .A2(n6084), .ZN(n5334) );
  INV_X1 U6455 ( .A(n5313), .ZN(n5285) );
  AOI22_X1 U6456 ( .A1(n6092), .A2(n5282), .B1(n6090), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5284) );
  AOI21_X1 U6457 ( .B1(n6094), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6053), 
        .ZN(n5283) );
  OAI211_X1 U6458 ( .C1(n5285), .C2(n6104), .A(n5284), .B(n5283), .ZN(n5288)
         );
  NOR3_X1 U6459 ( .A1(n5286), .A2(n5337), .A3(n5336), .ZN(n5287) );
  AOI211_X1 U6460 ( .C1(REIP_REG_8__SCAN_IN), .C2(n5334), .A(n5288), .B(n5287), 
        .ZN(n5289) );
  OAI21_X1 U6461 ( .B1(n5310), .B2(n5873), .A(n5289), .ZN(U2819) );
  OAI22_X1 U6462 ( .A1(n5291), .A2(n6019), .B1(n6104), .B2(n5290), .ZN(n5295)
         );
  NOR3_X1 U6463 ( .A1(n5336), .A2(REIP_REG_7__SCAN_IN), .A3(n6083), .ZN(n5292)
         );
  AOI21_X1 U6464 ( .B1(n6232), .B2(n6092), .A(n5292), .ZN(n5293) );
  OAI21_X1 U6465 ( .B1(n6932), .B2(n6080), .A(n5293), .ZN(n5294) );
  NOR3_X1 U6466 ( .A1(n5295), .A2(n6053), .A3(n5294), .ZN(n5298) );
  NOR2_X1 U6467 ( .A1(n6083), .A2(REIP_REG_6__SCAN_IN), .ZN(n5296) );
  OAI21_X1 U6468 ( .B1(n5324), .B2(n5296), .A(REIP_REG_7__SCAN_IN), .ZN(n5297)
         );
  OAI211_X1 U6469 ( .C1(n5299), .C2(n5873), .A(n5298), .B(n5297), .ZN(U2820)
         );
  AOI21_X1 U6470 ( .B1(n5301), .B2(n3147), .A(n5300), .ZN(n5302) );
  INV_X1 U6471 ( .A(n5302), .ZN(n5365) );
  XNOR2_X1 U6472 ( .A(n5303), .B(n6050), .ZN(n5340) );
  INV_X1 U6473 ( .A(n5340), .ZN(n6207) );
  AOI22_X1 U6474 ( .A1(n6113), .A2(n6207), .B1(n5588), .B2(EBX_REG_10__SCAN_IN), .ZN(n5304) );
  OAI21_X1 U6475 ( .B1(n5365), .B2(n5592), .A(n5304), .ZN(U2849) );
  INV_X1 U6476 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5306) );
  INV_X1 U6477 ( .A(DATAI_10_), .ZN(n5305) );
  OAI222_X1 U6478 ( .A1(n5365), .A2(n6135), .B1(n6134), .B2(n5306), .C1(n5305), 
        .C2(n6133), .ZN(U2881) );
  OAI21_X1 U6479 ( .B1(n3108), .B2(n5308), .A(n5307), .ZN(n6222) );
  OAI22_X1 U6480 ( .A1(n5686), .A2(n6782), .B1(n6253), .B2(n6619), .ZN(n5312)
         );
  NOR2_X1 U6481 ( .A1(n5310), .A2(n5696), .ZN(n5311) );
  AOI211_X1 U6482 ( .C1(n6168), .C2(n5313), .A(n5312), .B(n5311), .ZN(n5314)
         );
  OAI21_X1 U6483 ( .B1(n6172), .B2(n6222), .A(n5314), .ZN(U2978) );
  NAND2_X1 U6484 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  XNOR2_X1 U6485 ( .A(n5318), .B(n5317), .ZN(n6218) );
  NAND2_X1 U6486 ( .A1(n6218), .A2(n6191), .ZN(n5322) );
  INV_X1 U6487 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6488 ( .A1(n6197), .A2(REIP_REG_9__SCAN_IN), .ZN(n6214) );
  OAI21_X1 U6489 ( .B1(n5686), .B2(n5319), .A(n6214), .ZN(n5320) );
  AOI21_X1 U6490 ( .B1(n6168), .B2(n6055), .A(n5320), .ZN(n5321) );
  OAI211_X1 U6491 ( .C1(n5696), .C2(n6054), .A(n5322), .B(n5321), .ZN(U2977)
         );
  INV_X1 U6492 ( .A(n6178), .ZN(n5323) );
  NAND2_X1 U6493 ( .A1(n6071), .A2(n5323), .ZN(n5327) );
  NAND2_X1 U6494 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5326)
         );
  AOI22_X1 U6495 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6090), .B1(
        REIP_REG_6__SCAN_IN), .B2(n5324), .ZN(n5325) );
  NAND4_X1 U6496 ( .A1(n5327), .A2(n5326), .A3(n5325), .A4(n6027), .ZN(n5332)
         );
  NAND3_X1 U6497 ( .A1(n6063), .A2(n5328), .A3(n4527), .ZN(n5329) );
  OAI21_X1 U6498 ( .B1(n5330), .B2(n5871), .A(n5329), .ZN(n5331) );
  AOI211_X1 U6499 ( .C1(n6174), .C2(n6056), .A(n5332), .B(n5331), .ZN(n5333)
         );
  INV_X1 U6500 ( .A(n5333), .ZN(U2821) );
  INV_X1 U6501 ( .A(n5334), .ZN(n5335) );
  OAI21_X1 U6502 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6083), .A(n5335), .ZN(n6057)
         );
  AOI22_X1 U6503 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6090), .B1(
        REIP_REG_10__SCAN_IN), .B2(n6057), .ZN(n5344) );
  NOR4_X1 U6504 ( .A1(n6083), .A2(n5337), .A3(n6619), .A4(n5336), .ZN(n6058)
         );
  INV_X1 U6505 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6621) );
  NOR2_X1 U6506 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6621), .ZN(n5342) );
  NOR2_X1 U6507 ( .A1(n6019), .A2(n5360), .ZN(n5338) );
  AOI211_X1 U6508 ( .C1(n6071), .C2(n5362), .A(n6053), .B(n5338), .ZN(n5339)
         );
  OAI21_X1 U6509 ( .B1(n5340), .B2(n5871), .A(n5339), .ZN(n5341) );
  AOI21_X1 U6510 ( .B1(n6058), .B2(n5342), .A(n5341), .ZN(n5343) );
  OAI211_X1 U6511 ( .C1(n5365), .C2(n5873), .A(n5344), .B(n5343), .ZN(U2817)
         );
  NOR2_X1 U6512 ( .A1(n5300), .A2(n5345), .ZN(n5346) );
  OR2_X1 U6513 ( .A1(n5367), .A2(n5346), .ZN(n6046) );
  AOI22_X1 U6514 ( .A1(n5613), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6128), .ZN(n5347) );
  OAI21_X1 U6515 ( .B1(n6046), .B2(n6135), .A(n5347), .ZN(U2880) );
  INV_X1 U6516 ( .A(n5962), .ZN(n5355) );
  INV_X1 U6517 ( .A(n6187), .ZN(n5348) );
  AOI22_X1 U6518 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n6094), .B1(n6071), 
        .B2(n5348), .ZN(n5350) );
  NAND2_X1 U6519 ( .A1(n6090), .A2(EBX_REG_4__SCAN_IN), .ZN(n5349) );
  OAI211_X1 U6520 ( .C1(n6254), .C2(n5871), .A(n5350), .B(n5349), .ZN(n5354)
         );
  INV_X1 U6521 ( .A(n6084), .ZN(n6093) );
  OAI21_X1 U6522 ( .B1(n6093), .B2(n5351), .A(n6086), .ZN(n6075) );
  OAI221_X1 U6523 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5352), .C1(n6613), .C2(
        n6075), .A(n6027), .ZN(n5353) );
  AOI211_X1 U6524 ( .C1(n6095), .C2(n5355), .A(n5354), .B(n5353), .ZN(n5356)
         );
  OAI21_X1 U6525 ( .B1(n6064), .B2(n6183), .A(n5356), .ZN(U2823) );
  NAND2_X1 U6526 ( .A1(n6162), .A2(n5358), .ZN(n5359) );
  XNOR2_X1 U6527 ( .A(n5357), .B(n5359), .ZN(n6210) );
  NAND2_X1 U6528 ( .A1(n6210), .A2(n6191), .ZN(n5364) );
  NAND2_X1 U6529 ( .A1(n6197), .A2(REIP_REG_10__SCAN_IN), .ZN(n6205) );
  OAI21_X1 U6530 ( .B1(n5686), .B2(n5360), .A(n6205), .ZN(n5361) );
  AOI21_X1 U6531 ( .B1(n6168), .B2(n5362), .A(n5361), .ZN(n5363) );
  OAI211_X1 U6532 ( .C1(n5696), .C2(n5365), .A(n5364), .B(n5363), .ZN(U2976)
         );
  XNOR2_X1 U6533 ( .A(n5367), .B(n5366), .ZN(n5410) );
  OR2_X1 U6534 ( .A1(n5369), .A2(n5368), .ZN(n5370) );
  NAND2_X1 U6535 ( .A1(n5370), .A2(n5948), .ZN(n5398) );
  INV_X1 U6536 ( .A(n5398), .ZN(n5371) );
  AOI22_X1 U6537 ( .A1(n6113), .A2(n5371), .B1(n5588), .B2(EBX_REG_12__SCAN_IN), .ZN(n5372) );
  OAI21_X1 U6538 ( .B1(n5410), .B2(n5592), .A(n5372), .ZN(U2847) );
  INV_X1 U6539 ( .A(n5375), .ZN(n5374) );
  INV_X1 U6540 ( .A(n6086), .ZN(n5373) );
  AOI21_X1 U6541 ( .B1(n6084), .B2(n5374), .A(n5373), .ZN(n6043) );
  NOR3_X1 U6542 ( .A1(n6083), .A2(REIP_REG_12__SCAN_IN), .A3(n5375), .ZN(n6037) );
  INV_X1 U6543 ( .A(n6037), .ZN(n5380) );
  OAI22_X1 U6544 ( .A1(n5403), .A2(n6104), .B1(n6019), .B2(n5405), .ZN(n5378)
         );
  NOR2_X1 U6545 ( .A1(n5376), .A2(n6080), .ZN(n5377) );
  NOR3_X1 U6546 ( .A1(n5378), .A2(n6053), .A3(n5377), .ZN(n5379) );
  OAI211_X1 U6547 ( .C1(n5398), .C2(n5871), .A(n5380), .B(n5379), .ZN(n5381)
         );
  AOI21_X1 U6548 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6043), .A(n5381), .ZN(n5382) );
  OAI21_X1 U6549 ( .B1(n5410), .B2(n5873), .A(n5382), .ZN(U2815) );
  INV_X1 U6550 ( .A(DATAI_12_), .ZN(n5384) );
  OAI222_X1 U6551 ( .A1(n6133), .A2(n5384), .B1(n6135), .B2(n5410), .C1(n5383), 
        .C2(n6134), .ZN(U2879) );
  NAND2_X1 U6552 ( .A1(n3252), .A2(n5386), .ZN(n5387) );
  XNOR2_X1 U6553 ( .A(n5385), .B(n5387), .ZN(n5402) );
  NOR2_X1 U6554 ( .A1(n5937), .A2(n3649), .ZN(n5397) );
  INV_X1 U6555 ( .A(n5388), .ZN(n5390) );
  NOR2_X1 U6556 ( .A1(n5390), .A2(n5389), .ZN(n5392) );
  AOI211_X1 U6557 ( .C1(n6252), .C2(n6204), .A(n5392), .B(n5391), .ZN(n6238)
         );
  OAI21_X1 U6558 ( .B1(n5393), .B2(n6209), .A(n6238), .ZN(n6200) );
  AOI221_X1 U6559 ( .B1(n6252), .B2(n3649), .C1(n5394), .C2(n3649), .A(n6200), 
        .ZN(n5395) );
  INV_X1 U6560 ( .A(n5395), .ZN(n5396) );
  MUX2_X1 U6561 ( .A(n5397), .B(n5396), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n5400) );
  NAND2_X1 U6562 ( .A1(n6197), .A2(REIP_REG_12__SCAN_IN), .ZN(n5404) );
  OAI21_X1 U6563 ( .B1(n6255), .B2(n5398), .A(n5404), .ZN(n5399) );
  AOI211_X1 U6564 ( .C1(n5402), .C2(n6269), .A(n5400), .B(n5399), .ZN(n5401)
         );
  INV_X1 U6565 ( .A(n5401), .ZN(U3006) );
  NAND2_X1 U6566 ( .A1(n5402), .A2(n6191), .ZN(n5409) );
  INV_X1 U6567 ( .A(n5403), .ZN(n5407) );
  OAI21_X1 U6568 ( .B1(n5686), .B2(n5405), .A(n5404), .ZN(n5406) );
  AOI21_X1 U6569 ( .B1(n6168), .B2(n5407), .A(n5406), .ZN(n5408) );
  OAI211_X1 U6570 ( .C1(n5410), .C2(n5696), .A(n5409), .B(n5408), .ZN(U2974)
         );
  XNOR2_X1 U6571 ( .A(n6164), .B(n5421), .ZN(n5411) );
  XNOR2_X1 U6572 ( .A(n5412), .B(n5411), .ZN(n5703) );
  OAI22_X1 U6573 ( .A1(n5414), .A2(n5413), .B1(n5422), .B2(n5952), .ZN(n5415)
         );
  NOR2_X1 U6574 ( .A1(n6200), .A2(n5415), .ZN(n5954) );
  NOR3_X1 U6575 ( .A1(n5417), .A2(n5416), .A3(n5944), .ZN(n5419) );
  NOR2_X1 U6576 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5418), .ZN(n5946)
         );
  OAI21_X1 U6577 ( .B1(n5420), .B2(n5419), .A(n5946), .ZN(n5958) );
  INV_X1 U6578 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5421) );
  AOI21_X1 U6579 ( .B1(n5954), .B2(n5958), .A(n5421), .ZN(n5426) );
  INV_X1 U6580 ( .A(n5937), .ZN(n6199) );
  AND3_X1 U6581 ( .A1(n5422), .A2(n5421), .A3(n6199), .ZN(n5425) );
  XNOR2_X1 U6582 ( .A(n5423), .B(n5947), .ZN(n6014) );
  OAI22_X1 U6583 ( .A1(n6255), .A2(n6014), .B1(n6628), .B2(n6253), .ZN(n5424)
         );
  NOR3_X1 U6584 ( .A1(n5426), .A2(n5425), .A3(n5424), .ZN(n5427) );
  OAI21_X1 U6585 ( .B1(n5703), .B2(n6223), .A(n5427), .ZN(U3004) );
  NAND2_X1 U6586 ( .A1(n5429), .A2(n5430), .ZN(n5431) );
  INV_X1 U6587 ( .A(n6108), .ZN(n5433) );
  AOI22_X1 U6588 ( .A1(n5613), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n6128), .ZN(n5432) );
  OAI21_X1 U6589 ( .B1(n5433), .B2(n6135), .A(n5432), .ZN(U2878) );
  INV_X1 U6590 ( .A(n5434), .ZN(n5447) );
  NOR2_X2 U6591 ( .A1(n6128), .A2(n5435), .ZN(n6125) );
  AOI22_X1 U6592 ( .A1(n6125), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6128), .ZN(n5438) );
  NOR3_X1 U6593 ( .A1(n6128), .A2(n5593), .A3(n3119), .ZN(n5436) );
  NAND2_X1 U6594 ( .A1(n6129), .A2(DATAI_13_), .ZN(n5437) );
  OAI211_X1 U6595 ( .C1(n5447), .C2(n6135), .A(n5438), .B(n5437), .ZN(U2862)
         );
  INV_X1 U6596 ( .A(n5439), .ZN(n5440) );
  AOI22_X1 U6597 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6094), .B1(n6071), 
        .B2(n5440), .ZN(n5442) );
  NAND2_X1 U6598 ( .A1(n6090), .A2(EBX_REG_29__SCAN_IN), .ZN(n5441) );
  OAI211_X1 U6599 ( .C1(n5731), .C2(n5871), .A(n5442), .B(n5441), .ZN(n5443)
         );
  NOR2_X1 U6600 ( .A1(n5444), .A2(n5443), .ZN(n5446) );
  NAND2_X1 U6601 ( .A1(n5474), .A2(REIP_REG_29__SCAN_IN), .ZN(n5445) );
  OAI211_X1 U6602 ( .C1(n5447), .C2(n5873), .A(n5446), .B(n5445), .ZN(U2798)
         );
  AOI22_X1 U6603 ( .A1(n6125), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6128), .ZN(n5449) );
  NAND2_X1 U6604 ( .A1(n6129), .A2(DATAI_14_), .ZN(n5448) );
  OAI211_X1 U6605 ( .C1(n5450), .C2(n6135), .A(n5449), .B(n5448), .ZN(U2861)
         );
  INV_X1 U6606 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6754) );
  OAI222_X1 U6607 ( .A1(n5592), .A2(n5450), .B1(n5591), .B2(n5722), .C1(n6754), 
        .C2(n6117), .ZN(U2829) );
  OAI21_X1 U6608 ( .B1(n5451), .B2(n5454), .A(n5453), .ZN(n5698) );
  AOI22_X1 U6609 ( .A1(n5613), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6128), .ZN(n5455) );
  OAI21_X1 U6610 ( .B1(n5698), .B2(n6135), .A(n5455), .ZN(U2877) );
  AOI21_X1 U6611 ( .B1(n5458), .B2(n5456), .A(n5465), .ZN(n5466) );
  INV_X1 U6612 ( .A(n5457), .ZN(n5461) );
  NAND3_X1 U6613 ( .A1(n5458), .A2(n4582), .A3(n3194), .ZN(n5459) );
  OAI21_X1 U6614 ( .B1(n5461), .B2(n5460), .A(n5459), .ZN(n5462) );
  AOI21_X1 U6615 ( .B1(n5463), .B2(n6667), .A(n5462), .ZN(n5464) );
  OAI22_X1 U6616 ( .A1(n5466), .A2(n3194), .B1(n5465), .B2(n5464), .ZN(U3459)
         );
  OAI22_X1 U6617 ( .A1(n5468), .A2(n5591), .B1(n5467), .B2(n6117), .ZN(U2828)
         );
  NAND2_X1 U6618 ( .A1(n3143), .A2(n5469), .ZN(n5470) );
  NAND2_X1 U6619 ( .A1(n5471), .A2(n5470), .ZN(n5739) );
  AOI22_X1 U6620 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6094), .B1(n6071), 
        .B2(n5472), .ZN(n5473) );
  OAI21_X1 U6621 ( .B1(n5739), .B2(n5871), .A(n5473), .ZN(n5478) );
  INV_X1 U6622 ( .A(n5474), .ZN(n5476) );
  AOI21_X1 U6623 ( .B1(n5483), .B2(REIP_REG_27__SCAN_IN), .A(
        REIP_REG_28__SCAN_IN), .ZN(n5475) );
  NOR2_X1 U6624 ( .A1(n5476), .A2(n5475), .ZN(n5477) );
  AOI211_X1 U6625 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6090), .A(n5478), .B(n5477), 
        .ZN(n5479) );
  OAI21_X1 U6626 ( .B1(n3121), .B2(n5873), .A(n5479), .ZN(U2799) );
  AOI21_X1 U6627 ( .B1(n5481), .B2(n5480), .A(n4234), .ZN(n5621) );
  INV_X1 U6628 ( .A(n5621), .ZN(n5602) );
  INV_X1 U6629 ( .A(n5482), .ZN(n5500) );
  INV_X1 U6630 ( .A(n5483), .ZN(n5490) );
  OR2_X1 U6631 ( .A1(n5494), .A2(n5484), .ZN(n5485) );
  NAND2_X1 U6632 ( .A1(n3143), .A2(n5485), .ZN(n5749) );
  NOR2_X1 U6633 ( .A1(n5871), .A2(n5749), .ZN(n5488) );
  OAI22_X1 U6634 ( .A1(n5486), .A2(n6019), .B1(n6104), .B2(n5619), .ZN(n5487)
         );
  AOI211_X1 U6635 ( .C1(EBX_REG_27__SCAN_IN), .C2(n6090), .A(n5488), .B(n5487), 
        .ZN(n5489) );
  OAI21_X1 U6636 ( .B1(n5490), .B2(REIP_REG_27__SCAN_IN), .A(n5489), .ZN(n5491) );
  AOI21_X1 U6637 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5500), .A(n5491), .ZN(n5492) );
  OAI21_X1 U6638 ( .B1(n5602), .B2(n5873), .A(n5492), .ZN(U2800) );
  OAI21_X1 U6639 ( .B1(n4533), .B2(n5493), .A(n5480), .ZN(n5626) );
  AOI21_X1 U6640 ( .B1(n5496), .B2(n5495), .A(n5494), .ZN(n5765) );
  INV_X1 U6641 ( .A(n5765), .ZN(n5498) );
  AOI22_X1 U6642 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6094), .B1(n6071), 
        .B2(n5627), .ZN(n5497) );
  OAI21_X1 U6643 ( .B1(n5498), .B2(n5871), .A(n5497), .ZN(n5499) );
  AOI21_X1 U6644 ( .B1(n6090), .B2(EBX_REG_26__SCAN_IN), .A(n5499), .ZN(n5503)
         );
  INV_X1 U6645 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6643) );
  INV_X1 U6646 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5637) );
  NOR3_X1 U6647 ( .A1(n5511), .A2(n6643), .A3(n5637), .ZN(n5501) );
  OAI21_X1 U6648 ( .B1(REIP_REG_26__SCAN_IN), .B2(n5501), .A(n5500), .ZN(n5502) );
  OAI211_X1 U6649 ( .C1(n5626), .C2(n5873), .A(n5503), .B(n5502), .ZN(U2801)
         );
  AOI21_X1 U6650 ( .B1(n5504), .B2(n4473), .A(n4531), .ZN(n5652) );
  INV_X1 U6651 ( .A(n5652), .ZN(n5610) );
  INV_X1 U6652 ( .A(n5650), .ZN(n5509) );
  OAI22_X1 U6653 ( .A1(n6809), .A2(n6080), .B1(n5505), .B2(n6019), .ZN(n5508)
         );
  XNOR2_X1 U6654 ( .A(n4431), .B(n5506), .ZN(n5781) );
  NOR2_X1 U6655 ( .A1(n5871), .A2(n5781), .ZN(n5507) );
  AOI211_X1 U6656 ( .C1(n6071), .C2(n5509), .A(n5508), .B(n5507), .ZN(n5510)
         );
  OAI21_X1 U6657 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5511), .A(n5510), .ZN(n5512) );
  AOI21_X1 U6658 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5877), .A(n5512), .ZN(n5513) );
  OAI21_X1 U6659 ( .B1(n5610), .B2(n5873), .A(n5513), .ZN(U2803) );
  INV_X1 U6660 ( .A(n5515), .ZN(n5516) );
  NOR2_X1 U6661 ( .A1(n5516), .A2(n5517), .ZN(n5518) );
  OR2_X1 U6662 ( .A1(n5514), .A2(n5518), .ZN(n5664) );
  INV_X1 U6663 ( .A(n5664), .ZN(n5902) );
  OAI21_X1 U6664 ( .B1(n5520), .B2(n5519), .A(n3149), .ZN(n5797) );
  NAND2_X1 U6665 ( .A1(n6090), .A2(EBX_REG_21__SCAN_IN), .ZN(n5526) );
  INV_X1 U6666 ( .A(n5890), .ZN(n5521) );
  AOI22_X1 U6667 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6094), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5521), .ZN(n5523) );
  INV_X1 U6668 ( .A(n5870), .ZN(n5522) );
  OR2_X1 U6669 ( .A1(n5522), .A2(REIP_REG_21__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U6670 ( .A1(n5523), .A2(n5881), .ZN(n5524) );
  AOI21_X1 U6671 ( .B1(n6071), .B2(n5667), .A(n5524), .ZN(n5525) );
  OAI211_X1 U6672 ( .C1(n5871), .C2(n5797), .A(n5526), .B(n5525), .ZN(n5527)
         );
  AOI21_X1 U6673 ( .B1(n5902), .B2(n6056), .A(n5527), .ZN(n5528) );
  INV_X1 U6674 ( .A(n5528), .ZN(U2806) );
  AOI21_X1 U6675 ( .B1(n5532), .B2(n5529), .A(n5531), .ZN(n5908) );
  INV_X1 U6676 ( .A(n5908), .ZN(n5578) );
  INV_X1 U6677 ( .A(n5678), .ZN(n5537) );
  XNOR2_X1 U6678 ( .A(n5805), .B(n4297), .ZN(n5582) );
  NAND2_X1 U6679 ( .A1(n5809), .A2(n5582), .ZN(n5536) );
  INV_X1 U6680 ( .A(n5582), .ZN(n5534) );
  OAI21_X1 U6681 ( .B1(n5534), .B2(n5927), .A(n5533), .ZN(n5535) );
  NAND2_X1 U6682 ( .A1(n5536), .A2(n5535), .ZN(n5825) );
  OAI22_X1 U6683 ( .A1(n5537), .A2(n6104), .B1(n5871), .B2(n5825), .ZN(n5543)
         );
  OAI21_X1 U6684 ( .B1(n6093), .B2(n5538), .A(n6086), .ZN(n6003) );
  AOI21_X1 U6685 ( .B1(n6094), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6053), 
        .ZN(n5541) );
  NOR2_X1 U6686 ( .A1(n6083), .A2(n5538), .ZN(n5990) );
  OAI211_X1 U6687 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5990), .B(n5539), .ZN(n5540) );
  OAI211_X1 U6688 ( .C1(n6635), .C2(n6003), .A(n5541), .B(n5540), .ZN(n5542)
         );
  AOI211_X1 U6689 ( .C1(n6090), .C2(EBX_REG_19__SCAN_IN), .A(n5543), .B(n5542), 
        .ZN(n5544) );
  OAI21_X1 U6690 ( .B1(n5578), .B2(n5873), .A(n5544), .ZN(U2808) );
  OAI21_X1 U6691 ( .B1(n5545), .B2(n5547), .A(n5546), .ZN(n6124) );
  OAI21_X1 U6692 ( .B1(n5549), .B2(n5548), .A(n5929), .ZN(n5845) );
  INV_X1 U6693 ( .A(n5845), .ZN(n5559) );
  INV_X1 U6694 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U6695 ( .A1(n6071), .A2(n5689), .ZN(n5550) );
  OAI211_X1 U6696 ( .C1(n6019), .C2(n5685), .A(n5550), .B(n6027), .ZN(n5558)
         );
  INV_X1 U6697 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U6698 ( .A1(n6063), .A2(n5552), .ZN(n5551) );
  NOR2_X1 U6699 ( .A1(n6717), .A2(n5551), .ZN(n5997) );
  INV_X1 U6700 ( .A(n5997), .ZN(n5555) );
  NOR2_X1 U6701 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5551), .ZN(n6005) );
  INV_X1 U6702 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U6703 ( .A1(n6063), .A2(n5553), .ZN(n6017) );
  NAND2_X1 U6704 ( .A1(n6017), .A2(n6084), .ZN(n6016) );
  NOR2_X1 U6705 ( .A1(n6005), .A2(n6016), .ZN(n5554) );
  MUX2_X1 U6706 ( .A(n5555), .B(n5554), .S(REIP_REG_16__SCAN_IN), .Z(n5556) );
  OAI21_X1 U6707 ( .B1(n4341), .B2(n6080), .A(n5556), .ZN(n5557) );
  AOI211_X1 U6708 ( .C1(n5559), .C2(n6092), .A(n5558), .B(n5557), .ZN(n5560)
         );
  OAI21_X1 U6709 ( .B1(n6124), .B2(n5873), .A(n5560), .ZN(U2811) );
  OAI222_X1 U6710 ( .A1(n5562), .A2(n6117), .B1(n5591), .B2(n5739), .C1(n3121), 
        .C2(n5592), .ZN(U2831) );
  OAI222_X1 U6711 ( .A1(n5563), .A2(n6117), .B1(n5591), .B2(n5749), .C1(n5602), 
        .C2(n5592), .ZN(U2832) );
  AOI22_X1 U6712 ( .A1(n5765), .A2(n6113), .B1(n5588), .B2(EBX_REG_26__SCAN_IN), .ZN(n5564) );
  OAI21_X1 U6713 ( .B1(n5626), .B2(n5592), .A(n5564), .ZN(U2833) );
  INV_X1 U6714 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5565) );
  OAI222_X1 U6715 ( .A1(n5769), .A2(n5591), .B1(n5565), .B2(n6117), .C1(n5607), 
        .C2(n5592), .ZN(U2834) );
  INV_X1 U6716 ( .A(n5781), .ZN(n5566) );
  AOI22_X1 U6717 ( .A1(n6113), .A2(n5566), .B1(n5588), .B2(EBX_REG_24__SCAN_IN), .ZN(n5567) );
  OAI21_X1 U6718 ( .B1(n5610), .B2(n5592), .A(n5567), .ZN(U2835) );
  INV_X1 U6719 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6757) );
  INV_X1 U6720 ( .A(n5568), .ZN(n5872) );
  OAI222_X1 U6721 ( .A1(n5592), .A2(n5874), .B1(n6117), .B2(n6757), .C1(n5872), 
        .C2(n5591), .ZN(U2836) );
  OR2_X1 U6722 ( .A1(n5514), .A2(n5569), .ZN(n5570) );
  AND2_X1 U6723 ( .A1(n4474), .A2(n5570), .ZN(n5899) );
  INV_X1 U6724 ( .A(n5899), .ZN(n5575) );
  AND2_X1 U6725 ( .A1(n3149), .A2(n5571), .ZN(n5572) );
  NOR2_X1 U6726 ( .A1(n5573), .A2(n5572), .ZN(n5885) );
  AOI22_X1 U6727 ( .A1(n6113), .A2(n5885), .B1(EBX_REG_22__SCAN_IN), .B2(n5588), .ZN(n5574) );
  OAI21_X1 U6728 ( .B1(n5575), .B2(n5592), .A(n5574), .ZN(U2837) );
  INV_X1 U6729 ( .A(n5797), .ZN(n5576) );
  AOI22_X1 U6730 ( .A1(n6113), .A2(n5576), .B1(n5588), .B2(EBX_REG_21__SCAN_IN), .ZN(n5577) );
  OAI21_X1 U6731 ( .B1(n5664), .B2(n5592), .A(n5577), .ZN(U2838) );
  OAI222_X1 U6732 ( .A1(n5592), .A2(n5578), .B1(n6117), .B2(n4288), .C1(n5825), 
        .C2(n5591), .ZN(U2840) );
  NAND2_X1 U6733 ( .A1(n5579), .A2(n5580), .ZN(n5581) );
  AND2_X1 U6734 ( .A1(n5529), .A2(n5581), .ZN(n6118) );
  INV_X1 U6735 ( .A(n6118), .ZN(n5584) );
  XNOR2_X1 U6736 ( .A(n5582), .B(n5927), .ZN(n5993) );
  AOI22_X1 U6737 ( .A1(n6113), .A2(n5993), .B1(n5588), .B2(EBX_REG_18__SCAN_IN), .ZN(n5583) );
  OAI21_X1 U6738 ( .B1(n5584), .B2(n5592), .A(n5583), .ZN(U2841) );
  OAI222_X1 U6739 ( .A1(n5845), .A2(n5591), .B1(n6117), .B2(n4341), .C1(n5592), 
        .C2(n6124), .ZN(U2843) );
  AOI21_X1 U6740 ( .B1(n5585), .B2(n5453), .A(n5545), .ZN(n6008) );
  INV_X1 U6741 ( .A(n6008), .ZN(n5697) );
  AOI21_X1 U6742 ( .B1(n5587), .B2(n5586), .A(n5548), .ZN(n6009) );
  AOI22_X1 U6743 ( .A1(n6113), .A2(n6009), .B1(n5588), .B2(EBX_REG_15__SCAN_IN), .ZN(n5589) );
  OAI21_X1 U6744 ( .B1(n5697), .B2(n5592), .A(n5589), .ZN(U2844) );
  OAI222_X1 U6745 ( .A1(n5698), .A2(n5592), .B1(n5591), .B2(n6014), .C1(n6117), 
        .C2(n5590), .ZN(U2845) );
  AND2_X1 U6746 ( .A1(n6134), .A2(n5593), .ZN(n5594) );
  NAND2_X1 U6747 ( .A1(n5595), .A2(n5594), .ZN(n5597) );
  AOI22_X1 U6748 ( .A1(n6125), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6128), .ZN(n5596) );
  NAND2_X1 U6749 ( .A1(n5597), .A2(n5596), .ZN(U2860) );
  AOI22_X1 U6750 ( .A1(n6125), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6128), .ZN(n5599) );
  NAND2_X1 U6751 ( .A1(n6129), .A2(DATAI_12_), .ZN(n5598) );
  OAI211_X1 U6752 ( .C1(n3121), .C2(n6135), .A(n5599), .B(n5598), .ZN(U2863)
         );
  AOI22_X1 U6753 ( .A1(n6125), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6128), .ZN(n5601) );
  NAND2_X1 U6754 ( .A1(n6129), .A2(DATAI_11_), .ZN(n5600) );
  OAI211_X1 U6755 ( .C1(n5602), .C2(n6135), .A(n5601), .B(n5600), .ZN(U2864)
         );
  AOI22_X1 U6756 ( .A1(n6125), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6128), .ZN(n5604) );
  NAND2_X1 U6757 ( .A1(n6129), .A2(DATAI_10_), .ZN(n5603) );
  OAI211_X1 U6758 ( .C1(n5626), .C2(n6135), .A(n5604), .B(n5603), .ZN(U2865)
         );
  AOI22_X1 U6759 ( .A1(n6125), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6128), .ZN(n5606) );
  NAND2_X1 U6760 ( .A1(n6129), .A2(DATAI_9_), .ZN(n5605) );
  OAI211_X1 U6761 ( .C1(n5607), .C2(n6135), .A(n5606), .B(n5605), .ZN(U2866)
         );
  AOI22_X1 U6762 ( .A1(n6125), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6128), .ZN(n5609) );
  NAND2_X1 U6763 ( .A1(n6129), .A2(DATAI_8_), .ZN(n5608) );
  OAI211_X1 U6764 ( .C1(n5610), .C2(n6135), .A(n5609), .B(n5608), .ZN(U2867)
         );
  AOI22_X1 U6765 ( .A1(n6129), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6128), .ZN(n5612) );
  NAND2_X1 U6766 ( .A1(n6125), .A2(DATAI_23_), .ZN(n5611) );
  OAI211_X1 U6767 ( .C1(n5874), .C2(n6135), .A(n5612), .B(n5611), .ZN(U2868)
         );
  AOI22_X1 U6768 ( .A1(n5613), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6128), .ZN(n5614) );
  OAI21_X1 U6769 ( .B1(n5697), .B2(n6135), .A(n5614), .ZN(U2876) );
  NAND2_X1 U6770 ( .A1(n5616), .A2(n5615), .ZN(n5617) );
  XNOR2_X1 U6771 ( .A(n5617), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5758)
         );
  INV_X1 U6772 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6815) );
  NOR2_X1 U6773 ( .A1(n6253), .A2(n6815), .ZN(n5750) );
  AOI21_X1 U6774 ( .B1(n6188), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5750), 
        .ZN(n5618) );
  OAI21_X1 U6775 ( .B1(n6195), .B2(n5619), .A(n5618), .ZN(n5620) );
  AOI21_X1 U6776 ( .B1(n5621), .B2(n3103), .A(n5620), .ZN(n5622) );
  OAI21_X1 U6777 ( .B1(n5758), .B2(n6172), .A(n5622), .ZN(U2959) );
  NAND2_X1 U6778 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  XNOR2_X1 U6779 ( .A(n3139), .B(n5625), .ZN(n5768) );
  INV_X1 U6780 ( .A(n5626), .ZN(n5631) );
  INV_X1 U6781 ( .A(n5627), .ZN(n5629) );
  INV_X1 U6782 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6646) );
  NOR2_X1 U6783 ( .A1(n6253), .A2(n6646), .ZN(n5764) );
  AOI21_X1 U6784 ( .B1(n6188), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5764), 
        .ZN(n5628) );
  OAI21_X1 U6785 ( .B1(n6195), .B2(n5629), .A(n5628), .ZN(n5630) );
  AOI21_X1 U6786 ( .B1(n5631), .B2(n3103), .A(n5630), .ZN(n5632) );
  OAI21_X1 U6787 ( .B1(n5768), .B2(n6172), .A(n5632), .ZN(U2960) );
  OAI21_X1 U6788 ( .B1(n5635), .B2(n5634), .A(n5633), .ZN(n5636) );
  INV_X1 U6789 ( .A(n5636), .ZN(n5776) );
  NOR2_X1 U6790 ( .A1(n6253), .A2(n5637), .ZN(n5770) );
  AOI21_X1 U6791 ( .B1(n6188), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5770), 
        .ZN(n5638) );
  OAI21_X1 U6792 ( .B1(n6195), .B2(n5639), .A(n5638), .ZN(n5640) );
  AOI21_X1 U6793 ( .B1(n5641), .B2(n3103), .A(n5640), .ZN(n5642) );
  OAI21_X1 U6794 ( .B1(n5776), .B2(n6172), .A(n5642), .ZN(U2961) );
  NAND3_X1 U6795 ( .A1(n5655), .A2(n5643), .A3(n3253), .ZN(n5647) );
  NAND2_X1 U6796 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  XNOR2_X1 U6797 ( .A(n5648), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5786)
         );
  NAND2_X1 U6798 ( .A1(n6197), .A2(REIP_REG_24__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U6799 ( .A1(n6188), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5649)
         );
  OAI211_X1 U6800 ( .C1(n6195), .C2(n5650), .A(n5780), .B(n5649), .ZN(n5651)
         );
  AOI21_X1 U6801 ( .B1(n5652), .B2(n3103), .A(n5651), .ZN(n5653) );
  OAI21_X1 U6802 ( .B1(n5786), .B2(n6172), .A(n5653), .ZN(U2962) );
  AOI21_X1 U6803 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6164), .A(n5654), 
        .ZN(n5656) );
  XOR2_X1 U6804 ( .A(n5656), .B(n5655), .Z(n5794) );
  NAND2_X1 U6805 ( .A1(n6197), .A2(REIP_REG_22__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U6806 ( .A1(n6188), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5657)
         );
  OAI211_X1 U6807 ( .C1(n6195), .C2(n5888), .A(n5789), .B(n5657), .ZN(n5658)
         );
  AOI21_X1 U6808 ( .B1(n5899), .B2(n3103), .A(n5658), .ZN(n5659) );
  OAI21_X1 U6809 ( .B1(n5794), .B2(n6172), .A(n5659), .ZN(U2964) );
  AOI21_X1 U6810 ( .B1(n5662), .B2(n5661), .A(n5660), .ZN(n5803) );
  INV_X1 U6811 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U6812 ( .A1(n6197), .A2(REIP_REG_21__SCAN_IN), .ZN(n5796) );
  OAI21_X1 U6813 ( .B1(n5686), .B2(n5663), .A(n5796), .ZN(n5666) );
  NOR2_X1 U6814 ( .A1(n5664), .A2(n5696), .ZN(n5665) );
  AOI211_X1 U6815 ( .C1(n6168), .C2(n5667), .A(n5666), .B(n5665), .ZN(n5668)
         );
  OAI21_X1 U6816 ( .B1(n5803), .B2(n6172), .A(n5668), .ZN(U2965) );
  XNOR2_X1 U6817 ( .A(n5670), .B(n5669), .ZN(n5820) );
  INV_X1 U6818 ( .A(n5671), .ZN(n5673) );
  INV_X1 U6819 ( .A(n5531), .ZN(n5672) );
  AOI21_X1 U6820 ( .B1(n5673), .B2(n5672), .A(n5516), .ZN(n5905) );
  NAND2_X1 U6821 ( .A1(n6197), .A2(REIP_REG_20__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U6822 ( .A1(n6188), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5674)
         );
  OAI211_X1 U6823 ( .C1(n6195), .C2(n5896), .A(n5816), .B(n5674), .ZN(n5675)
         );
  AOI21_X1 U6824 ( .B1(n5905), .B2(n3103), .A(n5675), .ZN(n5676) );
  OAI21_X1 U6825 ( .B1(n5820), .B2(n6172), .A(n5676), .ZN(U2966) );
  XNOR2_X1 U6826 ( .A(n3107), .B(n3140), .ZN(n5829) );
  NAND2_X1 U6827 ( .A1(n6168), .A2(n5678), .ZN(n5679) );
  NAND2_X1 U6828 ( .A1(n6197), .A2(REIP_REG_19__SCAN_IN), .ZN(n5823) );
  OAI211_X1 U6829 ( .C1(n5686), .C2(n5680), .A(n5679), .B(n5823), .ZN(n5681)
         );
  AOI21_X1 U6830 ( .B1(n5908), .B2(n3103), .A(n5681), .ZN(n5682) );
  OAI21_X1 U6831 ( .B1(n5829), .B2(n6172), .A(n5682), .ZN(U2967) );
  XNOR2_X1 U6832 ( .A(n6164), .B(n5840), .ZN(n5684) );
  XNOR2_X1 U6833 ( .A(n5683), .B(n5684), .ZN(n5849) );
  NAND2_X1 U6834 ( .A1(n6197), .A2(REIP_REG_16__SCAN_IN), .ZN(n5844) );
  OAI21_X1 U6835 ( .B1(n5686), .B2(n5685), .A(n5844), .ZN(n5688) );
  NOR2_X1 U6836 ( .A1(n6124), .A2(n5696), .ZN(n5687) );
  AOI211_X1 U6837 ( .C1(n6168), .C2(n5689), .A(n5688), .B(n5687), .ZN(n5690)
         );
  OAI21_X1 U6838 ( .B1(n6172), .B2(n5849), .A(n5690), .ZN(U2970) );
  NOR2_X1 U6839 ( .A1(n6253), .A2(n6717), .ZN(n5935) );
  NOR2_X1 U6840 ( .A1(n6195), .A2(n6006), .ZN(n5691) );
  AOI211_X1 U6841 ( .C1(n6188), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5935), 
        .B(n5691), .ZN(n5695) );
  XNOR2_X1 U6842 ( .A(n6164), .B(n5942), .ZN(n5693) );
  XNOR2_X1 U6843 ( .A(n5692), .B(n5693), .ZN(n5939) );
  NAND2_X1 U6844 ( .A1(n5939), .A2(n6191), .ZN(n5694) );
  OAI211_X1 U6845 ( .C1(n5697), .C2(n5696), .A(n5695), .B(n5694), .ZN(U2971)
         );
  INV_X1 U6846 ( .A(n5698), .ZN(n6023) );
  INV_X1 U6847 ( .A(n6022), .ZN(n5700) );
  AOI22_X1 U6848 ( .A1(n6188), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6197), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5699) );
  OAI21_X1 U6849 ( .B1(n6195), .B2(n5700), .A(n5699), .ZN(n5701) );
  AOI21_X1 U6850 ( .B1(n6023), .B2(n3103), .A(n5701), .ZN(n5702) );
  OAI21_X1 U6851 ( .B1(n5703), .B2(n6172), .A(n5702), .ZN(U2972) );
  INV_X1 U6852 ( .A(n5704), .ZN(n5721) );
  INV_X1 U6853 ( .A(n5705), .ZN(n5713) );
  NAND2_X1 U6854 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5759) );
  NOR2_X1 U6855 ( .A1(n5773), .A2(n5759), .ZN(n5753) );
  NAND2_X1 U6856 ( .A1(n5753), .A2(n5706), .ZN(n5730) );
  INV_X1 U6857 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5707) );
  NOR4_X1 U6858 ( .A1(n5730), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6776), 
        .A4(n5707), .ZN(n5708) );
  AOI211_X1 U6859 ( .C1(n6266), .C2(n5710), .A(n5709), .B(n5708), .ZN(n5720)
         );
  NAND2_X1 U6860 ( .A1(n5712), .A2(n5711), .ZN(n5804) );
  NAND2_X1 U6861 ( .A1(n5804), .A2(n5713), .ZN(n5714) );
  NAND2_X1 U6862 ( .A1(n5787), .A2(n5714), .ZN(n5784) );
  AND2_X1 U6863 ( .A1(n5838), .A2(n5759), .ZN(n5715) );
  NOR2_X1 U6864 ( .A1(n5784), .A2(n5715), .ZN(n5754) );
  NAND2_X1 U6865 ( .A1(n5838), .A2(n5742), .ZN(n5716) );
  AND2_X1 U6866 ( .A1(n5754), .A2(n5716), .ZN(n5735) );
  NAND2_X1 U6867 ( .A1(n5838), .A2(n6776), .ZN(n5717) );
  AND2_X1 U6868 ( .A1(n5735), .A2(n5717), .ZN(n5725) );
  OAI21_X1 U6869 ( .B1(n6209), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5725), 
        .ZN(n5718) );
  NAND2_X1 U6870 ( .A1(n5718), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5719) );
  OAI211_X1 U6871 ( .C1(n5721), .C2(n6223), .A(n5720), .B(n5719), .ZN(U2987)
         );
  NOR3_X1 U6872 ( .A1(n5730), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6776), 
        .ZN(n5723) );
  AOI211_X1 U6873 ( .C1(n6266), .C2(n3208), .A(n5724), .B(n5723), .ZN(n5728)
         );
  INV_X1 U6874 ( .A(n5725), .ZN(n5726) );
  NAND2_X1 U6875 ( .A1(n5726), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5727) );
  OAI211_X1 U6876 ( .C1(n5729), .C2(n6223), .A(n5728), .B(n5727), .ZN(U2988)
         );
  INV_X1 U6877 ( .A(n5730), .ZN(n5734) );
  NOR2_X1 U6878 ( .A1(n5731), .A2(n6255), .ZN(n5733) );
  AOI211_X1 U6879 ( .C1(n5734), .C2(n6776), .A(n5733), .B(n5732), .ZN(n5737)
         );
  OR2_X1 U6880 ( .A1(n5735), .A2(n6776), .ZN(n5736) );
  OAI211_X1 U6881 ( .C1(n5738), .C2(n6223), .A(n5737), .B(n5736), .ZN(U2989)
         );
  INV_X1 U6882 ( .A(n5739), .ZN(n5741) );
  AOI21_X1 U6883 ( .B1(n5741), .B2(n6266), .A(n5740), .ZN(n5745) );
  NAND3_X1 U6884 ( .A1(n5753), .A2(n5743), .A3(n5742), .ZN(n5744) );
  OAI211_X1 U6885 ( .C1(n5754), .C2(n6983), .A(n5745), .B(n5744), .ZN(n5746)
         );
  INV_X1 U6886 ( .A(n5746), .ZN(n5747) );
  OAI21_X1 U6887 ( .B1(n5748), .B2(n6223), .A(n5747), .ZN(U2990) );
  NOR2_X1 U6888 ( .A1(n5749), .A2(n6255), .ZN(n5751) );
  AOI211_X1 U6889 ( .C1(n5753), .C2(n5752), .A(n5751), .B(n5750), .ZN(n5757)
         );
  INV_X1 U6890 ( .A(n5754), .ZN(n5755) );
  NAND2_X1 U6891 ( .A1(n5755), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5756) );
  OAI211_X1 U6892 ( .C1(n5758), .C2(n6223), .A(n5757), .B(n5756), .ZN(U2991)
         );
  INV_X1 U6893 ( .A(n5759), .ZN(n5760) );
  AOI211_X1 U6894 ( .C1(n5762), .C2(n5761), .A(n5760), .B(n5773), .ZN(n5763)
         );
  AOI211_X1 U6895 ( .C1(n6266), .C2(n5765), .A(n5764), .B(n5763), .ZN(n5767)
         );
  NAND2_X1 U6896 ( .A1(n5784), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5766) );
  OAI211_X1 U6897 ( .C1(n5768), .C2(n6223), .A(n5767), .B(n5766), .ZN(U2992)
         );
  INV_X1 U6898 ( .A(n5769), .ZN(n5771) );
  AOI21_X1 U6899 ( .B1(n6266), .B2(n5771), .A(n5770), .ZN(n5772) );
  OAI21_X1 U6900 ( .B1(n5773), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5772), 
        .ZN(n5774) );
  AOI21_X1 U6901 ( .B1(n5784), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5774), 
        .ZN(n5775) );
  OAI21_X1 U6902 ( .B1(n5776), .B2(n6223), .A(n5775), .ZN(U2993) );
  OAI21_X1 U6903 ( .B1(n5779), .B2(n5778), .A(n5777), .ZN(n5783) );
  OAI21_X1 U6904 ( .B1(n6255), .B2(n5781), .A(n5780), .ZN(n5782) );
  AOI21_X1 U6905 ( .B1(n5784), .B2(n5783), .A(n5782), .ZN(n5785) );
  OAI21_X1 U6906 ( .B1(n5786), .B2(n6223), .A(n5785), .ZN(U2994) );
  INV_X1 U6907 ( .A(n5787), .ZN(n5792) );
  NAND2_X1 U6908 ( .A1(n6266), .A2(n5885), .ZN(n5788) );
  OAI211_X1 U6909 ( .C1(n5790), .C2(n6723), .A(n5789), .B(n5788), .ZN(n5791)
         );
  AOI21_X1 U6910 ( .B1(n5792), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5791), 
        .ZN(n5793) );
  OAI21_X1 U6911 ( .B1(n5794), .B2(n6223), .A(n5793), .ZN(U2996) );
  INV_X1 U6912 ( .A(n5795), .ZN(n5801) );
  OAI21_X1 U6913 ( .B1(n6255), .B2(n5797), .A(n5796), .ZN(n5800) );
  NOR2_X1 U6914 ( .A1(n5798), .A2(n6723), .ZN(n5799) );
  AOI211_X1 U6915 ( .C1(n5801), .C2(n6723), .A(n5800), .B(n5799), .ZN(n5802)
         );
  OAI21_X1 U6916 ( .B1(n5803), .B2(n6223), .A(n5802), .ZN(U2997) );
  AOI21_X1 U6917 ( .B1(n5930), .B2(n5804), .A(n5925), .ZN(n5833) );
  OAI21_X1 U6918 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6209), .A(n5833), 
        .ZN(n5827) );
  INV_X1 U6919 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U6920 ( .A1(n5809), .A2(n5806), .ZN(n5807) );
  OAI21_X1 U6921 ( .B1(n5809), .B2(n5808), .A(n5807), .ZN(n5812) );
  INV_X1 U6922 ( .A(n5810), .ZN(n5811) );
  XNOR2_X1 U6923 ( .A(n5812), .B(n5811), .ZN(n5893) );
  INV_X1 U6924 ( .A(n5813), .ZN(n5815) );
  NAND3_X1 U6925 ( .A1(n5822), .A2(n5815), .A3(n5814), .ZN(n5817) );
  OAI211_X1 U6926 ( .C1(n5893), .C2(n6255), .A(n5817), .B(n5816), .ZN(n5818)
         );
  AOI21_X1 U6927 ( .B1(INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n5827), .A(n5818), 
        .ZN(n5819) );
  OAI21_X1 U6928 ( .B1(n5820), .B2(n6223), .A(n5819), .ZN(U2998) );
  NAND2_X1 U6929 ( .A1(n5822), .A2(n5821), .ZN(n5824) );
  OAI211_X1 U6930 ( .C1(n6255), .C2(n5825), .A(n5824), .B(n5823), .ZN(n5826)
         );
  AOI21_X1 U6931 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5827), .A(n5826), 
        .ZN(n5828) );
  OAI21_X1 U6932 ( .B1(n5829), .B2(n6223), .A(n5828), .ZN(U2999) );
  NAND3_X1 U6933 ( .A1(n5683), .A2(n3140), .A3(n5840), .ZN(n5914) );
  NOR3_X1 U6934 ( .A1(n5683), .A2(n3140), .A3(n5840), .ZN(n5916) );
  NAND2_X1 U6935 ( .A1(n5916), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5830) );
  OAI21_X1 U6936 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5914), .A(n5830), 
        .ZN(n5831) );
  XNOR2_X1 U6937 ( .A(n5831), .B(n5832), .ZN(n5911) );
  INV_X1 U6938 ( .A(n5911), .ZN(n5837) );
  OAI22_X1 U6939 ( .A1(n5833), .A2(n5832), .B1(n6253), .B2(n6633), .ZN(n5835)
         );
  NOR3_X1 U6940 ( .A1(n5926), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5930), 
        .ZN(n5834) );
  AOI211_X1 U6941 ( .C1(n6266), .C2(n5993), .A(n5835), .B(n5834), .ZN(n5836)
         );
  OAI21_X1 U6942 ( .B1(n5837), .B2(n6223), .A(n5836), .ZN(U3000) );
  AND2_X1 U6943 ( .A1(n5838), .A2(n5936), .ZN(n5839) );
  NOR2_X1 U6944 ( .A1(n6200), .A2(n5839), .ZN(n5943) );
  INV_X1 U6945 ( .A(n5943), .ZN(n5847) );
  AOI211_X1 U6946 ( .C1(n5942), .C2(n5840), .A(n5937), .B(n5936), .ZN(n5842)
         );
  NAND2_X1 U6947 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  OAI211_X1 U6948 ( .C1(n6255), .C2(n5845), .A(n5844), .B(n5843), .ZN(n5846)
         );
  AOI21_X1 U6949 ( .B1(n5847), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5846), 
        .ZN(n5848) );
  OAI21_X1 U6950 ( .B1(n5849), .B2(n6223), .A(n5848), .ZN(U3002) );
  INV_X1 U6951 ( .A(n5850), .ZN(n5858) );
  INV_X1 U6952 ( .A(n6515), .ZN(n5856) );
  OAI211_X1 U6953 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3129), .A(n5856), .B(
        n6409), .ZN(n5851) );
  OAI21_X1 U6954 ( .B1(n5858), .B2(n5852), .A(n5851), .ZN(n5853) );
  MUX2_X1 U6955 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5853), .S(n6275), 
        .Z(U3464) );
  INV_X1 U6956 ( .A(n4914), .ZN(n5859) );
  NAND2_X1 U6957 ( .A1(n5855), .A2(n5854), .ZN(n6312) );
  NOR2_X1 U6958 ( .A1(n6432), .A2(n5856), .ZN(n6483) );
  NOR2_X1 U6959 ( .A1(n6312), .A2(n6483), .ZN(n5857) );
  OAI222_X1 U6960 ( .A1(n5859), .A2(n6280), .B1(n5858), .B2(n6354), .C1(n6527), 
        .C2(n5857), .ZN(n5860) );
  MUX2_X1 U6961 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5860), .S(n6275), 
        .Z(U3462) );
  INV_X1 U6962 ( .A(n5861), .ZN(n5864) );
  OAI22_X1 U6963 ( .A1(n5864), .A2(n6673), .B1(n5863), .B2(n5862), .ZN(n5865)
         );
  MUX2_X1 U6964 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5865), .S(n6669), 
        .Z(U3456) );
  AOI21_X1 U6965 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5867), .A(n5866), .ZN(
        n5868) );
  INV_X1 U6966 ( .A(n5868), .ZN(U2788) );
  AOI22_X1 U6967 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6090), .B1(n5869), .B2(n6071), .ZN(n5879) );
  INV_X1 U6968 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U6969 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5870), .ZN(n5882) );
  OAI21_X1 U6970 ( .B1(n6640), .B2(n5882), .A(n4367), .ZN(n5876) );
  OAI22_X1 U6971 ( .A1(n5874), .A2(n5873), .B1(n5872), .B2(n5871), .ZN(n5875)
         );
  AOI21_X1 U6972 ( .B1(n5877), .B2(n5876), .A(n5875), .ZN(n5878) );
  OAI211_X1 U6973 ( .C1(n5880), .C2(n6019), .A(n5879), .B(n5878), .ZN(U2804)
         );
  AOI21_X1 U6974 ( .B1(n5890), .B2(n5881), .A(n6640), .ZN(n5884) );
  INV_X1 U6975 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6745) );
  OAI22_X1 U6976 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5882), .B1(n6745), .B2(
        n6019), .ZN(n5883) );
  AOI211_X1 U6977 ( .C1(n6090), .C2(EBX_REG_22__SCAN_IN), .A(n5884), .B(n5883), 
        .ZN(n5887) );
  AOI22_X1 U6978 ( .A1(n5899), .A2(n6056), .B1(n5885), .B2(n6092), .ZN(n5886)
         );
  OAI211_X1 U6979 ( .C1(n5888), .C2(n6104), .A(n5887), .B(n5886), .ZN(U2805)
         );
  AOI21_X1 U6980 ( .B1(n5889), .B2(n5990), .A(REIP_REG_20__SCAN_IN), .ZN(n5891) );
  INV_X1 U6981 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6899) );
  OAI22_X1 U6982 ( .A1(n5891), .A2(n5890), .B1(n6899), .B2(n6080), .ZN(n5892)
         );
  AOI21_X1 U6983 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6094), .A(n5892), 
        .ZN(n5895) );
  INV_X1 U6984 ( .A(n5893), .ZN(n5897) );
  AOI22_X1 U6985 ( .A1(n5905), .A2(n6056), .B1(n6092), .B2(n5897), .ZN(n5894)
         );
  OAI211_X1 U6986 ( .C1(n5896), .C2(n6104), .A(n5895), .B(n5894), .ZN(U2807)
         );
  AOI22_X1 U6987 ( .A1(n5905), .A2(n6114), .B1(n6113), .B2(n5897), .ZN(n5898)
         );
  OAI21_X1 U6988 ( .B1(n6899), .B2(n6117), .A(n5898), .ZN(U2839) );
  AOI22_X1 U6989 ( .A1(n5899), .A2(n6126), .B1(n6125), .B2(DATAI_22_), .ZN(
        n5901) );
  AOI22_X1 U6990 ( .A1(n6129), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6128), .ZN(n5900) );
  NAND2_X1 U6991 ( .A1(n5901), .A2(n5900), .ZN(U2869) );
  AOI22_X1 U6992 ( .A1(n5902), .A2(n6126), .B1(n6125), .B2(DATAI_21_), .ZN(
        n5904) );
  AOI22_X1 U6993 ( .A1(n6129), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6128), .ZN(n5903) );
  NAND2_X1 U6994 ( .A1(n5904), .A2(n5903), .ZN(U2870) );
  AOI22_X1 U6995 ( .A1(n5905), .A2(n6126), .B1(n6125), .B2(DATAI_20_), .ZN(
        n5907) );
  AOI22_X1 U6996 ( .A1(n6129), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6128), .ZN(n5906) );
  NAND2_X1 U6997 ( .A1(n5907), .A2(n5906), .ZN(U2871) );
  AOI22_X1 U6998 ( .A1(n5908), .A2(n6126), .B1(n6125), .B2(DATAI_19_), .ZN(
        n5910) );
  AOI22_X1 U6999 ( .A1(n6129), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6128), .ZN(n5909) );
  NAND2_X1 U7000 ( .A1(n5910), .A2(n5909), .ZN(U2872) );
  AOI22_X1 U7001 ( .A1(n6197), .A2(REIP_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6188), .ZN(n5913) );
  AOI22_X1 U7002 ( .A1(n5911), .A2(n6191), .B1(n3103), .B2(n6118), .ZN(n5912)
         );
  OAI211_X1 U7003 ( .C1(n5996), .C2(n6195), .A(n5913), .B(n5912), .ZN(U2968)
         );
  INV_X1 U7004 ( .A(n5914), .ZN(n5915) );
  NOR2_X1 U7005 ( .A1(n5916), .A2(n5915), .ZN(n5917) );
  XNOR2_X1 U7006 ( .A(n5917), .B(n5930), .ZN(n5934) );
  AOI22_X1 U7007 ( .A1(n6197), .A2(REIP_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6188), .ZN(n5920) );
  XOR2_X1 U7008 ( .A(n5918), .B(n5546), .Z(n6121) );
  AOI22_X1 U7009 ( .A1(n6121), .A2(n3103), .B1(n6168), .B2(n6000), .ZN(n5919)
         );
  OAI211_X1 U7010 ( .C1(n5934), .C2(n6172), .A(n5920), .B(n5919), .ZN(U2969)
         );
  AOI22_X1 U7011 ( .A1(n6197), .A2(REIP_REG_13__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n6188), .ZN(n5924) );
  XNOR2_X1 U7012 ( .A(n5922), .B(n5921), .ZN(n5956) );
  AOI22_X1 U7013 ( .A1(n5956), .A2(n6191), .B1(n3103), .B2(n6108), .ZN(n5923)
         );
  OAI211_X1 U7014 ( .C1(n6040), .C2(n6195), .A(n5924), .B(n5923), .ZN(U2973)
         );
  AOI22_X1 U7015 ( .A1(n6197), .A2(REIP_REG_17__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5925), .ZN(n5933) );
  INV_X1 U7016 ( .A(n5926), .ZN(n5931) );
  AOI21_X1 U7017 ( .B1(n5929), .B2(n5928), .A(n4348), .ZN(n6105) );
  AOI22_X1 U7018 ( .A1(n5931), .A2(n5930), .B1(n6105), .B2(n6266), .ZN(n5932)
         );
  OAI211_X1 U7019 ( .C1(n5934), .C2(n6223), .A(n5933), .B(n5932), .ZN(U3001)
         );
  AOI21_X1 U7020 ( .B1(n6266), .B2(n6009), .A(n5935), .ZN(n5941) );
  NOR2_X1 U7021 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  AOI22_X1 U7022 ( .A1(n5939), .A2(n6269), .B1(n5938), .B2(n5942), .ZN(n5940)
         );
  OAI211_X1 U7023 ( .C1(n5943), .C2(n5942), .A(n5941), .B(n5940), .ZN(U3003)
         );
  INV_X1 U7024 ( .A(n5944), .ZN(n5945) );
  NAND2_X1 U7025 ( .A1(n5946), .A2(n5945), .ZN(n5951) );
  AOI21_X1 U7026 ( .B1(n5949), .B2(n5948), .A(n5947), .ZN(n6107) );
  INV_X1 U7027 ( .A(n6107), .ZN(n5950) );
  OAI22_X1 U7028 ( .A1(n5952), .A2(n5951), .B1(n6255), .B2(n5950), .ZN(n5953)
         );
  INV_X1 U7029 ( .A(n5953), .ZN(n5960) );
  INV_X1 U7030 ( .A(n5954), .ZN(n5955) );
  AOI22_X1 U7031 ( .A1(n5956), .A2(n6269), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5955), .ZN(n5959) );
  NAND2_X1 U7032 ( .A1(n6197), .A2(REIP_REG_13__SCAN_IN), .ZN(n5957) );
  NAND4_X1 U7033 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(U3005)
         );
  OR4_X1 U7034 ( .A1(n5962), .A2(n5961), .A3(n6673), .A4(n4282), .ZN(n5963) );
  OAI21_X1 U7035 ( .B1(n6669), .B2(n5964), .A(n5963), .ZN(U3455) );
  AOI21_X1 U7036 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6608), .A(n6602), .ZN(n5971) );
  INV_X1 U7037 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5965) );
  AOI21_X1 U7038 ( .B1(n5971), .B2(n5965), .A(n6684), .ZN(U2789) );
  NAND2_X1 U7039 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5966), .ZN(n5969) );
  OAI21_X1 U7040 ( .B1(n5967), .B2(n6582), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5968) );
  OAI21_X1 U7041 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5969), .A(n5968), .ZN(
        U2790) );
  INV_X2 U7042 ( .A(n6684), .ZN(n6700) );
  NOR2_X1 U7043 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5972) );
  OAI21_X1 U7044 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5972), .A(n6700), .ZN(n5970)
         );
  OAI21_X1 U7045 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6700), .A(n5970), .ZN(
        U2791) );
  NOR2_X1 U7046 ( .A1(n6684), .A2(n5971), .ZN(n6661) );
  OAI21_X1 U7047 ( .B1(n5972), .B2(BS16_N), .A(n6661), .ZN(n6659) );
  OAI21_X1 U7048 ( .B1(n6661), .B2(n6703), .A(n6659), .ZN(U2792) );
  OAI21_X1 U7049 ( .B1(n5974), .B2(n5973), .A(n6172), .ZN(U2793) );
  NOR4_X1 U7050 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5978) );
  NOR4_X1 U7051 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(DATAWIDTH_REG_14__SCAN_IN), .ZN(n5977)
         );
  NOR4_X1 U7052 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n5976) );
  NOR4_X1 U7053 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n5975) );
  NAND4_X1 U7054 ( .A1(n5978), .A2(n5977), .A3(n5976), .A4(n5975), .ZN(n5984)
         );
  NOR4_X1 U7055 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_30__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5982) );
  AOI211_X1 U7056 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_18__SCAN_IN), .B(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5981) );
  NOR4_X1 U7057 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5980) );
  NOR4_X1 U7058 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n5979) );
  NAND4_X1 U7059 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n5983)
         );
  NOR2_X1 U7060 ( .A1(n5984), .A2(n5983), .ZN(n6678) );
  INV_X1 U7061 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5986) );
  NOR3_X1 U7062 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5987) );
  OAI21_X1 U7063 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5987), .A(n6678), .ZN(n5985)
         );
  OAI21_X1 U7064 ( .B1(n6678), .B2(n5986), .A(n5985), .ZN(U2794) );
  INV_X1 U7065 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6980) );
  INV_X1 U7066 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6660) );
  AOI21_X1 U7067 ( .B1(n6980), .B2(n6660), .A(n5987), .ZN(n5989) );
  INV_X1 U7068 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5988) );
  INV_X1 U7069 ( .A(n6678), .ZN(n6681) );
  AOI22_X1 U7070 ( .A1(n6678), .A2(n5989), .B1(n5988), .B2(n6681), .ZN(U2795)
         );
  AOI22_X1 U7071 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6090), .B1(n5990), .B2(n6633), .ZN(n5991) );
  OAI21_X1 U7072 ( .B1(n6633), .B2(n6003), .A(n5991), .ZN(n5992) );
  AOI211_X1 U7073 ( .C1(n6094), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6053), 
        .B(n5992), .ZN(n5995) );
  AOI22_X1 U7074 ( .A1(n6118), .A2(n6056), .B1(n6092), .B2(n5993), .ZN(n5994)
         );
  OAI211_X1 U7075 ( .C1(n5996), .C2(n6104), .A(n5995), .B(n5994), .ZN(U2809)
         );
  AOI21_X1 U7076 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5997), .A(
        REIP_REG_17__SCAN_IN), .ZN(n6004) );
  INV_X1 U7077 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6735) );
  OAI22_X1 U7078 ( .A1(n6735), .A2(n6080), .B1(n5998), .B2(n6019), .ZN(n5999)
         );
  AOI211_X1 U7079 ( .C1(n6071), .C2(n6000), .A(n6053), .B(n5999), .ZN(n6002)
         );
  AOI22_X1 U7080 ( .A1(n6121), .A2(n6056), .B1(n6092), .B2(n6105), .ZN(n6001)
         );
  OAI211_X1 U7081 ( .C1(n6004), .C2(n6003), .A(n6002), .B(n6001), .ZN(U2810)
         );
  AOI22_X1 U7082 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6090), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6016), .ZN(n6013) );
  AOI211_X1 U7083 ( .C1(n6094), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6053), 
        .B(n6005), .ZN(n6012) );
  INV_X1 U7084 ( .A(n6006), .ZN(n6007) );
  AOI22_X1 U7085 ( .A1(n6008), .A2(n6056), .B1(n6007), .B2(n6071), .ZN(n6011)
         );
  NAND2_X1 U7086 ( .A1(n6092), .A2(n6009), .ZN(n6010) );
  NAND4_X1 U7087 ( .A1(n6013), .A2(n6012), .A3(n6011), .A4(n6010), .ZN(U2812)
         );
  INV_X1 U7088 ( .A(n6014), .ZN(n6015) );
  AOI22_X1 U7089 ( .A1(n6016), .A2(REIP_REG_14__SCAN_IN), .B1(n6092), .B2(
        n6015), .ZN(n6026) );
  OAI22_X1 U7090 ( .A1(n6020), .A2(n6019), .B1(n6018), .B2(n6017), .ZN(n6021)
         );
  AOI211_X1 U7091 ( .C1(n6090), .C2(EBX_REG_14__SCAN_IN), .A(n6053), .B(n6021), 
        .ZN(n6025) );
  AOI22_X1 U7092 ( .A1(n6023), .A2(n6056), .B1(n6071), .B2(n6022), .ZN(n6024)
         );
  NAND3_X1 U7093 ( .A1(n6026), .A2(n6025), .A3(n6024), .ZN(U2813) );
  NAND2_X1 U7094 ( .A1(n6092), .A2(n6107), .ZN(n6035) );
  NAND2_X1 U7095 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6028)
         );
  AND2_X1 U7096 ( .A1(n6028), .A2(n6027), .ZN(n6034) );
  NAND2_X1 U7097 ( .A1(n6090), .A2(EBX_REG_13__SCAN_IN), .ZN(n6033) );
  INV_X1 U7098 ( .A(n6029), .ZN(n6030) );
  NOR2_X1 U7099 ( .A1(n6030), .A2(REIP_REG_13__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7100 ( .A1(n6063), .A2(n6031), .ZN(n6032) );
  NAND4_X1 U7101 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n6036)
         );
  AOI21_X1 U7102 ( .B1(n6108), .B2(n6056), .A(n6036), .ZN(n6039) );
  OAI21_X1 U7103 ( .B1(n6037), .B2(n6043), .A(REIP_REG_13__SCAN_IN), .ZN(n6038) );
  OAI211_X1 U7104 ( .C1(n6104), .C2(n6040), .A(n6039), .B(n6038), .ZN(U2814)
         );
  NAND3_X1 U7105 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n6058), .ZN(n6049) );
  INV_X1 U7106 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6112) );
  AOI21_X1 U7107 ( .B1(n6042), .B2(n6041), .A(n5368), .ZN(n6198) );
  AOI22_X1 U7108 ( .A1(n6043), .A2(REIP_REG_11__SCAN_IN), .B1(n6092), .B2(
        n6198), .ZN(n6044) );
  OAI21_X1 U7109 ( .B1(n6112), .B2(n6080), .A(n6044), .ZN(n6045) );
  AOI211_X1 U7110 ( .C1(n6094), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6053), 
        .B(n6045), .ZN(n6048) );
  AOI22_X1 U7111 ( .A1(n6169), .A2(n6056), .B1(n6071), .B2(n6167), .ZN(n6047)
         );
  OAI211_X1 U7112 ( .C1(REIP_REG_11__SCAN_IN), .C2(n6049), .A(n6048), .B(n6047), .ZN(U2816) );
  AOI22_X1 U7113 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6090), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n6094), .ZN(n6062) );
  AOI21_X1 U7114 ( .B1(n6052), .B2(n6051), .A(n6050), .ZN(n6216) );
  AOI21_X1 U7115 ( .B1(n6092), .B2(n6216), .A(n6053), .ZN(n6061) );
  INV_X1 U7116 ( .A(n6054), .ZN(n6115) );
  AOI22_X1 U7117 ( .A1(n6115), .A2(n6056), .B1(n6071), .B2(n6055), .ZN(n6060)
         );
  OAI21_X1 U7118 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6058), .A(n6057), .ZN(n6059)
         );
  NAND4_X1 U7119 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(U2818)
         );
  NAND2_X1 U7120 ( .A1(n6063), .A2(n6980), .ZN(n6096) );
  NAND3_X1 U7121 ( .A1(n6096), .A2(REIP_REG_2__SCAN_IN), .A3(n6084), .ZN(n6074) );
  INV_X1 U7122 ( .A(n6064), .ZN(n6101) );
  NAND2_X1 U7123 ( .A1(n6065), .A2(n6101), .ZN(n6069) );
  AOI22_X1 U7124 ( .A1(n6092), .A2(n6265), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n6094), .ZN(n6068) );
  NAND2_X1 U7125 ( .A1(n6095), .A2(n3118), .ZN(n6067) );
  NAND2_X1 U7126 ( .A1(n6090), .A2(EBX_REG_3__SCAN_IN), .ZN(n6066) );
  NAND4_X1 U7127 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n6070)
         );
  AOI21_X1 U7128 ( .B1(n6072), .B2(n6071), .A(n6070), .ZN(n6073) );
  OAI221_X1 U7129 ( .B1(n6075), .B2(n4829), .C1(n6075), .C2(n6074), .A(n6073), 
        .ZN(U2824) );
  INV_X1 U7130 ( .A(n6076), .ZN(n6077) );
  AOI22_X1 U7131 ( .A1(n6092), .A2(n6077), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6094), .ZN(n6079) );
  NAND2_X1 U7132 ( .A1(n6095), .A2(n4761), .ZN(n6078) );
  OAI211_X1 U7133 ( .C1(n6081), .C2(n6080), .A(n6079), .B(n6078), .ZN(n6082)
         );
  AOI21_X1 U7134 ( .B1(n6190), .B2(n6101), .A(n6082), .ZN(n6089) );
  NOR2_X1 U7135 ( .A1(n6083), .A2(n6980), .ZN(n6087) );
  NAND3_X1 U7136 ( .A1(n6084), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6085) );
  OAI211_X1 U7137 ( .C1(n6087), .C2(REIP_REG_2__SCAN_IN), .A(n6086), .B(n6085), 
        .ZN(n6088) );
  OAI211_X1 U7138 ( .C1(n6104), .C2(n6196), .A(n6089), .B(n6088), .ZN(U2825)
         );
  AOI22_X1 U7139 ( .A1(n6092), .A2(n6091), .B1(n6090), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n6099) );
  AOI22_X1 U7140 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6093), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7141 ( .A1(n6095), .A2(n4575), .ZN(n6097) );
  NAND4_X1 U7142 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), .ZN(n6100)
         );
  AOI21_X1 U7143 ( .B1(n6102), .B2(n6101), .A(n6100), .ZN(n6103) );
  OAI21_X1 U7144 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6104), .A(n6103), 
        .ZN(U2826) );
  AOI22_X1 U7145 ( .A1(n6121), .A2(n6114), .B1(n6113), .B2(n6105), .ZN(n6106)
         );
  OAI21_X1 U7146 ( .B1(n6735), .B2(n6117), .A(n6106), .ZN(U2842) );
  INV_X1 U7147 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6110) );
  AOI22_X1 U7148 ( .A1(n6108), .A2(n6114), .B1(n6113), .B2(n6107), .ZN(n6109)
         );
  OAI21_X1 U7149 ( .B1(n6110), .B2(n6117), .A(n6109), .ZN(U2846) );
  AOI22_X1 U7150 ( .A1(n6169), .A2(n6114), .B1(n6113), .B2(n6198), .ZN(n6111)
         );
  OAI21_X1 U7151 ( .B1(n6112), .B2(n6117), .A(n6111), .ZN(U2848) );
  AOI22_X1 U7152 ( .A1(n6115), .A2(n6114), .B1(n6113), .B2(n6216), .ZN(n6116)
         );
  OAI21_X1 U7153 ( .B1(n6732), .B2(n6117), .A(n6116), .ZN(U2850) );
  AOI22_X1 U7154 ( .A1(n6118), .A2(n6126), .B1(n6125), .B2(DATAI_18_), .ZN(
        n6120) );
  AOI22_X1 U7155 ( .A1(n6129), .A2(DATAI_2_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6128), .ZN(n6119) );
  NAND2_X1 U7156 ( .A1(n6120), .A2(n6119), .ZN(U2873) );
  AOI22_X1 U7157 ( .A1(n6121), .A2(n6126), .B1(n6125), .B2(DATAI_17_), .ZN(
        n6123) );
  AOI22_X1 U7158 ( .A1(n6129), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6128), .ZN(n6122) );
  NAND2_X1 U7159 ( .A1(n6123), .A2(n6122), .ZN(U2874) );
  INV_X1 U7160 ( .A(n6124), .ZN(n6127) );
  AOI22_X1 U7161 ( .A1(n6127), .A2(n6126), .B1(n6125), .B2(DATAI_16_), .ZN(
        n6131) );
  AOI22_X1 U7162 ( .A1(n6129), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6128), .ZN(n6130) );
  NAND2_X1 U7163 ( .A1(n6131), .A2(n6130), .ZN(U2875) );
  INV_X1 U7164 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6918) );
  OAI222_X1 U7165 ( .A1(n6136), .A2(n6135), .B1(n6134), .B2(n6918), .C1(n6133), 
        .C2(n6132), .ZN(U2891) );
  INV_X1 U7166 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6762) );
  AOI22_X1 U7167 ( .A1(n6140), .A2(DATAO_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6139), .ZN(n6137) );
  OAI21_X1 U7168 ( .B1(n6142), .B2(n6762), .A(n6137), .ZN(U2913) );
  INV_X1 U7169 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n6993) );
  AOI22_X1 U7170 ( .A1(n6140), .A2(DATAO_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6139), .ZN(n6138) );
  OAI21_X1 U7171 ( .B1(n6142), .B2(n6993), .A(n6138), .ZN(U2915) );
  INV_X1 U7172 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6884) );
  AOI22_X1 U7173 ( .A1(n6140), .A2(DATAO_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6139), .ZN(n6141) );
  OAI21_X1 U7174 ( .B1(n6142), .B2(n6884), .A(n6141), .ZN(U2917) );
  AOI22_X1 U7175 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7176 ( .A1(n6146), .A2(DATAI_8_), .ZN(n6148) );
  NAND2_X1 U7177 ( .A1(n6143), .A2(n6148), .ZN(U2932) );
  AOI22_X1 U7178 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7179 ( .A1(n6146), .A2(DATAI_9_), .ZN(n6150) );
  NAND2_X1 U7180 ( .A1(n6144), .A2(n6150), .ZN(U2933) );
  AOI22_X1 U7181 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7182 ( .A1(n6146), .A2(DATAI_11_), .ZN(n6154) );
  NAND2_X1 U7183 ( .A1(n6145), .A2(n6154), .ZN(U2935) );
  AOI22_X1 U7184 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7185 ( .A1(n6146), .A2(DATAI_12_), .ZN(n6156) );
  NAND2_X1 U7186 ( .A1(n6147), .A2(n6156), .ZN(U2936) );
  AOI22_X1 U7187 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7188 ( .A1(n6149), .A2(n6148), .ZN(U2947) );
  AOI22_X1 U7189 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7190 ( .A1(n6151), .A2(n6150), .ZN(U2948) );
  AOI22_X1 U7191 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7192 ( .A1(n6153), .A2(n6152), .ZN(U2949) );
  AOI22_X1 U7193 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7194 ( .A1(n6155), .A2(n6154), .ZN(U2950) );
  AOI22_X1 U7195 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7196 ( .A1(n6157), .A2(n6156), .ZN(U2951) );
  AOI22_X1 U7197 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6159), .B1(n6158), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7198 ( .A1(n6161), .A2(n6160), .ZN(U2952) );
  NAND2_X1 U7199 ( .A1(n6163), .A2(n6162), .ZN(n6166) );
  XNOR2_X1 U7200 ( .A(n6164), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6165)
         );
  XNOR2_X1 U7201 ( .A(n6166), .B(n6165), .ZN(n6203) );
  AOI22_X1 U7202 ( .A1(n6197), .A2(REIP_REG_11__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6188), .ZN(n6171) );
  AOI22_X1 U7203 ( .A1(n6169), .A2(n3103), .B1(n6168), .B2(n6167), .ZN(n6170)
         );
  OAI211_X1 U7204 ( .C1(n6203), .C2(n6172), .A(n6171), .B(n6170), .ZN(U2975)
         );
  AOI22_X1 U7205 ( .A1(n6197), .A2(REIP_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6188), .ZN(n6177) );
  INV_X1 U7206 ( .A(n6173), .ZN(n6175) );
  AOI22_X1 U7207 ( .A1(n6175), .A2(n6191), .B1(n6174), .B2(n3103), .ZN(n6176)
         );
  OAI211_X1 U7208 ( .C1(n6178), .C2(n6195), .A(n6177), .B(n6176), .ZN(U2980)
         );
  AOI22_X1 U7209 ( .A1(n6197), .A2(REIP_REG_4__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6188), .ZN(n6186) );
  OAI21_X1 U7210 ( .B1(n6181), .B2(n6180), .A(n6179), .ZN(n6182) );
  INV_X1 U7211 ( .A(n6182), .ZN(n6257) );
  INV_X1 U7212 ( .A(n6183), .ZN(n6184) );
  AOI22_X1 U7213 ( .A1(n6257), .A2(n6191), .B1(n3103), .B2(n6184), .ZN(n6185)
         );
  OAI211_X1 U7214 ( .C1(n6187), .C2(n6195), .A(n6186), .B(n6185), .ZN(U2982)
         );
  AOI22_X1 U7215 ( .A1(n6197), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6188), .ZN(n6194) );
  INV_X1 U7216 ( .A(n6189), .ZN(n6192) );
  AOI22_X1 U7217 ( .A1(n6192), .A2(n6191), .B1(n3103), .B2(n6190), .ZN(n6193)
         );
  OAI211_X1 U7218 ( .C1(n6196), .C2(n6195), .A(n6194), .B(n6193), .ZN(U2984)
         );
  AOI22_X1 U7219 ( .A1(n6266), .A2(n6198), .B1(n6197), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6202) );
  AOI22_X1 U7220 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6200), .B1(n6199), .B2(n3649), .ZN(n6201) );
  OAI211_X1 U7221 ( .C1(n6203), .C2(n6223), .A(n6202), .B(n6201), .ZN(U3007)
         );
  NOR2_X1 U7222 ( .A1(n6258), .A2(n6204), .ZN(n6234) );
  NAND2_X1 U7223 ( .A1(n6208), .A2(n6234), .ZN(n6221) );
  AOI22_X1 U7224 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n3648), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6967), .ZN(n6213) );
  INV_X1 U7225 ( .A(n6205), .ZN(n6206) );
  AOI21_X1 U7226 ( .B1(n6266), .B2(n6207), .A(n6206), .ZN(n6212) );
  OAI21_X1 U7227 ( .B1(n6209), .B2(n6208), .A(n6238), .ZN(n6217) );
  AOI22_X1 U7228 ( .A1(n6210), .A2(n6269), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6217), .ZN(n6211) );
  OAI211_X1 U7229 ( .C1(n6221), .C2(n6213), .A(n6212), .B(n6211), .ZN(U3008)
         );
  INV_X1 U7230 ( .A(n6214), .ZN(n6215) );
  AOI21_X1 U7231 ( .B1(n6266), .B2(n6216), .A(n6215), .ZN(n6220) );
  AOI22_X1 U7232 ( .A1(n6218), .A2(n6269), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6217), .ZN(n6219) );
  OAI211_X1 U7233 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6221), .A(n6220), 
        .B(n6219), .ZN(U3009) );
  OAI222_X1 U7234 ( .A1(n6224), .A2(n6255), .B1(n6253), .B2(n6619), .C1(n6223), 
        .C2(n6222), .ZN(n6225) );
  INV_X1 U7235 ( .A(n6225), .ZN(n6228) );
  OAI211_X1 U7236 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6234), .B(n6226), .ZN(n6227) );
  OAI211_X1 U7237 ( .C1(n6238), .C2(n6229), .A(n6228), .B(n6227), .ZN(U3010)
         );
  INV_X1 U7238 ( .A(n6230), .ZN(n6231) );
  AOI21_X1 U7239 ( .B1(n6266), .B2(n6232), .A(n6231), .ZN(n6237) );
  INV_X1 U7240 ( .A(n6233), .ZN(n6235) );
  AOI22_X1 U7241 ( .A1(n6235), .A2(n6269), .B1(n6234), .B2(n6913), .ZN(n6236)
         );
  OAI211_X1 U7242 ( .C1(n6238), .C2(n6913), .A(n6237), .B(n6236), .ZN(U3011)
         );
  AOI21_X1 U7243 ( .B1(n6252), .B2(n6239), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6249) );
  INV_X1 U7244 ( .A(n6240), .ZN(n6241) );
  AOI21_X1 U7245 ( .B1(n6266), .B2(n6242), .A(n6241), .ZN(n6248) );
  INV_X1 U7246 ( .A(n6243), .ZN(n6246) );
  NOR2_X1 U7247 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6260), .ZN(n6245)
         );
  AOI22_X1 U7248 ( .A1(n6246), .A2(n6269), .B1(n6245), .B2(n6244), .ZN(n6247)
         );
  OAI211_X1 U7249 ( .C1(n6250), .C2(n6249), .A(n6248), .B(n6247), .ZN(U3013)
         );
  AOI21_X1 U7250 ( .B1(n6252), .B2(n6259), .A(n6251), .ZN(n6274) );
  OAI22_X1 U7251 ( .A1(n6255), .A2(n6254), .B1(n6613), .B2(n6253), .ZN(n6256)
         );
  AOI21_X1 U7252 ( .B1(n6257), .B2(n6269), .A(n6256), .ZN(n6262) );
  NOR2_X1 U7253 ( .A1(n6259), .A2(n6258), .ZN(n6270) );
  OAI211_X1 U7254 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6270), .B(n6260), .ZN(n6261) );
  OAI211_X1 U7255 ( .C1(n6274), .C2(n6263), .A(n6262), .B(n6261), .ZN(U3014)
         );
  AOI21_X1 U7256 ( .B1(n6266), .B2(n6265), .A(n6264), .ZN(n6272) );
  INV_X1 U7257 ( .A(n6267), .ZN(n6268) );
  AOI22_X1 U7258 ( .A1(n6270), .A2(n6273), .B1(n6269), .B2(n6268), .ZN(n6271)
         );
  OAI211_X1 U7259 ( .C1(n6274), .C2(n6273), .A(n6272), .B(n6271), .ZN(U3015)
         );
  NOR2_X1 U7260 ( .A1(n6276), .A2(n6275), .ZN(U3019) );
  NAND2_X1 U7261 ( .A1(n6354), .A2(n6277), .ZN(n6313) );
  NAND2_X1 U7262 ( .A1(n6278), .A2(n6359), .ZN(n6433) );
  OAI22_X1 U7263 ( .A1(n6313), .A2(n6527), .B1(n6444), .B2(n6433), .ZN(n6300)
         );
  NAND3_X1 U7264 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6359), .A3(n6279), .ZN(n6317) );
  NOR2_X1 U7265 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6317), .ZN(n6299)
         );
  AOI22_X1 U7266 ( .A1(n6437), .A2(n6300), .B1(n6522), .B2(n6299), .ZN(n6286)
         );
  INV_X1 U7267 ( .A(n6348), .ZN(n6281) );
  OAI21_X1 U7268 ( .B1(n6281), .B2(n6301), .A(n6280), .ZN(n6282) );
  AOI21_X1 U7269 ( .B1(n6282), .B2(n6313), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6284) );
  AOI22_X1 U7270 ( .A1(n6302), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6531), 
        .B2(n6301), .ZN(n6285) );
  OAI211_X1 U7271 ( .C1(n6449), .C2(n6348), .A(n6286), .B(n6285), .ZN(U3036)
         );
  AOI22_X1 U7272 ( .A1(n6450), .A2(n6300), .B1(n6535), .B2(n6299), .ZN(n6288)
         );
  AOI22_X1 U7273 ( .A1(n6302), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6537), 
        .B2(n6301), .ZN(n6287) );
  OAI211_X1 U7274 ( .C1(n6348), .C2(n6453), .A(n6288), .B(n6287), .ZN(U3037)
         );
  AOI22_X1 U7275 ( .A1(n6454), .A2(n6300), .B1(n6541), .B2(n6299), .ZN(n6290)
         );
  AOI22_X1 U7276 ( .A1(n6302), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6542), 
        .B2(n6301), .ZN(n6289) );
  OAI211_X1 U7277 ( .C1(n6348), .C2(n6457), .A(n6290), .B(n6289), .ZN(U3038)
         );
  AOI22_X1 U7278 ( .A1(n6458), .A2(n6300), .B1(n6547), .B2(n6299), .ZN(n6292)
         );
  AOI22_X1 U7279 ( .A1(n6302), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6549), 
        .B2(n6301), .ZN(n6291) );
  OAI211_X1 U7280 ( .C1(n6348), .C2(n6461), .A(n6292), .B(n6291), .ZN(U3039)
         );
  AOI22_X1 U7281 ( .A1(n6462), .A2(n6300), .B1(n6553), .B2(n6299), .ZN(n6294)
         );
  AOI22_X1 U7282 ( .A1(n6302), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6554), 
        .B2(n6301), .ZN(n6293) );
  OAI211_X1 U7283 ( .C1(n6348), .C2(n6465), .A(n6294), .B(n6293), .ZN(U3040)
         );
  AOI22_X1 U7284 ( .A1(n6466), .A2(n6300), .B1(n6559), .B2(n6299), .ZN(n6296)
         );
  AOI22_X1 U7285 ( .A1(n6302), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6560), 
        .B2(n6301), .ZN(n6295) );
  OAI211_X1 U7286 ( .C1(n6348), .C2(n6469), .A(n6296), .B(n6295), .ZN(U3041)
         );
  AOI22_X1 U7287 ( .A1(n6470), .A2(n6300), .B1(n6565), .B2(n6299), .ZN(n6298)
         );
  AOI22_X1 U7288 ( .A1(n6302), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6567), 
        .B2(n6301), .ZN(n6297) );
  OAI211_X1 U7289 ( .C1(n6348), .C2(n6473), .A(n6298), .B(n6297), .ZN(U3042)
         );
  AOI22_X1 U7290 ( .A1(n6476), .A2(n6300), .B1(n6572), .B2(n6299), .ZN(n6304)
         );
  AOI22_X1 U7291 ( .A1(n6302), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6573), 
        .B2(n6301), .ZN(n6303) );
  OAI211_X1 U7292 ( .C1(n6348), .C2(n6482), .A(n6304), .B(n6303), .ZN(U3043)
         );
  INV_X1 U7293 ( .A(n6305), .ZN(n6306) );
  INV_X1 U7294 ( .A(n6308), .ZN(n6518) );
  NAND2_X1 U7295 ( .A1(n6518), .A2(n6359), .ZN(n6346) );
  OAI22_X1 U7296 ( .A1(n6348), .A2(n6371), .B1(n6309), .B2(n6346), .ZN(n6310)
         );
  INV_X1 U7297 ( .A(n6310), .ZN(n6321) );
  NAND2_X1 U7298 ( .A1(n6515), .A2(n4782), .ZN(n6311) );
  OAI21_X1 U7299 ( .B1(n6312), .B2(n6311), .A(n6409), .ZN(n6319) );
  OR2_X1 U7300 ( .A1(n6313), .A2(n6484), .ZN(n6314) );
  AND2_X1 U7301 ( .A1(n6314), .A2(n6346), .ZN(n6318) );
  INV_X1 U7302 ( .A(n6318), .ZN(n6316) );
  AOI21_X1 U7303 ( .B1(n6527), .B2(n6317), .A(n6525), .ZN(n6315) );
  OAI21_X1 U7304 ( .B1(n6319), .B2(n6316), .A(n6315), .ZN(n6351) );
  OAI22_X1 U7305 ( .A1(n6319), .A2(n6318), .B1(n6317), .B2(n6695), .ZN(n6350)
         );
  AOI22_X1 U7306 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6351), .B1(n6437), 
        .B2(n6350), .ZN(n6320) );
  OAI211_X1 U7307 ( .C1(n6449), .C2(n6395), .A(n6321), .B(n6320), .ZN(U3044)
         );
  OAI22_X1 U7308 ( .A1(n6348), .A2(n6374), .B1(n6322), .B2(n6346), .ZN(n6323)
         );
  INV_X1 U7309 ( .A(n6323), .ZN(n6325) );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6351), .B1(n6450), 
        .B2(n6350), .ZN(n6324) );
  OAI211_X1 U7311 ( .C1(n6453), .C2(n6395), .A(n6325), .B(n6324), .ZN(U3045)
         );
  OAI22_X1 U7312 ( .A1(n6348), .A2(n6377), .B1(n6326), .B2(n6346), .ZN(n6327)
         );
  INV_X1 U7313 ( .A(n6327), .ZN(n6329) );
  AOI22_X1 U7314 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6351), .B1(n6454), 
        .B2(n6350), .ZN(n6328) );
  OAI211_X1 U7315 ( .C1(n6457), .C2(n6395), .A(n6329), .B(n6328), .ZN(U3046)
         );
  OAI22_X1 U7316 ( .A1(n6348), .A2(n6380), .B1(n6330), .B2(n6346), .ZN(n6331)
         );
  INV_X1 U7317 ( .A(n6331), .ZN(n6333) );
  AOI22_X1 U7318 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6351), .B1(n6458), 
        .B2(n6350), .ZN(n6332) );
  OAI211_X1 U7319 ( .C1(n6461), .C2(n6395), .A(n6333), .B(n6332), .ZN(U3047)
         );
  OAI22_X1 U7320 ( .A1(n6348), .A2(n6383), .B1(n6334), .B2(n6346), .ZN(n6335)
         );
  INV_X1 U7321 ( .A(n6335), .ZN(n6337) );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6351), .B1(n6462), 
        .B2(n6350), .ZN(n6336) );
  OAI211_X1 U7323 ( .C1(n6465), .C2(n6395), .A(n6337), .B(n6336), .ZN(U3048)
         );
  OAI22_X1 U7324 ( .A1(n6348), .A2(n6386), .B1(n6338), .B2(n6346), .ZN(n6339)
         );
  INV_X1 U7325 ( .A(n6339), .ZN(n6341) );
  AOI22_X1 U7326 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6351), .B1(n6466), 
        .B2(n6350), .ZN(n6340) );
  OAI211_X1 U7327 ( .C1(n6469), .C2(n6395), .A(n6341), .B(n6340), .ZN(U3049)
         );
  OAI22_X1 U7328 ( .A1(n6348), .A2(n6389), .B1(n6342), .B2(n6346), .ZN(n6343)
         );
  INV_X1 U7329 ( .A(n6343), .ZN(n6345) );
  AOI22_X1 U7330 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6351), .B1(n6470), 
        .B2(n6350), .ZN(n6344) );
  OAI211_X1 U7331 ( .C1(n6473), .C2(n6395), .A(n6345), .B(n6344), .ZN(U3050)
         );
  OAI22_X1 U7332 ( .A1(n6348), .A2(n6396), .B1(n6347), .B2(n6346), .ZN(n6349)
         );
  INV_X1 U7333 ( .A(n6349), .ZN(n6353) );
  AOI22_X1 U7334 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6351), .B1(n6476), 
        .B2(n6350), .ZN(n6352) );
  OAI211_X1 U7335 ( .C1(n6482), .C2(n6395), .A(n6353), .B(n6352), .ZN(U3051)
         );
  NAND2_X1 U7336 ( .A1(n6354), .A2(n6409), .ZN(n6436) );
  INV_X1 U7337 ( .A(n6362), .ZN(n6357) );
  INV_X1 U7338 ( .A(n6355), .ZN(n6434) );
  OAI22_X1 U7339 ( .A1(n6436), .A2(n6357), .B1(n6434), .B2(n6356), .ZN(n6391)
         );
  NAND3_X1 U7340 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6359), .A3(n6358), .ZN(n6401) );
  NOR2_X1 U7341 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6401), .ZN(n6390)
         );
  AOI22_X1 U7342 ( .A1(n6437), .A2(n6391), .B1(n6522), .B2(n6390), .ZN(n6370)
         );
  INV_X1 U7343 ( .A(n6432), .ZN(n6361) );
  AOI21_X1 U7344 ( .B1(n6361), .B2(n6360), .A(n6527), .ZN(n6405) );
  NAND2_X1 U7345 ( .A1(n6362), .A2(n6438), .ZN(n6397) );
  OAI211_X1 U7346 ( .C1(n6395), .C2(n6440), .A(n6405), .B(n6397), .ZN(n6367)
         );
  INV_X1 U7347 ( .A(n6390), .ZN(n6365) );
  AOI211_X1 U7348 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6365), .A(n6364), .B(
        n6363), .ZN(n6366) );
  NAND2_X1 U7349 ( .A1(n6367), .A2(n6366), .ZN(n6392) );
  NOR2_X2 U7350 ( .A1(n6432), .A2(n6368), .ZN(n6425) );
  AOI22_X1 U7351 ( .A1(n6392), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6523), 
        .B2(n6425), .ZN(n6369) );
  OAI211_X1 U7352 ( .C1(n6371), .C2(n6395), .A(n6370), .B(n6369), .ZN(U3052)
         );
  AOI22_X1 U7353 ( .A1(n6450), .A2(n6391), .B1(n6535), .B2(n6390), .ZN(n6373)
         );
  AOI22_X1 U7354 ( .A1(n6392), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6536), 
        .B2(n6425), .ZN(n6372) );
  OAI211_X1 U7355 ( .C1(n6374), .C2(n6395), .A(n6373), .B(n6372), .ZN(U3053)
         );
  AOI22_X1 U7356 ( .A1(n6454), .A2(n6391), .B1(n6541), .B2(n6390), .ZN(n6376)
         );
  AOI22_X1 U7357 ( .A1(n6392), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6543), 
        .B2(n6425), .ZN(n6375) );
  OAI211_X1 U7358 ( .C1(n6377), .C2(n6395), .A(n6376), .B(n6375), .ZN(U3054)
         );
  AOI22_X1 U7359 ( .A1(n6458), .A2(n6391), .B1(n6547), .B2(n6390), .ZN(n6379)
         );
  AOI22_X1 U7360 ( .A1(n6392), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6548), 
        .B2(n6425), .ZN(n6378) );
  OAI211_X1 U7361 ( .C1(n6380), .C2(n6395), .A(n6379), .B(n6378), .ZN(U3055)
         );
  AOI22_X1 U7362 ( .A1(n6462), .A2(n6391), .B1(n6553), .B2(n6390), .ZN(n6382)
         );
  AOI22_X1 U7363 ( .A1(n6392), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6555), 
        .B2(n6425), .ZN(n6381) );
  OAI211_X1 U7364 ( .C1(n6383), .C2(n6395), .A(n6382), .B(n6381), .ZN(U3056)
         );
  AOI22_X1 U7365 ( .A1(n6466), .A2(n6391), .B1(n6559), .B2(n6390), .ZN(n6385)
         );
  AOI22_X1 U7366 ( .A1(n6392), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6561), 
        .B2(n6425), .ZN(n6384) );
  OAI211_X1 U7367 ( .C1(n6386), .C2(n6395), .A(n6385), .B(n6384), .ZN(U3057)
         );
  AOI22_X1 U7368 ( .A1(n6470), .A2(n6391), .B1(n6565), .B2(n6390), .ZN(n6388)
         );
  AOI22_X1 U7369 ( .A1(n6392), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6566), 
        .B2(n6425), .ZN(n6387) );
  OAI211_X1 U7370 ( .C1(n6389), .C2(n6395), .A(n6388), .B(n6387), .ZN(U3058)
         );
  AOI22_X1 U7371 ( .A1(n6476), .A2(n6391), .B1(n6572), .B2(n6390), .ZN(n6394)
         );
  AOI22_X1 U7372 ( .A1(n6392), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6576), 
        .B2(n6425), .ZN(n6393) );
  OAI211_X1 U7373 ( .C1(n6396), .C2(n6395), .A(n6394), .B(n6393), .ZN(U3059)
         );
  OR2_X1 U7374 ( .A1(n6397), .A2(n6484), .ZN(n6400) );
  NOR2_X1 U7375 ( .A1(n6398), .A2(n6401), .ZN(n6424) );
  INV_X1 U7376 ( .A(n6424), .ZN(n6399) );
  INV_X1 U7377 ( .A(n6404), .ZN(n6402) );
  INV_X1 U7378 ( .A(n6401), .ZN(n6408) );
  AOI22_X1 U7379 ( .A1(n6477), .A2(n6523), .B1(n6522), .B2(n6424), .ZN(n6411)
         );
  NAND2_X1 U7380 ( .A1(n6405), .A2(n6404), .ZN(n6407) );
  OAI211_X1 U7381 ( .C1(n6409), .C2(n6408), .A(n6407), .B(n6406), .ZN(n6426)
         );
  AOI22_X1 U7382 ( .A1(n6426), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n6531), 
        .B2(n6425), .ZN(n6410) );
  OAI211_X1 U7383 ( .C1(n6429), .C2(n6534), .A(n6411), .B(n6410), .ZN(U3060)
         );
  AOI22_X1 U7384 ( .A1(n6477), .A2(n6536), .B1(n6535), .B2(n6424), .ZN(n6413)
         );
  AOI22_X1 U7385 ( .A1(n6426), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n6537), 
        .B2(n6425), .ZN(n6412) );
  OAI211_X1 U7386 ( .C1(n6429), .C2(n6540), .A(n6413), .B(n6412), .ZN(U3061)
         );
  AOI22_X1 U7387 ( .A1(n6477), .A2(n6543), .B1(n6541), .B2(n6424), .ZN(n6415)
         );
  AOI22_X1 U7388 ( .A1(n6426), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n6542), 
        .B2(n6425), .ZN(n6414) );
  OAI211_X1 U7389 ( .C1(n6429), .C2(n6546), .A(n6415), .B(n6414), .ZN(U3062)
         );
  AOI22_X1 U7390 ( .A1(n6477), .A2(n6548), .B1(n6547), .B2(n6424), .ZN(n6417)
         );
  AOI22_X1 U7391 ( .A1(n6426), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n6549), 
        .B2(n6425), .ZN(n6416) );
  OAI211_X1 U7392 ( .C1(n6429), .C2(n6552), .A(n6417), .B(n6416), .ZN(U3063)
         );
  AOI22_X1 U7393 ( .A1(n6477), .A2(n6555), .B1(n6553), .B2(n6424), .ZN(n6419)
         );
  AOI22_X1 U7394 ( .A1(n6426), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n6554), 
        .B2(n6425), .ZN(n6418) );
  OAI211_X1 U7395 ( .C1(n6429), .C2(n6558), .A(n6419), .B(n6418), .ZN(U3064)
         );
  AOI22_X1 U7396 ( .A1(n6477), .A2(n6561), .B1(n6559), .B2(n6424), .ZN(n6421)
         );
  AOI22_X1 U7397 ( .A1(n6426), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n6560), 
        .B2(n6425), .ZN(n6420) );
  OAI211_X1 U7398 ( .C1(n6429), .C2(n6564), .A(n6421), .B(n6420), .ZN(U3065)
         );
  AOI22_X1 U7399 ( .A1(n6477), .A2(n6566), .B1(n6565), .B2(n6424), .ZN(n6423)
         );
  AOI22_X1 U7400 ( .A1(n6426), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n6567), 
        .B2(n6425), .ZN(n6422) );
  OAI211_X1 U7401 ( .C1(n6429), .C2(n6570), .A(n6423), .B(n6422), .ZN(U3066)
         );
  AOI22_X1 U7402 ( .A1(n6477), .A2(n6576), .B1(n6572), .B2(n6424), .ZN(n6428)
         );
  AOI22_X1 U7403 ( .A1(n6426), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n6573), 
        .B2(n6425), .ZN(n6427) );
  OAI211_X1 U7404 ( .C1(n6429), .C2(n6580), .A(n6428), .B(n6427), .ZN(U3067)
         );
  INV_X1 U7405 ( .A(n6430), .ZN(n6431) );
  OAI22_X1 U7406 ( .A1(n6436), .A2(n6435), .B1(n6434), .B2(n6433), .ZN(n6475)
         );
  NOR2_X1 U7407 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6490), .ZN(n6474)
         );
  AOI22_X1 U7408 ( .A1(n6437), .A2(n6475), .B1(n6522), .B2(n6474), .ZN(n6448)
         );
  NOR3_X1 U7409 ( .A1(n6510), .A2(n6477), .A3(n6527), .ZN(n6441) );
  NAND2_X1 U7410 ( .A1(n6439), .A2(n6438), .ZN(n6485) );
  OAI21_X1 U7411 ( .B1(n6441), .B2(n6440), .A(n6485), .ZN(n6446) );
  INV_X1 U7412 ( .A(n6474), .ZN(n6443) );
  AOI211_X1 U7413 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6443), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6442), .ZN(n6445) );
  NAND3_X1 U7414 ( .A1(n6446), .A2(n6445), .A3(n6444), .ZN(n6478) );
  AOI22_X1 U7415 ( .A1(n6478), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6531), 
        .B2(n6477), .ZN(n6447) );
  OAI211_X1 U7416 ( .C1(n6449), .C2(n6481), .A(n6448), .B(n6447), .ZN(U3068)
         );
  AOI22_X1 U7417 ( .A1(n6450), .A2(n6475), .B1(n6535), .B2(n6474), .ZN(n6452)
         );
  AOI22_X1 U7418 ( .A1(n6478), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6537), 
        .B2(n6477), .ZN(n6451) );
  OAI211_X1 U7419 ( .C1(n6453), .C2(n6481), .A(n6452), .B(n6451), .ZN(U3069)
         );
  AOI22_X1 U7420 ( .A1(n6454), .A2(n6475), .B1(n6541), .B2(n6474), .ZN(n6456)
         );
  AOI22_X1 U7421 ( .A1(n6478), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6542), 
        .B2(n6477), .ZN(n6455) );
  OAI211_X1 U7422 ( .C1(n6457), .C2(n6481), .A(n6456), .B(n6455), .ZN(U3070)
         );
  AOI22_X1 U7423 ( .A1(n6458), .A2(n6475), .B1(n6547), .B2(n6474), .ZN(n6460)
         );
  AOI22_X1 U7424 ( .A1(n6478), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6549), 
        .B2(n6477), .ZN(n6459) );
  OAI211_X1 U7425 ( .C1(n6461), .C2(n6481), .A(n6460), .B(n6459), .ZN(U3071)
         );
  AOI22_X1 U7426 ( .A1(n6462), .A2(n6475), .B1(n6553), .B2(n6474), .ZN(n6464)
         );
  AOI22_X1 U7427 ( .A1(n6478), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6554), 
        .B2(n6477), .ZN(n6463) );
  OAI211_X1 U7428 ( .C1(n6465), .C2(n6481), .A(n6464), .B(n6463), .ZN(U3072)
         );
  AOI22_X1 U7429 ( .A1(n6466), .A2(n6475), .B1(n6559), .B2(n6474), .ZN(n6468)
         );
  AOI22_X1 U7430 ( .A1(n6478), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6560), 
        .B2(n6477), .ZN(n6467) );
  OAI211_X1 U7431 ( .C1(n6469), .C2(n6481), .A(n6468), .B(n6467), .ZN(U3073)
         );
  AOI22_X1 U7432 ( .A1(n6470), .A2(n6475), .B1(n6565), .B2(n6474), .ZN(n6472)
         );
  AOI22_X1 U7433 ( .A1(n6478), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6567), 
        .B2(n6477), .ZN(n6471) );
  OAI211_X1 U7434 ( .C1(n6473), .C2(n6481), .A(n6472), .B(n6471), .ZN(U3074)
         );
  AOI22_X1 U7435 ( .A1(n6476), .A2(n6475), .B1(n6572), .B2(n6474), .ZN(n6480)
         );
  AOI22_X1 U7436 ( .A1(n6478), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6573), 
        .B2(n6477), .ZN(n6479) );
  OAI211_X1 U7437 ( .C1(n6482), .C2(n6481), .A(n6480), .B(n6479), .ZN(U3075)
         );
  NOR2_X1 U7438 ( .A1(n6483), .A2(n6527), .ZN(n6489) );
  OR2_X1 U7439 ( .A1(n6485), .A2(n6484), .ZN(n6486) );
  NAND2_X1 U7440 ( .A1(n6486), .A2(n6488), .ZN(n6492) );
  INV_X1 U7441 ( .A(n6488), .ZN(n6508) );
  AOI22_X1 U7442 ( .A1(n6509), .A2(n6523), .B1(n6522), .B2(n6508), .ZN(n6495)
         );
  INV_X1 U7443 ( .A(n6489), .ZN(n6493) );
  AOI21_X1 U7444 ( .B1(n6527), .B2(n6490), .A(n6525), .ZN(n6491) );
  AOI22_X1 U7445 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6511), .B1(n6531), 
        .B2(n6510), .ZN(n6494) );
  OAI211_X1 U7446 ( .C1(n6514), .C2(n6534), .A(n6495), .B(n6494), .ZN(U3076)
         );
  AOI22_X1 U7447 ( .A1(n6509), .A2(n6536), .B1(n6535), .B2(n6508), .ZN(n6497)
         );
  AOI22_X1 U7448 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6511), .B1(n6537), 
        .B2(n6510), .ZN(n6496) );
  OAI211_X1 U7449 ( .C1(n6514), .C2(n6540), .A(n6497), .B(n6496), .ZN(U3077)
         );
  AOI22_X1 U7450 ( .A1(n6509), .A2(n6543), .B1(n6541), .B2(n6508), .ZN(n6499)
         );
  AOI22_X1 U7451 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6511), .B1(n6542), 
        .B2(n6510), .ZN(n6498) );
  OAI211_X1 U7452 ( .C1(n6514), .C2(n6546), .A(n6499), .B(n6498), .ZN(U3078)
         );
  AOI22_X1 U7453 ( .A1(n6510), .A2(n6549), .B1(n6547), .B2(n6508), .ZN(n6501)
         );
  AOI22_X1 U7454 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6511), .B1(n6548), 
        .B2(n6509), .ZN(n6500) );
  OAI211_X1 U7455 ( .C1(n6514), .C2(n6552), .A(n6501), .B(n6500), .ZN(U3079)
         );
  AOI22_X1 U7456 ( .A1(n6510), .A2(n6554), .B1(n6553), .B2(n6508), .ZN(n6503)
         );
  AOI22_X1 U7457 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6511), .B1(n6555), 
        .B2(n6509), .ZN(n6502) );
  OAI211_X1 U7458 ( .C1(n6514), .C2(n6558), .A(n6503), .B(n6502), .ZN(U3080)
         );
  AOI22_X1 U7459 ( .A1(n6509), .A2(n6561), .B1(n6559), .B2(n6508), .ZN(n6505)
         );
  AOI22_X1 U7460 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6511), .B1(n6560), 
        .B2(n6510), .ZN(n6504) );
  OAI211_X1 U7461 ( .C1(n6514), .C2(n6564), .A(n6505), .B(n6504), .ZN(U3081)
         );
  AOI22_X1 U7462 ( .A1(n6510), .A2(n6567), .B1(n6565), .B2(n6508), .ZN(n6507)
         );
  AOI22_X1 U7463 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6511), .B1(n6566), 
        .B2(n6509), .ZN(n6506) );
  OAI211_X1 U7464 ( .C1(n6514), .C2(n6570), .A(n6507), .B(n6506), .ZN(U3082)
         );
  AOI22_X1 U7465 ( .A1(n6509), .A2(n6576), .B1(n6572), .B2(n6508), .ZN(n6513)
         );
  AOI22_X1 U7466 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6511), .B1(n6573), 
        .B2(n6510), .ZN(n6512) );
  OAI211_X1 U7467 ( .C1(n6514), .C2(n6580), .A(n6513), .B(n6512), .ZN(U3083)
         );
  AOI21_X1 U7468 ( .B1(n6516), .B2(n6515), .A(n6527), .ZN(n6524) );
  NAND2_X1 U7469 ( .A1(n6517), .A2(n3130), .ZN(n6519) );
  NAND2_X1 U7470 ( .A1(n6518), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U7471 ( .A1(n6519), .A2(n6521), .ZN(n6529) );
  INV_X1 U7472 ( .A(n6526), .ZN(n6520) );
  INV_X1 U7473 ( .A(n6521), .ZN(n6571) );
  AOI22_X1 U7474 ( .A1(n6575), .A2(n6523), .B1(n6522), .B2(n6571), .ZN(n6533)
         );
  INV_X1 U7475 ( .A(n6524), .ZN(n6530) );
  AOI21_X1 U7476 ( .B1(n6527), .B2(n6526), .A(n6525), .ZN(n6528) );
  AOI22_X1 U7477 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6577), .B1(n6531), 
        .B2(n6574), .ZN(n6532) );
  OAI211_X1 U7478 ( .C1(n6581), .C2(n6534), .A(n6533), .B(n6532), .ZN(U3108)
         );
  AOI22_X1 U7479 ( .A1(n6575), .A2(n6536), .B1(n6535), .B2(n6571), .ZN(n6539)
         );
  AOI22_X1 U7480 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6577), .B1(n6537), 
        .B2(n6574), .ZN(n6538) );
  OAI211_X1 U7481 ( .C1(n6581), .C2(n6540), .A(n6539), .B(n6538), .ZN(U3109)
         );
  AOI22_X1 U7482 ( .A1(n6574), .A2(n6542), .B1(n6541), .B2(n6571), .ZN(n6545)
         );
  AOI22_X1 U7483 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6577), .B1(n6543), 
        .B2(n6575), .ZN(n6544) );
  OAI211_X1 U7484 ( .C1(n6581), .C2(n6546), .A(n6545), .B(n6544), .ZN(U3110)
         );
  AOI22_X1 U7485 ( .A1(n6575), .A2(n6548), .B1(n6547), .B2(n6571), .ZN(n6551)
         );
  AOI22_X1 U7486 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6577), .B1(n6549), 
        .B2(n6574), .ZN(n6550) );
  OAI211_X1 U7487 ( .C1(n6581), .C2(n6552), .A(n6551), .B(n6550), .ZN(U3111)
         );
  AOI22_X1 U7488 ( .A1(n6574), .A2(n6554), .B1(n6553), .B2(n6571), .ZN(n6557)
         );
  AOI22_X1 U7489 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6577), .B1(n6555), 
        .B2(n6575), .ZN(n6556) );
  OAI211_X1 U7490 ( .C1(n6581), .C2(n6558), .A(n6557), .B(n6556), .ZN(U3112)
         );
  AOI22_X1 U7491 ( .A1(n6574), .A2(n6560), .B1(n6559), .B2(n6571), .ZN(n6563)
         );
  AOI22_X1 U7492 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6577), .B1(n6561), 
        .B2(n6575), .ZN(n6562) );
  OAI211_X1 U7493 ( .C1(n6581), .C2(n6564), .A(n6563), .B(n6562), .ZN(U3113)
         );
  AOI22_X1 U7494 ( .A1(n6575), .A2(n6566), .B1(n6565), .B2(n6571), .ZN(n6569)
         );
  AOI22_X1 U7495 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6577), .B1(n6567), 
        .B2(n6574), .ZN(n6568) );
  OAI211_X1 U7496 ( .C1(n6581), .C2(n6570), .A(n6569), .B(n6568), .ZN(U3114)
         );
  AOI22_X1 U7497 ( .A1(n6574), .A2(n6573), .B1(n6572), .B2(n6571), .ZN(n6579)
         );
  AOI22_X1 U7498 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6577), .B1(n6576), 
        .B2(n6575), .ZN(n6578) );
  OAI211_X1 U7499 ( .C1(n6581), .C2(n6580), .A(n6579), .B(n6578), .ZN(U3115)
         );
  OAI21_X1 U7500 ( .B1(READY_N), .B2(n6583), .A(n6582), .ZN(n6586) );
  AOI211_X1 U7501 ( .C1(n6664), .C2(n6588), .A(n6591), .B(n6981), .ZN(n6584)
         );
  AOI211_X1 U7502 ( .C1(n6664), .C2(n6586), .A(n6585), .B(n6584), .ZN(n6587)
         );
  INV_X1 U7503 ( .A(n6587), .ZN(U3149) );
  NAND3_X1 U7504 ( .A1(n6589), .A2(n6588), .A3(n6662), .ZN(n6590) );
  OAI22_X1 U7505 ( .A1(n6591), .A2(n6590), .B1(n6694), .B2(n6703), .ZN(U3150)
         );
  AND2_X1 U7506 ( .A1(n6592), .A2(DATAWIDTH_REG_31__SCAN_IN), .ZN(U3151) );
  AND2_X1 U7507 ( .A1(n6592), .A2(DATAWIDTH_REG_30__SCAN_IN), .ZN(U3152) );
  AND2_X1 U7508 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6592), .ZN(U3153) );
  AND2_X1 U7509 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6592), .ZN(U3154) );
  AND2_X1 U7510 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6592), .ZN(U3155) );
  AND2_X1 U7511 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6592), .ZN(U3156) );
  AND2_X1 U7512 ( .A1(n6592), .A2(DATAWIDTH_REG_25__SCAN_IN), .ZN(U3157) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6592), .ZN(U3158) );
  AND2_X1 U7514 ( .A1(n6592), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7515 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6592), .ZN(U3160) );
  AND2_X1 U7516 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6592), .ZN(U3161) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6592), .ZN(U3162) );
  AND2_X1 U7518 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6592), .ZN(U3163) );
  AND2_X1 U7519 ( .A1(n6592), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  AND2_X1 U7520 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6592), .ZN(U3165) );
  AND2_X1 U7521 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6592), .ZN(U3166) );
  AND2_X1 U7522 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6592), .ZN(U3167) );
  AND2_X1 U7523 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6592), .ZN(U3168) );
  AND2_X1 U7524 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6592), .ZN(U3169) );
  AND2_X1 U7525 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6592), .ZN(U3170) );
  AND2_X1 U7526 ( .A1(n6592), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(U3171) );
  AND2_X1 U7527 ( .A1(n6592), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  AND2_X1 U7528 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6592), .ZN(U3173) );
  AND2_X1 U7529 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6592), .ZN(U3174) );
  AND2_X1 U7530 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6592), .ZN(U3175) );
  AND2_X1 U7531 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6592), .ZN(U3176) );
  AND2_X1 U7532 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6592), .ZN(U3177) );
  AND2_X1 U7533 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6592), .ZN(U3178) );
  AND2_X1 U7534 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6592), .ZN(U3179) );
  AND2_X1 U7535 ( .A1(n6592), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  INV_X1 U7536 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6598) );
  NOR2_X1 U7537 ( .A1(n6608), .A2(n6598), .ZN(n6599) );
  AOI22_X1 U7538 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6607) );
  AND2_X1 U7539 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6596) );
  INV_X1 U7540 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6594) );
  INV_X1 U7541 ( .A(NA_N), .ZN(n6600) );
  AOI221_X1 U7542 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6600), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6604) );
  AOI221_X1 U7543 ( .B1(n6596), .B2(n6700), .C1(n6594), .C2(n6700), .A(n6604), 
        .ZN(n6593) );
  OAI21_X1 U7544 ( .B1(n6599), .B2(n6607), .A(n6593), .ZN(U3181) );
  NOR2_X1 U7545 ( .A1(n6602), .A2(n6594), .ZN(n6601) );
  NAND2_X1 U7546 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6595) );
  OAI21_X1 U7547 ( .B1(n6601), .B2(n6596), .A(n6595), .ZN(n6597) );
  OAI211_X1 U7548 ( .C1(n6598), .C2(n6690), .A(n6689), .B(n6597), .ZN(U3182)
         );
  AOI21_X1 U7549 ( .B1(n6601), .B2(n6600), .A(n6599), .ZN(n6606) );
  AOI221_X1 U7550 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6690), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6603) );
  AOI221_X1 U7551 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6603), .C2(HOLD), .A(n6602), .ZN(n6605) );
  OAI22_X1 U7552 ( .A1(n6607), .A2(n6606), .B1(n6605), .B2(n6604), .ZN(U3183)
         );
  NOR2_X2 U7553 ( .A1(n6608), .A2(n6700), .ZN(n6650) );
  NAND2_X1 U7554 ( .A1(n6608), .A2(n6684), .ZN(n6652) );
  INV_X1 U7555 ( .A(n6652), .ZN(n6653) );
  AOI22_X1 U7556 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6700), .ZN(n6609) );
  OAI21_X1 U7557 ( .B1(n6980), .B2(n6655), .A(n6609), .ZN(U3184) );
  AOI22_X1 U7558 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6650), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6700), .ZN(n6610) );
  OAI21_X1 U7559 ( .B1(n4829), .B2(n6652), .A(n6610), .ZN(U3185) );
  AOI222_X1 U7560 ( .A1(n6650), .A2(REIP_REG_3__SCAN_IN), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6700), .C1(REIP_REG_4__SCAN_IN), .C2(
        n6653), .ZN(n6611) );
  INV_X1 U7561 ( .A(n6611), .ZN(U3186) );
  AOI22_X1 U7562 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6700), .ZN(n6612) );
  OAI21_X1 U7563 ( .B1(n6613), .B2(n6655), .A(n6612), .ZN(U3187) );
  AOI22_X1 U7564 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6700), .ZN(n6614) );
  OAI21_X1 U7565 ( .B1(n6615), .B2(n6655), .A(n6614), .ZN(U3188) );
  AOI222_X1 U7566 ( .A1(n6650), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6700), .C1(REIP_REG_7__SCAN_IN), .C2(
        n6653), .ZN(n6616) );
  INV_X1 U7567 ( .A(n6616), .ZN(U3189) );
  AOI222_X1 U7568 ( .A1(n6650), .A2(REIP_REG_7__SCAN_IN), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6700), .C1(REIP_REG_8__SCAN_IN), .C2(
        n6653), .ZN(n6617) );
  INV_X1 U7569 ( .A(n6617), .ZN(U3190) );
  AOI22_X1 U7570 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6700), .ZN(n6618) );
  OAI21_X1 U7571 ( .B1(n6619), .B2(n6655), .A(n6618), .ZN(U3191) );
  AOI22_X1 U7572 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6700), .ZN(n6620) );
  OAI21_X1 U7573 ( .B1(n6621), .B2(n6655), .A(n6620), .ZN(U3192) );
  INV_X1 U7574 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6623) );
  AOI22_X1 U7575 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6700), .ZN(n6622) );
  OAI21_X1 U7576 ( .B1(n6623), .B2(n6655), .A(n6622), .ZN(U3193) );
  AOI22_X1 U7577 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6650), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6700), .ZN(n6624) );
  OAI21_X1 U7578 ( .B1(n6626), .B2(n6652), .A(n6624), .ZN(U3194) );
  AOI22_X1 U7579 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6700), .ZN(n6625) );
  OAI21_X1 U7580 ( .B1(n6626), .B2(n6655), .A(n6625), .ZN(U3195) );
  AOI22_X1 U7581 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6650), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6700), .ZN(n6627) );
  OAI21_X1 U7582 ( .B1(n6628), .B2(n6652), .A(n6627), .ZN(U3196) );
  AOI22_X1 U7583 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6650), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6700), .ZN(n6629) );
  OAI21_X1 U7584 ( .B1(n6717), .B2(n6652), .A(n6629), .ZN(U3197) );
  INV_X1 U7585 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6631) );
  INV_X1 U7586 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6969) );
  OAI222_X1 U7587 ( .A1(n6652), .A2(n6631), .B1(n6969), .B2(n6684), .C1(n6717), 
        .C2(n6655), .ZN(U3198) );
  AOI22_X1 U7588 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6700), .ZN(n6630) );
  OAI21_X1 U7589 ( .B1(n6631), .B2(n6655), .A(n6630), .ZN(U3199) );
  AOI22_X1 U7590 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6650), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6700), .ZN(n6632) );
  OAI21_X1 U7591 ( .B1(n6633), .B2(n6652), .A(n6632), .ZN(U3200) );
  AOI22_X1 U7592 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6650), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6700), .ZN(n6634) );
  OAI21_X1 U7593 ( .B1(n6635), .B2(n6652), .A(n6634), .ZN(U3201) );
  AOI222_X1 U7594 ( .A1(n6650), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6700), .C1(REIP_REG_20__SCAN_IN), .C2(
        n6653), .ZN(n6636) );
  INV_X1 U7595 ( .A(n6636), .ZN(U3202) );
  AOI22_X1 U7596 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6700), .ZN(n6637) );
  OAI21_X1 U7597 ( .B1(n6739), .B2(n6655), .A(n6637), .ZN(U3203) );
  AOI222_X1 U7598 ( .A1(n6650), .A2(REIP_REG_21__SCAN_IN), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6700), .C1(REIP_REG_22__SCAN_IN), .C2(
        n6653), .ZN(n6638) );
  INV_X1 U7599 ( .A(n6638), .ZN(U3204) );
  AOI22_X1 U7600 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6700), .ZN(n6639) );
  OAI21_X1 U7601 ( .B1(n6640), .B2(n6655), .A(n6639), .ZN(U3205) );
  AOI222_X1 U7602 ( .A1(n6650), .A2(REIP_REG_23__SCAN_IN), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6700), .C1(REIP_REG_24__SCAN_IN), .C2(
        n6653), .ZN(n6641) );
  INV_X1 U7603 ( .A(n6641), .ZN(U3206) );
  AOI22_X1 U7604 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6700), .ZN(n6642) );
  OAI21_X1 U7605 ( .B1(n6643), .B2(n6655), .A(n6642), .ZN(U3207) );
  AOI22_X1 U7606 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6650), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6700), .ZN(n6644) );
  OAI21_X1 U7607 ( .B1(n6646), .B2(n6652), .A(n6644), .ZN(U3208) );
  AOI22_X1 U7608 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6700), .ZN(n6645) );
  OAI21_X1 U7609 ( .B1(n6646), .B2(n6655), .A(n6645), .ZN(U3209) );
  AOI22_X1 U7610 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6700), .ZN(n6647) );
  OAI21_X1 U7611 ( .B1(n6815), .B2(n6655), .A(n6647), .ZN(U3210) );
  AOI22_X1 U7612 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6700), .ZN(n6648) );
  OAI21_X1 U7613 ( .B1(n6649), .B2(n6655), .A(n6648), .ZN(U3211) );
  AOI22_X1 U7614 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6650), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6700), .ZN(n6651) );
  OAI21_X1 U7615 ( .B1(n6656), .B2(n6652), .A(n6651), .ZN(U3212) );
  AOI22_X1 U7616 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6700), .ZN(n6654) );
  OAI21_X1 U7617 ( .B1(n6656), .B2(n6655), .A(n6654), .ZN(U3213) );
  OAI22_X1 U7618 ( .A1(n6700), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6684), .ZN(n6657) );
  INV_X1 U7619 ( .A(n6657), .ZN(U3445) );
  MUX2_X1 U7620 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6700), .Z(U3446) );
  MUX2_X1 U7621 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6700), .Z(U3447) );
  MUX2_X1 U7622 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6700), .Z(U3448) );
  OAI21_X1 U7623 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6661), .A(n6659), .ZN(
        n6658) );
  INV_X1 U7624 ( .A(n6658), .ZN(U3451) );
  OAI21_X1 U7625 ( .B1(n6661), .B2(n6660), .A(n6659), .ZN(U3452) );
  OAI211_X1 U7626 ( .C1(n6665), .C2(n6664), .A(n6663), .B(n6662), .ZN(U3453)
         );
  OAI211_X1 U7627 ( .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n6981), .A(n6669), 
        .B(n6666), .ZN(n6671) );
  AND2_X1 U7628 ( .A1(n6668), .A2(n6667), .ZN(n6670) );
  OAI22_X1 U7629 ( .A1(n6671), .A2(n6670), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6669), .ZN(n6672) );
  OAI21_X1 U7630 ( .B1(n6674), .B2(n6673), .A(n6672), .ZN(U3461) );
  AOI21_X1 U7631 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6675) );
  AOI22_X1 U7632 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6675), .B2(n6980), .ZN(n6677) );
  INV_X1 U7633 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6676) );
  AOI22_X1 U7634 ( .A1(n6678), .A2(n6677), .B1(n6676), .B2(n6681), .ZN(U3468)
         );
  INV_X1 U7635 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6682) );
  NOR2_X1 U7636 ( .A1(n6681), .A2(REIP_REG_1__SCAN_IN), .ZN(n6679) );
  AOI22_X1 U7637 ( .A1(n6682), .A2(n6681), .B1(n6680), .B2(n6679), .ZN(U3469)
         );
  INV_X1 U7638 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6683) );
  AOI22_X1 U7639 ( .A1(n6684), .A2(READREQUEST_REG_SCAN_IN), .B1(n6683), .B2(
        n6700), .ZN(U3470) );
  AOI211_X1 U7640 ( .C1(n6687), .C2(n6690), .A(n6686), .B(n6685), .ZN(n6699)
         );
  INV_X1 U7641 ( .A(n6688), .ZN(n6693) );
  OAI21_X1 U7642 ( .B1(n6689), .B2(n6703), .A(n3406), .ZN(n6691) );
  OAI211_X1 U7643 ( .C1(n6693), .C2(n6692), .A(n6691), .B(n6690), .ZN(n6696)
         );
  AOI22_X1 U7644 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6696), .B1(n6695), .B2(
        n6694), .ZN(n6698) );
  NAND2_X1 U7645 ( .A1(n6699), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6697) );
  OAI21_X1 U7646 ( .B1(n6699), .B2(n6698), .A(n6697), .ZN(U3472) );
  MUX2_X1 U7647 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6700), .Z(U3473) );
  INV_X1 U7648 ( .A(DATAI_19_), .ZN(n6702) );
  AOI22_X1 U7649 ( .A1(n6703), .A2(keyinput118), .B1(keyinput115), .B2(n6702), 
        .ZN(n6701) );
  OAI221_X1 U7650 ( .B1(n6703), .B2(keyinput118), .C1(n6702), .C2(keyinput115), 
        .A(n6701), .ZN(n6715) );
  INV_X1 U7651 ( .A(keyinput17), .ZN(n6862) );
  AOI22_X1 U7652 ( .A1(n6705), .A2(keyinput55), .B1(ADDRESS_REG_15__SCAN_IN), 
        .B2(n6862), .ZN(n6704) );
  OAI221_X1 U7653 ( .B1(n6705), .B2(keyinput55), .C1(n6862), .C2(
        ADDRESS_REG_15__SCAN_IN), .A(n6704), .ZN(n6714) );
  INV_X1 U7654 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6708) );
  INV_X1 U7655 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6707) );
  AOI22_X1 U7656 ( .A1(n6708), .A2(keyinput88), .B1(n6707), .B2(keyinput78), 
        .ZN(n6706) );
  OAI221_X1 U7657 ( .B1(n6708), .B2(keyinput88), .C1(n6707), .C2(keyinput78), 
        .A(n6706), .ZN(n6713) );
  INV_X1 U7658 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6709) );
  XOR2_X1 U7659 ( .A(n6709), .B(keyinput39), .Z(n6711) );
  XNOR2_X1 U7660 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .B(keyinput53), .ZN(n6710)
         );
  NAND2_X1 U7661 ( .A1(n6711), .A2(n6710), .ZN(n6712) );
  NOR4_X1 U7662 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n7016)
         );
  AOI22_X1 U7663 ( .A1(n6718), .A2(keyinput33), .B1(keyinput0), .B2(n6717), 
        .ZN(n6716) );
  OAI221_X1 U7664 ( .B1(n6718), .B2(keyinput33), .C1(n6717), .C2(keyinput0), 
        .A(n6716), .ZN(n6730) );
  INV_X1 U7665 ( .A(keyinput3), .ZN(n6720) );
  AOI22_X1 U7666 ( .A1(n6721), .A2(keyinput112), .B1(ADDRESS_REG_18__SCAN_IN), 
        .B2(n6720), .ZN(n6719) );
  OAI221_X1 U7667 ( .B1(n6721), .B2(keyinput112), .C1(n6720), .C2(
        ADDRESS_REG_18__SCAN_IN), .A(n6719), .ZN(n6729) );
  AOI22_X1 U7668 ( .A1(n6723), .A2(keyinput81), .B1(keyinput105), .B2(n4288), 
        .ZN(n6722) );
  OAI221_X1 U7669 ( .B1(n6723), .B2(keyinput81), .C1(n4288), .C2(keyinput105), 
        .A(n6722), .ZN(n6728) );
  INV_X1 U7670 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6725) );
  AOI22_X1 U7671 ( .A1(n6726), .A2(keyinput80), .B1(n6725), .B2(keyinput19), 
        .ZN(n6724) );
  OAI221_X1 U7672 ( .B1(n6726), .B2(keyinput80), .C1(n6725), .C2(keyinput19), 
        .A(n6724), .ZN(n6727) );
  NOR4_X1 U7673 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n7015)
         );
  INV_X1 U7674 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6733) );
  AOI22_X1 U7675 ( .A1(n6733), .A2(keyinput103), .B1(n6732), .B2(keyinput108), 
        .ZN(n6731) );
  OAI221_X1 U7676 ( .B1(n6733), .B2(keyinput103), .C1(n6732), .C2(keyinput108), 
        .A(n6731), .ZN(n6752) );
  INV_X1 U7677 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6736) );
  AOI22_X1 U7678 ( .A1(n6736), .A2(keyinput34), .B1(keyinput119), .B2(n6735), 
        .ZN(n6734) );
  OAI221_X1 U7679 ( .B1(n6736), .B2(keyinput34), .C1(n6735), .C2(keyinput119), 
        .A(n6734), .ZN(n6751) );
  AOI22_X1 U7680 ( .A1(n6738), .A2(keyinput110), .B1(n5118), .B2(keyinput41), 
        .ZN(n6737) );
  OAI221_X1 U7681 ( .B1(n6738), .B2(keyinput110), .C1(n5118), .C2(keyinput41), 
        .A(n6737), .ZN(n6750) );
  XOR2_X1 U7682 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput10), .Z(n6743)
         );
  XOR2_X1 U7683 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput97), .Z(n6742)
         );
  XOR2_X1 U7684 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .B(keyinput37), .Z(n6741)
         );
  XNOR2_X1 U7685 ( .A(keyinput15), .B(n6739), .ZN(n6740) );
  NOR4_X1 U7686 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6748)
         );
  XOR2_X1 U7687 ( .A(n6744), .B(keyinput126), .Z(n6747) );
  XOR2_X1 U7688 ( .A(n6745), .B(keyinput74), .Z(n6746) );
  NAND3_X1 U7689 ( .A1(n6748), .A2(n6747), .A3(n6746), .ZN(n6749) );
  OR4_X1 U7690 ( .A1(n6752), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(n6792) );
  OAI22_X1 U7691 ( .A1(n6754), .A2(keyinput38), .B1(n4625), .B2(keyinput77), 
        .ZN(n6753) );
  AOI221_X1 U7692 ( .B1(n6754), .B2(keyinput38), .C1(keyinput77), .C2(n4625), 
        .A(n6753), .ZN(n6773) );
  INV_X1 U7693 ( .A(keyinput64), .ZN(n6756) );
  OAI22_X1 U7694 ( .A1(n6757), .A2(keyinput70), .B1(n6756), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n6755) );
  AOI221_X1 U7695 ( .B1(n6757), .B2(keyinput70), .C1(ADDRESS_REG_22__SCAN_IN), 
        .C2(n6756), .A(n6755), .ZN(n6772) );
  INV_X1 U7696 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6760) );
  INV_X1 U7697 ( .A(keyinput87), .ZN(n6759) );
  AOI22_X1 U7698 ( .A1(n6760), .A2(keyinput47), .B1(ADDRESS_REG_2__SCAN_IN), 
        .B2(n6759), .ZN(n6758) );
  OAI221_X1 U7699 ( .B1(n6760), .B2(keyinput47), .C1(n6759), .C2(
        ADDRESS_REG_2__SCAN_IN), .A(n6758), .ZN(n6770) );
  AOI22_X1 U7700 ( .A1(n4341), .A2(keyinput25), .B1(keyinput71), .B2(n6762), 
        .ZN(n6761) );
  OAI221_X1 U7701 ( .B1(n4341), .B2(keyinput25), .C1(n6762), .C2(keyinput71), 
        .A(n6761), .ZN(n6769) );
  INV_X1 U7702 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6765) );
  AOI22_X1 U7703 ( .A1(n6765), .A2(keyinput120), .B1(keyinput46), .B2(n6764), 
        .ZN(n6763) );
  OAI221_X1 U7704 ( .B1(n6765), .B2(keyinput120), .C1(n6764), .C2(keyinput46), 
        .A(n6763), .ZN(n6768) );
  AOI22_X1 U7705 ( .A1(n4620), .A2(keyinput5), .B1(n5134), .B2(keyinput73), 
        .ZN(n6766) );
  OAI221_X1 U7706 ( .B1(n4620), .B2(keyinput5), .C1(n5134), .C2(keyinput73), 
        .A(n6766), .ZN(n6767) );
  NOR4_X1 U7707 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n6771)
         );
  NAND3_X1 U7708 ( .A1(n6773), .A2(n6772), .A3(n6771), .ZN(n6791) );
  INV_X1 U7709 ( .A(keyinput51), .ZN(n6775) );
  AOI22_X1 U7710 ( .A1(n6776), .A2(keyinput11), .B1(CODEFETCH_REG_SCAN_IN), 
        .B2(n6775), .ZN(n6774) );
  OAI221_X1 U7711 ( .B1(n6776), .B2(keyinput11), .C1(n6775), .C2(
        CODEFETCH_REG_SCAN_IN), .A(n6774), .ZN(n6789) );
  INV_X1 U7712 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6779) );
  INV_X1 U7713 ( .A(keyinput75), .ZN(n6778) );
  AOI22_X1 U7714 ( .A1(n6779), .A2(keyinput121), .B1(BE_N_REG_3__SCAN_IN), 
        .B2(n6778), .ZN(n6777) );
  OAI221_X1 U7715 ( .B1(n6779), .B2(keyinput121), .C1(n6778), .C2(
        BE_N_REG_3__SCAN_IN), .A(n6777), .ZN(n6788) );
  INV_X1 U7716 ( .A(keyinput117), .ZN(n6781) );
  AOI22_X1 U7717 ( .A1(n6782), .A2(keyinput99), .B1(DATAWIDTH_REG_25__SCAN_IN), 
        .B2(n6781), .ZN(n6780) );
  OAI221_X1 U7718 ( .B1(n6782), .B2(keyinput99), .C1(n6781), .C2(
        DATAWIDTH_REG_25__SCAN_IN), .A(n6780), .ZN(n6787) );
  INV_X1 U7719 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6784) );
  AOI22_X1 U7720 ( .A1(n6785), .A2(keyinput12), .B1(n6784), .B2(keyinput116), 
        .ZN(n6783) );
  OAI221_X1 U7721 ( .B1(n6785), .B2(keyinput12), .C1(n6784), .C2(keyinput116), 
        .A(n6783), .ZN(n6786) );
  OR4_X1 U7722 ( .A1(n6789), .A2(n6788), .A3(n6787), .A4(n6786), .ZN(n6790) );
  NOR3_X1 U7723 ( .A1(n6792), .A2(n6791), .A3(n6790), .ZN(n6825) );
  INV_X1 U7724 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6794) );
  AOI22_X1 U7725 ( .A1(n6795), .A2(keyinput57), .B1(n6794), .B2(keyinput14), 
        .ZN(n6793) );
  OAI221_X1 U7726 ( .B1(n6795), .B2(keyinput57), .C1(n6794), .C2(keyinput14), 
        .A(n6793), .ZN(n6807) );
  INV_X1 U7727 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6798) );
  AOI22_X1 U7728 ( .A1(n6798), .A2(keyinput9), .B1(keyinput67), .B2(n6797), 
        .ZN(n6796) );
  OAI221_X1 U7729 ( .B1(n6798), .B2(keyinput9), .C1(n6797), .C2(keyinput67), 
        .A(n6796), .ZN(n6806) );
  AOI22_X1 U7730 ( .A1(n3779), .A2(keyinput30), .B1(n6800), .B2(keyinput54), 
        .ZN(n6799) );
  OAI221_X1 U7731 ( .B1(n3779), .B2(keyinput30), .C1(n6800), .C2(keyinput54), 
        .A(n6799), .ZN(n6805) );
  INV_X1 U7732 ( .A(DATAI_25_), .ZN(n6802) );
  AOI22_X1 U7733 ( .A1(n6803), .A2(keyinput107), .B1(keyinput20), .B2(n6802), 
        .ZN(n6801) );
  OAI221_X1 U7734 ( .B1(n6803), .B2(keyinput107), .C1(n6802), .C2(keyinput20), 
        .A(n6801), .ZN(n6804) );
  NOR4_X1 U7735 ( .A1(n6807), .A2(n6806), .A3(n6805), .A4(n6804), .ZN(n6824)
         );
  AOI22_X1 U7736 ( .A1(n6810), .A2(keyinput76), .B1(n6809), .B2(keyinput2), 
        .ZN(n6808) );
  OAI221_X1 U7737 ( .B1(n6810), .B2(keyinput76), .C1(n6809), .C2(keyinput2), 
        .A(n6808), .ZN(n6822) );
  INV_X1 U7738 ( .A(keyinput52), .ZN(n6831) );
  AOI22_X1 U7739 ( .A1(n6812), .A2(keyinput45), .B1(BYTEENABLE_REG_0__SCAN_IN), 
        .B2(n6831), .ZN(n6811) );
  OAI221_X1 U7740 ( .B1(n6812), .B2(keyinput45), .C1(n6831), .C2(
        BYTEENABLE_REG_0__SCAN_IN), .A(n6811), .ZN(n6821) );
  INV_X1 U7741 ( .A(keyinput32), .ZN(n6814) );
  AOI22_X1 U7742 ( .A1(n6815), .A2(keyinput65), .B1(DATAO_REG_14__SCAN_IN), 
        .B2(n6814), .ZN(n6813) );
  OAI221_X1 U7743 ( .B1(n6815), .B2(keyinput65), .C1(n6814), .C2(
        DATAO_REG_14__SCAN_IN), .A(n6813), .ZN(n6820) );
  INV_X1 U7744 ( .A(keyinput123), .ZN(n6817) );
  AOI22_X1 U7745 ( .A1(n6818), .A2(keyinput89), .B1(ADDRESS_REG_5__SCAN_IN), 
        .B2(n6817), .ZN(n6816) );
  OAI221_X1 U7746 ( .B1(n6818), .B2(keyinput89), .C1(n6817), .C2(
        ADDRESS_REG_5__SCAN_IN), .A(n6816), .ZN(n6819) );
  NOR4_X1 U7747 ( .A1(n6822), .A2(n6821), .A3(n6820), .A4(n6819), .ZN(n6823)
         );
  AND3_X1 U7748 ( .A1(n6825), .A2(n6824), .A3(n6823), .ZN(n7014) );
  NOR2_X1 U7749 ( .A1(keyinput57), .A2(keyinput20), .ZN(n6826) );
  NAND3_X1 U7750 ( .A1(keyinput14), .A2(keyinput107), .A3(n6826), .ZN(n6827)
         );
  NOR3_X1 U7751 ( .A1(keyinput30), .A2(keyinput54), .A3(n6827), .ZN(n6828) );
  NAND3_X1 U7752 ( .A1(keyinput9), .A2(keyinput67), .A3(n6828), .ZN(n6850) );
  NOR2_X1 U7753 ( .A1(keyinput11), .A2(keyinput108), .ZN(n6829) );
  NAND3_X1 U7754 ( .A1(keyinput51), .A2(keyinput103), .A3(n6829), .ZN(n6830)
         );
  NOR3_X1 U7755 ( .A1(keyinput15), .A2(keyinput37), .A3(n6830), .ZN(n6838) );
  NAND4_X1 U7756 ( .A1(keyinput89), .A2(keyinput123), .A3(keyinput32), .A4(
        keyinput65), .ZN(n6836) );
  NAND4_X1 U7757 ( .A1(keyinput45), .A2(keyinput76), .A3(keyinput2), .A4(n6831), .ZN(n6835) );
  NAND4_X1 U7758 ( .A1(keyinput34), .A2(keyinput119), .A3(keyinput74), .A4(
        keyinput10), .ZN(n6834) );
  NOR2_X1 U7759 ( .A1(keyinput99), .A2(keyinput41), .ZN(n6832) );
  NAND3_X1 U7760 ( .A1(keyinput110), .A2(keyinput117), .A3(n6832), .ZN(n6833)
         );
  NOR4_X1 U7761 ( .A1(n6836), .A2(n6835), .A3(n6834), .A4(n6833), .ZN(n6837)
         );
  NAND4_X1 U7762 ( .A1(keyinput121), .A2(keyinput75), .A3(n6838), .A4(n6837), 
        .ZN(n6849) );
  NOR4_X1 U7763 ( .A1(keyinput109), .A2(keyinput113), .A3(keyinput85), .A4(
        keyinput8), .ZN(n6842) );
  NOR4_X1 U7764 ( .A1(keyinput27), .A2(keyinput22), .A3(keyinput18), .A4(
        keyinput7), .ZN(n6841) );
  NOR4_X1 U7765 ( .A1(keyinput56), .A2(keyinput61), .A3(keyinput29), .A4(
        keyinput124), .ZN(n6840) );
  NOR4_X1 U7766 ( .A1(keyinput28), .A2(keyinput36), .A3(keyinput60), .A4(
        keyinput48), .ZN(n6839) );
  NAND4_X1 U7767 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .ZN(n6848)
         );
  NOR4_X1 U7768 ( .A1(keyinput90), .A2(keyinput86), .A3(keyinput83), .A4(
        keyinput79), .ZN(n6846) );
  NOR4_X1 U7769 ( .A1(keyinput44), .A2(keyinput111), .A3(keyinput102), .A4(
        keyinput94), .ZN(n6845) );
  NOR4_X1 U7770 ( .A1(keyinput59), .A2(keyinput50), .A3(keyinput43), .A4(
        keyinput31), .ZN(n6844) );
  NOR4_X1 U7771 ( .A1(keyinput66), .A2(keyinput62), .A3(keyinput63), .A4(
        keyinput58), .ZN(n6843) );
  NAND4_X1 U7772 ( .A1(n6846), .A2(n6845), .A3(n6844), .A4(n6843), .ZN(n6847)
         );
  NOR4_X1 U7773 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n7012)
         );
  NAND4_X1 U7774 ( .A1(keyinput39), .A2(keyinput53), .A3(keyinput118), .A4(
        keyinput115), .ZN(n6851) );
  NOR3_X1 U7775 ( .A1(keyinput88), .A2(keyinput78), .A3(n6851), .ZN(n6864) );
  NAND2_X1 U7776 ( .A1(keyinput64), .A2(keyinput97), .ZN(n6852) );
  NOR3_X1 U7777 ( .A1(keyinput126), .A2(keyinput70), .A3(n6852), .ZN(n6853) );
  NAND3_X1 U7778 ( .A1(keyinput38), .A2(keyinput77), .A3(n6853), .ZN(n6861) );
  NAND3_X1 U7779 ( .A1(keyinput80), .A2(keyinput33), .A3(keyinput0), .ZN(n6854) );
  NOR2_X1 U7780 ( .A1(keyinput19), .A2(n6854), .ZN(n6859) );
  NOR4_X1 U7781 ( .A1(keyinput112), .A2(keyinput3), .A3(keyinput81), .A4(
        keyinput105), .ZN(n6858) );
  NAND2_X1 U7782 ( .A1(keyinput5), .A2(keyinput47), .ZN(n6855) );
  NOR3_X1 U7783 ( .A1(keyinput87), .A2(keyinput73), .A3(n6855), .ZN(n6857) );
  NOR4_X1 U7784 ( .A1(keyinput25), .A2(keyinput71), .A3(keyinput120), .A4(
        keyinput46), .ZN(n6856) );
  NAND4_X1 U7785 ( .A1(n6859), .A2(n6858), .A3(n6857), .A4(n6856), .ZN(n6860)
         );
  NOR4_X1 U7786 ( .A1(keyinput12), .A2(keyinput116), .A3(n6861), .A4(n6860), 
        .ZN(n6863) );
  NAND4_X1 U7787 ( .A1(keyinput55), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(
        n6875) );
  NAND4_X1 U7788 ( .A1(keyinput23), .A2(keyinput26), .A3(keyinput6), .A4(
        keyinput101), .ZN(n6874) );
  NAND4_X1 U7789 ( .A1(keyinput95), .A2(keyinput82), .A3(keyinput42), .A4(
        keyinput35), .ZN(n6873) );
  NAND4_X1 U7790 ( .A1(keyinput114), .A2(keyinput106), .A3(keyinput98), .A4(
        keyinput91), .ZN(n6865) );
  NOR3_X1 U7791 ( .A1(keyinput104), .A2(keyinput96), .A3(n6865), .ZN(n6871) );
  NAND4_X1 U7792 ( .A1(keyinput4), .A2(keyinput40), .A3(keyinput16), .A4(
        keyinput68), .ZN(n6869) );
  NAND4_X1 U7793 ( .A1(keyinput125), .A2(keyinput69), .A3(keyinput93), .A4(
        keyinput24), .ZN(n6868) );
  NAND4_X1 U7794 ( .A1(keyinput92), .A2(keyinput84), .A3(keyinput72), .A4(
        keyinput100), .ZN(n6867) );
  NAND4_X1 U7795 ( .A1(keyinput49), .A2(keyinput1), .A3(keyinput13), .A4(
        keyinput21), .ZN(n6866) );
  NOR4_X1 U7796 ( .A1(n6869), .A2(n6868), .A3(n6867), .A4(n6866), .ZN(n6870)
         );
  NAND4_X1 U7797 ( .A1(keyinput122), .A2(keyinput127), .A3(n6871), .A4(n6870), 
        .ZN(n6872) );
  NOR4_X1 U7798 ( .A1(n6875), .A2(n6874), .A3(n6873), .A4(n6872), .ZN(n7011)
         );
  INV_X1 U7799 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6878) );
  AOI22_X1 U7800 ( .A1(n6878), .A2(keyinput66), .B1(n6877), .B2(keyinput82), 
        .ZN(n6876) );
  OAI221_X1 U7801 ( .B1(n6878), .B2(keyinput66), .C1(n6877), .C2(keyinput82), 
        .A(n6876), .ZN(n6891) );
  INV_X1 U7802 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6881) );
  INV_X1 U7803 ( .A(keyinput31), .ZN(n6880) );
  AOI22_X1 U7804 ( .A1(n6881), .A2(keyinput69), .B1(DATAWIDTH_REG_18__SCAN_IN), 
        .B2(n6880), .ZN(n6879) );
  OAI221_X1 U7805 ( .B1(n6881), .B2(keyinput69), .C1(n6880), .C2(
        DATAWIDTH_REG_18__SCAN_IN), .A(n6879), .ZN(n6890) );
  INV_X1 U7806 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6883) );
  AOI22_X1 U7807 ( .A1(n6884), .A2(keyinput124), .B1(n6883), .B2(keyinput23), 
        .ZN(n6882) );
  OAI221_X1 U7808 ( .B1(n6884), .B2(keyinput124), .C1(n6883), .C2(keyinput23), 
        .A(n6882), .ZN(n6889) );
  INV_X1 U7809 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6886) );
  AOI22_X1 U7810 ( .A1(n6887), .A2(keyinput85), .B1(n6886), .B2(keyinput8), 
        .ZN(n6885) );
  OAI221_X1 U7811 ( .B1(n6887), .B2(keyinput85), .C1(n6886), .C2(keyinput8), 
        .A(n6885), .ZN(n6888) );
  NOR4_X1 U7812 ( .A1(n6891), .A2(n6890), .A3(n6889), .A4(n6888), .ZN(n6943)
         );
  INV_X1 U7813 ( .A(keyinput84), .ZN(n6893) );
  AOI22_X1 U7814 ( .A1(n6894), .A2(keyinput86), .B1(BYTEENABLE_REG_1__SCAN_IN), 
        .B2(n6893), .ZN(n6892) );
  OAI221_X1 U7815 ( .B1(n6894), .B2(keyinput86), .C1(n6893), .C2(
        BYTEENABLE_REG_1__SCAN_IN), .A(n6892), .ZN(n6907) );
  INV_X1 U7816 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6897) );
  INV_X1 U7817 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6896) );
  AOI22_X1 U7818 ( .A1(n6897), .A2(keyinput102), .B1(n6896), .B2(keyinput90), 
        .ZN(n6895) );
  OAI221_X1 U7819 ( .B1(n6897), .B2(keyinput102), .C1(n6896), .C2(keyinput90), 
        .A(n6895), .ZN(n6906) );
  INV_X1 U7820 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6900) );
  AOI22_X1 U7821 ( .A1(n6900), .A2(keyinput36), .B1(keyinput35), .B2(n6899), 
        .ZN(n6898) );
  OAI221_X1 U7822 ( .B1(n6900), .B2(keyinput36), .C1(n6899), .C2(keyinput35), 
        .A(n6898), .ZN(n6905) );
  INV_X1 U7823 ( .A(keyinput16), .ZN(n6902) );
  AOI22_X1 U7824 ( .A1(n6903), .A2(keyinput26), .B1(BYTEENABLE_REG_3__SCAN_IN), 
        .B2(n6902), .ZN(n6901) );
  OAI221_X1 U7825 ( .B1(n6903), .B2(keyinput26), .C1(n6902), .C2(
        BYTEENABLE_REG_3__SCAN_IN), .A(n6901), .ZN(n6904) );
  NOR4_X1 U7826 ( .A1(n6907), .A2(n6906), .A3(n6905), .A4(n6904), .ZN(n6942)
         );
  INV_X1 U7827 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U7828 ( .A1(n6910), .A2(keyinput40), .B1(keyinput100), .B2(n6909), 
        .ZN(n6908) );
  OAI221_X1 U7829 ( .B1(n6910), .B2(keyinput40), .C1(n6909), .C2(keyinput100), 
        .A(n6908), .ZN(n6923) );
  INV_X1 U7830 ( .A(keyinput79), .ZN(n6912) );
  AOI22_X1 U7831 ( .A1(n6913), .A2(keyinput59), .B1(DATAO_REG_11__SCAN_IN), 
        .B2(n6912), .ZN(n6911) );
  OAI221_X1 U7832 ( .B1(n6913), .B2(keyinput59), .C1(n6912), .C2(
        DATAO_REG_11__SCAN_IN), .A(n6911), .ZN(n6922) );
  INV_X1 U7833 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6915) );
  AOI22_X1 U7834 ( .A1(n6916), .A2(keyinput58), .B1(n6915), .B2(keyinput42), 
        .ZN(n6914) );
  OAI221_X1 U7835 ( .B1(n6916), .B2(keyinput58), .C1(n6915), .C2(keyinput42), 
        .A(n6914), .ZN(n6921) );
  INV_X1 U7836 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6919) );
  AOI22_X1 U7837 ( .A1(n6919), .A2(keyinput94), .B1(keyinput56), .B2(n6918), 
        .ZN(n6917) );
  OAI221_X1 U7838 ( .B1(n6919), .B2(keyinput94), .C1(n6918), .C2(keyinput56), 
        .A(n6917), .ZN(n6920) );
  NOR4_X1 U7839 ( .A1(n6923), .A2(n6922), .A3(n6921), .A4(n6920), .ZN(n6941)
         );
  INV_X1 U7840 ( .A(keyinput60), .ZN(n6926) );
  INV_X1 U7841 ( .A(keyinput91), .ZN(n6925) );
  AOI22_X1 U7842 ( .A1(n6926), .A2(ADDRESS_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6925), .ZN(n6924) );
  OAI221_X1 U7843 ( .B1(n6926), .B2(ADDRESS_REG_20__SCAN_IN), .C1(n6925), .C2(
        ADDRESS_REG_6__SCAN_IN), .A(n6924), .ZN(n6939) );
  INV_X1 U7844 ( .A(keyinput43), .ZN(n6928) );
  AOI22_X1 U7845 ( .A1(n6929), .A2(keyinput125), .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(n6928), .ZN(n6927) );
  OAI221_X1 U7846 ( .B1(n6929), .B2(keyinput125), .C1(n6928), .C2(
        DATAWIDTH_REG_23__SCAN_IN), .A(n6927), .ZN(n6938) );
  INV_X1 U7847 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U7848 ( .A1(n6932), .A2(keyinput111), .B1(n6931), .B2(keyinput127), 
        .ZN(n6930) );
  OAI221_X1 U7849 ( .B1(n6932), .B2(keyinput111), .C1(n6931), .C2(keyinput127), 
        .A(n6930), .ZN(n6937) );
  INV_X1 U7850 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U7851 ( .A1(n6935), .A2(keyinput114), .B1(n6934), .B2(keyinput6), 
        .ZN(n6933) );
  OAI221_X1 U7852 ( .B1(n6935), .B2(keyinput114), .C1(n6934), .C2(keyinput6), 
        .A(n6933), .ZN(n6936) );
  NOR4_X1 U7853 ( .A1(n6939), .A2(n6938), .A3(n6937), .A4(n6936), .ZN(n6940)
         );
  NAND4_X1 U7854 ( .A1(n6943), .A2(n6942), .A3(n6941), .A4(n6940), .ZN(n7010)
         );
  INV_X1 U7855 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6946) );
  INV_X1 U7856 ( .A(keyinput27), .ZN(n6945) );
  AOI22_X1 U7857 ( .A1(n6946), .A2(keyinput93), .B1(BYTEENABLE_REG_2__SCAN_IN), 
        .B2(n6945), .ZN(n6944) );
  OAI221_X1 U7858 ( .B1(n6946), .B2(keyinput93), .C1(n6945), .C2(
        BYTEENABLE_REG_2__SCAN_IN), .A(n6944), .ZN(n6959) );
  INV_X1 U7859 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6949) );
  INV_X1 U7860 ( .A(keyinput104), .ZN(n6948) );
  AOI22_X1 U7861 ( .A1(n6949), .A2(keyinput72), .B1(ADS_N_REG_SCAN_IN), .B2(
        n6948), .ZN(n6947) );
  OAI221_X1 U7862 ( .B1(n6949), .B2(keyinput72), .C1(n6948), .C2(
        ADS_N_REG_SCAN_IN), .A(n6947), .ZN(n6958) );
  INV_X1 U7863 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6951) );
  AOI22_X1 U7864 ( .A1(n6952), .A2(keyinput50), .B1(keyinput61), .B2(n6951), 
        .ZN(n6950) );
  OAI221_X1 U7865 ( .B1(n6952), .B2(keyinput50), .C1(n6951), .C2(keyinput61), 
        .A(n6950), .ZN(n6957) );
  INV_X1 U7866 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6955) );
  INV_X1 U7867 ( .A(keyinput106), .ZN(n6954) );
  AOI22_X1 U7868 ( .A1(n6955), .A2(keyinput96), .B1(DATAWIDTH_REG_30__SCAN_IN), 
        .B2(n6954), .ZN(n6953) );
  OAI221_X1 U7869 ( .B1(n6955), .B2(keyinput96), .C1(n6954), .C2(
        DATAWIDTH_REG_30__SCAN_IN), .A(n6953), .ZN(n6956) );
  NOR4_X1 U7870 ( .A1(n6959), .A2(n6958), .A3(n6957), .A4(n6956), .ZN(n7008)
         );
  INV_X1 U7871 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6962) );
  INV_X1 U7872 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n6961) );
  AOI22_X1 U7873 ( .A1(n6962), .A2(keyinput95), .B1(keyinput101), .B2(n6961), 
        .ZN(n6960) );
  OAI221_X1 U7874 ( .B1(n6962), .B2(keyinput95), .C1(n6961), .C2(keyinput101), 
        .A(n6960), .ZN(n6974) );
  INV_X1 U7875 ( .A(keyinput122), .ZN(n6964) );
  AOI22_X1 U7876 ( .A1(n4367), .A2(keyinput29), .B1(W_R_N_REG_SCAN_IN), .B2(
        n6964), .ZN(n6963) );
  OAI221_X1 U7877 ( .B1(n4367), .B2(keyinput29), .C1(n6964), .C2(
        W_R_N_REG_SCAN_IN), .A(n6963), .ZN(n6973) );
  INV_X1 U7878 ( .A(keyinput7), .ZN(n6966) );
  AOI22_X1 U7879 ( .A1(n6967), .A2(keyinput109), .B1(DATAWIDTH_REG_11__SCAN_IN), .B2(n6966), .ZN(n6965) );
  OAI221_X1 U7880 ( .B1(n6967), .B2(keyinput109), .C1(n6966), .C2(
        DATAWIDTH_REG_11__SCAN_IN), .A(n6965), .ZN(n6972) );
  INV_X1 U7881 ( .A(keyinput44), .ZN(n6970) );
  AOI22_X1 U7882 ( .A1(n6970), .A2(DATAWIDTH_REG_31__SCAN_IN), .B1(keyinput48), 
        .B2(n6969), .ZN(n6968) );
  OAI221_X1 U7883 ( .B1(n6970), .B2(DATAWIDTH_REG_31__SCAN_IN), .C1(n6969), 
        .C2(keyinput48), .A(n6968), .ZN(n6971) );
  NOR4_X1 U7884 ( .A1(n6974), .A2(n6973), .A3(n6972), .A4(n6971), .ZN(n7007)
         );
  INV_X1 U7885 ( .A(keyinput68), .ZN(n6976) );
  AOI22_X1 U7886 ( .A1(n4527), .A2(keyinput24), .B1(DATAWIDTH_REG_10__SCAN_IN), 
        .B2(n6976), .ZN(n6975) );
  OAI221_X1 U7887 ( .B1(n4527), .B2(keyinput24), .C1(n6976), .C2(
        DATAWIDTH_REG_10__SCAN_IN), .A(n6975), .ZN(n6988) );
  INV_X1 U7888 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6978) );
  AOI22_X1 U7889 ( .A1(n6978), .A2(keyinput4), .B1(keyinput92), .B2(n4309), 
        .ZN(n6977) );
  OAI221_X1 U7890 ( .B1(n6978), .B2(keyinput4), .C1(n4309), .C2(keyinput92), 
        .A(n6977), .ZN(n6987) );
  AOI22_X1 U7891 ( .A1(n6981), .A2(keyinput63), .B1(keyinput13), .B2(n6980), 
        .ZN(n6979) );
  OAI221_X1 U7892 ( .B1(n6981), .B2(keyinput63), .C1(n6980), .C2(keyinput13), 
        .A(n6979), .ZN(n6986) );
  INV_X1 U7893 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6984) );
  AOI22_X1 U7894 ( .A1(n6984), .A2(keyinput62), .B1(keyinput22), .B2(n6983), 
        .ZN(n6982) );
  OAI221_X1 U7895 ( .B1(n6984), .B2(keyinput62), .C1(n6983), .C2(keyinput22), 
        .A(n6982), .ZN(n6985) );
  NOR4_X1 U7896 ( .A1(n6988), .A2(n6987), .A3(n6986), .A4(n6985), .ZN(n7006)
         );
  INV_X1 U7897 ( .A(keyinput28), .ZN(n6990) );
  AOI22_X1 U7898 ( .A1(n6991), .A2(keyinput113), .B1(ADDRESS_REG_12__SCAN_IN), 
        .B2(n6990), .ZN(n6989) );
  OAI221_X1 U7899 ( .B1(n6991), .B2(keyinput113), .C1(n6990), .C2(
        ADDRESS_REG_12__SCAN_IN), .A(n6989), .ZN(n7004) );
  INV_X1 U7900 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6994) );
  AOI22_X1 U7901 ( .A1(n6994), .A2(keyinput83), .B1(keyinput98), .B2(n6993), 
        .ZN(n6992) );
  OAI221_X1 U7902 ( .B1(n6994), .B2(keyinput83), .C1(n6993), .C2(keyinput98), 
        .A(n6992), .ZN(n7003) );
  INV_X1 U7903 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n6997) );
  INV_X1 U7904 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6996) );
  AOI22_X1 U7905 ( .A1(n6997), .A2(keyinput18), .B1(n6996), .B2(keyinput21), 
        .ZN(n6995) );
  OAI221_X1 U7906 ( .B1(n6997), .B2(keyinput18), .C1(n6996), .C2(keyinput21), 
        .A(n6995), .ZN(n7002) );
  INV_X1 U7907 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n7000) );
  INV_X1 U7908 ( .A(keyinput49), .ZN(n6999) );
  AOI22_X1 U7909 ( .A1(n7000), .A2(keyinput1), .B1(DATAWIDTH_REG_2__SCAN_IN), 
        .B2(n6999), .ZN(n6998) );
  OAI221_X1 U7910 ( .B1(n7000), .B2(keyinput1), .C1(n6999), .C2(
        DATAWIDTH_REG_2__SCAN_IN), .A(n6998), .ZN(n7001) );
  NOR4_X1 U7911 ( .A1(n7004), .A2(n7003), .A3(n7002), .A4(n7001), .ZN(n7005)
         );
  NAND4_X1 U7912 ( .A1(n7008), .A2(n7007), .A3(n7006), .A4(n7005), .ZN(n7009)
         );
  AOI211_X1 U7913 ( .C1(n7012), .C2(n7011), .A(n7010), .B(n7009), .ZN(n7013)
         );
  NAND4_X1 U7914 ( .A1(n7016), .A2(n7015), .A3(n7014), .A4(n7013), .ZN(n7018)
         );
  NAND2_X1 U7915 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n6140), .ZN(n7017) );
  XOR2_X1 U7916 ( .A(n7018), .B(n7017), .Z(U2892) );
  CLKBUF_X1 U3563 ( .A(n3356), .Z(n3116) );
  CLKBUF_X2 U3587 ( .A(n3134), .Z(n3135) );
  CLKBUF_X1 U3604 ( .A(n4317), .Z(n4676) );
  CLKBUF_X1 U3605 ( .A(n4742), .Z(n3118) );
endmodule

