

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944;

  BUF_X1 U2307 ( .A(n2507), .Z(n2837) );
  CLKBUF_X2 U2308 ( .A(n2510), .Z(n3169) );
  CLKBUF_X2 U2309 ( .A(n2533), .Z(n3102) );
  CLKBUF_X2 U2310 ( .A(n2531), .Z(n2273) );
  NAND4_X2 U2311 ( .A1(n2537), .A2(n2536), .A3(n2535), .A4(n2534), .ZN(n3985)
         );
  XNOR2_X1 U2312 ( .A(n2488), .B(IR_REG_22__SCAN_IN), .ZN(n3962) );
  INV_X1 U2313 ( .A(n3050), .ZN(n3158) );
  NAND2_X1 U2314 ( .A1(n2916), .A2(IR_REG_31__SCAN_IN), .ZN(n2433) );
  NAND4_X2 U2315 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n3049)
         );
  NAND2_X1 U2316 ( .A1(n3004), .A2(n2481), .ZN(n2482) );
  NOR4_X1 U2317 ( .A1(n3927), .A2(n3926), .A3(n4050), .A4(n3925), .ZN(n3937)
         );
  INV_X1 U2318 ( .A(n3985), .ZN(n3110) );
  INV_X2 U2319 ( .A(n2510), .ZN(n2538) );
  OAI21_X1 U2320 ( .B1(n2555), .B2(n2522), .A(n2521), .ZN(n3356) );
  XOR2_X1 U2321 ( .A(n2991), .B(n4939), .Z(n4781) );
  NAND2_X1 U2322 ( .A1(n3144), .A2(n3871), .ZN(n4050) );
  OR2_X1 U2323 ( .A1(n3329), .A2(n2596), .ZN(n2272) );
  MUX2_X2 U2324 ( .A(IR_REG_31__SCAN_IN), .B(n2502), .S(IR_REG_1__SCAN_IN), 
        .Z(n2503) );
  NAND2_X2 U2325 ( .A1(n3684), .A2(n2789), .ZN(n3696) );
  OR2_X2 U2326 ( .A1(n3407), .A2(n3943), .ZN(n3408) );
  NOR2_X2 U2327 ( .A1(n2766), .A2(n3793), .ZN(n2777) );
  NAND2_X2 U2328 ( .A1(n2457), .A2(IR_REG_31__SCAN_IN), .ZN(n2454) );
  NOR2_X1 U2329 ( .A1(n3285), .A2(n2562), .ZN(n3287) );
  OAI22_X2 U2330 ( .A1(n4739), .A2(n2408), .B1(REG1_REG_11__SCAN_IN), .B2(
        n4737), .ZN(n2985) );
  NAND2_X2 U2331 ( .A1(n4727), .A2(n2984), .ZN(n4739) );
  INV_X2 U2332 ( .A(n3049), .ZN(n2509) );
  OAI21_X2 U2333 ( .B1(n3709), .B2(n2288), .A(n2372), .ZN(n3802) );
  NAND2_X2 U2334 ( .A1(n3747), .A2(n2864), .ZN(n3709) );
  OAI22_X2 U2335 ( .A1(n3279), .A2(n3280), .B1(n2514), .B2(n2513), .ZN(n3273)
         );
  AND2_X2 U2336 ( .A1(n2496), .A2(n2495), .ZN(n3279) );
  NOR2_X2 U2337 ( .A1(n4100), .A2(n3866), .ZN(n4081) );
  NOR2_X2 U2338 ( .A1(n4119), .A2(n3896), .ZN(n4100) );
  XNOR2_X2 U2339 ( .A(n2433), .B(n2435), .ZN(n3212) );
  XNOR2_X2 U2340 ( .A(n2454), .B(n3630), .ZN(n2460) );
  NOR2_X2 U2341 ( .A1(n2978), .A2(n3249), .ZN(n4719) );
  AOI22_X2 U2342 ( .A1(n2690), .A2(n3621), .B1(n2689), .B2(n2688), .ZN(n3766)
         );
  NAND2_X1 U2343 ( .A1(n4239), .A2(n4233), .ZN(n4232) );
  AND2_X1 U2344 ( .A1(n3329), .A2(n2596), .ZN(n2598) );
  NAND2_X1 U2345 ( .A1(n3813), .A2(n3816), .ZN(n3407) );
  CLKBUF_X2 U2346 ( .A(U4043), .Z(n4683) );
  NAND2_X1 U2347 ( .A1(n2930), .A2(n3190), .ZN(n2556) );
  CLKBUF_X2 U2348 ( .A(n2497), .Z(n2844) );
  AND2_X1 U2349 ( .A1(n3217), .A2(n2460), .ZN(n2533) );
  NAND2_X1 U2350 ( .A1(n2455), .A2(n2453), .ZN(n2457) );
  AOI21_X1 U2351 ( .B1(n2899), .B2(n2898), .A(n2897), .ZN(n3177) );
  NAND2_X1 U2352 ( .A1(n3885), .A2(n3550), .ZN(n4281) );
  OR2_X2 U2353 ( .A1(n4232), .A2(n4212), .ZN(n4369) );
  AND2_X2 U2354 ( .A1(n3389), .A2(n4909), .ZN(n4944) );
  NOR2_X1 U2355 ( .A1(n2975), .A2(n3252), .ZN(n2978) );
  NAND2_X1 U2356 ( .A1(n2490), .A2(n2489), .ZN(n2839) );
  OAI22_X1 U2357 ( .A1(n4711), .A2(n4709), .B1(n4703), .B2(REG1_REG_7__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U2358 ( .A1(n2974), .A2(n4698), .ZN(n4711) );
  NOR2_X1 U2359 ( .A1(n3190), .A2(n3960), .ZN(U4043) );
  NAND4_X1 U2360 ( .A1(n2464), .A2(n2463), .A3(n2462), .A4(n2461), .ZN(n3987)
         );
  NOR2_X1 U2361 ( .A1(n3962), .A2(n3814), .ZN(n4788) );
  INV_X1 U2362 ( .A(n3950), .ZN(n3814) );
  AND2_X1 U2363 ( .A1(n3217), .A2(n3219), .ZN(n2531) );
  AND2_X1 U2364 ( .A1(n3219), .A2(n2459), .ZN(n2515) );
  INV_X1 U2365 ( .A(n2459), .ZN(n3217) );
  OR2_X2 U2366 ( .A1(n3004), .A2(n2414), .ZN(n2483) );
  OAI22_X1 U2367 ( .A1(n3258), .A2(n2971), .B1(n2970), .B2(n2969), .ZN(n3239)
         );
  NAND2_X1 U2368 ( .A1(n2458), .A2(n2457), .ZN(n2459) );
  OR2_X1 U2369 ( .A1(n2718), .A2(n2717), .ZN(n2731) );
  XNOR2_X1 U2370 ( .A(n2970), .B(n2969), .ZN(n3258) );
  MUX2_X1 U2371 ( .A(IR_REG_31__SCAN_IN), .B(n2456), .S(IR_REG_29__SCAN_IN), 
        .Z(n2458) );
  OAI21_X1 U2372 ( .B1(n2494), .B2(IR_REG_19__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2471) );
  XNOR2_X1 U2373 ( .A(n2448), .B(IR_REG_26__SCAN_IN), .ZN(n2913) );
  AOI22_X1 U2374 ( .A1(n3228), .A2(REG1_REG_3__SCAN_IN), .B1(n4467), .B2(n2968), .ZN(n2970) );
  AND2_X1 U2375 ( .A1(n2544), .A2(n2553), .ZN(n4467) );
  AND2_X1 U2376 ( .A1(n2405), .A2(n2423), .ZN(n2404) );
  NOR2_X1 U2377 ( .A1(n2276), .A2(n2737), .ZN(n2358) );
  AND2_X1 U2378 ( .A1(n2424), .A2(n2406), .ZN(n2405) );
  AND3_X1 U2379 ( .A1(n2322), .A2(n2321), .A3(n2320), .ZN(n2424) );
  INV_X1 U2380 ( .A(IR_REG_0__SCAN_IN), .ZN(n2318) );
  NOR2_X1 U2381 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2441)
         );
  INV_X1 U2382 ( .A(IR_REG_18__SCAN_IN), .ZN(n2772) );
  INV_X1 U2383 ( .A(IR_REG_23__SCAN_IN), .ZN(n2918) );
  NOR2_X1 U2384 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2440)
         );
  NOR2_X1 U2385 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2442)
         );
  INV_X1 U2386 ( .A(IR_REG_7__SCAN_IN), .ZN(n4676) );
  INV_X1 U2387 ( .A(IR_REG_8__SCAN_IN), .ZN(n2621) );
  INV_X1 U2388 ( .A(IR_REG_2__SCAN_IN), .ZN(n2539) );
  INV_X1 U2389 ( .A(IR_REG_17__SCAN_IN), .ZN(n2757) );
  INV_X1 U2390 ( .A(IR_REG_5__SCAN_IN), .ZN(n2419) );
  INV_X1 U2391 ( .A(IR_REG_6__SCAN_IN), .ZN(n2421) );
  INV_X2 U2392 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U2393 ( .A1(n3159), .A2(n3312), .ZN(n3376) );
  INV_X1 U2394 ( .A(n3397), .ZN(n3159) );
  NAND2_X1 U2395 ( .A1(n3674), .A2(n2411), .ZN(n3562) );
  NOR2_X4 U2396 ( .A1(n4321), .A2(n3655), .ZN(n4293) );
  NOR2_X4 U2397 ( .A1(n4328), .A2(n4332), .ZN(n4327) );
  NAND2_X2 U2398 ( .A1(n4045), .A2(n3874), .ZN(n4328) );
  AOI21_X2 U2399 ( .B1(n2272), .B2(n2599), .A(n2598), .ZN(n3461) );
  NOR2_X4 U2400 ( .A1(n4072), .A2(n3179), .ZN(n4045) );
  NAND2_X2 U2401 ( .A1(n4291), .A2(n3582), .ZN(n4383) );
  AND2_X2 U2402 ( .A1(n4293), .A2(n4294), .ZN(n4291) );
  OAI21_X2 U2403 ( .B1(n3461), .B2(n3462), .A(n2612), .ZN(n3476) );
  NOR2_X2 U2404 ( .A1(n2731), .A2(n4539), .ZN(n2752) );
  AOI21_X2 U2405 ( .B1(n3300), .B2(n3296), .A(n3297), .ZN(n3329) );
  NOR2_X2 U2406 ( .A1(n3287), .A2(n2565), .ZN(n3300) );
  INV_X2 U2407 ( .A(n3391), .ZN(n3398) );
  AOI21_X2 U2408 ( .B1(n3562), .B2(n3564), .A(n3563), .ZN(n3619) );
  NOR2_X4 U2409 ( .A1(n4273), .A2(n4244), .ZN(n4239) );
  OR2_X2 U2410 ( .A1(n4383), .A2(n4271), .ZN(n4273) );
  NAND2_X1 U2411 ( .A1(n2353), .A2(n2352), .ZN(n2351) );
  NOR2_X1 U2412 ( .A1(n4167), .A2(n4137), .ZN(n2356) );
  INV_X1 U2413 ( .A(n3086), .ZN(n2352) );
  AOI21_X1 U2414 ( .B1(n2349), .B2(n2354), .A(n4139), .ZN(n2348) );
  AOI21_X1 U2415 ( .B1(n2385), .B2(n2383), .A(n3778), .ZN(n2381) );
  INV_X1 U2416 ( .A(n2383), .ZN(n2382) );
  INV_X1 U2417 ( .A(n2394), .ZN(n2393) );
  OAI21_X1 U2418 ( .B1(n2293), .B2(n2397), .A(n2395), .ZN(n2394) );
  NAND2_X1 U2419 ( .A1(n2399), .A2(n2396), .ZN(n2395) );
  NAND2_X1 U2420 ( .A1(n3200), .A2(n3009), .ZN(n3010) );
  AOI21_X1 U2421 ( .B1(n3448), .B2(n2361), .A(n2359), .ZN(n3548) );
  AND2_X1 U2422 ( .A1(n3073), .A2(n2274), .ZN(n2361) );
  OAI21_X1 U2423 ( .B1(n2275), .B2(n2360), .A(n2292), .ZN(n2359) );
  NOR2_X1 U2424 ( .A1(n2335), .A2(n3063), .ZN(n2333) );
  NAND2_X1 U2425 ( .A1(n3448), .A2(n2274), .ZN(n2363) );
  NAND2_X1 U2426 ( .A1(n2465), .A2(n2426), .ZN(n2439) );
  NAND2_X1 U2427 ( .A1(n2765), .A2(n2291), .ZN(n2371) );
  NAND2_X1 U2428 ( .A1(n2538), .A2(n3987), .ZN(n2367) );
  OAI211_X1 U2429 ( .C1(n4762), .C2(n2303), .A(n2301), .B(n2300), .ZN(n3588)
         );
  INV_X1 U2430 ( .A(n2305), .ZN(n2303) );
  AOI22_X1 U2431 ( .A1(n2305), .A2(n2302), .B1(n2304), .B2(n4759), .ZN(n2301)
         );
  AND2_X1 U2432 ( .A1(n3190), .A2(n3225), .ZN(n3269) );
  AOI21_X1 U2433 ( .B1(n3769), .B2(n2403), .A(n2402), .ZN(n2401) );
  INV_X1 U2434 ( .A(n3652), .ZN(n2402) );
  NOR2_X1 U2435 ( .A1(n3769), .A2(n2403), .ZN(n2399) );
  INV_X1 U2436 ( .A(n3979), .ZN(n3120) );
  AND2_X1 U2437 ( .A1(n2675), .A2(n2674), .ZN(n2676) );
  AOI22_X1 U2438 ( .A1(n3199), .A2(n3198), .B1(n3007), .B2(REG1_REG_2__SCAN_IN), .ZN(n2967) );
  NOR2_X1 U2439 ( .A1(n3229), .A2(n2418), .ZN(n3011) );
  INV_X1 U2440 ( .A(n3930), .ZN(n2362) );
  INV_X1 U2441 ( .A(n3980), .ZN(n3495) );
  INV_X1 U2442 ( .A(n3063), .ZN(n2332) );
  NAND2_X1 U2443 ( .A1(n3061), .A2(n2337), .ZN(n2336) );
  INV_X1 U2444 ( .A(n3060), .ZN(n2337) );
  AOI21_X1 U2445 ( .B1(n2274), .B2(n3069), .A(n2365), .ZN(n2364) );
  NOR2_X1 U2446 ( .A1(n3120), .A2(n3535), .ZN(n2365) );
  AND2_X1 U2447 ( .A1(n3516), .A2(n3518), .ZN(n3930) );
  INV_X1 U2448 ( .A(IR_REG_16__SCAN_IN), .ZN(n2425) );
  INV_X1 U2449 ( .A(IR_REG_13__SCAN_IN), .ZN(n2406) );
  INV_X1 U2450 ( .A(n3634), .ZN(n3098) );
  INV_X1 U2451 ( .A(n2555), .ZN(n2504) );
  INV_X1 U2452 ( .A(n2751), .ZN(n2390) );
  INV_X1 U2453 ( .A(n2287), .ZN(n2389) );
  NOR2_X1 U2454 ( .A1(n3686), .A2(n2370), .ZN(n2369) );
  INV_X1 U2455 ( .A(n2776), .ZN(n2370) );
  AND2_X1 U2456 ( .A1(n2708), .A2(n2707), .ZN(n3769) );
  INV_X1 U2457 ( .A(n3758), .ZN(n2386) );
  OR2_X1 U2458 ( .A1(n2820), .A2(n2821), .ZN(n2383) );
  BUF_X1 U2459 ( .A(n3103), .Z(n3635) );
  INV_X1 U2460 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2316) );
  INV_X1 U2461 ( .A(n3241), .ZN(n2314) );
  XNOR2_X1 U2462 ( .A(n3011), .B(n4466), .ZN(n3257) );
  NAND2_X1 U2463 ( .A1(n4743), .A2(n3024), .ZN(n3025) );
  OR2_X1 U2464 ( .A1(n4762), .A2(n4759), .ZN(n2299) );
  NAND2_X1 U2465 ( .A1(n4773), .A2(n3033), .ZN(n4014) );
  NAND2_X1 U2466 ( .A1(n4014), .A2(n4016), .ZN(n4015) );
  AOI21_X1 U2467 ( .B1(n2343), .B2(n2342), .A(n2294), .ZN(n2341) );
  AND2_X1 U2468 ( .A1(n3869), .A2(n4048), .ZN(n4069) );
  NAND2_X1 U2469 ( .A1(n4104), .A2(n4090), .ZN(n3092) );
  AOI21_X1 U2470 ( .B1(n2346), .B2(n2347), .A(n2295), .ZN(n2344) );
  AND2_X1 U2471 ( .A1(n2846), .A2(n2832), .ZN(n4158) );
  AOI21_X1 U2472 ( .B1(n3490), .B2(n3067), .A(n2412), .ZN(n3448) );
  INV_X1 U2473 ( .A(n3061), .ZN(n2338) );
  AND4_X1 U2474 ( .A1(n2519), .A2(n2518), .A3(n2517), .A4(n2516), .ZN(n3344)
         );
  OAI21_X1 U2475 ( .B1(n2917), .B2(n2436), .A(IR_REG_31__SCAN_IN), .ZN(n2438)
         );
  INV_X1 U2476 ( .A(IR_REG_25__SCAN_IN), .ZN(n2437) );
  INV_X1 U2477 ( .A(n2908), .ZN(n2450) );
  INV_X1 U2478 ( .A(n3212), .ZN(n2451) );
  INV_X1 U2479 ( .A(n3802), .ZN(n2899) );
  NAND2_X1 U2480 ( .A1(n2878), .A2(n2366), .ZN(n2495) );
  AND2_X1 U2481 ( .A1(n2367), .A2(n2368), .ZN(n2366) );
  NAND2_X1 U2482 ( .A1(n2555), .A2(n3007), .ZN(n2521) );
  NAND2_X1 U2483 ( .A1(n4744), .A2(n4745), .ZN(n4743) );
  INV_X1 U2484 ( .A(n2401), .ZN(n2397) );
  NAND2_X1 U2485 ( .A1(n4918), .A2(n4760), .ZN(n2306) );
  AND2_X1 U2486 ( .A1(n2802), .A2(REG3_REG_21__SCAN_IN), .ZN(n2822) );
  AND2_X1 U2487 ( .A1(n2790), .A2(REG3_REG_20__SCAN_IN), .ZN(n2802) );
  INV_X1 U2488 ( .A(n3073), .ZN(n2360) );
  INV_X1 U2489 ( .A(n2443), .ZN(n2429) );
  INV_X1 U2490 ( .A(n3160), .ZN(n2489) );
  OR2_X1 U2491 ( .A1(n4693), .A2(n3015), .ZN(n2307) );
  INV_X1 U2492 ( .A(n2306), .ZN(n2302) );
  AOI21_X1 U2493 ( .B1(n4759), .B2(n2306), .A(n3209), .ZN(n2305) );
  AND2_X1 U2494 ( .A1(n2306), .A2(n3209), .ZN(n2304) );
  INV_X1 U2495 ( .A(n3092), .ZN(n2342) );
  AOI21_X1 U2496 ( .B1(n2348), .B2(n2350), .A(n2298), .ZN(n2346) );
  INV_X1 U2497 ( .A(n2348), .ZN(n2347) );
  OAI21_X1 U2498 ( .B1(n3053), .B2(n2326), .A(n3055), .ZN(n2324) );
  NAND2_X1 U2499 ( .A1(n3158), .A2(n3049), .ZN(n3813) );
  AND2_X1 U2500 ( .A1(n3814), .A2(n3962), .ZN(n3107) );
  AND2_X1 U2501 ( .A1(n2358), .A2(n2285), .ZN(n2357) );
  INV_X1 U2502 ( .A(IR_REG_12__SCAN_IN), .ZN(n2320) );
  INV_X1 U2503 ( .A(IR_REG_9__SCAN_IN), .ZN(n2423) );
  AOI21_X1 U2504 ( .B1(n2381), .B2(n2382), .A(n2379), .ZN(n2378) );
  INV_X1 U2505 ( .A(n2859), .ZN(n2379) );
  AND2_X1 U2506 ( .A1(n3098), .A2(DATAI_20_), .ZN(n4212) );
  AND2_X1 U2507 ( .A1(n2691), .A2(REG3_REG_13__SCAN_IN), .ZN(n2709) );
  AND2_X1 U2508 ( .A1(n3675), .A2(n3673), .ZN(n2658) );
  NAND2_X1 U2509 ( .A1(n2392), .A2(n2287), .ZN(n2391) );
  INV_X1 U2510 ( .A(n3766), .ZN(n2392) );
  AND4_X1 U2511 ( .A1(n2607), .A2(n2606), .A3(n2605), .A4(n2604), .ZN(n3369)
         );
  XNOR2_X1 U2512 ( .A(n3010), .B(n4467), .ZN(n3230) );
  NOR2_X1 U2513 ( .A1(n3230), .A2(n3231), .ZN(n3229) );
  AND2_X1 U2514 ( .A1(n2575), .A2(n2419), .ZN(n2373) );
  NAND2_X1 U2515 ( .A1(n2977), .A2(n2976), .ZN(n3250) );
  NAND2_X1 U2516 ( .A1(n4722), .A2(n3020), .ZN(n3022) );
  NAND2_X1 U2517 ( .A1(n2982), .A2(n2981), .ZN(n2983) );
  NAND2_X1 U2518 ( .A1(n2980), .A2(REG1_REG_9__SCAN_IN), .ZN(n2981) );
  NAND2_X1 U2519 ( .A1(n2979), .A2(n4716), .ZN(n2982) );
  NAND2_X1 U2520 ( .A1(n4001), .A2(n3029), .ZN(n4002) );
  INV_X1 U2521 ( .A(n4004), .ZN(n3029) );
  AND2_X1 U2522 ( .A1(n4002), .A2(n3030), .ZN(n3032) );
  NAND2_X1 U2523 ( .A1(n4015), .A2(n3035), .ZN(n4028) );
  INV_X1 U2524 ( .A(n4069), .ZN(n4062) );
  AND4_X1 U2525 ( .A1(n2888), .A2(n2887), .A3(n2886), .A4(n2885), .ZN(n4085)
         );
  AOI21_X1 U2526 ( .B1(n3089), .B2(n3088), .A(n3087), .ZN(n4097) );
  NAND2_X1 U2527 ( .A1(n4151), .A2(n4128), .ZN(n3088) );
  AND2_X1 U2528 ( .A1(n3141), .A2(n4122), .ZN(n3087) );
  INV_X1 U2529 ( .A(n4187), .ZN(n4149) );
  OR2_X1 U2530 ( .A1(n4183), .A2(n4141), .ZN(n4143) );
  AND4_X1 U2531 ( .A1(n2836), .A2(n2835), .A3(n2834), .A4(n2833), .ZN(n4171)
         );
  AND2_X1 U2532 ( .A1(n2355), .A2(n2281), .ZN(n4182) );
  NAND2_X1 U2533 ( .A1(n4207), .A2(n3086), .ZN(n2355) );
  AOI21_X1 U2534 ( .B1(n3572), .B2(n3081), .A(n2417), .ZN(n4254) );
  AND4_X1 U2535 ( .A1(n2770), .A2(n2769), .A3(n2768), .A4(n2767), .ZN(n4270)
         );
  AND4_X1 U2536 ( .A1(n2756), .A2(n2755), .A3(n2754), .A4(n2753), .ZN(n4247)
         );
  AOI21_X1 U2537 ( .B1(n3548), .B2(n3077), .A(n3076), .ZN(n3573) );
  OR2_X1 U2538 ( .A1(n3078), .A2(n3886), .ZN(n3574) );
  NAND2_X1 U2539 ( .A1(n2709), .A2(REG3_REG_14__SCAN_IN), .ZN(n2718) );
  AND4_X1 U2540 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), .ZN(n4311)
         );
  AND4_X1 U2541 ( .A1(n2669), .A2(n2668), .A3(n2667), .A4(n2666), .ZN(n3536)
         );
  NOR2_X1 U2542 ( .A1(n2663), .A2(n2662), .ZN(n2678) );
  INV_X1 U2543 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4528) );
  OR2_X1 U2544 ( .A1(n2630), .A2(n2629), .ZN(n2644) );
  AND2_X1 U2545 ( .A1(n2331), .A2(n2330), .ZN(n2329) );
  OR2_X1 U2546 ( .A1(n3982), .A2(n3375), .ZN(n2330) );
  AND2_X1 U2547 ( .A1(n3114), .A2(n3838), .ZN(n4847) );
  INV_X1 U2548 ( .A(n3463), .ZN(n4856) );
  AND4_X1 U2549 ( .A1(n2552), .A2(n2551), .A3(n2550), .A4(n2549), .ZN(n3313)
         );
  AND2_X1 U2550 ( .A1(n3147), .A2(n3146), .ZN(n4863) );
  AND4_X1 U2551 ( .A1(n2573), .A2(n2572), .A3(n2571), .A4(n2570), .ZN(n3393)
         );
  AND2_X1 U2552 ( .A1(n3823), .A2(n3826), .ZN(n3929) );
  AND2_X1 U2553 ( .A1(n3817), .A2(n3820), .ZN(n3928) );
  AOI21_X1 U2554 ( .B1(n3223), .B2(n3227), .A(n3226), .ZN(n3163) );
  AND2_X1 U2555 ( .A1(n4462), .A2(n4788), .ZN(n4331) );
  INV_X1 U2556 ( .A(n3143), .ZN(n4073) );
  INV_X1 U2557 ( .A(n4122), .ZN(n4128) );
  CLKBUF_X1 U2558 ( .A(n4154), .Z(n4359) );
  NOR2_X2 U2559 ( .A1(n4369), .A2(n3703), .ZN(n4190) );
  INV_X1 U2560 ( .A(n4919), .ZN(n4294) );
  INV_X1 U2561 ( .A(n3623), .ZN(n3522) );
  NAND2_X1 U2562 ( .A1(n2363), .A2(n2364), .ZN(n3601) );
  INV_X1 U2563 ( .A(n3677), .ZN(n3535) );
  AND2_X1 U2564 ( .A1(n4842), .A2(n4856), .ZN(n4843) );
  NOR2_X2 U2565 ( .A1(n3376), .A2(n3375), .ZN(n4842) );
  NAND2_X1 U2566 ( .A1(n3399), .A2(n3398), .ZN(n3397) );
  AND3_X1 U2567 ( .A1(n3156), .A2(n3155), .A3(n3154), .ZN(n3164) );
  INV_X1 U2568 ( .A(n2475), .ZN(n2472) );
  NOR2_X1 U2569 ( .A1(n2467), .A2(n2375), .ZN(n2374) );
  INV_X1 U2570 ( .A(n2466), .ZN(n2375) );
  INV_X1 U2571 ( .A(IR_REG_15__SCAN_IN), .ZN(n2726) );
  AND2_X1 U2572 ( .A1(n2685), .A2(n2672), .ZN(n4737) );
  NAND2_X1 U2573 ( .A1(n2621), .A2(n4676), .ZN(n2422) );
  INV_X1 U2574 ( .A(IR_REG_31__SCAN_IN), .ZN(n2650) );
  NAND2_X1 U2575 ( .A1(n2503), .A2(n2319), .ZN(n3988) );
  INV_X1 U2576 ( .A(n3769), .ZN(n2398) );
  NAND2_X1 U2577 ( .A1(n3766), .A2(n3768), .ZN(n2400) );
  AOI21_X1 U2578 ( .B1(n2278), .B2(n2389), .A(n2297), .ZN(n2388) );
  INV_X1 U2579 ( .A(n3286), .ZN(n2560) );
  CLKBUF_X1 U2580 ( .A(n3766), .Z(n3767) );
  NAND2_X1 U2581 ( .A1(n3696), .A2(n2384), .ZN(n2380) );
  CLKBUF_X1 U2582 ( .A(n3806), .Z(n4924) );
  INV_X1 U2583 ( .A(n3688), .ZN(n4920) );
  OR2_X1 U2584 ( .A1(n3710), .A2(n3711), .ZN(n2372) );
  AND2_X1 U2585 ( .A1(n2935), .A2(n2934), .ZN(n4938) );
  INV_X1 U2586 ( .A(n4123), .ZN(n3971) );
  NAND4_X1 U2587 ( .A1(n2649), .A2(n2648), .A3(n2647), .A4(n2646), .ZN(n3979)
         );
  INV_X1 U2588 ( .A(n3450), .ZN(n4860) );
  INV_X1 U2589 ( .A(n3369), .ZN(n3981) );
  INV_X1 U2590 ( .A(n3393), .ZN(n3983) );
  INV_X1 U2591 ( .A(n3313), .ZN(n3984) );
  INV_X1 U2592 ( .A(n3344), .ZN(n3986) );
  NAND2_X1 U2593 ( .A1(n2515), .A2(REG2_REG_0__SCAN_IN), .ZN(n2463) );
  AND2_X1 U2594 ( .A1(n3257), .A2(REG2_REG_4__SCAN_IN), .ZN(n3263) );
  NAND2_X1 U2595 ( .A1(n3257), .A2(n2315), .ZN(n2313) );
  NOR2_X1 U2596 ( .A1(n3241), .A2(n2316), .ZN(n2315) );
  NOR2_X1 U2597 ( .A1(n3263), .A2(n2413), .ZN(n3242) );
  NOR2_X1 U2598 ( .A1(n4694), .A2(n4695), .ZN(n4693) );
  NAND2_X1 U2599 ( .A1(n4723), .A2(n4724), .ZN(n4722) );
  XNOR2_X1 U2600 ( .A(n2983), .B(n4890), .ZN(n4728) );
  NAND2_X1 U2601 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4728), .ZN(n4727) );
  NAND2_X1 U2602 ( .A1(n3026), .A2(n4753), .ZN(n4762) );
  XNOR2_X1 U2603 ( .A(n3032), .B(n3031), .ZN(n4776) );
  AND2_X1 U2604 ( .A1(n3043), .A2(n3042), .ZN(n4779) );
  AND2_X1 U2605 ( .A1(n4689), .A2(n3958), .ZN(n4780) );
  XNOR2_X1 U2606 ( .A(n2309), .B(n3039), .ZN(n2308) );
  NAND2_X1 U2607 ( .A1(n2311), .A2(n2310), .ZN(n2309) );
  NAND2_X1 U2608 ( .A1(n3214), .A2(REG2_REG_18__SCAN_IN), .ZN(n2310) );
  AND2_X1 U2609 ( .A1(n2950), .A2(n2884), .ZN(n4068) );
  AOI21_X1 U2610 ( .B1(n2339), .B2(n3092), .A(n3091), .ZN(n4070) );
  OAI21_X1 U2611 ( .B1(n3448), .B2(n3069), .A(n3068), .ZN(n3533) );
  OAI21_X1 U2612 ( .B1(n3383), .B2(n2338), .A(n2334), .ZN(n3366) );
  NAND2_X1 U2613 ( .A1(n4849), .A2(n3417), .ZN(n4905) );
  NAND2_X1 U2614 ( .A1(n3352), .A2(n3054), .ZN(n3337) );
  NAND2_X1 U2615 ( .A1(n3153), .A2(n3269), .ZN(n4909) );
  INV_X1 U2616 ( .A(n4905), .ZN(n4940) );
  INV_X1 U2617 ( .A(n4875), .ZN(n4873) );
  AND2_X2 U2618 ( .A1(n3164), .A2(n3163), .ZN(n4875) );
  INV_X2 U2619 ( .A(n4876), .ZN(n4879) );
  AND2_X1 U2620 ( .A1(n3002), .A2(STATE_REG_SCAN_IN), .ZN(n3225) );
  NAND2_X1 U2621 ( .A1(n3224), .A2(n3269), .ZN(n4470) );
  NOR2_X1 U2622 ( .A1(n2480), .A2(n2445), .ZN(n2446) );
  NOR2_X1 U2623 ( .A1(IR_REG_25__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2445)
         );
  INV_X1 U2624 ( .A(n3031), .ZN(n4939) );
  NAND2_X1 U2625 ( .A1(n2319), .A2(IR_REG_31__SCAN_IN), .ZN(n2520) );
  INV_X1 U2626 ( .A(n3988), .ZN(n4468) );
  AND4_X1 U2627 ( .A1(n4680), .A2(n4679), .A3(n4678), .A4(n4677), .ZN(n4685)
         );
  OR2_X1 U2628 ( .A1(n4037), .A2(n4406), .ZN(n3161) );
  OR2_X1 U2629 ( .A1(n4037), .A2(n4459), .ZN(n3167) );
  BUF_X1 U2630 ( .A(n2839), .Z(n3170) );
  INV_X2 U2631 ( .A(n2839), .ZN(n2491) );
  AND2_X4 U2632 ( .A1(n2460), .A2(n2459), .ZN(n2497) );
  AND2_X1 U2633 ( .A1(n2296), .A2(n3068), .ZN(n2274) );
  NAND2_X1 U2634 ( .A1(n2477), .A2(n3190), .ZN(n2510) );
  AND2_X1 U2635 ( .A1(n2364), .A2(n2362), .ZN(n2275) );
  NAND2_X1 U2636 ( .A1(n2371), .A2(n2776), .ZN(n3683) );
  INV_X1 U2637 ( .A(n2354), .ZN(n2353) );
  NAND2_X1 U2638 ( .A1(n2281), .A2(n4136), .ZN(n2354) );
  OR2_X1 U2639 ( .A1(n2444), .A2(n2443), .ZN(n2276) );
  INV_X1 U2640 ( .A(n2350), .ZN(n2349) );
  NAND2_X1 U2641 ( .A1(n2356), .A2(n2351), .ZN(n2350) );
  AND2_X1 U2642 ( .A1(n2374), .A2(n2284), .ZN(n2277) );
  AND2_X1 U2643 ( .A1(n2393), .A2(n2390), .ZN(n2278) );
  OR2_X1 U2644 ( .A1(n3046), .A2(n3045), .ZN(n2279) );
  INV_X1 U2646 ( .A(IR_REG_3__SCAN_IN), .ZN(n2542) );
  NAND2_X1 U2647 ( .A1(n2391), .A2(n2393), .ZN(n3720) );
  NAND2_X1 U2648 ( .A1(n4776), .A2(n4775), .ZN(n4773) );
  NAND2_X1 U2649 ( .A1(n2373), .A2(n2574), .ZN(n2579) );
  NAND2_X1 U2650 ( .A1(n2387), .A2(n2388), .ZN(n3737) );
  AND2_X1 U2651 ( .A1(n2400), .A2(n2398), .ZN(n2280) );
  NAND2_X1 U2652 ( .A1(n3972), .A2(n4212), .ZN(n2281) );
  OR2_X1 U2653 ( .A1(n3190), .A2(n2964), .ZN(n2282) );
  INV_X1 U2654 ( .A(n3312), .ZN(n3307) );
  AND2_X1 U2655 ( .A1(n2380), .A2(n2383), .ZN(n2283) );
  INV_X2 U2656 ( .A(n2319), .ZN(n2575) );
  NAND2_X1 U2657 ( .A1(n2465), .A2(n2358), .ZN(n2478) );
  NAND2_X1 U2658 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2284) );
  INV_X1 U2659 ( .A(n2335), .ZN(n2334) );
  NAND2_X1 U2660 ( .A1(n3062), .A2(n2336), .ZN(n2335) );
  INV_X1 U2661 ( .A(n2737), .ZN(n2426) );
  NAND2_X1 U2662 ( .A1(n2726), .A2(n2425), .ZN(n2737) );
  INV_X1 U2663 ( .A(n2507), .ZN(n2878) );
  NOR2_X1 U2664 ( .A1(IR_REG_26__SCAN_IN), .A2(n2452), .ZN(n2285) );
  AND2_X1 U2665 ( .A1(n2299), .A2(n2304), .ZN(n2286) );
  NAND2_X1 U2666 ( .A1(n2715), .A2(n2466), .ZN(n2725) );
  NAND2_X1 U2667 ( .A1(n2363), .A2(n2275), .ZN(n3526) );
  INV_X1 U2668 ( .A(n3651), .ZN(n2403) );
  AND2_X1 U2669 ( .A1(n2637), .A2(n2423), .ZN(n2639) );
  OR2_X1 U2670 ( .A1(n2401), .A2(n2399), .ZN(n2287) );
  NAND2_X1 U2671 ( .A1(n2345), .A2(n2344), .ZN(n4116) );
  AOI21_X1 U2672 ( .B1(n4230), .B2(n3085), .A(n3084), .ZN(n4207) );
  NAND2_X1 U2673 ( .A1(n2700), .A2(IR_REG_31__SCAN_IN), .ZN(n2715) );
  AND2_X1 U2674 ( .A1(n3710), .A2(n3711), .ZN(n2288) );
  NAND2_X1 U2675 ( .A1(n2639), .A2(n2424), .ZN(n2697) );
  OR2_X1 U2676 ( .A1(n3788), .A2(n3789), .ZN(n2289) );
  INV_X1 U2677 ( .A(n3054), .ZN(n2326) );
  NOR2_X1 U2678 ( .A1(n3970), .A2(n3143), .ZN(n2290) );
  AND2_X1 U2679 ( .A1(n2289), .A2(n3735), .ZN(n2291) );
  OR2_X1 U2680 ( .A1(n3072), .A2(n4301), .ZN(n2292) );
  AND2_X1 U2681 ( .A1(n3768), .A2(n2403), .ZN(n2293) );
  NOR2_X1 U2682 ( .A1(n4085), .A2(n4073), .ZN(n2294) );
  NOR2_X1 U2683 ( .A1(n4171), .A2(n4148), .ZN(n2295) );
  OR2_X1 U2684 ( .A1(n3979), .A2(n3677), .ZN(n2296) );
  NAND2_X1 U2685 ( .A1(n2750), .A2(n3724), .ZN(n2297) );
  NOR2_X1 U2686 ( .A1(n4125), .A2(n4155), .ZN(n2298) );
  INV_X1 U2687 ( .A(n2385), .ZN(n2384) );
  OR2_X1 U2688 ( .A1(n2820), .A2(n2386), .ZN(n2385) );
  AND2_X1 U2689 ( .A1(n3142), .A2(n4084), .ZN(n3091) );
  NOR2_X1 U2690 ( .A1(n3091), .A2(n2290), .ZN(n2343) );
  INV_X1 U2691 ( .A(n3785), .ZN(n4933) );
  NOR2_X1 U2692 ( .A1(n3319), .A2(n3318), .ZN(n3285) );
  INV_X1 U2693 ( .A(IR_REG_11__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U2694 ( .A1(n3383), .A2(n3060), .ZN(n3309) );
  INV_X1 U2695 ( .A(n3768), .ZN(n2396) );
  NAND2_X1 U2696 ( .A1(n2715), .A2(n2374), .ZN(n2376) );
  INV_X1 U2697 ( .A(IR_REG_10__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U2698 ( .A1(n2327), .A2(n3053), .ZN(n3352) );
  AND2_X2 U2699 ( .A1(n2922), .A2(n4788), .ZN(n3160) );
  INV_X1 U2700 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2629) );
  NAND3_X1 U2701 ( .A1(n2451), .A2(n2450), .A3(n2449), .ZN(n3190) );
  OR2_X4 U2702 ( .A1(n3531), .A2(n3677), .ZN(n3599) );
  AOI21_X2 U2704 ( .B1(n4035), .B2(n4871), .A(n4039), .ZN(n3165) );
  OAI21_X2 U2705 ( .B1(n4061), .B2(n3881), .A(n3871), .ZN(n3145) );
  AOI21_X1 U2706 ( .B1(n4183), .B2(n3894), .A(n3892), .ZN(n4119) );
  NAND2_X1 U2707 ( .A1(n3115), .A2(n3838), .ZN(n3493) );
  NAND2_X1 U2708 ( .A1(n3131), .A2(n3835), .ZN(n3575) );
  NOR2_X2 U2709 ( .A1(n4063), .A2(n4062), .ZN(n4061) );
  NOR2_X2 U2710 ( .A1(n3137), .A2(n3136), .ZN(n4183) );
  NAND2_X1 U2711 ( .A1(n3128), .A2(n3852), .ZN(n3885) );
  NAND2_X1 U2712 ( .A1(n3339), .A2(n3340), .ZN(n3338) );
  NAND2_X1 U2713 ( .A1(n3121), .A2(n3850), .ZN(n3603) );
  OR2_X2 U2714 ( .A1(n3390), .A2(n3112), .ZN(n3113) );
  NAND2_X1 U2715 ( .A1(n4190), .A2(n4177), .ZN(n4154) );
  NAND2_X1 U2716 ( .A1(n2480), .A2(n2479), .ZN(n2939) );
  INV_X2 U2717 ( .A(n2700), .ZN(n2465) );
  NAND2_X1 U2718 ( .A1(n4762), .A2(n2304), .ZN(n2300) );
  INV_X1 U2719 ( .A(n2307), .ZN(n4706) );
  NOR2_X1 U2720 ( .A1(n2307), .A2(REG2_REG_7__SCAN_IN), .ZN(n3016) );
  XNOR2_X1 U2721 ( .A(n3014), .B(n4833), .ZN(n4694) );
  AOI21_X1 U2722 ( .B1(n2308), .B2(n4754), .A(n2279), .ZN(n3047) );
  INV_X1 U2723 ( .A(n4027), .ZN(n2311) );
  NAND2_X1 U2724 ( .A1(n2413), .A2(n2314), .ZN(n2312) );
  NAND2_X1 U2725 ( .A1(n2313), .A2(n2312), .ZN(n3240) );
  NAND2_X2 U2726 ( .A1(n2318), .A2(n2317), .ZN(n2319) );
  INV_X2 U2727 ( .A(IR_REG_1__SCAN_IN), .ZN(n2317) );
  INV_X1 U2728 ( .A(n3354), .ZN(n2327) );
  NAND2_X1 U2729 ( .A1(n2325), .A2(n2323), .ZN(n3057) );
  INV_X1 U2730 ( .A(n2324), .ZN(n2323) );
  NAND2_X1 U2731 ( .A1(n3354), .A2(n3054), .ZN(n2325) );
  NAND2_X1 U2732 ( .A1(n3383), .A2(n2333), .ZN(n2328) );
  NAND2_X1 U2733 ( .A1(n2329), .A2(n2328), .ZN(n4846) );
  NAND3_X1 U2734 ( .A1(n2332), .A2(n2334), .A3(n2338), .ZN(n2331) );
  NAND2_X1 U2735 ( .A1(n4078), .A2(n2343), .ZN(n2340) );
  INV_X1 U2736 ( .A(n4078), .ZN(n2339) );
  NAND2_X1 U2737 ( .A1(n2340), .A2(n2341), .ZN(n4043) );
  NAND2_X1 U2738 ( .A1(n4207), .A2(n2346), .ZN(n2345) );
  AND2_X2 U2739 ( .A1(n2465), .A2(n2357), .ZN(n2455) );
  NAND3_X1 U2740 ( .A1(n2367), .A2(n2368), .A3(n2282), .ZN(n3192) );
  NAND2_X1 U2741 ( .A1(n2490), .A2(n3419), .ZN(n2368) );
  NAND2_X1 U2742 ( .A1(n2371), .A2(n2369), .ZN(n3684) );
  NAND2_X1 U2743 ( .A1(n2765), .A2(n3735), .ZN(n3787) );
  NAND4_X2 U2744 ( .A1(n2574), .A2(n2575), .A3(n2419), .A4(n2421), .ZN(n2608)
         );
  NAND2_X1 U2745 ( .A1(n2715), .A2(n2277), .ZN(n2771) );
  INV_X1 U2746 ( .A(n2771), .ZN(n2469) );
  NAND2_X1 U2747 ( .A1(n3696), .A2(n2381), .ZN(n2377) );
  OAI21_X1 U2748 ( .B1(n3696), .B2(n2382), .A(n2381), .ZN(n3663) );
  NAND2_X1 U2749 ( .A1(n2377), .A2(n2378), .ZN(n3666) );
  NAND2_X1 U2750 ( .A1(n3766), .A2(n2278), .ZN(n2387) );
  NAND2_X1 U2751 ( .A1(n2637), .A2(n2404), .ZN(n2700) );
  NAND2_X1 U2752 ( .A1(n2561), .A2(n2560), .ZN(n2562) );
  NAND2_X1 U2753 ( .A1(n3405), .A2(n3052), .ZN(n3354) );
  NAND2_X1 U2754 ( .A1(n2515), .A2(REG2_REG_1__SCAN_IN), .ZN(n2498) );
  INV_X1 U2755 ( .A(n2460), .ZN(n3219) );
  OAI21_X2 U2756 ( .B1(n4081), .B2(n3880), .A(n3940), .ZN(n4063) );
  AOI211_X2 U2757 ( .C1(n3639), .C2(n3968), .A(n3150), .B(n3149), .ZN(n3151)
         );
  AND2_X1 U2758 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  OAI21_X2 U2759 ( .B1(n3476), .B2(n3477), .A(n3478), .ZN(n3507) );
  NOR2_X2 U2760 ( .A1(n3273), .A2(n3275), .ZN(n3274) );
  AND2_X1 U2761 ( .A1(n2427), .A2(n2470), .ZN(n2407) );
  AND2_X1 U2762 ( .A1(n4737), .A2(REG1_REG_11__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U2763 ( .A1(n3526), .A2(n4300), .ZN(n2409) );
  AND2_X1 U2764 ( .A1(n3175), .A2(n2415), .ZN(n2410) );
  INV_X1 U2765 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2600) );
  INV_X1 U2766 ( .A(n4888), .ZN(n4716) );
  OR2_X1 U2767 ( .A1(n2661), .A2(n2660), .ZN(n2411) );
  INV_X1 U2768 ( .A(DATAI_0_), .ZN(n2485) );
  AND2_X1 U2769 ( .A1(n3450), .A2(n3494), .ZN(n2412) );
  AND2_X1 U2770 ( .A1(n3012), .A2(n4466), .ZN(n2413) );
  NAND2_X1 U2771 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2414) );
  AND2_X1 U2772 ( .A1(n3180), .A2(n4933), .ZN(n2415) );
  AND2_X1 U2773 ( .A1(n2925), .A2(n2924), .ZN(n2416) );
  NOR2_X1 U2774 ( .A1(n4257), .A2(n4252), .ZN(n2417) );
  AND2_X1 U2775 ( .A1(n3010), .A2(n4467), .ZN(n2418) );
  INV_X1 U2776 ( .A(n3327), .ZN(n2599) );
  INV_X1 U2777 ( .A(IR_REG_4__SCAN_IN), .ZN(n2420) );
  INV_X1 U2778 ( .A(n3890), .ZN(n3136) );
  NAND2_X1 U2779 ( .A1(n2407), .A2(n2429), .ZN(n2430) );
  AND2_X1 U2780 ( .A1(n2862), .A2(n2861), .ZN(n2857) );
  OR2_X1 U2781 ( .A1(n3344), .A2(n2839), .ZN(n2525) );
  NOR2_X1 U2782 ( .A1(n2831), .A2(n4571), .ZN(n2845) );
  INV_X1 U2783 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3034) );
  AND2_X1 U2784 ( .A1(REG3_REG_19__SCAN_IN), .A2(n2777), .ZN(n2790) );
  NAND2_X1 U2785 ( .A1(n3118), .A2(n3117), .ZN(n3119) );
  INV_X1 U2786 ( .A(n4847), .ZN(n3064) );
  INV_X1 U2787 ( .A(IR_REG_26__SCAN_IN), .ZN(n2479) );
  INV_X1 U2788 ( .A(n2817), .ZN(n2821) );
  NAND2_X1 U2789 ( .A1(n2822), .A2(REG3_REG_22__SCAN_IN), .ZN(n2831) );
  INV_X1 U2790 ( .A(n4466), .ZN(n2969) );
  NAND2_X1 U2791 ( .A1(n4020), .A2(n3034), .ZN(n3035) );
  AND2_X1 U2792 ( .A1(n2678), .A2(REG3_REG_12__SCAN_IN), .ZN(n2691) );
  AND3_X1 U2793 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2589) );
  INV_X1 U2794 ( .A(n4192), .ZN(n3703) );
  INV_X1 U2795 ( .A(n3356), .ZN(n3362) );
  INV_X1 U2796 ( .A(n3799), .ZN(n2898) );
  NAND2_X1 U2797 ( .A1(n2555), .A2(IR_REG_0__SCAN_IN), .ZN(n2484) );
  OR2_X1 U2798 ( .A1(n2527), .A2(n2526), .ZN(n2528) );
  AND2_X1 U2799 ( .A1(n4144), .A2(n3139), .ZN(n4167) );
  OR2_X1 U2800 ( .A1(n2644), .A2(n4528), .ZN(n2663) );
  OR2_X1 U2801 ( .A1(n3959), .A2(n3108), .ZN(n4857) );
  INV_X1 U2802 ( .A(n4331), .ZN(n4855) );
  AND2_X1 U2803 ( .A1(n4222), .A2(n4223), .ZN(n4257) );
  AND2_X1 U2804 ( .A1(n2910), .A2(n2449), .ZN(n3223) );
  INV_X1 U2805 ( .A(n2913), .ZN(n2449) );
  AND2_X1 U2806 ( .A1(n3098), .A2(DATAI_23_), .ZN(n4155) );
  NOR2_X1 U2807 ( .A1(n2947), .A2(n3221), .ZN(n3806) );
  AND4_X1 U2808 ( .A1(n2955), .A2(n2954), .A3(n2953), .A4(n2952), .ZN(n4064)
         );
  AND4_X1 U2809 ( .A1(n2868), .A2(n2867), .A3(n2866), .A4(n2865), .ZN(n4123)
         );
  AND4_X1 U2810 ( .A1(n2796), .A2(n2795), .A3(n2794), .A4(n2793), .ZN(n4226)
         );
  AND4_X1 U2811 ( .A1(n2618), .A2(n2617), .A3(n2616), .A4(n2615), .ZN(n3450)
         );
  AND2_X1 U2812 ( .A1(n4689), .A2(n3040), .ZN(n4754) );
  AND2_X1 U2813 ( .A1(n3043), .A2(n3041), .ZN(n4689) );
  AND2_X1 U2814 ( .A1(n4036), .A2(n2951), .ZN(n4044) );
  INV_X1 U2815 ( .A(n4794), .ZN(n4861) );
  NOR2_X1 U2816 ( .A1(n2601), .A2(n2600), .ZN(n2613) );
  INV_X1 U2817 ( .A(n4863), .ZN(n4791) );
  AND2_X1 U2818 ( .A1(n3987), .A2(n3419), .ZN(n3406) );
  OR2_X1 U2819 ( .A1(n4798), .A2(n3962), .ZN(n4804) );
  NAND2_X1 U2820 ( .A1(n4316), .A2(n4804), .ZN(n4871) );
  AND2_X1 U2821 ( .A1(n2739), .A2(n2738), .ZN(n3031) );
  OR2_X1 U2822 ( .A1(n2936), .A2(n2923), .ZN(n3785) );
  INV_X1 U2823 ( .A(n4064), .ZN(n3969) );
  INV_X1 U2824 ( .A(n4226), .ZN(n3972) );
  NAND4_X1 U2825 ( .A1(n2696), .A2(n2695), .A3(n2694), .A4(n2693), .ZN(n3976)
         );
  INV_X1 U2826 ( .A(n4754), .ZN(n4774) );
  INV_X1 U2827 ( .A(n4780), .ZN(n4768) );
  NAND2_X1 U2828 ( .A1(n3160), .A2(n4875), .ZN(n4406) );
  NAND2_X1 U2829 ( .A1(n4879), .A2(n3160), .ZN(n4459) );
  NAND2_X1 U2830 ( .A1(n3164), .A2(n3388), .ZN(n4876) );
  INV_X1 U2831 ( .A(n2782), .ZN(n4851) );
  INV_X1 U2832 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2964) );
  AND3_X2 U2833 ( .A1(n2539), .A2(n2420), .A3(n2542), .ZN(n2574) );
  NOR2_X2 U2834 ( .A1(n2608), .A2(n2422), .ZN(n2637) );
  INV_X1 U2835 ( .A(IR_REG_19__SCAN_IN), .ZN(n2427) );
  INV_X1 U2836 ( .A(IR_REG_20__SCAN_IN), .ZN(n2470) );
  INV_X1 U2837 ( .A(IR_REG_14__SCAN_IN), .ZN(n2428) );
  NAND3_X1 U2838 ( .A1(n2772), .A2(n2428), .A3(n2757), .ZN(n2443) );
  NOR2_X2 U2839 ( .A1(n2439), .A2(n2430), .ZN(n2475) );
  INV_X1 U2840 ( .A(IR_REG_22__SCAN_IN), .ZN(n2431) );
  INV_X1 U2841 ( .A(IR_REG_21__SCAN_IN), .ZN(n2474) );
  AND2_X1 U2842 ( .A1(n2431), .A2(n2474), .ZN(n2434) );
  AND2_X1 U2843 ( .A1(n2434), .A2(n2918), .ZN(n2432) );
  NAND2_X1 U2844 ( .A1(n2475), .A2(n2432), .ZN(n2916) );
  INV_X1 U2845 ( .A(IR_REG_24__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U2846 ( .A1(n2475), .A2(n2434), .ZN(n2917) );
  NAND2_X1 U2847 ( .A1(n2918), .A2(n2435), .ZN(n2436) );
  OR2_X1 U2848 ( .A1(n2438), .A2(n2437), .ZN(n2447) );
  NAND4_X1 U2849 ( .A1(n2442), .A2(n2441), .A3(n2440), .A4(n2918), .ZN(n2444)
         );
  NAND2_X1 U2850 ( .A1(n2447), .A2(n2446), .ZN(n2908) );
  AND2_X1 U2851 ( .A1(n2478), .A2(IR_REG_31__SCAN_IN), .ZN(n2448) );
  NOR2_X1 U2852 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2481)
         );
  INV_X1 U2853 ( .A(n2481), .ZN(n2452) );
  INV_X1 U2854 ( .A(IR_REG_29__SCAN_IN), .ZN(n2453) );
  INV_X1 U2855 ( .A(IR_REG_30__SCAN_IN), .ZN(n3630) );
  INV_X1 U2856 ( .A(n2455), .ZN(n2945) );
  NAND2_X1 U2857 ( .A1(n2945), .A2(IR_REG_31__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U2858 ( .A1(n2497), .A2(REG0_REG_0__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U2859 ( .A1(n2531), .A2(REG3_REG_0__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U2860 ( .A1(n2533), .A2(REG1_REG_0__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U2861 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2466) );
  AND2_X1 U2862 ( .A1(n2737), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U2863 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U2864 ( .A1(n2469), .A2(n2468), .ZN(n2494) );
  XNOR2_X1 U2865 ( .A(n2471), .B(n2470), .ZN(n2486) );
  NAND2_X1 U2866 ( .A1(n2472), .A2(IR_REG_31__SCAN_IN), .ZN(n2473) );
  MUX2_X1 U2867 ( .A(IR_REG_31__SCAN_IN), .B(n2473), .S(IR_REG_21__SCAN_IN), 
        .Z(n2476) );
  NAND2_X1 U2868 ( .A1(n2475), .A2(n2474), .ZN(n2487) );
  NAND2_X1 U2869 ( .A1(n2476), .A2(n2487), .ZN(n3950) );
  NAND2_X1 U2870 ( .A1(n2486), .A2(n3814), .ZN(n2930) );
  INV_X1 U2871 ( .A(n2930), .ZN(n2477) );
  INV_X2 U2872 ( .A(n2556), .ZN(n2490) );
  INV_X1 U2873 ( .A(n2478), .ZN(n2480) );
  NAND2_X2 U2874 ( .A1(n2939), .A2(IR_REG_31__SCAN_IN), .ZN(n3004) );
  NAND2_X4 U2875 ( .A1(n2483), .A2(n2482), .ZN(n2555) );
  OAI21_X2 U2876 ( .B1(n2555), .B2(n2485), .A(n2484), .ZN(n3419) );
  BUF_X1 U2877 ( .A(n2486), .Z(n2922) );
  NAND2_X1 U2878 ( .A1(n2487), .A2(IR_REG_31__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U2879 ( .A1(n3987), .A2(n2491), .ZN(n2493) );
  INV_X1 U2880 ( .A(n3190), .ZN(n2929) );
  AOI22_X1 U2881 ( .A1(n2538), .A2(n3419), .B1(IR_REG_0__SCAN_IN), .B2(n2929), 
        .ZN(n2492) );
  NAND2_X1 U2882 ( .A1(n2493), .A2(n2492), .ZN(n3193) );
  NAND2_X1 U2883 ( .A1(n3192), .A2(n3193), .ZN(n2496) );
  XNOR2_X2 U2884 ( .A(n2494), .B(IR_REG_19__SCAN_IN), .ZN(n2782) );
  NAND2_X1 U2885 ( .A1(n2782), .A2(n3962), .ZN(n2931) );
  NAND2_X1 U2886 ( .A1(n2931), .A2(n2930), .ZN(n2507) );
  NAND2_X1 U2887 ( .A1(n2531), .A2(REG3_REG_1__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U2888 ( .A1(n2533), .A2(REG1_REG_1__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U2889 ( .A1(n2497), .A2(REG0_REG_1__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U2890 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2502)
         );
  NAND2_X1 U2891 ( .A1(n2555), .A2(n4468), .ZN(n2506) );
  NAND2_X1 U2892 ( .A1(n2504), .A2(DATAI_1_), .ZN(n2505) );
  NAND2_X1 U2893 ( .A1(n2506), .A2(n2505), .ZN(n3050) );
  OAI22_X1 U2894 ( .A1(n2509), .A2(n2510), .B1(n3158), .B2(n2556), .ZN(n2508)
         );
  XNOR2_X1 U2895 ( .A(n2508), .B(n2507), .ZN(n2512) );
  OAI22_X1 U2896 ( .A1(n2509), .A2(n2839), .B1(n3158), .B2(n2510), .ZN(n2511)
         );
  XNOR2_X1 U2897 ( .A(n2512), .B(n2511), .ZN(n3280) );
  INV_X1 U2898 ( .A(n2511), .ZN(n2514) );
  INV_X1 U2899 ( .A(n2512), .ZN(n2513) );
  NAND2_X1 U2900 ( .A1(n2497), .A2(REG0_REG_2__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U2901 ( .A1(n2515), .A2(REG2_REG_2__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U2902 ( .A1(n2531), .A2(REG3_REG_2__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U2903 ( .A1(n2533), .A2(REG1_REG_2__SCAN_IN), .ZN(n2516) );
  INV_X1 U2904 ( .A(DATAI_2_), .ZN(n2522) );
  XNOR2_X2 U2905 ( .A(n2520), .B(IR_REG_2__SCAN_IN), .ZN(n3007) );
  OAI22_X1 U2906 ( .A1(n3344), .A2(n2510), .B1(n3362), .B2(n2556), .ZN(n2523)
         );
  XNOR2_X1 U2907 ( .A(n2523), .B(n2878), .ZN(n2527) );
  NAND2_X1 U2908 ( .A1(n2538), .A2(n3356), .ZN(n2524) );
  AND2_X1 U2909 ( .A1(n2525), .A2(n2524), .ZN(n2526) );
  NAND2_X1 U2910 ( .A1(n2527), .A2(n2526), .ZN(n2529) );
  NAND2_X1 U2911 ( .A1(n2528), .A2(n2529), .ZN(n3275) );
  INV_X1 U2912 ( .A(n2529), .ZN(n2530) );
  NOR2_X1 U2913 ( .A1(n3274), .A2(n2530), .ZN(n3319) );
  NAND2_X1 U2914 ( .A1(n2844), .A2(REG0_REG_3__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U2916 ( .A1(n3103), .A2(REG2_REG_3__SCAN_IN), .ZN(n2536) );
  INV_X1 U2917 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U2918 ( .A1(n2531), .A2(n2532), .ZN(n2535) );
  NAND2_X1 U2919 ( .A1(n2533), .A2(REG1_REG_3__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U2920 ( .A1(n3985), .A2(n2538), .ZN(n2546) );
  AND2_X1 U2921 ( .A1(n2575), .A2(n2539), .ZN(n2540) );
  NOR2_X1 U2922 ( .A1(n2540), .A2(n2650), .ZN(n2541) );
  NAND2_X1 U2923 ( .A1(n2541), .A2(IR_REG_3__SCAN_IN), .ZN(n2544) );
  INV_X1 U2924 ( .A(n2541), .ZN(n2543) );
  NAND2_X1 U2925 ( .A1(n2543), .A2(n2542), .ZN(n2553) );
  MUX2_X1 U2926 ( .A(DATAI_3_), .B(n4467), .S(n2555), .Z(n3347) );
  NAND2_X1 U2927 ( .A1(n2490), .A2(n3347), .ZN(n2545) );
  NAND2_X1 U2928 ( .A1(n2546), .A2(n2545), .ZN(n2547) );
  XNOR2_X1 U2929 ( .A(n2547), .B(n2837), .ZN(n2559) );
  INV_X1 U2930 ( .A(n3347), .ZN(n3111) );
  OAI22_X1 U2931 ( .A1(n3110), .A2(n3170), .B1(n3111), .B2(n3169), .ZN(n2558)
         );
  XNOR2_X1 U2932 ( .A(n2559), .B(n2558), .ZN(n3318) );
  NAND2_X1 U2933 ( .A1(n2844), .A2(REG0_REG_4__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U2934 ( .A1(n3103), .A2(REG2_REG_4__SCAN_IN), .ZN(n2551) );
  INV_X1 U2935 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2548) );
  XNOR2_X1 U2936 ( .A(n2548), .B(REG3_REG_3__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U2937 ( .A1(n2273), .A2(n3290), .ZN(n2550) );
  NAND2_X1 U2938 ( .A1(n3102), .A2(REG1_REG_4__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U2939 ( .A1(n2553), .A2(IR_REG_31__SCAN_IN), .ZN(n2554) );
  XNOR2_X1 U2940 ( .A(n2554), .B(IR_REG_4__SCAN_IN), .ZN(n4466) );
  MUX2_X1 U2941 ( .A(DATAI_4_), .B(n4466), .S(n3634), .Z(n3391) );
  OAI22_X1 U2942 ( .A1(n3313), .A2(n3169), .B1(n3398), .B2(n3172), .ZN(n2557)
         );
  XNOR2_X1 U2943 ( .A(n2557), .B(n2837), .ZN(n2564) );
  OAI22_X1 U2944 ( .A1(n3313), .A2(n3170), .B1(n3398), .B2(n3169), .ZN(n2563)
         );
  XNOR2_X1 U2945 ( .A(n2564), .B(n2563), .ZN(n3289) );
  INV_X1 U2946 ( .A(n3289), .ZN(n2561) );
  NOR2_X1 U2947 ( .A1(n2559), .A2(n2558), .ZN(n3286) );
  NAND2_X1 U2948 ( .A1(n2844), .A2(REG0_REG_5__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U2949 ( .A1(n3103), .A2(REG2_REG_5__SCAN_IN), .ZN(n2572) );
  INV_X1 U2950 ( .A(n2589), .ZN(n2588) );
  INV_X1 U2951 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U2952 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2566) );
  NAND2_X1 U2953 ( .A1(n2567), .A2(n2566), .ZN(n2568) );
  NAND2_X1 U2954 ( .A1(n2588), .A2(n2568), .ZN(n3424) );
  INV_X1 U2955 ( .A(n3424), .ZN(n2569) );
  NAND2_X1 U2956 ( .A1(n2273), .A2(n2569), .ZN(n2571) );
  NAND2_X1 U2957 ( .A1(n3102), .A2(REG1_REG_5__SCAN_IN), .ZN(n2570) );
  OR2_X1 U2958 ( .A1(n3393), .A2(n3170), .ZN(n2582) );
  INV_X1 U2959 ( .A(DATAI_5_), .ZN(n4621) );
  AND2_X1 U2960 ( .A1(n2575), .A2(n2574), .ZN(n2576) );
  NOR2_X1 U2961 ( .A1(n2576), .A2(n2650), .ZN(n2577) );
  MUX2_X1 U2962 ( .A(n2650), .B(n2577), .S(IR_REG_5__SCAN_IN), .Z(n2578) );
  INV_X1 U2963 ( .A(n2578), .ZN(n2580) );
  NAND2_X1 U2964 ( .A1(n2580), .A2(n2579), .ZN(n3246) );
  MUX2_X1 U2965 ( .A(n4621), .B(n3246), .S(n3634), .Z(n3312) );
  NAND2_X1 U2966 ( .A1(n2538), .A2(n3307), .ZN(n2581) );
  AND2_X1 U2967 ( .A1(n2582), .A2(n2581), .ZN(n2586) );
  INV_X1 U2968 ( .A(n2586), .ZN(n2585) );
  OAI22_X1 U2969 ( .A1(n3393), .A2(n3169), .B1(n3312), .B2(n3172), .ZN(n2583)
         );
  XNOR2_X1 U2970 ( .A(n2583), .B(n2878), .ZN(n2587) );
  INV_X1 U2971 ( .A(n2587), .ZN(n2584) );
  NAND2_X1 U2972 ( .A1(n2585), .A2(n2584), .ZN(n3296) );
  AND2_X1 U2973 ( .A1(n2587), .A2(n2586), .ZN(n3297) );
  NAND2_X1 U2974 ( .A1(n2844), .A2(REG0_REG_6__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U2975 ( .A1(n3635), .A2(REG2_REG_6__SCAN_IN), .ZN(n2593) );
  INV_X1 U2976 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U2977 ( .A1(n2588), .A2(n3330), .ZN(n2590) );
  NAND2_X1 U2978 ( .A1(n2589), .A2(REG3_REG_6__SCAN_IN), .ZN(n2601) );
  AND2_X1 U2979 ( .A1(n2590), .A2(n2601), .ZN(n4834) );
  NAND2_X1 U2980 ( .A1(n2273), .A2(n4834), .ZN(n2592) );
  NAND2_X1 U2981 ( .A1(n3102), .A2(REG1_REG_6__SCAN_IN), .ZN(n2591) );
  NAND4_X1 U2982 ( .A1(n2594), .A2(n2593), .A3(n2592), .A4(n2591), .ZN(n3982)
         );
  NAND2_X1 U2983 ( .A1(n2579), .A2(IR_REG_31__SCAN_IN), .ZN(n2595) );
  XNOR2_X1 U2984 ( .A(n2595), .B(IR_REG_6__SCAN_IN), .ZN(n3013) );
  MUX2_X1 U2985 ( .A(DATAI_6_), .B(n3013), .S(n3634), .Z(n3375) );
  AOI22_X1 U2986 ( .A1(n3982), .A2(n2491), .B1(n3375), .B2(n2538), .ZN(n3326)
         );
  INV_X1 U2987 ( .A(n3326), .ZN(n2596) );
  INV_X1 U2988 ( .A(n3982), .ZN(n4858) );
  INV_X1 U2989 ( .A(n3375), .ZN(n3368) );
  OAI22_X1 U2990 ( .A1(n4858), .A2(n3169), .B1(n3368), .B2(n3172), .ZN(n2597)
         );
  XOR2_X1 U2991 ( .A(n2837), .B(n2597), .Z(n3327) );
  NAND2_X1 U2992 ( .A1(n2844), .A2(REG0_REG_7__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U2993 ( .A1(n3103), .A2(REG2_REG_7__SCAN_IN), .ZN(n2606) );
  AND2_X1 U2994 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  OR2_X1 U2995 ( .A1(n2602), .A2(n2613), .ZN(n4867) );
  INV_X1 U2996 ( .A(n4867), .ZN(n2603) );
  NAND2_X1 U2997 ( .A1(n2273), .A2(n2603), .ZN(n2605) );
  NAND2_X1 U2998 ( .A1(n3102), .A2(REG1_REG_7__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U2999 ( .A1(n2608), .A2(IR_REG_31__SCAN_IN), .ZN(n2619) );
  XNOR2_X1 U3000 ( .A(n2619), .B(IR_REG_7__SCAN_IN), .ZN(n4703) );
  MUX2_X1 U3001 ( .A(DATAI_7_), .B(n4703), .S(n3634), .Z(n3463) );
  OAI22_X1 U3002 ( .A1(n3369), .A2(n3169), .B1(n4856), .B2(n3172), .ZN(n2609)
         );
  XNOR2_X1 U3003 ( .A(n2609), .B(n2837), .ZN(n2610) );
  OAI22_X1 U3004 ( .A1(n3369), .A2(n3170), .B1(n4856), .B2(n3169), .ZN(n2611)
         );
  XNOR2_X1 U3005 ( .A(n2610), .B(n2611), .ZN(n3462) );
  NAND2_X1 U3006 ( .A1(n2610), .A2(n2611), .ZN(n2612) );
  NAND2_X1 U3007 ( .A1(n2844), .A2(REG0_REG_8__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U3008 ( .A1(n3103), .A2(REG2_REG_8__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U3009 ( .A1(n2613), .A2(REG3_REG_8__SCAN_IN), .ZN(n2630) );
  OR2_X1 U3010 ( .A1(n2613), .A2(REG3_REG_8__SCAN_IN), .ZN(n2614) );
  AND2_X1 U3011 ( .A1(n2630), .A2(n2614), .ZN(n4880) );
  NAND2_X1 U3012 ( .A1(n2273), .A2(n4880), .ZN(n2616) );
  NAND2_X1 U3013 ( .A1(n3102), .A2(REG1_REG_8__SCAN_IN), .ZN(n2615) );
  INV_X1 U3014 ( .A(DATAI_8_), .ZN(n2623) );
  NAND2_X1 U3015 ( .A1(n2619), .A2(n4676), .ZN(n2620) );
  NAND2_X1 U3016 ( .A1(n2620), .A2(IR_REG_31__SCAN_IN), .ZN(n2622) );
  XNOR2_X1 U3017 ( .A(n2622), .B(n2621), .ZN(n3252) );
  MUX2_X1 U3018 ( .A(n2623), .B(n3252), .S(n3634), .Z(n3494) );
  OAI22_X1 U3019 ( .A1(n3450), .A2(n3169), .B1(n3494), .B2(n3172), .ZN(n2624)
         );
  XNOR2_X1 U3020 ( .A(n2624), .B(n2878), .ZN(n2628) );
  OR2_X1 U3021 ( .A1(n3450), .A2(n3170), .ZN(n2626) );
  INV_X1 U3022 ( .A(n3494), .ZN(n3481) );
  NAND2_X1 U3023 ( .A1(n2538), .A2(n3481), .ZN(n2625) );
  AND2_X1 U3024 ( .A1(n2626), .A2(n2625), .ZN(n2627) );
  NOR2_X1 U3025 ( .A1(n2628), .A2(n2627), .ZN(n3477) );
  NAND2_X1 U3026 ( .A1(n2628), .A2(n2627), .ZN(n3478) );
  NAND2_X1 U3027 ( .A1(n2844), .A2(REG0_REG_9__SCAN_IN), .ZN(n2636) );
  NAND2_X1 U3028 ( .A1(n3103), .A2(REG2_REG_9__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U3029 ( .A1(n2630), .A2(n2629), .ZN(n2631) );
  NAND2_X1 U3030 ( .A1(n2644), .A2(n2631), .ZN(n3512) );
  INV_X1 U3031 ( .A(n3512), .ZN(n2632) );
  NAND2_X1 U3032 ( .A1(n2273), .A2(n2632), .ZN(n2634) );
  NAND2_X1 U3033 ( .A1(n3102), .A2(REG1_REG_9__SCAN_IN), .ZN(n2633) );
  NAND4_X1 U3034 ( .A1(n2636), .A2(n2635), .A3(n2634), .A4(n2633), .ZN(n3980)
         );
  NOR2_X1 U3035 ( .A1(n2637), .A2(n2650), .ZN(n2638) );
  MUX2_X1 U3036 ( .A(n2650), .B(n2638), .S(IR_REG_9__SCAN_IN), .Z(n2640) );
  OR2_X1 U3037 ( .A1(n2640), .A2(n2639), .ZN(n4888) );
  MUX2_X1 U3038 ( .A(DATAI_9_), .B(n4716), .S(n3634), .Z(n3509) );
  INV_X1 U3039 ( .A(n3509), .ZN(n3454) );
  OAI22_X1 U3040 ( .A1(n3495), .A2(n3170), .B1(n3454), .B2(n3169), .ZN(n2655)
         );
  NAND2_X1 U3041 ( .A1(n3980), .A2(n2538), .ZN(n2642) );
  NAND2_X1 U3042 ( .A1(n2490), .A2(n3509), .ZN(n2641) );
  NAND2_X1 U3043 ( .A1(n2642), .A2(n2641), .ZN(n2643) );
  XNOR2_X1 U3044 ( .A(n2643), .B(n2837), .ZN(n2654) );
  XOR2_X1 U3045 ( .A(n2655), .B(n2654), .Z(n3508) );
  NAND2_X1 U3046 ( .A1(n3507), .A2(n3508), .ZN(n3506) );
  NAND2_X1 U3047 ( .A1(n2497), .A2(REG0_REG_10__SCAN_IN), .ZN(n2649) );
  NAND2_X1 U3048 ( .A1(n3103), .A2(REG2_REG_10__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3049 ( .A1(n2644), .A2(n4528), .ZN(n2645) );
  AND2_X1 U3050 ( .A1(n2663), .A2(n2645), .ZN(n4892) );
  NAND2_X1 U3051 ( .A1(n2273), .A2(n4892), .ZN(n2647) );
  NAND2_X1 U3052 ( .A1(n3102), .A2(REG1_REG_10__SCAN_IN), .ZN(n2646) );
  OR2_X1 U3053 ( .A1(n2639), .A2(n2650), .ZN(n2651) );
  XNOR2_X1 U3054 ( .A(n2651), .B(IR_REG_10__SCAN_IN), .ZN(n3021) );
  MUX2_X1 U3055 ( .A(DATAI_10_), .B(n3021), .S(n3634), .Z(n3677) );
  OAI22_X1 U3056 ( .A1(n3120), .A2(n3169), .B1(n3535), .B2(n3172), .ZN(n2652)
         );
  XNOR2_X1 U3057 ( .A(n2652), .B(n2837), .ZN(n2659) );
  NOR2_X1 U3058 ( .A1(n3169), .A2(n3535), .ZN(n2653) );
  AOI21_X1 U3059 ( .B1(n3979), .B2(n2491), .A(n2653), .ZN(n2660) );
  XNOR2_X1 U3060 ( .A(n2659), .B(n2660), .ZN(n3675) );
  INV_X1 U3061 ( .A(n2654), .ZN(n2657) );
  INV_X1 U3062 ( .A(n2655), .ZN(n2656) );
  NAND2_X1 U3063 ( .A1(n2657), .A2(n2656), .ZN(n3673) );
  NAND2_X1 U3064 ( .A1(n3506), .A2(n2658), .ZN(n3674) );
  INV_X1 U3065 ( .A(n2659), .ZN(n2661) );
  NAND2_X1 U3066 ( .A1(n2844), .A2(REG0_REG_11__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3067 ( .A1(n3103), .A2(REG2_REG_11__SCAN_IN), .ZN(n2668) );
  INV_X1 U3068 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2662) );
  AND2_X1 U3069 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  OR2_X1 U3070 ( .A1(n2664), .A2(n2678), .ZN(n4910) );
  INV_X1 U3071 ( .A(n4910), .ZN(n2665) );
  NAND2_X1 U3072 ( .A1(n2273), .A2(n2665), .ZN(n2667) );
  NAND2_X1 U3073 ( .A1(n3102), .A2(REG1_REG_11__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3074 ( .A1(n2639), .A2(n2322), .ZN(n2670) );
  NAND2_X1 U3075 ( .A1(n2670), .A2(IR_REG_31__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U3076 ( .A1(n2671), .A2(n2321), .ZN(n2685) );
  OR2_X1 U3077 ( .A1(n2671), .A2(n2321), .ZN(n2672) );
  MUX2_X1 U3078 ( .A(DATAI_11_), .B(n4737), .S(n3634), .Z(n3600) );
  INV_X1 U3079 ( .A(n3600), .ZN(n3606) );
  OAI22_X1 U3080 ( .A1(n3536), .A2(n3169), .B1(n3606), .B2(n3172), .ZN(n2673)
         );
  XNOR2_X1 U3081 ( .A(n2673), .B(n2878), .ZN(n2677) );
  OR2_X1 U3082 ( .A1(n3536), .A2(n2839), .ZN(n2675) );
  NAND2_X1 U3083 ( .A1(n2538), .A2(n3600), .ZN(n2674) );
  NAND2_X1 U3084 ( .A1(n2677), .A2(n2676), .ZN(n3564) );
  NOR2_X1 U3085 ( .A1(n2677), .A2(n2676), .ZN(n3563) );
  NAND2_X1 U3086 ( .A1(n2844), .A2(REG0_REG_12__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3087 ( .A1(n3635), .A2(REG2_REG_12__SCAN_IN), .ZN(n2683) );
  NOR2_X1 U3088 ( .A1(n2678), .A2(REG3_REG_12__SCAN_IN), .ZN(n2679) );
  OR2_X1 U3089 ( .A1(n2691), .A2(n2679), .ZN(n3626) );
  INV_X1 U3090 ( .A(n3626), .ZN(n2680) );
  NAND2_X1 U3091 ( .A1(n2273), .A2(n2680), .ZN(n2682) );
  NAND2_X1 U3092 ( .A1(n3102), .A2(REG1_REG_12__SCAN_IN), .ZN(n2681) );
  NAND4_X1 U3093 ( .A1(n2684), .A2(n2683), .A3(n2682), .A4(n2681), .ZN(n3977)
         );
  NAND2_X1 U3094 ( .A1(n2685), .A2(IR_REG_31__SCAN_IN), .ZN(n2686) );
  XNOR2_X1 U3095 ( .A(n2686), .B(IR_REG_12__SCAN_IN), .ZN(n4915) );
  MUX2_X1 U3096 ( .A(DATAI_12_), .B(n4915), .S(n3634), .Z(n3623) );
  AOI22_X1 U3097 ( .A1(n3977), .A2(n2491), .B1(n3623), .B2(n2538), .ZN(n3620)
         );
  NAND2_X1 U3098 ( .A1(n3619), .A2(n3620), .ZN(n2690) );
  INV_X1 U3099 ( .A(n3977), .ZN(n4309) );
  OAI22_X1 U3100 ( .A1(n4309), .A2(n3169), .B1(n3522), .B2(n3172), .ZN(n2687)
         );
  XNOR2_X1 U3101 ( .A(n2687), .B(n2837), .ZN(n3621) );
  INV_X1 U3102 ( .A(n3620), .ZN(n2689) );
  INV_X1 U3103 ( .A(n3619), .ZN(n2688) );
  NAND2_X1 U3104 ( .A1(n2497), .A2(REG0_REG_13__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3105 ( .A1(n3635), .A2(REG2_REG_13__SCAN_IN), .ZN(n2695) );
  NOR2_X1 U3106 ( .A1(n2691), .A2(REG3_REG_13__SCAN_IN), .ZN(n2692) );
  OR2_X1 U3107 ( .A1(n2709), .A2(n2692), .ZN(n3773) );
  INV_X1 U3108 ( .A(n3773), .ZN(n4322) );
  NAND2_X1 U3109 ( .A1(n2273), .A2(n4322), .ZN(n2694) );
  NAND2_X1 U3110 ( .A1(n3102), .A2(REG1_REG_13__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3111 ( .A1(n3976), .A2(n2538), .ZN(n2702) );
  NAND2_X1 U3112 ( .A1(n2697), .A2(IR_REG_31__SCAN_IN), .ZN(n2698) );
  MUX2_X1 U3113 ( .A(IR_REG_31__SCAN_IN), .B(n2698), .S(IR_REG_13__SCAN_IN), 
        .Z(n2699) );
  AND2_X1 U3114 ( .A1(n2700), .A2(n2699), .ZN(n3027) );
  MUX2_X1 U3115 ( .A(DATAI_13_), .B(n3027), .S(n3634), .Z(n4318) );
  NAND2_X1 U3116 ( .A1(n2490), .A2(n4318), .ZN(n2701) );
  NAND2_X1 U3117 ( .A1(n2702), .A2(n2701), .ZN(n2703) );
  XNOR2_X1 U3118 ( .A(n2703), .B(n2878), .ZN(n2708) );
  INV_X1 U3119 ( .A(n2708), .ZN(n2706) );
  INV_X1 U3120 ( .A(n4318), .ZN(n4310) );
  NOR2_X1 U3121 ( .A1(n3169), .A2(n4310), .ZN(n2704) );
  AOI21_X1 U3122 ( .B1(n3976), .B2(n2491), .A(n2704), .ZN(n2707) );
  INV_X1 U3123 ( .A(n2707), .ZN(n2705) );
  NAND2_X1 U3124 ( .A1(n2706), .A2(n2705), .ZN(n3768) );
  NAND2_X1 U3125 ( .A1(n2497), .A2(REG0_REG_14__SCAN_IN), .ZN(n2714) );
  NAND2_X1 U3126 ( .A1(n3103), .A2(REG2_REG_14__SCAN_IN), .ZN(n2713) );
  OR2_X1 U3127 ( .A1(n2709), .A2(REG3_REG_14__SCAN_IN), .ZN(n2710) );
  AND2_X1 U3128 ( .A1(n2710), .A2(n2718), .ZN(n3654) );
  NAND2_X1 U3129 ( .A1(n2273), .A2(n3654), .ZN(n2712) );
  NAND2_X1 U3130 ( .A1(n3102), .A2(REG1_REG_14__SCAN_IN), .ZN(n2711) );
  XNOR2_X1 U3131 ( .A(n2715), .B(IR_REG_14__SCAN_IN), .ZN(n3209) );
  MUX2_X1 U3132 ( .A(DATAI_14_), .B(n3209), .S(n3634), .Z(n3655) );
  INV_X1 U3133 ( .A(n3655), .ZN(n3556) );
  OAI22_X1 U3134 ( .A1(n4311), .A2(n3170), .B1(n3556), .B2(n3169), .ZN(n3651)
         );
  OAI22_X1 U3135 ( .A1(n4311), .A2(n3169), .B1(n3556), .B2(n3172), .ZN(n2716)
         );
  XNOR2_X1 U3136 ( .A(n2716), .B(n2837), .ZN(n3652) );
  NAND2_X1 U3137 ( .A1(n2497), .A2(REG0_REG_15__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U3138 ( .A1(n3635), .A2(REG2_REG_15__SCAN_IN), .ZN(n2723) );
  INV_X1 U3139 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2717) );
  NAND2_X1 U3140 ( .A1(n2718), .A2(n2717), .ZN(n2719) );
  NAND2_X1 U3141 ( .A1(n2731), .A2(n2719), .ZN(n4937) );
  INV_X1 U3142 ( .A(n4937), .ZN(n2720) );
  NAND2_X1 U3143 ( .A1(n2273), .A2(n2720), .ZN(n2722) );
  NAND2_X1 U3144 ( .A1(n3102), .A2(REG1_REG_15__SCAN_IN), .ZN(n2721) );
  NAND4_X1 U3145 ( .A1(n2724), .A2(n2723), .A3(n2722), .A4(n2721), .ZN(n3975)
         );
  NAND2_X1 U3146 ( .A1(n3975), .A2(n2538), .ZN(n2728) );
  XNOR2_X1 U3147 ( .A(n2725), .B(n2726), .ZN(n4464) );
  MUX2_X1 U31480 ( .A(DATAI_15_), .B(n4464), .S(n3634), .Z(n4919) );
  NAND2_X1 U31490 ( .A1(n2490), .A2(n4919), .ZN(n2727) );
  NAND2_X1 U3150 ( .A1(n2728), .A2(n2727), .ZN(n2729) );
  XNOR2_X1 U3151 ( .A(n2729), .B(n2878), .ZN(n4931) );
  NOR2_X1 U3152 ( .A1(n3169), .A2(n4294), .ZN(n2730) );
  AOI21_X1 U3153 ( .B1(n3975), .B2(n2491), .A(n2730), .ZN(n4930) );
  NAND2_X1 U3154 ( .A1(n2497), .A2(REG0_REG_16__SCAN_IN), .ZN(n2735) );
  NAND2_X1 U3155 ( .A1(n3103), .A2(REG2_REG_16__SCAN_IN), .ZN(n2734) );
  INV_X1 U3156 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4539) );
  AOI21_X1 U3157 ( .B1(n2731), .B2(n4539), .A(n2752), .ZN(n3580) );
  NAND2_X1 U3158 ( .A1(n2273), .A2(n3580), .ZN(n2733) );
  NAND2_X1 U3159 ( .A1(n3102), .A2(REG1_REG_16__SCAN_IN), .ZN(n2732) );
  NAND4_X1 U3160 ( .A1(n2735), .A2(n2734), .A3(n2733), .A4(n2732), .ZN(n4923)
         );
  NAND2_X1 U3161 ( .A1(n4923), .A2(n2538), .ZN(n2742) );
  INV_X1 U3162 ( .A(DATAI_16_), .ZN(n2740) );
  OAI21_X1 U3163 ( .B1(n2725), .B2(IR_REG_15__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2736) );
  MUX2_X1 U3164 ( .A(IR_REG_31__SCAN_IN), .B(n2736), .S(IR_REG_16__SCAN_IN), 
        .Z(n2739) );
  OR2_X1 U3165 ( .A1(n2725), .A2(n2737), .ZN(n2738) );
  MUX2_X1 U3166 ( .A(n2740), .B(n4939), .S(n3634), .Z(n3582) );
  INV_X1 U3167 ( .A(n3582), .ZN(n3728) );
  NAND2_X1 U3168 ( .A1(n2490), .A2(n3728), .ZN(n2741) );
  NAND2_X1 U3169 ( .A1(n2742), .A2(n2741), .ZN(n2743) );
  XNOR2_X1 U3170 ( .A(n2743), .B(n2837), .ZN(n2746) );
  NAND2_X1 U3171 ( .A1(n4923), .A2(n2491), .ZN(n2745) );
  NAND2_X1 U3172 ( .A1(n2538), .A2(n3728), .ZN(n2744) );
  NAND2_X1 U3173 ( .A1(n2745), .A2(n2744), .ZN(n2747) );
  NAND2_X1 U3174 ( .A1(n2746), .A2(n2747), .ZN(n3725) );
  OAI21_X1 U3175 ( .B1(n4931), .B2(n4930), .A(n3725), .ZN(n2751) );
  NAND3_X1 U3176 ( .A1(n3725), .A2(n4930), .A3(n4931), .ZN(n2750) );
  INV_X1 U3177 ( .A(n2746), .ZN(n2749) );
  INV_X1 U3178 ( .A(n2747), .ZN(n2748) );
  NAND2_X1 U3179 ( .A1(n2749), .A2(n2748), .ZN(n3724) );
  NAND2_X1 U3180 ( .A1(n2844), .A2(REG0_REG_17__SCAN_IN), .ZN(n2756) );
  NAND2_X1 U3181 ( .A1(n3103), .A2(REG2_REG_17__SCAN_IN), .ZN(n2755) );
  NAND2_X1 U3182 ( .A1(n2752), .A2(REG3_REG_17__SCAN_IN), .ZN(n2766) );
  OAI21_X1 U3183 ( .B1(REG3_REG_17__SCAN_IN), .B2(n2752), .A(n2766), .ZN(n3741) );
  INV_X1 U3184 ( .A(n3741), .ZN(n4274) );
  NAND2_X1 U3185 ( .A1(n2273), .A2(n4274), .ZN(n2754) );
  NAND2_X1 U3186 ( .A1(n3102), .A2(REG1_REG_17__SCAN_IN), .ZN(n2753) );
  XNOR2_X1 U3187 ( .A(n2376), .B(n2757), .ZN(n4463) );
  MUX2_X1 U3188 ( .A(DATAI_17_), .B(n4463), .S(n3634), .Z(n4271) );
  INV_X1 U3189 ( .A(n4271), .ZN(n3080) );
  OAI22_X1 U3190 ( .A1(n4247), .A2(n3169), .B1(n3080), .B2(n3172), .ZN(n2758)
         );
  XNOR2_X1 U3191 ( .A(n2758), .B(n2837), .ZN(n2761) );
  OR2_X1 U3192 ( .A1(n4247), .A2(n2839), .ZN(n2760) );
  NAND2_X1 U3193 ( .A1(n2538), .A2(n4271), .ZN(n2759) );
  NAND2_X1 U3194 ( .A1(n2760), .A2(n2759), .ZN(n2762) );
  NAND2_X1 U3195 ( .A1(n2761), .A2(n2762), .ZN(n3736) );
  NAND2_X1 U3196 ( .A1(n3737), .A2(n3736), .ZN(n2765) );
  INV_X1 U3197 ( .A(n2761), .ZN(n2764) );
  INV_X1 U3198 ( .A(n2762), .ZN(n2763) );
  NAND2_X1 U3199 ( .A1(n2764), .A2(n2763), .ZN(n3735) );
  NAND2_X1 U3200 ( .A1(n2844), .A2(REG0_REG_18__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U3201 ( .A1(n3635), .A2(REG2_REG_18__SCAN_IN), .ZN(n2769) );
  INV_X1 U3202 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3793) );
  AOI21_X1 U3203 ( .B1(n3793), .B2(n2766), .A(n2777), .ZN(n3791) );
  NAND2_X1 U3204 ( .A1(n2273), .A2(n3791), .ZN(n2768) );
  NAND2_X1 U3205 ( .A1(n3102), .A2(REG1_REG_18__SCAN_IN), .ZN(n2767) );
  XNOR2_X1 U3206 ( .A(n2771), .B(n2772), .ZN(n3214) );
  MUX2_X1 U3207 ( .A(DATAI_18_), .B(n3214), .S(n3634), .Z(n4244) );
  INV_X1 U3208 ( .A(n4244), .ZN(n4241) );
  OAI22_X1 U3209 ( .A1(n4270), .A2(n3169), .B1(n4241), .B2(n3172), .ZN(n2773)
         );
  XNOR2_X1 U32100 ( .A(n2773), .B(n2837), .ZN(n3788) );
  OR2_X1 U32110 ( .A1(n4270), .A2(n3170), .ZN(n2775) );
  NAND2_X1 U32120 ( .A1(n2538), .A2(n4244), .ZN(n2774) );
  NAND2_X1 U32130 ( .A1(n2775), .A2(n2774), .ZN(n3789) );
  NAND2_X1 U32140 ( .A1(n3788), .A2(n3789), .ZN(n2776) );
  NAND2_X1 U32150 ( .A1(n2844), .A2(REG0_REG_19__SCAN_IN), .ZN(n2781) );
  NAND2_X1 U32160 ( .A1(n3103), .A2(REG2_REG_19__SCAN_IN), .ZN(n2780) );
  INV_X1 U32170 ( .A(n2790), .ZN(n2791) );
  OAI21_X1 U32180 ( .B1(REG3_REG_19__SCAN_IN), .B2(n2777), .A(n2791), .ZN(
        n4234) );
  INV_X1 U32190 ( .A(n4234), .ZN(n3691) );
  NAND2_X1 U32200 ( .A1(n2273), .A2(n3691), .ZN(n2779) );
  NAND2_X1 U32210 ( .A1(n3102), .A2(REG1_REG_19__SCAN_IN), .ZN(n2778) );
  NAND4_X1 U32220 ( .A1(n2781), .A2(n2780), .A3(n2779), .A4(n2778), .ZN(n4245)
         );
  NAND2_X1 U32230 ( .A1(n4245), .A2(n2538), .ZN(n2784) );
  INV_X1 U32240 ( .A(DATAI_19_), .ZN(n4497) );
  MUX2_X1 U32250 ( .A(n4497), .B(n2782), .S(n3634), .Z(n4233) );
  INV_X1 U32260 ( .A(n4233), .ZN(n3083) );
  NAND2_X1 U32270 ( .A1(n2490), .A2(n3083), .ZN(n2783) );
  NAND2_X1 U32280 ( .A1(n2784), .A2(n2783), .ZN(n2785) );
  XNOR2_X1 U32290 ( .A(n2785), .B(n2878), .ZN(n2788) );
  NOR2_X1 U32300 ( .A1(n3169), .A2(n4233), .ZN(n2786) );
  AOI21_X1 U32310 ( .B1(n4245), .B2(n2491), .A(n2786), .ZN(n2787) );
  NAND2_X1 U32320 ( .A1(n2788), .A2(n2787), .ZN(n2789) );
  OAI21_X1 U32330 ( .B1(n2788), .B2(n2787), .A(n2789), .ZN(n3686) );
  NAND2_X1 U32340 ( .A1(n2844), .A2(REG0_REG_20__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U32350 ( .A1(n3635), .A2(REG2_REG_20__SCAN_IN), .ZN(n2795) );
  INV_X1 U32360 ( .A(n2802), .ZN(n2804) );
  INV_X1 U32370 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4552) );
  NAND2_X1 U32380 ( .A1(n4552), .A2(n2791), .ZN(n2792) );
  AND2_X1 U32390 ( .A1(n2804), .A2(n2792), .ZN(n3760) );
  NAND2_X1 U32400 ( .A1(n2273), .A2(n3760), .ZN(n2794) );
  NAND2_X1 U32410 ( .A1(n3102), .A2(REG1_REG_20__SCAN_IN), .ZN(n2793) );
  INV_X1 U32420 ( .A(n4212), .ZN(n3133) );
  OAI22_X1 U32430 ( .A1(n4226), .A2(n3169), .B1(n3133), .B2(n3172), .ZN(n2797)
         );
  XNOR2_X1 U32440 ( .A(n2797), .B(n2878), .ZN(n2816) );
  INV_X1 U32450 ( .A(n2816), .ZN(n2801) );
  OR2_X1 U32460 ( .A1(n4226), .A2(n2839), .ZN(n2799) );
  NAND2_X1 U32470 ( .A1(n2538), .A2(n4212), .ZN(n2798) );
  AND2_X1 U32480 ( .A1(n2799), .A2(n2798), .ZN(n2815) );
  INV_X1 U32490 ( .A(n2815), .ZN(n2800) );
  NAND2_X1 U32500 ( .A1(n2801), .A2(n2800), .ZN(n3758) );
  NAND2_X1 U32510 ( .A1(n2844), .A2(REG0_REG_21__SCAN_IN), .ZN(n2809) );
  NAND2_X1 U32520 ( .A1(n3635), .A2(REG2_REG_21__SCAN_IN), .ZN(n2808) );
  INV_X1 U32530 ( .A(n2822), .ZN(n2824) );
  INV_X1 U32540 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U32550 ( .A1(n2804), .A2(n2803), .ZN(n2805) );
  AND2_X1 U32560 ( .A1(n2824), .A2(n2805), .ZN(n3702) );
  NAND2_X1 U32570 ( .A1(n2273), .A2(n3702), .ZN(n2807) );
  NAND2_X1 U32580 ( .A1(n3102), .A2(REG1_REG_21__SCAN_IN), .ZN(n2806) );
  NAND4_X1 U32590 ( .A1(n2809), .A2(n2808), .A3(n2807), .A4(n2806), .ZN(n4204)
         );
  NAND2_X1 U32600 ( .A1(n4204), .A2(n2491), .ZN(n2811) );
  NAND2_X1 U32610 ( .A1(n3098), .A2(DATAI_21_), .ZN(n4192) );
  NAND2_X1 U32620 ( .A1(n2538), .A2(n3703), .ZN(n2810) );
  NAND2_X1 U32630 ( .A1(n2811), .A2(n2810), .ZN(n3698) );
  NAND2_X1 U32640 ( .A1(n4204), .A2(n2538), .ZN(n2813) );
  NAND2_X1 U32650 ( .A1(n2490), .A2(n3703), .ZN(n2812) );
  NAND2_X1 U32660 ( .A1(n2813), .A2(n2812), .ZN(n2814) );
  XNOR2_X1 U32670 ( .A(n2814), .B(n2837), .ZN(n3699) );
  NAND2_X1 U32680 ( .A1(n2816), .A2(n2815), .ZN(n3757) );
  OAI21_X1 U32690 ( .B1(n3698), .B2(n3699), .A(n3757), .ZN(n2817) );
  INV_X1 U32700 ( .A(n3699), .ZN(n2819) );
  INV_X1 U32710 ( .A(n3698), .ZN(n2818) );
  NOR2_X1 U32720 ( .A1(n2819), .A2(n2818), .ZN(n2820) );
  NAND2_X1 U32730 ( .A1(n3635), .A2(REG2_REG_22__SCAN_IN), .ZN(n2829) );
  NAND2_X1 U32740 ( .A1(n3102), .A2(REG1_REG_22__SCAN_IN), .ZN(n2828) );
  INV_X1 U32750 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2823) );
  NAND2_X1 U32760 ( .A1(n2824), .A2(n2823), .ZN(n2825) );
  AND2_X1 U32770 ( .A1(n2831), .A2(n2825), .ZN(n3779) );
  NAND2_X1 U32780 ( .A1(n2273), .A2(n3779), .ZN(n2827) );
  NAND2_X1 U32790 ( .A1(n2844), .A2(REG0_REG_22__SCAN_IN), .ZN(n2826) );
  NAND4_X1 U32800 ( .A1(n2829), .A2(n2828), .A3(n2827), .A4(n2826), .ZN(n4187)
         );
  NAND2_X1 U32810 ( .A1(n3098), .A2(DATAI_22_), .ZN(n4177) );
  OAI22_X1 U32820 ( .A1(n4149), .A2(n3169), .B1(n4177), .B2(n3172), .ZN(n2830)
         );
  XNOR2_X1 U32830 ( .A(n2837), .B(n2830), .ZN(n2843) );
  OAI22_X1 U32840 ( .A1(n4149), .A2(n3170), .B1(n4177), .B2(n3169), .ZN(n2842)
         );
  XNOR2_X1 U32850 ( .A(n2843), .B(n2842), .ZN(n3778) );
  NAND2_X1 U32860 ( .A1(n2844), .A2(REG0_REG_23__SCAN_IN), .ZN(n2836) );
  NAND2_X1 U32870 ( .A1(n3635), .A2(REG2_REG_23__SCAN_IN), .ZN(n2835) );
  INV_X1 U32880 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4571) );
  INV_X1 U32890 ( .A(n2845), .ZN(n2846) );
  NAND2_X1 U32900 ( .A1(n2831), .A2(n4571), .ZN(n2832) );
  NAND2_X1 U32910 ( .A1(n2273), .A2(n4158), .ZN(n2834) );
  NAND2_X1 U32920 ( .A1(n3102), .A2(REG1_REG_23__SCAN_IN), .ZN(n2833) );
  INV_X1 U32930 ( .A(n4155), .ZN(n4148) );
  OAI22_X1 U32940 ( .A1(n4171), .A2(n3169), .B1(n3172), .B2(n4148), .ZN(n2838)
         );
  XNOR2_X1 U32950 ( .A(n2838), .B(n2837), .ZN(n2856) );
  OR2_X1 U32960 ( .A1(n4171), .A2(n2839), .ZN(n2841) );
  NAND2_X1 U32970 ( .A1(n2538), .A2(n4155), .ZN(n2840) );
  NAND2_X1 U32980 ( .A1(n2841), .A2(n2840), .ZN(n2855) );
  XNOR2_X1 U32990 ( .A(n2856), .B(n2855), .ZN(n3664) );
  NOR2_X1 U33000 ( .A1(n2843), .A2(n2842), .ZN(n3665) );
  NOR2_X1 U33010 ( .A1(n3664), .A2(n3665), .ZN(n2859) );
  NAND2_X1 U33020 ( .A1(n2844), .A2(REG0_REG_24__SCAN_IN), .ZN(n2851) );
  NAND2_X1 U33030 ( .A1(n3635), .A2(REG2_REG_24__SCAN_IN), .ZN(n2850) );
  NAND2_X1 U33040 ( .A1(n2845), .A2(REG3_REG_24__SCAN_IN), .ZN(n2870) );
  INV_X1 U33050 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4472) );
  NAND2_X1 U33060 ( .A1(n2846), .A2(n4472), .ZN(n2847) );
  AND2_X1 U33070 ( .A1(n2870), .A2(n2847), .ZN(n4131) );
  NAND2_X1 U33080 ( .A1(n2273), .A2(n4131), .ZN(n2849) );
  NAND2_X1 U33090 ( .A1(n3102), .A2(REG1_REG_24__SCAN_IN), .ZN(n2848) );
  NAND4_X1 U33100 ( .A1(n2851), .A2(n2850), .A3(n2849), .A4(n2848), .ZN(n4151)
         );
  NAND2_X1 U33110 ( .A1(n4151), .A2(n2538), .ZN(n2853) );
  NAND2_X1 U33120 ( .A1(n3098), .A2(DATAI_24_), .ZN(n4122) );
  NAND2_X1 U33130 ( .A1(n2490), .A2(n4128), .ZN(n2852) );
  NAND2_X1 U33140 ( .A1(n2853), .A2(n2852), .ZN(n2854) );
  XNOR2_X1 U33150 ( .A(n2854), .B(n2837), .ZN(n2858) );
  INV_X1 U33160 ( .A(n2858), .ZN(n2862) );
  NAND2_X1 U33170 ( .A1(n2856), .A2(n2855), .ZN(n2861) );
  NAND2_X1 U33180 ( .A1(n3666), .A2(n2857), .ZN(n3747) );
  AND2_X1 U33190 ( .A1(n2859), .A2(n2858), .ZN(n2860) );
  NAND2_X1 U33200 ( .A1(n3663), .A2(n2860), .ZN(n3746) );
  OR2_X1 U33210 ( .A1(n2862), .A2(n2861), .ZN(n3745) );
  AOI22_X1 U33220 ( .A1(n4151), .A2(n2491), .B1(n4128), .B2(n2538), .ZN(n3750)
         );
  AND2_X1 U33230 ( .A1(n3745), .A2(n3750), .ZN(n2863) );
  NAND2_X1 U33240 ( .A1(n3746), .A2(n2863), .ZN(n2864) );
  NAND2_X1 U33250 ( .A1(n3635), .A2(REG2_REG_25__SCAN_IN), .ZN(n2868) );
  NAND2_X1 U33260 ( .A1(n3102), .A2(REG1_REG_25__SCAN_IN), .ZN(n2867) );
  XNOR2_X1 U33270 ( .A(n2870), .B(REG3_REG_25__SCAN_IN), .ZN(n4111) );
  NAND2_X1 U33280 ( .A1(n2273), .A2(n4111), .ZN(n2866) );
  NAND2_X1 U33290 ( .A1(n2497), .A2(REG0_REG_25__SCAN_IN), .ZN(n2865) );
  AND2_X1 U33300 ( .A1(n3098), .A2(DATAI_25_), .ZN(n3713) );
  INV_X1 U33310 ( .A(n3713), .ZN(n4109) );
  OAI22_X1 U33320 ( .A1(n4123), .A2(n3169), .B1(n3172), .B2(n4109), .ZN(n2869)
         );
  XOR2_X1 U33330 ( .A(n2837), .B(n2869), .Z(n3710) );
  AOI22_X1 U33340 ( .A1(n3971), .A2(n2491), .B1(n2538), .B2(n3713), .ZN(n3711)
         );
  NAND2_X1 U33350 ( .A1(n2497), .A2(REG0_REG_26__SCAN_IN), .ZN(n2875) );
  NAND2_X1 U33360 ( .A1(n3635), .A2(REG2_REG_26__SCAN_IN), .ZN(n2874) );
  INV_X1 U33370 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4648) );
  INV_X1 U33380 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3804) );
  OAI21_X1 U33390 ( .B1(n2870), .B2(n4648), .A(n3804), .ZN(n2871) );
  OR3_X2 U33400 ( .A1(n2870), .A2(n4648), .A3(n3804), .ZN(n2883) );
  AND2_X1 U33410 ( .A1(n2871), .A2(n2883), .ZN(n3803) );
  NAND2_X1 U33420 ( .A1(n2273), .A2(n3803), .ZN(n2873) );
  NAND2_X1 U33430 ( .A1(n3102), .A2(REG1_REG_26__SCAN_IN), .ZN(n2872) );
  NAND4_X1 U33440 ( .A1(n2875), .A2(n2874), .A3(n2873), .A4(n2872), .ZN(n4104)
         );
  NAND2_X1 U33450 ( .A1(n4104), .A2(n2538), .ZN(n2877) );
  NAND2_X1 U33460 ( .A1(n3098), .A2(DATAI_26_), .ZN(n4084) );
  INV_X1 U33470 ( .A(n4084), .ZN(n4090) );
  NAND2_X1 U33480 ( .A1(n2490), .A2(n4090), .ZN(n2876) );
  NAND2_X1 U33490 ( .A1(n2877), .A2(n2876), .ZN(n2879) );
  XNOR2_X1 U33500 ( .A(n2879), .B(n2878), .ZN(n2895) );
  NOR2_X1 U33510 ( .A1(n3169), .A2(n4084), .ZN(n2880) );
  AOI21_X1 U33520 ( .B1(n4104), .B2(n2491), .A(n2880), .ZN(n2894) );
  NOR2_X1 U3353 ( .A1(n2895), .A2(n2894), .ZN(n3799) );
  NAND2_X1 U33540 ( .A1(n3635), .A2(REG2_REG_27__SCAN_IN), .ZN(n2888) );
  NAND2_X1 U3355 ( .A1(n3102), .A2(REG1_REG_27__SCAN_IN), .ZN(n2887) );
  INV_X1 U3356 ( .A(n2883), .ZN(n2881) );
  NAND2_X1 U3357 ( .A1(n2881), .A2(REG3_REG_27__SCAN_IN), .ZN(n2950) );
  INV_X1 U3358 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U3359 ( .A1(n2883), .A2(n2882), .ZN(n2884) );
  NAND2_X1 U3360 ( .A1(n2273), .A2(n4068), .ZN(n2886) );
  NAND2_X1 U3361 ( .A1(n2497), .A2(REG0_REG_27__SCAN_IN), .ZN(n2885) );
  AND2_X1 U3362 ( .A1(n3098), .A2(DATAI_27_), .ZN(n3143) );
  OAI22_X1 U3363 ( .A1(n4085), .A2(n3169), .B1(n3172), .B2(n4073), .ZN(n2889)
         );
  XNOR2_X1 U3364 ( .A(n2889), .B(n2837), .ZN(n2893) );
  OR2_X1 U3365 ( .A1(n4085), .A2(n3170), .ZN(n2891) );
  NAND2_X1 U3366 ( .A1(n2538), .A2(n3143), .ZN(n2890) );
  NAND2_X1 U3367 ( .A1(n2891), .A2(n2890), .ZN(n2892) );
  NAND2_X1 U3368 ( .A1(n2893), .A2(n2892), .ZN(n3180) );
  OAI21_X1 U3369 ( .B1(n2893), .B2(n2892), .A(n3180), .ZN(n2924) );
  INV_X1 U3370 ( .A(n2924), .ZN(n2896) );
  NAND2_X1 U3371 ( .A1(n2895), .A2(n2894), .ZN(n3800) );
  NAND2_X1 U3372 ( .A1(n2896), .A2(n3800), .ZN(n2897) );
  INV_X1 U3373 ( .A(n3177), .ZN(n3176) );
  NOR4_X1 U3374 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2903) );
  NOR4_X1 U3375 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2902) );
  NOR4_X1 U3376 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2901) );
  NOR4_X1 U3377 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2900) );
  NAND4_X1 U3378 ( .A1(n2903), .A2(n2902), .A3(n2901), .A4(n2900), .ZN(n2912)
         );
  NOR2_X1 U3379 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_30__SCAN_IN), .ZN(n2907)
         );
  NOR4_X1 U3380 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2906) );
  NOR4_X1 U3381 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2905) );
  NOR4_X1 U3382 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2904) );
  NAND4_X1 U3383 ( .A1(n2907), .A2(n2906), .A3(n2905), .A4(n2904), .ZN(n2911)
         );
  NAND2_X1 U3384 ( .A1(n3212), .A2(n2908), .ZN(n2909) );
  MUX2_X1 U3385 ( .A(n3212), .B(n2909), .S(B_REG_SCAN_IN), .Z(n2910) );
  OAI21_X1 U3386 ( .B1(n2912), .B2(n2911), .A(n3223), .ZN(n3154) );
  NAND2_X1 U3387 ( .A1(n2908), .A2(n2913), .ZN(n4461) );
  AND2_X1 U3388 ( .A1(n3154), .A2(n4461), .ZN(n3386) );
  INV_X1 U3389 ( .A(D_REG_0__SCAN_IN), .ZN(n3227) );
  AND2_X1 U3390 ( .A1(n3212), .A2(n2913), .ZN(n3226) );
  INV_X1 U3391 ( .A(D_REG_1__SCAN_IN), .ZN(n2914) );
  NAND2_X1 U3392 ( .A1(n3223), .A2(n2914), .ZN(n3385) );
  NAND3_X1 U3393 ( .A1(n3386), .A2(n3163), .A3(n3385), .ZN(n2938) );
  OR2_X1 U3394 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2915)
         );
  AND2_X1 U3395 ( .A1(n2916), .A2(n2915), .ZN(n2921) );
  NAND2_X1 U3396 ( .A1(n2917), .A2(IR_REG_31__SCAN_IN), .ZN(n2919) );
  OR2_X1 U3397 ( .A1(n2919), .A2(n2918), .ZN(n2920) );
  NAND2_X1 U3398 ( .A1(n2921), .A2(n2920), .ZN(n3002) );
  INV_X1 U3399 ( .A(n3269), .ZN(n3001) );
  OR2_X1 U3400 ( .A1(n2938), .A2(n3001), .ZN(n2936) );
  NAND2_X1 U3401 ( .A1(n2922), .A2(n2782), .ZN(n2927) );
  AOI21_X1 U3402 ( .B1(n2927), .B2(n4788), .A(n3107), .ZN(n2926) );
  INV_X1 U3403 ( .A(n2926), .ZN(n2923) );
  NAND2_X1 U3404 ( .A1(n3176), .A2(n4933), .ZN(n2961) );
  OAI21_X1 U3405 ( .B1(n3802), .B2(n3799), .A(n3800), .ZN(n2925) );
  NAND2_X1 U3406 ( .A1(n2938), .A2(n2926), .ZN(n2928) );
  NAND2_X1 U3407 ( .A1(n2927), .A2(n3107), .ZN(n3152) );
  NAND2_X1 U3408 ( .A1(n2928), .A2(n3152), .ZN(n3267) );
  OAI21_X1 U3409 ( .B1(n3267), .B2(n2929), .A(STATE_REG_SCAN_IN), .ZN(n2935)
         );
  INV_X1 U3410 ( .A(n2922), .ZN(n4462) );
  NOR2_X1 U3411 ( .A1(n2930), .A2(n2931), .ZN(n2932) );
  NAND2_X1 U3412 ( .A1(n3269), .A2(n2932), .ZN(n2937) );
  OAI21_X1 U3413 ( .B1(U3149), .B2(n4855), .A(n2937), .ZN(n2933) );
  NAND2_X1 U3414 ( .A1(n2938), .A2(n2933), .ZN(n3268) );
  OR2_X1 U3415 ( .A1(n3002), .A2(U3149), .ZN(n4469) );
  AND2_X1 U3416 ( .A1(n3268), .A2(n4469), .ZN(n2934) );
  INV_X1 U3417 ( .A(n4068), .ZN(n2958) );
  NAND2_X1 U3418 ( .A1(n2922), .A2(n4851), .ZN(n4798) );
  NOR2_X1 U3419 ( .A1(n4804), .A2(n3814), .ZN(n3153) );
  OAI21_X1 U3420 ( .B1(n2936), .B2(n4855), .A(n4909), .ZN(n3792) );
  INV_X1 U3421 ( .A(n3792), .ZN(n3688) );
  OR2_X1 U3422 ( .A1(n2938), .A2(n2937), .ZN(n2947) );
  INV_X1 U3423 ( .A(n2939), .ZN(n2941) );
  INV_X1 U3424 ( .A(IR_REG_27__SCAN_IN), .ZN(n2940) );
  AND2_X1 U3425 ( .A1(n2941), .A2(n2940), .ZN(n2942) );
  NOR2_X1 U3426 ( .A1(n2942), .A2(n2650), .ZN(n2943) );
  MUX2_X1 U3427 ( .A(n2650), .B(n2943), .S(IR_REG_28__SCAN_IN), .Z(n2944) );
  INV_X1 U3428 ( .A(n2944), .ZN(n2946) );
  NAND2_X1 U3429 ( .A1(n2946), .A2(n2945), .ZN(n3959) );
  OR2_X1 U3430 ( .A1(n2947), .A2(n3959), .ZN(n3687) );
  INV_X2 U3431 ( .A(n3687), .ZN(n4922) );
  AOI22_X1 U3432 ( .A1(n3143), .A2(n4920), .B1(n4922), .B2(n4104), .ZN(n2957)
         );
  INV_X1 U3433 ( .A(n3959), .ZN(n3221) );
  NAND2_X1 U3434 ( .A1(n2497), .A2(REG0_REG_28__SCAN_IN), .ZN(n2955) );
  NAND2_X1 U3435 ( .A1(n3635), .A2(REG2_REG_28__SCAN_IN), .ZN(n2954) );
  INV_X1 U3436 ( .A(n2950), .ZN(n2948) );
  NAND2_X1 U3437 ( .A1(n2948), .A2(REG3_REG_28__SCAN_IN), .ZN(n4036) );
  INV_X1 U3438 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2949) );
  NAND2_X1 U3439 ( .A1(n2950), .A2(n2949), .ZN(n2951) );
  NAND2_X1 U3440 ( .A1(n2273), .A2(n4044), .ZN(n2953) );
  NAND2_X1 U3441 ( .A1(n3102), .A2(REG1_REG_28__SCAN_IN), .ZN(n2952) );
  AOI22_X1 U3442 ( .A1(n4924), .A2(n3969), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n2956) );
  OAI211_X1 U3443 ( .C1(n4938), .C2(n2958), .A(n2957), .B(n2956), .ZN(n2959)
         );
  INV_X1 U3444 ( .A(n2959), .ZN(n2960) );
  OAI21_X1 U3445 ( .B1(n2961), .B2(n2416), .A(n2960), .ZN(U3211) );
  XNOR2_X1 U3446 ( .A(n3214), .B(REG1_REG_18__SCAN_IN), .ZN(n4025) );
  INV_X1 U3447 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4392) );
  XNOR2_X1 U3448 ( .A(n4464), .B(n4392), .ZN(n4000) );
  INV_X1 U3449 ( .A(n3246), .ZN(n4465) );
  NAND2_X1 U3450 ( .A1(n4465), .A2(REG1_REG_5__SCAN_IN), .ZN(n2972) );
  INV_X1 U3451 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2962) );
  MUX2_X1 U3452 ( .A(REG1_REG_5__SCAN_IN), .B(n2962), .S(n3246), .Z(n2963) );
  INV_X1 U3453 ( .A(n2963), .ZN(n3238) );
  INV_X1 U3454 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4809) );
  INV_X1 U3455 ( .A(IR_REG_0__SCAN_IN), .ZN(n4786) );
  AOI211_X1 U3456 ( .C1(n3988), .C2(n4809), .A(n4786), .B(n2964), .ZN(n2965)
         );
  NAND2_X1 U3457 ( .A1(n4468), .A2(REG1_REG_1__SCAN_IN), .ZN(n2966) );
  NAND2_X1 U34580 ( .A1(n2965), .A2(n2966), .ZN(n3989) );
  NAND2_X1 U34590 ( .A1(n3989), .A2(n2966), .ZN(n3199) );
  INV_X1 U3460 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3363) );
  XNOR2_X1 U3461 ( .A(n3007), .B(n3363), .ZN(n3198) );
  XNOR2_X1 U3462 ( .A(n2967), .B(n4467), .ZN(n3228) );
  INV_X1 U3463 ( .A(n2967), .ZN(n2968) );
  INV_X1 U3464 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U3465 ( .A1(n3238), .A2(n3239), .ZN(n3237) );
  NAND2_X1 U3466 ( .A1(n2972), .A2(n3237), .ZN(n2973) );
  NAND2_X1 U34670 ( .A1(n3013), .A2(n2973), .ZN(n2974) );
  INV_X1 U3468 ( .A(n3013), .ZN(n4833) );
  XNOR2_X1 U34690 ( .A(n2973), .B(n4833), .ZN(n4699) );
  NAND2_X1 U3470 ( .A1(REG1_REG_6__SCAN_IN), .A2(n4699), .ZN(n4698) );
  INV_X1 U34710 ( .A(n4703), .ZN(n4841) );
  INV_X1 U3472 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4874) );
  NOR2_X1 U34730 ( .A1(n4841), .A2(n4874), .ZN(n4709) );
  INV_X1 U3474 ( .A(n2978), .ZN(n2977) );
  NAND2_X1 U34750 ( .A1(n2975), .A2(n3252), .ZN(n2976) );
  INV_X1 U3476 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3504) );
  NOR2_X1 U34770 ( .A1(n3250), .A2(n3504), .ZN(n3249) );
  INV_X1 U3478 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U34790 ( .A1(n4719), .A2(n4715), .ZN(n2979) );
  INV_X1 U3480 ( .A(n4719), .ZN(n2980) );
  INV_X1 U34810 ( .A(n3021), .ZN(n4890) );
  NAND2_X1 U3482 ( .A1(n3021), .A2(n2983), .ZN(n2984) );
  INV_X1 U34830 ( .A(n4915), .ZN(n4758) );
  NOR2_X1 U3484 ( .A1(n2985), .A2(n4758), .ZN(n2986) );
  INV_X1 U34850 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4750) );
  XOR2_X1 U3486 ( .A(n2985), .B(n4915), .Z(n4749) );
  NOR2_X1 U34870 ( .A1(n4750), .A2(n4749), .ZN(n4748) );
  NOR2_X1 U3488 ( .A1(n2986), .A2(n4748), .ZN(n4766) );
  NAND2_X1 U34890 ( .A1(n3027), .A2(REG1_REG_13__SCAN_IN), .ZN(n4764) );
  INV_X1 U3490 ( .A(n3027), .ZN(n4918) );
  INV_X1 U34910 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U3492 ( .A1(n4918), .A2(n4400), .ZN(n4763) );
  INV_X1 U34930 ( .A(n4763), .ZN(n2987) );
  AOI21_X1 U3494 ( .B1(n4766), .B2(n4764), .A(n2987), .ZN(n2988) );
  NAND2_X1 U34950 ( .A1(n3209), .A2(n2988), .ZN(n2989) );
  INV_X1 U3496 ( .A(n3209), .ZN(n3591) );
  XNOR2_X1 U34970 ( .A(n2988), .B(n3591), .ZN(n3595) );
  NAND2_X1 U3498 ( .A1(REG1_REG_14__SCAN_IN), .A2(n3595), .ZN(n3594) );
  NAND2_X1 U34990 ( .A1(n2989), .A2(n3594), .ZN(n3999) );
  AOI22_X1 U3500 ( .A1(n4000), .A2(n3999), .B1(REG1_REG_15__SCAN_IN), .B2(
        n4464), .ZN(n2990) );
  INV_X1 U35010 ( .A(n2990), .ZN(n2991) );
  NOR2_X1 U3502 ( .A1(n3031), .A2(n2991), .ZN(n2992) );
  NOR2_X1 U35030 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4781), .ZN(n4782) );
  NOR2_X1 U3504 ( .A1(n2992), .A2(n4782), .ZN(n4013) );
  INV_X1 U35050 ( .A(n4463), .ZN(n4020) );
  INV_X1 U35060 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2994) );
  NOR2_X1 U35070 ( .A1(n4463), .A2(REG1_REG_17__SCAN_IN), .ZN(n2995) );
  INV_X1 U35080 ( .A(n2995), .ZN(n2993) );
  OAI21_X1 U35090 ( .B1(n4020), .B2(n2994), .A(n2993), .ZN(n4012) );
  NOR2_X1 U35100 ( .A1(n4013), .A2(n4012), .ZN(n4011) );
  NOR2_X2 U35110 ( .A1(n4011), .A2(n2995), .ZN(n4024) );
  INV_X1 U35120 ( .A(n4024), .ZN(n2997) );
  INV_X1 U35130 ( .A(n3214), .ZN(n4034) );
  INV_X1 U35140 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2996) );
  OAI22_X1 U35150 ( .A1(n4025), .A2(n2997), .B1(n4034), .B2(n2996), .ZN(n3000)
         );
  INV_X1 U35160 ( .A(REG1_REG_19__SCAN_IN), .ZN(n2998) );
  MUX2_X1 U35170 ( .A(REG1_REG_19__SCAN_IN), .B(n2998), .S(n2782), .Z(n2999)
         );
  XNOR2_X1 U35180 ( .A(n3000), .B(n2999), .ZN(n3005) );
  NAND2_X1 U35190 ( .A1(n3001), .A2(n4469), .ZN(n3043) );
  NAND2_X1 U35200 ( .A1(n3107), .A2(n3002), .ZN(n3003) );
  AND2_X1 U35210 ( .A1(n3003), .A2(n3098), .ZN(n3041) );
  XNOR2_X1 U35220 ( .A(n3004), .B(IR_REG_27__SCAN_IN), .ZN(n4687) );
  INV_X1 U35230 ( .A(n4687), .ZN(n3958) );
  NAND2_X1 U35240 ( .A1(n3005), .A2(n4780), .ZN(n3048) );
  INV_X1 U35250 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3589) );
  XNOR2_X1 U35260 ( .A(n3988), .B(REG2_REG_1__SCAN_IN), .ZN(n3994) );
  INV_X1 U35270 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4802) );
  NOR2_X1 U35280 ( .A1(n4786), .A2(n4802), .ZN(n3993) );
  NAND2_X1 U35290 ( .A1(n3994), .A2(n3993), .ZN(n3992) );
  NAND2_X1 U35300 ( .A1(n4468), .A2(REG2_REG_1__SCAN_IN), .ZN(n3006) );
  NAND2_X1 U35310 ( .A1(n3992), .A2(n3006), .ZN(n3201) );
  INV_X1 U35320 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3008) );
  MUX2_X1 U35330 ( .A(REG2_REG_2__SCAN_IN), .B(n3008), .S(n3007), .Z(n3202) );
  NAND2_X1 U35340 ( .A1(n3201), .A2(n3202), .ZN(n3200) );
  NAND2_X1 U35350 ( .A1(n3007), .A2(REG2_REG_2__SCAN_IN), .ZN(n3009) );
  INV_X1 U35360 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3231) );
  INV_X1 U35370 ( .A(n3011), .ZN(n3012) );
  XOR2_X1 U35380 ( .A(REG2_REG_5__SCAN_IN), .B(n3246), .Z(n3241) );
  AOI21_X1 U35390 ( .B1(REG2_REG_5__SCAN_IN), .B2(n4465), .A(n3240), .ZN(n3014) );
  NOR2_X1 U35400 ( .A1(n3014), .A2(n4833), .ZN(n3015) );
  INV_X1 U35410 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4695) );
  INV_X1 U35420 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4702) );
  OAI22_X1 U35430 ( .A1(n3016), .A2(n4841), .B1(n4706), .B2(n4702), .ZN(n3018)
         );
  INV_X1 U35440 ( .A(n3252), .ZN(n3017) );
  NAND2_X1 U35450 ( .A1(n3018), .A2(n3017), .ZN(n3019) );
  XNOR2_X1 U35460 ( .A(n3018), .B(n3252), .ZN(n3248) );
  NAND2_X1 U35470 ( .A1(n3248), .A2(REG2_REG_8__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U35480 ( .A1(n3019), .A2(n3247), .ZN(n4723) );
  INV_X1 U35490 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U35500 ( .A1(n4716), .A2(REG2_REG_9__SCAN_IN), .B1(n3456), .B2(
        n4888), .ZN(n4724) );
  NAND2_X1 U35510 ( .A1(n4716), .A2(REG2_REG_9__SCAN_IN), .ZN(n3020) );
  NAND2_X1 U35520 ( .A1(n3021), .A2(n3022), .ZN(n3023) );
  XNOR2_X1 U35530 ( .A(n3022), .B(n4890), .ZN(n4730) );
  NAND2_X1 U35540 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4730), .ZN(n4729) );
  NAND2_X1 U35550 ( .A1(n3023), .A2(n4729), .ZN(n4744) );
  INV_X1 U35560 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4908) );
  INV_X1 U35570 ( .A(n4737), .ZN(n4901) );
  AOI22_X1 U35580 ( .A1(n4737), .A2(REG2_REG_11__SCAN_IN), .B1(n4908), .B2(
        n4901), .ZN(n4745) );
  NAND2_X1 U35590 ( .A1(n4737), .A2(REG2_REG_11__SCAN_IN), .ZN(n3024) );
  NAND2_X1 U35600 ( .A1(n4915), .A2(n3025), .ZN(n3026) );
  XNOR2_X1 U35610 ( .A(n3025), .B(n4758), .ZN(n4755) );
  NAND2_X1 U35620 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4755), .ZN(n4753) );
  INV_X1 U35630 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4760) );
  NOR2_X1 U35640 ( .A1(n4918), .A2(n4760), .ZN(n4759) );
  NOR2_X1 U35650 ( .A1(n3589), .A2(n3588), .ZN(n3587) );
  OR2_X1 U35660 ( .A1(n3587), .A2(n2286), .ZN(n4001) );
  NAND2_X1 U35670 ( .A1(n4464), .A2(REG2_REG_15__SCAN_IN), .ZN(n3030) );
  OR2_X1 U35680 ( .A1(n4464), .A2(REG2_REG_15__SCAN_IN), .ZN(n3028) );
  NAND2_X1 U35690 ( .A1(n3030), .A2(n3028), .ZN(n4004) );
  NAND2_X1 U35700 ( .A1(n3032), .A2(n4939), .ZN(n3033) );
  INV_X1 U35710 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4775) );
  XNOR2_X1 U35720 ( .A(n4020), .B(REG2_REG_17__SCAN_IN), .ZN(n4016) );
  INV_X1 U35730 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3037) );
  NOR2_X1 U35740 ( .A1(n3214), .A2(n3037), .ZN(n3036) );
  AOI21_X1 U35750 ( .B1(n3037), .B2(n3214), .A(n3036), .ZN(n4029) );
  NOR2_X1 U35760 ( .A1(n4028), .A2(n4029), .ZN(n4027) );
  INV_X1 U35770 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3038) );
  MUX2_X1 U35780 ( .A(REG2_REG_19__SCAN_IN), .B(n3038), .S(n2782), .Z(n3039)
         );
  NOR2_X1 U35790 ( .A1(n3959), .A2(n3958), .ZN(n3040) );
  INV_X1 U35800 ( .A(n3041), .ZN(n3042) );
  INV_X1 U35810 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4638) );
  NOR2_X1 U3582 ( .A1(STATE_REG_SCAN_IN), .A2(n4638), .ZN(n3690) );
  AOI21_X1 U3583 ( .B1(n4779), .B2(ADDR_REG_19__SCAN_IN), .A(n3690), .ZN(n3044) );
  INV_X1 U3584 ( .A(n3044), .ZN(n3046) );
  NAND2_X1 U3585 ( .A1(n4689), .A2(n3959), .ZN(n4785) );
  NOR2_X1 U3586 ( .A1(n4785), .A2(n2782), .ZN(n3045) );
  NAND2_X1 U3587 ( .A1(n3048), .A2(n3047), .ZN(U3259) );
  INV_X1 U3588 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3157) );
  NAND2_X2 U3590 ( .A1(n2509), .A2(n3051), .ZN(n3816) );
  NAND2_X1 U3591 ( .A1(n3407), .A2(n3406), .ZN(n3405) );
  NAND2_X1 U3592 ( .A1(n3049), .A2(n3051), .ZN(n3052) );
  NAND2_X1 U3593 ( .A1(n3344), .A2(n3356), .ZN(n3817) );
  NAND2_X1 U3594 ( .A1(n3986), .A2(n3362), .ZN(n3820) );
  INV_X1 U3595 ( .A(n3928), .ZN(n3053) );
  NAND2_X1 U3596 ( .A1(n3344), .A2(n3362), .ZN(n3054) );
  NAND2_X1 U3597 ( .A1(n3985), .A2(n3347), .ZN(n3055) );
  NAND2_X1 U3598 ( .A1(n3110), .A2(n3111), .ZN(n3056) );
  NAND2_X1 U3599 ( .A1(n3057), .A2(n3056), .ZN(n3381) );
  INV_X1 U3600 ( .A(n3381), .ZN(n3059) );
  NAND2_X1 U3601 ( .A1(n3313), .A2(n3391), .ZN(n3823) );
  NAND2_X1 U3602 ( .A1(n3984), .A2(n3398), .ZN(n3826) );
  INV_X1 U3603 ( .A(n3929), .ZN(n3058) );
  NAND2_X1 U3604 ( .A1(n3059), .A2(n3058), .ZN(n3383) );
  NAND2_X1 U3605 ( .A1(n3984), .A2(n3391), .ZN(n3060) );
  NAND2_X1 U3606 ( .A1(n3393), .A2(n3312), .ZN(n3061) );
  NAND2_X1 U3607 ( .A1(n3983), .A2(n3307), .ZN(n3062) );
  AND2_X1 U3608 ( .A1(n3982), .A2(n3375), .ZN(n3063) );
  INV_X1 U3609 ( .A(n4846), .ZN(n3065) );
  NAND2_X1 U3610 ( .A1(n3369), .A2(n3463), .ZN(n3114) );
  NAND2_X1 U3611 ( .A1(n3981), .A2(n4856), .ZN(n3838) );
  NAND2_X1 U3612 ( .A1(n3065), .A2(n3064), .ZN(n3490) );
  NAND2_X1 U3613 ( .A1(n3981), .A2(n3463), .ZN(n3491) );
  NAND2_X1 U3614 ( .A1(n4860), .A2(n3481), .ZN(n3066) );
  AND2_X1 U3615 ( .A1(n3491), .A2(n3066), .ZN(n3067) );
  AND2_X1 U3616 ( .A1(n3980), .A2(n3509), .ZN(n3069) );
  NAND2_X1 U3617 ( .A1(n3495), .A2(n3454), .ZN(n3068) );
  NAND2_X1 U3618 ( .A1(n3536), .A2(n3600), .ZN(n3516) );
  INV_X1 U3619 ( .A(n3536), .ZN(n3978) );
  NAND2_X1 U3620 ( .A1(n3978), .A2(n3606), .ZN(n3518) );
  NAND2_X1 U3621 ( .A1(n3536), .A2(n3606), .ZN(n3527) );
  NAND2_X1 U3622 ( .A1(n4309), .A2(n3522), .ZN(n3070) );
  AND2_X1 U3623 ( .A1(n3527), .A2(n3070), .ZN(n4300) );
  NOR2_X1 U3624 ( .A1(n3976), .A2(n4318), .ZN(n3072) );
  INV_X1 U3625 ( .A(n3072), .ZN(n3071) );
  AND2_X1 U3626 ( .A1(n4300), .A2(n3071), .ZN(n3073) );
  NAND2_X1 U3627 ( .A1(n3977), .A2(n3623), .ZN(n4301) );
  NAND2_X1 U3628 ( .A1(n4311), .A2(n3655), .ZN(n4280) );
  INV_X1 U3629 ( .A(n4311), .ZN(n4921) );
  NAND2_X1 U3630 ( .A1(n4921), .A2(n3556), .ZN(n3834) );
  NAND2_X1 U3631 ( .A1(n4280), .A2(n3834), .ZN(n3924) );
  NAND2_X1 U3632 ( .A1(n3975), .A2(n4919), .ZN(n3074) );
  NAND2_X1 U3633 ( .A1(n3976), .A2(n4318), .ZN(n3547) );
  AND3_X1 U3634 ( .A1(n3924), .A2(n3074), .A3(n3547), .ZN(n3077) );
  NAND2_X1 U3635 ( .A1(n4311), .A2(n3556), .ZN(n4286) );
  INV_X1 U3636 ( .A(n3074), .ZN(n3075) );
  OAI22_X1 U3637 ( .A1(n4286), .A2(n3075), .B1(n3975), .B2(n4919), .ZN(n3076)
         );
  NAND2_X1 U3638 ( .A1(n4923), .A2(n3582), .ZN(n3883) );
  INV_X1 U3639 ( .A(n3883), .ZN(n3078) );
  NOR2_X1 U3640 ( .A1(n4923), .A2(n3582), .ZN(n3886) );
  NAND2_X1 U3641 ( .A1(n3573), .A2(n3574), .ZN(n3572) );
  NAND2_X1 U3642 ( .A1(n4923), .A2(n3728), .ZN(n4262) );
  INV_X1 U3643 ( .A(n4247), .ZN(n3974) );
  NAND2_X1 U3644 ( .A1(n3974), .A2(n4271), .ZN(n3079) );
  AND2_X1 U3645 ( .A1(n4262), .A2(n3079), .ZN(n4251) );
  NAND2_X1 U3646 ( .A1(n4270), .A2(n4244), .ZN(n4222) );
  INV_X1 U3647 ( .A(n4270), .ZN(n3973) );
  NAND2_X1 U3648 ( .A1(n3973), .A2(n4241), .ZN(n4223) );
  INV_X1 U3649 ( .A(n4257), .ZN(n3927) );
  AND2_X1 U3650 ( .A1(n4251), .A2(n3927), .ZN(n3081) );
  NAND2_X1 U3651 ( .A1(n4247), .A2(n3080), .ZN(n4252) );
  NAND2_X1 U3652 ( .A1(n4270), .A2(n4241), .ZN(n3082) );
  NAND2_X1 U3653 ( .A1(n4254), .A2(n3082), .ZN(n4230) );
  NAND2_X1 U3654 ( .A1(n4245), .A2(n3083), .ZN(n3085) );
  NOR2_X1 U3655 ( .A1(n4245), .A2(n3083), .ZN(n3084) );
  NAND2_X1 U3656 ( .A1(n4226), .A2(n3133), .ZN(n3086) );
  NAND2_X1 U3657 ( .A1(n4204), .A2(n3703), .ZN(n4136) );
  INV_X1 U3658 ( .A(n4177), .ZN(n3780) );
  NAND2_X1 U3659 ( .A1(n4149), .A2(n3780), .ZN(n4144) );
  NAND2_X1 U3660 ( .A1(n4187), .A2(n4177), .ZN(n3139) );
  NOR2_X1 U3661 ( .A1(n4204), .A2(n3703), .ZN(n4137) );
  NOR2_X1 U3662 ( .A1(n4149), .A2(n4177), .ZN(n4139) );
  INV_X1 U3663 ( .A(n4171), .ZN(n4125) );
  INV_X1 U3664 ( .A(n4116), .ZN(n3089) );
  INV_X1 U3665 ( .A(n4151), .ZN(n3141) );
  OAI21_X1 U3666 ( .B1(n3713), .B2(n3971), .A(n4097), .ZN(n3090) );
  OAI21_X1 U3667 ( .B1(n4123), .B2(n4109), .A(n3090), .ZN(n4078) );
  INV_X1 U3668 ( .A(n4104), .ZN(n3142) );
  INV_X1 U3669 ( .A(n4085), .ZN(n3970) );
  AND2_X1 U3670 ( .A1(n3098), .A2(DATAI_28_), .ZN(n3179) );
  NAND2_X1 U3671 ( .A1(n4064), .A2(n3179), .ZN(n3144) );
  INV_X1 U3672 ( .A(n3179), .ZN(n4052) );
  NAND2_X1 U3673 ( .A1(n3969), .A2(n4052), .ZN(n3871) );
  AOI22_X1 U3674 ( .A1(n4043), .A2(n4050), .B1(n3179), .B2(n3969), .ZN(n3099)
         );
  NAND2_X1 U3675 ( .A1(n2497), .A2(REG0_REG_29__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3676 ( .A1(n3103), .A2(REG2_REG_29__SCAN_IN), .ZN(n3096) );
  INV_X1 U3677 ( .A(n4036), .ZN(n3093) );
  NAND2_X1 U3678 ( .A1(n2273), .A2(n3093), .ZN(n3095) );
  NAND2_X1 U3679 ( .A1(n3102), .A2(REG1_REG_29__SCAN_IN), .ZN(n3094) );
  NAND4_X1 U3680 ( .A1(n3097), .A2(n3096), .A3(n3095), .A4(n3094), .ZN(n4054)
         );
  NAND2_X1 U3681 ( .A1(n3098), .A2(DATAI_29_), .ZN(n3874) );
  XNOR2_X1 U3682 ( .A(n4054), .B(n3874), .ZN(n3947) );
  XNOR2_X1 U3683 ( .A(n3099), .B(n3947), .ZN(n4035) );
  XNOR2_X1 U3684 ( .A(n3962), .B(n2930), .ZN(n3100) );
  NAND2_X1 U3685 ( .A1(n3100), .A2(n2782), .ZN(n4316) );
  NAND2_X1 U3686 ( .A1(n3959), .A2(n3107), .ZN(n4794) );
  AND2_X1 U3687 ( .A1(n4687), .A2(B_REG_SCAN_IN), .ZN(n3101) );
  NOR2_X1 U3688 ( .A1(n4794), .A2(n3101), .ZN(n3639) );
  NAND2_X1 U3689 ( .A1(n3102), .A2(REG1_REG_30__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U3690 ( .A1(n3103), .A2(REG2_REG_30__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U3691 ( .A1(n2497), .A2(REG0_REG_30__SCAN_IN), .ZN(n3104) );
  NAND3_X1 U3692 ( .A1(n3106), .A2(n3105), .A3(n3104), .ZN(n3968) );
  INV_X1 U3693 ( .A(n3107), .ZN(n3108) );
  OAI22_X1 U3694 ( .A1(n4064), .A2(n4857), .B1(n3874), .B2(n4855), .ZN(n3150)
         );
  INV_X1 U3695 ( .A(n3987), .ZN(n3410) );
  NAND2_X1 U3696 ( .A1(n3410), .A2(n3419), .ZN(n3943) );
  NAND2_X1 U3697 ( .A1(n3408), .A2(n3816), .ZN(n3355) );
  NAND2_X1 U3698 ( .A1(n3355), .A2(n3928), .ZN(n3109) );
  NAND2_X1 U3699 ( .A1(n3109), .A2(n3817), .ZN(n3339) );
  NAND2_X1 U3700 ( .A1(n3110), .A2(n3347), .ZN(n3822) );
  NAND2_X1 U3701 ( .A1(n3985), .A2(n3111), .ZN(n3819) );
  AND2_X1 U3702 ( .A1(n3822), .A2(n3819), .ZN(n3340) );
  NAND2_X1 U3703 ( .A1(n3338), .A2(n3822), .ZN(n3390) );
  INV_X1 U3704 ( .A(n3823), .ZN(n3112) );
  NAND2_X1 U3705 ( .A1(n3113), .A2(n3826), .ZN(n3311) );
  AND2_X1 U3706 ( .A1(n3983), .A2(n3312), .ZN(n3310) );
  NAND2_X1 U3707 ( .A1(n3393), .A2(n3307), .ZN(n3840) );
  OAI21_X2 U3708 ( .B1(n3311), .B2(n3310), .A(n3840), .ZN(n3367) );
  NAND2_X1 U3709 ( .A1(n3982), .A2(n3368), .ZN(n3839) );
  NAND2_X1 U3710 ( .A1(n3367), .A2(n3839), .ZN(n4853) );
  NAND2_X1 U3711 ( .A1(n4858), .A2(n3375), .ZN(n4852) );
  AND2_X1 U3712 ( .A1(n4852), .A2(n3114), .ZN(n3828) );
  NAND2_X1 U3713 ( .A1(n4853), .A2(n3828), .ZN(n3115) );
  NAND2_X1 U3714 ( .A1(n3450), .A2(n3481), .ZN(n3831) );
  NAND2_X1 U3715 ( .A1(n3493), .A2(n3831), .ZN(n3116) );
  NAND2_X1 U3716 ( .A1(n4860), .A2(n3494), .ZN(n3837) );
  NAND2_X1 U3717 ( .A1(n3116), .A2(n3837), .ZN(n3449) );
  INV_X1 U3718 ( .A(n3449), .ZN(n3118) );
  AND2_X1 U3719 ( .A1(n3980), .A2(n3454), .ZN(n3836) );
  INV_X1 U3720 ( .A(n3836), .ZN(n3117) );
  NAND2_X1 U3721 ( .A1(n3495), .A2(n3509), .ZN(n3832) );
  NAND2_X1 U3722 ( .A1(n3119), .A2(n3832), .ZN(n3534) );
  NAND2_X1 U3723 ( .A1(n3979), .A2(n3535), .ZN(n3848) );
  NAND2_X1 U3724 ( .A1(n3534), .A2(n3848), .ZN(n3121) );
  NAND2_X1 U3725 ( .A1(n3120), .A2(n3677), .ZN(n3850) );
  NAND2_X1 U3726 ( .A1(n3977), .A2(n3522), .ZN(n4303) );
  NAND2_X1 U3727 ( .A1(n3976), .A2(n4310), .ZN(n3122) );
  NAND2_X1 U3728 ( .A1(n4303), .A2(n3122), .ZN(n3124) );
  INV_X1 U3729 ( .A(n3518), .ZN(n3123) );
  NOR2_X1 U3730 ( .A1(n3124), .A2(n3123), .ZN(n3849) );
  NAND2_X1 U3731 ( .A1(n3603), .A2(n3849), .ZN(n3128) );
  NAND2_X1 U3732 ( .A1(n4309), .A2(n3623), .ZN(n4305) );
  NAND2_X1 U3733 ( .A1(n3516), .A2(n4305), .ZN(n3127) );
  INV_X1 U3734 ( .A(n3124), .ZN(n3126) );
  NOR2_X1 U3735 ( .A1(n3976), .A2(n4310), .ZN(n3125) );
  AOI21_X1 U3736 ( .B1(n3127), .B2(n3126), .A(n3125), .ZN(n3852) );
  INV_X1 U3737 ( .A(n3924), .ZN(n3550) );
  INV_X1 U3738 ( .A(n3975), .ZN(n3554) );
  NAND2_X1 U3739 ( .A1(n3554), .A2(n4919), .ZN(n3851) );
  NAND2_X1 U3740 ( .A1(n3975), .A2(n4294), .ZN(n3835) );
  NAND2_X1 U3741 ( .A1(n3851), .A2(n3835), .ZN(n4288) );
  INV_X1 U3742 ( .A(n4280), .ZN(n3129) );
  NOR2_X1 U3743 ( .A1(n4288), .A2(n3129), .ZN(n3130) );
  NAND2_X1 U3744 ( .A1(n4281), .A2(n3130), .ZN(n3131) );
  INV_X1 U3745 ( .A(n3574), .ZN(n3916) );
  NAND2_X1 U3746 ( .A1(n3575), .A2(n3916), .ZN(n3132) );
  NAND2_X2 U3747 ( .A1(n3132), .A2(n3883), .ZN(n4265) );
  NAND2_X1 U3748 ( .A1(n4245), .A2(n4233), .ZN(n3918) );
  AND2_X1 U3749 ( .A1(n4223), .A2(n3918), .ZN(n4200) );
  NAND2_X1 U3750 ( .A1(n3972), .A2(n3133), .ZN(n3911) );
  OR2_X1 U3751 ( .A1(n4247), .A2(n4271), .ZN(n4219) );
  AND3_X1 U3752 ( .A1(n4200), .A2(n3911), .A3(n4219), .ZN(n3860) );
  INV_X1 U3753 ( .A(n3860), .ZN(n3887) );
  NOR2_X2 U3754 ( .A1(n4265), .A2(n3887), .ZN(n3137) );
  NAND2_X1 U3755 ( .A1(n4247), .A2(n4271), .ZN(n4220) );
  NAND2_X1 U3756 ( .A1(n4222), .A2(n4220), .ZN(n3134) );
  NOR2_X1 U3757 ( .A1(n4245), .A2(n4233), .ZN(n3917) );
  AOI21_X1 U3758 ( .B1(n3134), .B2(n4200), .A(n3917), .ZN(n4201) );
  NAND2_X1 U3759 ( .A1(n4226), .A2(n4212), .ZN(n3912) );
  NAND2_X1 U3760 ( .A1(n4201), .A2(n3912), .ZN(n3135) );
  NAND2_X1 U3761 ( .A1(n3135), .A2(n3911), .ZN(n3890) );
  INV_X1 U3762 ( .A(n4204), .ZN(n3138) );
  NAND2_X1 U3763 ( .A1(n3138), .A2(n3703), .ZN(n4142) );
  AND2_X1 U3764 ( .A1(n4144), .A2(n4142), .ZN(n3894) );
  OR2_X1 U3765 ( .A1(n4171), .A2(n4155), .ZN(n3910) );
  AND2_X1 U3766 ( .A1(n3910), .A2(n3139), .ZN(n3864) );
  AND2_X1 U3767 ( .A1(n4204), .A2(n4192), .ZN(n4141) );
  NAND2_X1 U3768 ( .A1(n4144), .A2(n4141), .ZN(n3140) );
  NAND2_X1 U3769 ( .A1(n3864), .A2(n3140), .ZN(n3892) );
  NAND2_X1 U3770 ( .A1(n4171), .A2(n4155), .ZN(n4117) );
  NAND2_X1 U3771 ( .A1(n3141), .A2(n4128), .ZN(n3909) );
  NAND2_X1 U3772 ( .A1(n4117), .A2(n3909), .ZN(n3896) );
  OR2_X1 U3773 ( .A1(n4123), .A2(n3713), .ZN(n3908) );
  NAND2_X1 U3774 ( .A1(n4151), .A2(n4122), .ZN(n4098) );
  AND2_X1 U3775 ( .A1(n3908), .A2(n4098), .ZN(n3895) );
  INV_X1 U3776 ( .A(n3895), .ZN(n3866) );
  NAND2_X1 U3777 ( .A1(n4123), .A2(n3713), .ZN(n4079) );
  NAND2_X1 U3778 ( .A1(n3142), .A2(n4090), .ZN(n3941) );
  NAND2_X1 U3779 ( .A1(n4079), .A2(n3941), .ZN(n3880) );
  NAND2_X1 U3780 ( .A1(n4104), .A2(n4084), .ZN(n3940) );
  OR2_X1 U3781 ( .A1(n4085), .A2(n3143), .ZN(n3869) );
  NAND2_X1 U3782 ( .A1(n4085), .A2(n3143), .ZN(n4048) );
  NAND2_X1 U3783 ( .A1(n4048), .A2(n3144), .ZN(n3881) );
  XOR2_X1 U3784 ( .A(n3947), .B(n3145), .Z(n3148) );
  NAND2_X1 U3785 ( .A1(n4462), .A2(n3814), .ZN(n3147) );
  NAND2_X1 U3786 ( .A1(n4851), .A2(n3962), .ZN(n3146) );
  NOR2_X1 U3787 ( .A1(n3148), .A2(n4863), .ZN(n3149) );
  INV_X1 U3788 ( .A(n3151), .ZN(n4039) );
  NAND2_X1 U3789 ( .A1(n3385), .A2(n4461), .ZN(n3156) );
  NAND2_X1 U3790 ( .A1(n3269), .A2(n3152), .ZN(n3384) );
  NOR2_X1 U3791 ( .A1(n3153), .A2(n3384), .ZN(n3155) );
  MUX2_X1 U3792 ( .A(n3157), .B(n3165), .S(n4875), .Z(n3162) );
  INV_X2 U3793 ( .A(n3419), .ZN(n4790) );
  AND2_X2 U3794 ( .A1(n3158), .A2(n4790), .ZN(n3418) );
  NAND2_X1 U3795 ( .A1(n3418), .A2(n3362), .ZN(n3361) );
  NOR2_X2 U3796 ( .A1(n3361), .A2(n3347), .ZN(n3399) );
  NAND2_X1 U3797 ( .A1(n4843), .A2(n3494), .ZN(n3489) );
  OR2_X2 U3798 ( .A1(n3489), .A2(n3509), .ZN(n3531) );
  NOR2_X4 U3799 ( .A1(n3599), .A2(n3600), .ZN(n3598) );
  NAND2_X1 U3800 ( .A1(n3598), .A2(n3522), .ZN(n4319) );
  OR2_X2 U3801 ( .A1(n4319), .A2(n4318), .ZN(n4321) );
  OR2_X2 U3802 ( .A1(n4154), .A2(n4155), .ZN(n4157) );
  OR2_X2 U3803 ( .A1(n4157), .A2(n4128), .ZN(n4130) );
  NOR2_X2 U3804 ( .A1(n4130), .A2(n3713), .ZN(n4089) );
  AND2_X2 U3805 ( .A1(n4089), .A2(n4084), .ZN(n4071) );
  NAND2_X2 U3806 ( .A1(n4071), .A2(n4073), .ZN(n4072) );
  OAI21_X1 U3807 ( .B1(n4045), .B2(n3874), .A(n4328), .ZN(n4037) );
  NAND2_X1 U3808 ( .A1(n3162), .A2(n3161), .ZN(U3547) );
  INV_X1 U3809 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3166) );
  INV_X1 U3810 ( .A(n3163), .ZN(n3388) );
  MUX2_X1 U3811 ( .A(n3166), .B(n3165), .S(n4879), .Z(n3168) );
  NAND2_X1 U3812 ( .A1(n3168), .A2(n3167), .ZN(U3515) );
  OAI22_X1 U3813 ( .A1(n4064), .A2(n3170), .B1(n4052), .B2(n3169), .ZN(n3171)
         );
  XNOR2_X1 U3814 ( .A(n3171), .B(n2837), .ZN(n3174) );
  OAI22_X1 U3815 ( .A1(n4064), .A2(n3169), .B1(n4052), .B2(n3172), .ZN(n3173)
         );
  XNOR2_X1 U3816 ( .A(n3174), .B(n3173), .ZN(n3182) );
  INV_X1 U3817 ( .A(n3182), .ZN(n3175) );
  NAND2_X1 U3818 ( .A1(n3176), .A2(n2410), .ZN(n3189) );
  NAND3_X1 U3819 ( .A1(n3177), .A2(n4933), .A3(n3182), .ZN(n3188) );
  INV_X1 U3820 ( .A(n4044), .ZN(n3178) );
  OR2_X1 U3821 ( .A1(n4938), .A2(n3178), .ZN(n3186) );
  AOI22_X1 U3822 ( .A1(n3179), .A2(n4920), .B1(n3806), .B2(n4054), .ZN(n3185)
         );
  AOI22_X1 U3823 ( .A1(n4922), .A2(n3970), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3184) );
  INV_X1 U3824 ( .A(n3180), .ZN(n3181) );
  NAND3_X1 U3825 ( .A1(n3182), .A2(n4933), .A3(n3181), .ZN(n3183) );
  AND4_X1 U3826 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3187)
         );
  NAND3_X1 U3827 ( .A1(n3189), .A2(n3188), .A3(n3187), .ZN(U3217) );
  INV_X1 U3828 ( .A(n3225), .ZN(n3960) );
  AND2_X1 U3829 ( .A1(n4687), .A2(n4802), .ZN(n3191) );
  OR2_X1 U3830 ( .A1(n3959), .A2(n3191), .ZN(n4688) );
  INV_X1 U3831 ( .A(n4688), .ZN(n4686) );
  XOR2_X1 U3832 ( .A(n3192), .B(n3193), .Z(n3266) );
  NAND2_X1 U3833 ( .A1(n3266), .A2(n3958), .ZN(n3194) );
  OAI211_X1 U3834 ( .C1(n3993), .C2(n3958), .A(n3194), .B(n3221), .ZN(n3195)
         );
  OAI211_X1 U3835 ( .C1(IR_REG_0__SCAN_IN), .C2(n4686), .A(n3195), .B(n4683), 
        .ZN(n3260) );
  INV_X1 U3836 ( .A(n3260), .ZN(n3207) );
  INV_X1 U3837 ( .A(n3007), .ZN(n3197) );
  AOI22_X1 U3838 ( .A1(n4779), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3196) );
  OAI21_X1 U3839 ( .B1(n4785), .B2(n3197), .A(n3196), .ZN(n3206) );
  XNOR2_X1 U3840 ( .A(n3199), .B(n3198), .ZN(n3204) );
  OAI211_X1 U3841 ( .C1(n3202), .C2(n3201), .A(n4754), .B(n3200), .ZN(n3203)
         );
  OAI21_X1 U3842 ( .B1(n4768), .B2(n3204), .A(n3203), .ZN(n3205) );
  OR3_X1 U3843 ( .A1(n3207), .A2(n3206), .A3(n3205), .ZN(U3242) );
  MUX2_X1 U3844 ( .A(n3252), .B(n2623), .S(U3149), .Z(n3208) );
  INV_X1 U3845 ( .A(n3208), .ZN(U3344) );
  INV_X1 U3846 ( .A(DATAI_14_), .ZN(n4607) );
  NAND2_X1 U3847 ( .A1(n3209), .A2(STATE_REG_SCAN_IN), .ZN(n3210) );
  OAI21_X1 U3848 ( .B1(STATE_REG_SCAN_IN), .B2(n4607), .A(n3210), .ZN(U3338)
         );
  INV_X1 U3849 ( .A(DATAI_21_), .ZN(n4598) );
  NAND2_X1 U3850 ( .A1(n3814), .A2(STATE_REG_SCAN_IN), .ZN(n3211) );
  OAI21_X1 U3851 ( .B1(STATE_REG_SCAN_IN), .B2(n4598), .A(n3211), .ZN(U3331)
         );
  INV_X1 U3852 ( .A(DATAI_24_), .ZN(n4481) );
  MUX2_X1 U3853 ( .A(n4481), .B(n3212), .S(STATE_REG_SCAN_IN), .Z(n3213) );
  INV_X1 U3854 ( .A(n3213), .ZN(U3328) );
  INV_X1 U3855 ( .A(DATAI_18_), .ZN(n4600) );
  NAND2_X1 U3856 ( .A1(n3214), .A2(STATE_REG_SCAN_IN), .ZN(n3215) );
  OAI21_X1 U3857 ( .B1(STATE_REG_SCAN_IN), .B2(n4600), .A(n3215), .ZN(U3334)
         );
  INV_X1 U3858 ( .A(DATAI_22_), .ZN(n4596) );
  NAND2_X1 U3859 ( .A1(n3962), .A2(STATE_REG_SCAN_IN), .ZN(n3216) );
  OAI21_X1 U3860 ( .B1(STATE_REG_SCAN_IN), .B2(n4596), .A(n3216), .ZN(U3330)
         );
  INV_X1 U3861 ( .A(DATAI_29_), .ZN(n4588) );
  NAND2_X1 U3862 ( .A1(n3217), .A2(STATE_REG_SCAN_IN), .ZN(n3218) );
  OAI21_X1 U3863 ( .B1(STATE_REG_SCAN_IN), .B2(n4588), .A(n3218), .ZN(U3323)
         );
  INV_X1 U3864 ( .A(DATAI_30_), .ZN(n3633) );
  NAND2_X1 U3865 ( .A1(n3219), .A2(STATE_REG_SCAN_IN), .ZN(n3220) );
  OAI21_X1 U3866 ( .B1(STATE_REG_SCAN_IN), .B2(n3633), .A(n3220), .ZN(U3322)
         );
  INV_X1 U3867 ( .A(DATAI_28_), .ZN(n4591) );
  NAND2_X1 U3868 ( .A1(n3221), .A2(STATE_REG_SCAN_IN), .ZN(n3222) );
  OAI21_X1 U3869 ( .B1(STATE_REG_SCAN_IN), .B2(n4591), .A(n3222), .ZN(U3324)
         );
  INV_X1 U3870 ( .A(n3223), .ZN(n3224) );
  AOI22_X1 U3871 ( .A1(n4470), .A2(n3227), .B1(n3226), .B2(n3225), .ZN(U3458)
         );
  NOR2_X1 U3872 ( .A1(n4779), .A2(n4683), .ZN(U3148) );
  INV_X1 U3873 ( .A(n4467), .ZN(n3236) );
  INV_X1 U3874 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3349) );
  XNOR2_X1 U3875 ( .A(n3228), .B(n3349), .ZN(n3233) );
  AOI211_X1 U3876 ( .C1(n3231), .C2(n3230), .A(n3229), .B(n4774), .ZN(n3232)
         );
  AOI21_X1 U3877 ( .B1(n4780), .B2(n3233), .A(n3232), .ZN(n3235) );
  NOR2_X1 U3878 ( .A1(STATE_REG_SCAN_IN), .A2(n2532), .ZN(n3320) );
  AOI21_X1 U3879 ( .B1(n4779), .B2(ADDR_REG_3__SCAN_IN), .A(n3320), .ZN(n3234)
         );
  OAI211_X1 U3880 ( .C1(n3236), .C2(n4785), .A(n3235), .B(n3234), .ZN(U3243)
         );
  OAI211_X1 U3881 ( .C1(n3239), .C2(n3238), .A(n4780), .B(n3237), .ZN(n3245)
         );
  NOR2_X1 U3882 ( .A1(STATE_REG_SCAN_IN), .A2(n2567), .ZN(n3301) );
  AOI211_X1 U3883 ( .C1(n3242), .C2(n3241), .A(n3240), .B(n4774), .ZN(n3243)
         );
  AOI211_X1 U3884 ( .C1(n4779), .C2(ADDR_REG_5__SCAN_IN), .A(n3301), .B(n3243), 
        .ZN(n3244) );
  OAI211_X1 U3885 ( .C1(n4785), .C2(n3246), .A(n3245), .B(n3244), .ZN(U3245)
         );
  OAI211_X1 U3886 ( .C1(n3248), .C2(REG2_REG_8__SCAN_IN), .A(n4754), .B(n3247), 
        .ZN(n3256) );
  AOI211_X1 U3887 ( .C1(n3504), .C2(n3250), .A(n3249), .B(n4768), .ZN(n3254)
         );
  INV_X1 U3888 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4641) );
  NOR2_X1 U3889 ( .A1(STATE_REG_SCAN_IN), .A2(n4641), .ZN(n3482) );
  AOI21_X1 U3890 ( .B1(n4779), .B2(ADDR_REG_8__SCAN_IN), .A(n3482), .ZN(n3251)
         );
  OAI21_X1 U3891 ( .B1(n4785), .B2(n3252), .A(n3251), .ZN(n3253) );
  NOR2_X1 U3892 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  NAND2_X1 U3893 ( .A1(n3256), .A2(n3255), .ZN(U3248) );
  AND2_X1 U3894 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3291) );
  OAI21_X1 U3895 ( .B1(REG2_REG_4__SCAN_IN), .B2(n3257), .A(n4754), .ZN(n3262)
         );
  XNOR2_X1 U3896 ( .A(REG1_REG_4__SCAN_IN), .B(n3258), .ZN(n3259) );
  NAND2_X1 U3897 ( .A1(n4780), .A2(n3259), .ZN(n3261) );
  OAI211_X1 U3898 ( .C1(n3263), .C2(n3262), .A(n3261), .B(n3260), .ZN(n3264)
         );
  AOI211_X1 U3899 ( .C1(n4779), .C2(ADDR_REG_4__SCAN_IN), .A(n3291), .B(n3264), 
        .ZN(n3265) );
  OAI21_X1 U3900 ( .B1(n2969), .B2(n4785), .A(n3265), .ZN(U3244) );
  AOI22_X1 U3901 ( .A1(n3266), .A2(n4933), .B1(n4924), .B2(n3049), .ZN(n3272)
         );
  INV_X1 U3902 ( .A(n3267), .ZN(n3270) );
  NAND3_X1 U3903 ( .A1(n3270), .A2(n3269), .A3(n3268), .ZN(n3281) );
  AOI22_X1 U3904 ( .A1(n3281), .A2(REG3_REG_0__SCAN_IN), .B1(n4920), .B2(n3419), .ZN(n3271) );
  NAND2_X1 U3905 ( .A1(n3272), .A2(n3271), .ZN(U3229) );
  AOI21_X1 U3906 ( .B1(n3273), .B2(n3275), .A(n3274), .ZN(n3278) );
  AOI22_X1 U3907 ( .A1(n4924), .A2(n3985), .B1(n4922), .B2(n3049), .ZN(n3277)
         );
  AOI22_X1 U3908 ( .A1(n3281), .A2(REG3_REG_2__SCAN_IN), .B1(n4920), .B2(n3356), .ZN(n3276) );
  OAI211_X1 U3909 ( .C1(n3278), .C2(n3785), .A(n3277), .B(n3276), .ZN(U3234)
         );
  XNOR2_X1 U3910 ( .A(n3279), .B(n3280), .ZN(n3284) );
  AOI22_X1 U3911 ( .A1(n4922), .A2(n3987), .B1(n4924), .B2(n3986), .ZN(n3283)
         );
  AOI22_X1 U3912 ( .A1(n3281), .A2(REG3_REG_1__SCAN_IN), .B1(n4920), .B2(n3051), .ZN(n3282) );
  OAI211_X1 U3913 ( .C1(n3284), .C2(n3785), .A(n3283), .B(n3282), .ZN(U3219)
         );
  OR2_X1 U3914 ( .A1(n3285), .A2(n3286), .ZN(n3288) );
  AOI211_X1 U3915 ( .C1(n3289), .C2(n3288), .A(n3785), .B(n3287), .ZN(n3295)
         );
  INV_X1 U3916 ( .A(n3290), .ZN(n3400) );
  AOI22_X1 U3917 ( .A1(n3391), .A2(n4920), .B1(n4924), .B2(n3983), .ZN(n3293)
         );
  AOI21_X1 U3918 ( .B1(n4922), .B2(n3985), .A(n3291), .ZN(n3292) );
  OAI211_X1 U3919 ( .C1(n4938), .C2(n3400), .A(n3293), .B(n3292), .ZN(n3294)
         );
  OR2_X1 U3920 ( .A1(n3295), .A2(n3294), .ZN(U3227) );
  INV_X1 U3921 ( .A(n3296), .ZN(n3298) );
  NOR2_X1 U3922 ( .A1(n3298), .A2(n3297), .ZN(n3299) );
  XNOR2_X1 U3923 ( .A(n3300), .B(n3299), .ZN(n3305) );
  AOI22_X1 U3924 ( .A1(n3307), .A2(n3792), .B1(n4924), .B2(n3982), .ZN(n3303)
         );
  AOI21_X1 U3925 ( .B1(n4922), .B2(n3984), .A(n3301), .ZN(n3302) );
  OAI211_X1 U3926 ( .C1(n4938), .C2(n3424), .A(n3303), .B(n3302), .ZN(n3304)
         );
  AOI21_X1 U3927 ( .B1(n3305), .B2(n4933), .A(n3304), .ZN(n3306) );
  INV_X1 U3928 ( .A(n3306), .ZN(U3224) );
  NAND2_X1 U3929 ( .A1(n3397), .A2(n3307), .ZN(n3308) );
  NAND2_X1 U3930 ( .A1(n3376), .A2(n3308), .ZN(n3432) );
  INV_X1 U3931 ( .A(n3310), .ZN(n3825) );
  NAND2_X1 U3932 ( .A1(n3825), .A2(n3840), .ZN(n3926) );
  XOR2_X1 U3933 ( .A(n3309), .B(n3926), .Z(n3428) );
  XOR2_X1 U3934 ( .A(n3926), .B(n3311), .Z(n3316) );
  OAI22_X1 U3935 ( .A1(n3313), .A2(n4857), .B1(n4855), .B2(n3312), .ZN(n3314)
         );
  AOI21_X1 U3936 ( .B1(n4861), .B2(n3982), .A(n3314), .ZN(n3315) );
  OAI21_X1 U3937 ( .B1(n3316), .B2(n4863), .A(n3315), .ZN(n3422) );
  AOI21_X1 U3938 ( .B1(n3428), .B2(n4871), .A(n3422), .ZN(n3435) );
  MUX2_X1 U3939 ( .A(n2962), .B(n3435), .S(n4875), .Z(n3317) );
  OAI21_X1 U3940 ( .B1(n4406), .B2(n3432), .A(n3317), .ZN(U3523) );
  AOI21_X1 U3941 ( .B1(n3319), .B2(n3318), .A(n3285), .ZN(n3325) );
  AOI22_X1 U3942 ( .A1(n3347), .A2(n4920), .B1(n4924), .B2(n3984), .ZN(n3322)
         );
  AOI21_X1 U3943 ( .B1(n4922), .B2(n3986), .A(n3320), .ZN(n3321) );
  OAI211_X1 U3944 ( .C1(n4938), .C2(REG3_REG_3__SCAN_IN), .A(n3322), .B(n3321), 
        .ZN(n3323) );
  INV_X1 U3945 ( .A(n3323), .ZN(n3324) );
  OAI21_X1 U3946 ( .B1(n3325), .B2(n3785), .A(n3324), .ZN(U3215) );
  XNOR2_X1 U3947 ( .A(n3327), .B(n3326), .ZN(n3328) );
  XNOR2_X1 U3948 ( .A(n3329), .B(n3328), .ZN(n3335) );
  INV_X1 U3949 ( .A(n4834), .ZN(n3333) );
  AOI22_X1 U3950 ( .A1(n3375), .A2(n3792), .B1(n4922), .B2(n3983), .ZN(n3332)
         );
  NOR2_X1 U3951 ( .A1(STATE_REG_SCAN_IN), .A2(n3330), .ZN(n4696) );
  AOI21_X1 U3952 ( .B1(n3806), .B2(n3981), .A(n4696), .ZN(n3331) );
  OAI211_X1 U3953 ( .C1(n4938), .C2(n3333), .A(n3332), .B(n3331), .ZN(n3334)
         );
  AOI21_X1 U3954 ( .B1(n3335), .B2(n4933), .A(n3334), .ZN(n3336) );
  INV_X1 U3955 ( .A(n3336), .ZN(U3236) );
  INV_X1 U3956 ( .A(n3340), .ZN(n3934) );
  XNOR2_X1 U3957 ( .A(n3337), .B(n3934), .ZN(n4821) );
  INV_X1 U3958 ( .A(n4821), .ZN(n3346) );
  INV_X1 U3959 ( .A(n4316), .ZN(n4792) );
  OAI21_X1 U3960 ( .B1(n3340), .B2(n3339), .A(n3338), .ZN(n3341) );
  NAND2_X1 U3961 ( .A1(n3341), .A2(n4791), .ZN(n3343) );
  AOI22_X1 U3962 ( .A1(n3984), .A2(n4861), .B1(n4331), .B2(n3347), .ZN(n3342)
         );
  OAI211_X1 U3963 ( .C1(n3344), .C2(n4857), .A(n3343), .B(n3342), .ZN(n3345)
         );
  AOI21_X1 U3964 ( .B1(n4792), .B2(n4821), .A(n3345), .ZN(n4824) );
  OAI21_X1 U3965 ( .B1(n3346), .B2(n4804), .A(n4824), .ZN(n3438) );
  AND2_X1 U3966 ( .A1(n3361), .A2(n3347), .ZN(n3348) );
  OR2_X1 U3967 ( .A1(n3348), .A2(n3399), .ZN(n4819) );
  OAI22_X1 U3968 ( .A1(n4406), .A2(n4819), .B1(n4875), .B2(n3349), .ZN(n3350)
         );
  AOI21_X1 U3969 ( .B1(n3438), .B2(n4875), .A(n3350), .ZN(n3351) );
  INV_X1 U3970 ( .A(n3351), .ZN(U3521) );
  INV_X1 U3971 ( .A(n3352), .ZN(n3353) );
  AOI21_X1 U3972 ( .B1(n3928), .B2(n3354), .A(n3353), .ZN(n4812) );
  XNOR2_X1 U3973 ( .A(n3355), .B(n3928), .ZN(n3360) );
  AOI22_X1 U3974 ( .A1(n3985), .A2(n4861), .B1(n3356), .B2(n4331), .ZN(n3357)
         );
  OAI21_X1 U3975 ( .B1(n2509), .B2(n4857), .A(n3357), .ZN(n3359) );
  NOR2_X1 U3976 ( .A1(n4812), .A2(n4316), .ZN(n3358) );
  AOI211_X1 U3977 ( .C1(n3360), .C2(n4791), .A(n3359), .B(n3358), .ZN(n4818)
         );
  OAI21_X1 U3978 ( .B1(n4812), .B2(n4804), .A(n4818), .ZN(n3442) );
  OAI21_X1 U3979 ( .B1(n3418), .B2(n3362), .A(n3361), .ZN(n4813) );
  OAI22_X1 U3980 ( .A1(n4406), .A2(n4813), .B1(n4875), .B2(n3363), .ZN(n3364)
         );
  AOI21_X1 U3981 ( .B1(n3442), .B2(n4875), .A(n3364), .ZN(n3365) );
  INV_X1 U3982 ( .A(n3365), .ZN(U3520) );
  INV_X1 U3983 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3380) );
  NAND2_X1 U3984 ( .A1(n4852), .A2(n3839), .ZN(n3923) );
  XOR2_X1 U3985 ( .A(n3366), .B(n3923), .Z(n4836) );
  INV_X1 U3986 ( .A(n4836), .ZN(n3374) );
  XNOR2_X1 U3987 ( .A(n3367), .B(n3923), .ZN(n3372) );
  INV_X1 U3988 ( .A(n4857), .ZN(n4267) );
  OAI22_X1 U3989 ( .A1(n3369), .A2(n4794), .B1(n4855), .B2(n3368), .ZN(n3370)
         );
  AOI21_X1 U3990 ( .B1(n4267), .B2(n3983), .A(n3370), .ZN(n3371) );
  OAI21_X1 U3991 ( .B1(n3372), .B2(n4863), .A(n3371), .ZN(n3373) );
  AOI21_X1 U3992 ( .B1(n4836), .B2(n4792), .A(n3373), .ZN(n4839) );
  OAI21_X1 U3993 ( .B1(n4804), .B2(n3374), .A(n4839), .ZN(n3444) );
  NAND2_X1 U3994 ( .A1(n3444), .A2(n4875), .ZN(n3379) );
  AND2_X1 U3995 ( .A1(n3376), .A2(n3375), .ZN(n3377) );
  NOR2_X1 U3996 ( .A1(n4842), .A2(n3377), .ZN(n4835) );
  INV_X1 U3997 ( .A(n4406), .ZN(n3617) );
  NAND2_X1 U3998 ( .A1(n4835), .A2(n3617), .ZN(n3378) );
  OAI211_X1 U3999 ( .C1(n4875), .C2(n3380), .A(n3379), .B(n3378), .ZN(U3524)
         );
  NAND2_X1 U4000 ( .A1(n3381), .A2(n3929), .ZN(n3382) );
  AND2_X1 U4001 ( .A1(n3383), .A2(n3382), .ZN(n4829) );
  INV_X1 U4002 ( .A(n4829), .ZN(n3404) );
  INV_X1 U4003 ( .A(n3384), .ZN(n3387) );
  NAND4_X1 U4004 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), .ZN(n3389)
         );
  OR2_X1 U4005 ( .A1(n2930), .A2(n2782), .ZN(n3423) );
  NOR2_X1 U4006 ( .A1(n4944), .A2(n3423), .ZN(n4895) );
  INV_X1 U4007 ( .A(n4895), .ZN(n4906) );
  XOR2_X1 U4008 ( .A(n3929), .B(n3390), .Z(n3396) );
  AOI22_X1 U4009 ( .A1(n3985), .A2(n4267), .B1(n3391), .B2(n4331), .ZN(n3392)
         );
  OAI21_X1 U4010 ( .B1(n3393), .B2(n4794), .A(n3392), .ZN(n3394) );
  AOI21_X1 U4011 ( .B1(n4829), .B2(n4792), .A(n3394), .ZN(n3395) );
  OAI21_X1 U4012 ( .B1(n3396), .B2(n4863), .A(n3395), .ZN(n4826) );
  OAI211_X1 U4013 ( .C1(n3399), .C2(n3398), .A(n3397), .B(n3160), .ZN(n4825)
         );
  OAI22_X1 U4014 ( .A1(n4825), .A2(n4851), .B1(n3400), .B2(n4909), .ZN(n3401)
         );
  INV_X2 U4015 ( .A(n4944), .ZN(n4849) );
  OAI21_X1 U4016 ( .B1(n4826), .B2(n3401), .A(n4849), .ZN(n3403) );
  NAND2_X1 U4017 ( .A1(n4944), .A2(REG2_REG_4__SCAN_IN), .ZN(n3402) );
  OAI211_X1 U4018 ( .C1(n3404), .C2(n4906), .A(n3403), .B(n3402), .ZN(U3286)
         );
  OAI21_X1 U4019 ( .B1(n3407), .B2(n3406), .A(n3405), .ZN(n4805) );
  INV_X1 U4020 ( .A(n3407), .ZN(n3931) );
  INV_X1 U4021 ( .A(n3943), .ZN(n3815) );
  OAI21_X1 U4022 ( .B1(n3931), .B2(n3815), .A(n3408), .ZN(n3412) );
  AOI22_X1 U4023 ( .A1(n3986), .A2(n4861), .B1(n4331), .B2(n3051), .ZN(n3409)
         );
  OAI21_X1 U4024 ( .B1(n3410), .B2(n4857), .A(n3409), .ZN(n3411) );
  AOI21_X1 U4025 ( .B1(n3412), .B2(n4791), .A(n3411), .ZN(n3413) );
  OAI21_X1 U4026 ( .B1(n4316), .B2(n4805), .A(n3413), .ZN(n4806) );
  INV_X1 U4027 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3415) );
  INV_X1 U4028 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3414) );
  OAI22_X1 U4029 ( .A1(n4849), .A2(n3415), .B1(n3414), .B2(n4909), .ZN(n3416)
         );
  AOI21_X1 U4030 ( .B1(n4806), .B2(n4849), .A(n3416), .ZN(n3421) );
  AND2_X1 U4031 ( .A1(n3160), .A2(n2782), .ZN(n3417) );
  AOI21_X1 U4032 ( .B1(n3419), .B2(n3051), .A(n3418), .ZN(n4808) );
  NAND2_X1 U4033 ( .A1(n4940), .A2(n4808), .ZN(n3420) );
  OAI211_X1 U4034 ( .C1(n4805), .C2(n4906), .A(n3421), .B(n3420), .ZN(U3289)
         );
  INV_X1 U4035 ( .A(n3422), .ZN(n3430) );
  NAND2_X1 U4036 ( .A1(n4316), .A2(n3423), .ZN(n4848) );
  NAND2_X1 U4037 ( .A1(n4849), .A2(n4848), .ZN(n4278) );
  INV_X1 U4038 ( .A(n4278), .ZN(n4290) );
  NOR2_X1 U4039 ( .A1(n3424), .A2(n4909), .ZN(n3425) );
  AOI21_X1 U4040 ( .B1(n4944), .B2(REG2_REG_5__SCAN_IN), .A(n3425), .ZN(n3426)
         );
  OAI21_X1 U4041 ( .B1(n4905), .B2(n3432), .A(n3426), .ZN(n3427) );
  AOI21_X1 U4042 ( .B1(n3428), .B2(n4290), .A(n3427), .ZN(n3429) );
  OAI21_X1 U40430 ( .B1(n3430), .B2(n4944), .A(n3429), .ZN(U3285) );
  INV_X1 U4044 ( .A(REG0_REG_5__SCAN_IN), .ZN(n3431) );
  OAI22_X1 U4045 ( .A1(n4459), .A2(n3432), .B1(n4879), .B2(n3431), .ZN(n3433)
         );
  INV_X1 U4046 ( .A(n3433), .ZN(n3434) );
  OAI21_X1 U4047 ( .B1(n3435), .B2(n4876), .A(n3434), .ZN(U3477) );
  INV_X1 U4048 ( .A(REG0_REG_3__SCAN_IN), .ZN(n3436) );
  OAI22_X1 U4049 ( .A1(n4459), .A2(n4819), .B1(n4879), .B2(n3436), .ZN(n3437)
         );
  AOI21_X1 U4050 ( .B1(n3438), .B2(n4879), .A(n3437), .ZN(n3439) );
  INV_X1 U4051 ( .A(n3439), .ZN(U3473) );
  INV_X1 U4052 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3440) );
  OAI22_X1 U4053 ( .A1(n4459), .A2(n4813), .B1(n4879), .B2(n3440), .ZN(n3441)
         );
  AOI21_X1 U4054 ( .B1(n3442), .B2(n4879), .A(n3441), .ZN(n3443) );
  INV_X1 U4055 ( .A(n3443), .ZN(U3471) );
  INV_X1 U4056 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U4057 ( .A1(n3444), .A2(n4879), .ZN(n3446) );
  INV_X1 U4058 ( .A(n4459), .ZN(n3613) );
  NAND2_X1 U4059 ( .A1(n4835), .A2(n3613), .ZN(n3445) );
  OAI211_X1 U4060 ( .C1(n4879), .C2(n3447), .A(n3446), .B(n3445), .ZN(U3479)
         );
  NAND2_X1 U4061 ( .A1(n3117), .A2(n3832), .ZN(n3933) );
  XOR2_X1 U4062 ( .A(n3448), .B(n3933), .Z(n3470) );
  INV_X1 U4063 ( .A(n3470), .ZN(n3460) );
  XOR2_X1 U4064 ( .A(n3933), .B(n3449), .Z(n3453) );
  OAI22_X1 U4065 ( .A1(n3450), .A2(n4857), .B1(n3454), .B2(n4855), .ZN(n3451)
         );
  AOI21_X1 U4066 ( .B1(n4861), .B2(n3979), .A(n3451), .ZN(n3452) );
  OAI21_X1 U4067 ( .B1(n3453), .B2(n4863), .A(n3452), .ZN(n3469) );
  INV_X1 U4068 ( .A(n3489), .ZN(n3455) );
  OAI21_X1 U4069 ( .B1(n3455), .B2(n3454), .A(n3531), .ZN(n3475) );
  NOR2_X1 U4070 ( .A1(n3475), .A2(n4905), .ZN(n3458) );
  OAI22_X1 U4071 ( .A1(n3512), .A2(n4909), .B1(n3456), .B2(n4849), .ZN(n3457)
         );
  AOI211_X1 U4072 ( .C1(n3469), .C2(n4849), .A(n3458), .B(n3457), .ZN(n3459)
         );
  OAI21_X1 U4073 ( .B1(n4278), .B2(n3460), .A(n3459), .ZN(U3281) );
  XOR2_X1 U4074 ( .A(n3461), .B(n3462), .Z(n3467) );
  AOI22_X1 U4075 ( .A1(n3463), .A2(n4920), .B1(n4922), .B2(n3982), .ZN(n3465)
         );
  NOR2_X1 U4076 ( .A1(STATE_REG_SCAN_IN), .A2(n2600), .ZN(n4707) );
  AOI21_X1 U4077 ( .B1(n4924), .B2(n4860), .A(n4707), .ZN(n3464) );
  OAI211_X1 U4078 ( .C1(n4938), .C2(n4867), .A(n3465), .B(n3464), .ZN(n3466)
         );
  AOI21_X1 U4079 ( .B1(n3467), .B2(n4933), .A(n3466), .ZN(n3468) );
  INV_X1 U4080 ( .A(n3468), .ZN(U3210) );
  INV_X1 U4081 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3471) );
  AOI21_X1 U4082 ( .B1(n3470), .B2(n4871), .A(n3469), .ZN(n3473) );
  MUX2_X1 U4083 ( .A(n3471), .B(n3473), .S(n4879), .Z(n3472) );
  OAI21_X1 U4084 ( .B1(n3475), .B2(n4459), .A(n3472), .ZN(U3485) );
  MUX2_X1 U4085 ( .A(n4715), .B(n3473), .S(n4875), .Z(n3474) );
  OAI21_X1 U4086 ( .B1(n4406), .B2(n3475), .A(n3474), .ZN(U3527) );
  INV_X1 U4087 ( .A(n3477), .ZN(n3479) );
  NAND2_X1 U4088 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  XNOR2_X1 U4089 ( .A(n3476), .B(n3480), .ZN(n3487) );
  INV_X1 U4090 ( .A(n4880), .ZN(n3485) );
  AOI22_X1 U4091 ( .A1(n3481), .A2(n4920), .B1(n4924), .B2(n3980), .ZN(n3484)
         );
  AOI21_X1 U4092 ( .B1(n4922), .B2(n3981), .A(n3482), .ZN(n3483) );
  OAI211_X1 U4093 ( .C1(n4938), .C2(n3485), .A(n3484), .B(n3483), .ZN(n3486)
         );
  AOI21_X1 U4094 ( .B1(n3487), .B2(n4933), .A(n3486), .ZN(n3488) );
  INV_X1 U4095 ( .A(n3488), .ZN(U3218) );
  OAI21_X1 U4096 ( .B1(n4843), .B2(n3494), .A(n3489), .ZN(n4881) );
  INV_X1 U4097 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3501) );
  INV_X1 U4098 ( .A(n4804), .ZN(n4828) );
  NAND2_X1 U4099 ( .A1(n3831), .A2(n3837), .ZN(n3932) );
  NAND2_X1 U4100 ( .A1(n3490), .A2(n3491), .ZN(n3492) );
  XOR2_X1 U4101 ( .A(n3932), .B(n3492), .Z(n4883) );
  XOR2_X1 U4102 ( .A(n3493), .B(n3932), .Z(n3498) );
  OAI22_X1 U4103 ( .A1(n3495), .A2(n4794), .B1(n4855), .B2(n3494), .ZN(n3496)
         );
  AOI21_X1 U4104 ( .B1(n4267), .B2(n3981), .A(n3496), .ZN(n3497) );
  OAI21_X1 U4105 ( .B1(n3498), .B2(n4863), .A(n3497), .ZN(n3499) );
  AOI21_X1 U4106 ( .B1(n4883), .B2(n4792), .A(n3499), .ZN(n4886) );
  INV_X1 U4107 ( .A(n4886), .ZN(n3500) );
  AOI21_X1 U4108 ( .B1(n4828), .B2(n4883), .A(n3500), .ZN(n3503) );
  MUX2_X1 U4109 ( .A(n3501), .B(n3503), .S(n4879), .Z(n3502) );
  OAI21_X1 U4110 ( .B1(n4881), .B2(n4459), .A(n3502), .ZN(U3483) );
  MUX2_X1 U4111 ( .A(n3504), .B(n3503), .S(n4875), .Z(n3505) );
  OAI21_X1 U4112 ( .B1(n4881), .B2(n4406), .A(n3505), .ZN(U3526) );
  OAI21_X1 U4113 ( .B1(n3508), .B2(n3507), .A(n3506), .ZN(n3514) );
  AOI22_X1 U4114 ( .A1(n3509), .A2(n3792), .B1(n4922), .B2(n4860), .ZN(n3511)
         );
  NOR2_X1 U4115 ( .A1(STATE_REG_SCAN_IN), .A2(n2629), .ZN(n4720) );
  AOI21_X1 U4116 ( .B1(n3806), .B2(n3979), .A(n4720), .ZN(n3510) );
  OAI211_X1 U4117 ( .C1(n4938), .C2(n3512), .A(n3511), .B(n3510), .ZN(n3513)
         );
  AOI21_X1 U4118 ( .B1(n3514), .B2(n4933), .A(n3513), .ZN(n3515) );
  INV_X1 U4119 ( .A(n3515), .ZN(U3228) );
  OAI22_X1 U4120 ( .A1(n3536), .A2(n4857), .B1(n4855), .B2(n3522), .ZN(n3521)
         );
  INV_X1 U4121 ( .A(n3516), .ZN(n3517) );
  AOI21_X1 U4122 ( .B1(n3603), .B2(n3518), .A(n3517), .ZN(n4306) );
  AND2_X1 U4123 ( .A1(n4305), .A2(n4303), .ZN(n3913) );
  XNOR2_X1 U4124 ( .A(n4306), .B(n3913), .ZN(n3519) );
  NOR2_X1 U4125 ( .A1(n3519), .A2(n4863), .ZN(n3520) );
  AOI211_X1 U4126 ( .C1(n4861), .C2(n3976), .A(n3521), .B(n3520), .ZN(n4402)
         );
  OAI21_X1 U4127 ( .B1(n3598), .B2(n3522), .A(n4319), .ZN(n4460) );
  INV_X1 U4128 ( .A(n4460), .ZN(n3525) );
  INV_X1 U4129 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3523) );
  OAI22_X1 U4130 ( .A1(n4849), .A2(n3523), .B1(n3626), .B2(n4909), .ZN(n3524)
         );
  AOI21_X1 U4131 ( .B1(n3525), .B2(n4940), .A(n3524), .ZN(n3530) );
  NAND2_X1 U4132 ( .A1(n3526), .A2(n3527), .ZN(n3528) );
  XOR2_X1 U4133 ( .A(n3913), .B(n3528), .Z(n4404) );
  NAND2_X1 U4134 ( .A1(n4404), .A2(n4290), .ZN(n3529) );
  OAI211_X1 U4135 ( .C1(n4402), .C2(n4944), .A(n3530), .B(n3529), .ZN(U3278)
         );
  INV_X1 U4136 ( .A(n3531), .ZN(n3532) );
  OAI21_X1 U4137 ( .B1(n3532), .B2(n3535), .A(n3599), .ZN(n4893) );
  INV_X1 U4138 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3542) );
  NAND2_X1 U4139 ( .A1(n3850), .A2(n3848), .ZN(n3925) );
  XNOR2_X1 U4140 ( .A(n3533), .B(n3925), .ZN(n4896) );
  XNOR2_X1 U4141 ( .A(n3534), .B(n3925), .ZN(n3539) );
  OAI22_X1 U4142 ( .A1(n3536), .A2(n4794), .B1(n4855), .B2(n3535), .ZN(n3537)
         );
  AOI21_X1 U4143 ( .B1(n4267), .B2(n3980), .A(n3537), .ZN(n3538) );
  OAI21_X1 U4144 ( .B1(n3539), .B2(n4863), .A(n3538), .ZN(n3540) );
  AOI21_X1 U4145 ( .B1(n4792), .B2(n4896), .A(n3540), .ZN(n4899) );
  INV_X1 U4146 ( .A(n4899), .ZN(n3541) );
  AOI21_X1 U4147 ( .B1(n4828), .B2(n4896), .A(n3541), .ZN(n3544) );
  MUX2_X1 U4148 ( .A(n3542), .B(n3544), .S(n4875), .Z(n3543) );
  OAI21_X1 U4149 ( .B1(n4893), .B2(n4406), .A(n3543), .ZN(U3528) );
  INV_X1 U4150 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3545) );
  MUX2_X1 U4151 ( .A(n3545), .B(n3544), .S(n4879), .Z(n3546) );
  OAI21_X1 U4152 ( .B1(n4893), .B2(n4459), .A(n3546), .ZN(U3487) );
  AND2_X1 U4153 ( .A1(n3548), .A2(n3547), .ZN(n3549) );
  NAND2_X1 U4154 ( .A1(n3549), .A2(n3924), .ZN(n4287) );
  OAI21_X1 U4155 ( .B1(n3549), .B2(n3924), .A(n4287), .ZN(n4395) );
  INV_X1 U4156 ( .A(n4395), .ZN(n3561) );
  OAI21_X1 U4157 ( .B1(n3550), .B2(n3885), .A(n4281), .ZN(n3551) );
  NAND2_X1 U4158 ( .A1(n3551), .A2(n4791), .ZN(n3553) );
  AOI22_X1 U4159 ( .A1(n3976), .A2(n4267), .B1(n4331), .B2(n3655), .ZN(n3552)
         );
  OAI211_X1 U4160 ( .C1(n3554), .C2(n4794), .A(n3553), .B(n3552), .ZN(n4394)
         );
  INV_X1 U4161 ( .A(n4321), .ZN(n3557) );
  INV_X1 U4162 ( .A(n4293), .ZN(n3555) );
  OAI21_X1 U4163 ( .B1(n3557), .B2(n3556), .A(n3555), .ZN(n4451) );
  INV_X1 U4164 ( .A(n4909), .ZN(n4891) );
  AOI22_X1 U4165 ( .A1(n4944), .A2(REG2_REG_14__SCAN_IN), .B1(n3654), .B2(
        n4891), .ZN(n3558) );
  OAI21_X1 U4166 ( .B1(n4451), .B2(n4905), .A(n3558), .ZN(n3559) );
  AOI21_X1 U4167 ( .B1(n4394), .B2(n4849), .A(n3559), .ZN(n3560) );
  OAI21_X1 U4168 ( .B1(n3561), .B2(n4278), .A(n3560), .ZN(U3276) );
  INV_X1 U4169 ( .A(n3563), .ZN(n3565) );
  NAND2_X1 U4170 ( .A1(n3565), .A2(n3564), .ZN(n3566) );
  XNOR2_X1 U4171 ( .A(n3562), .B(n3566), .ZN(n3570) );
  AOI22_X1 U4172 ( .A1(n3600), .A2(n3792), .B1(n4922), .B2(n3979), .ZN(n3568)
         );
  AND2_X1 U4173 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4741) );
  AOI21_X1 U4174 ( .B1(n3806), .B2(n3977), .A(n4741), .ZN(n3567) );
  OAI211_X1 U4175 ( .C1(n4938), .C2(n4910), .A(n3568), .B(n3567), .ZN(n3569)
         );
  AOI21_X1 U4176 ( .B1(n3570), .B2(n4933), .A(n3569), .ZN(n3571) );
  INV_X1 U4177 ( .A(n3571), .ZN(U3233) );
  OAI21_X1 U4178 ( .B1(n3573), .B2(n3574), .A(n3572), .ZN(n4388) );
  XNOR2_X1 U4179 ( .A(n3575), .B(n3574), .ZN(n3579) );
  NOR2_X1 U4180 ( .A1(n3582), .A2(n4855), .ZN(n3576) );
  AOI21_X1 U4181 ( .B1(n3975), .B2(n4267), .A(n3576), .ZN(n3577) );
  OAI21_X1 U4182 ( .B1(n4247), .B2(n4794), .A(n3577), .ZN(n3578) );
  AOI21_X1 U4183 ( .B1(n3579), .B2(n4791), .A(n3578), .ZN(n4386) );
  INV_X1 U4184 ( .A(n3580), .ZN(n3731) );
  OAI22_X1 U4185 ( .A1(n4849), .A2(n4775), .B1(n3731), .B2(n4909), .ZN(n3581)
         );
  INV_X1 U4186 ( .A(n3581), .ZN(n3584) );
  OR2_X1 U4187 ( .A1(n4291), .A2(n3582), .ZN(n4384) );
  NAND3_X1 U4188 ( .A1(n4384), .A2(n4383), .A3(n4940), .ZN(n3583) );
  OAI211_X1 U4189 ( .C1(n4386), .C2(n4944), .A(n3584), .B(n3583), .ZN(n3585)
         );
  INV_X1 U4190 ( .A(n3585), .ZN(n3586) );
  OAI21_X1 U4191 ( .B1(n4388), .B2(n4278), .A(n3586), .ZN(U3274) );
  AOI211_X1 U4192 ( .C1(n3589), .C2(n3588), .A(n3587), .B(n4774), .ZN(n3593)
         );
  AND2_X1 U4193 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n3656) );
  AOI21_X1 U4194 ( .B1(n4779), .B2(ADDR_REG_14__SCAN_IN), .A(n3656), .ZN(n3590) );
  OAI21_X1 U4195 ( .B1(n4785), .B2(n3591), .A(n3590), .ZN(n3592) );
  NOR2_X1 U4196 ( .A1(n3593), .A2(n3592), .ZN(n3597) );
  OAI211_X1 U4197 ( .C1(n3595), .C2(REG1_REG_14__SCAN_IN), .A(n4780), .B(n3594), .ZN(n3596) );
  NAND2_X1 U4198 ( .A1(n3597), .A2(n3596), .ZN(U3254) );
  AOI21_X1 U4199 ( .B1(n3600), .B2(n3599), .A(n3598), .ZN(n4903) );
  NAND2_X1 U4200 ( .A1(n3601), .A2(n3930), .ZN(n3602) );
  NAND2_X1 U4201 ( .A1(n3526), .A2(n3602), .ZN(n4902) );
  NAND2_X1 U4202 ( .A1(n4902), .A2(n4792), .ZN(n3610) );
  XNOR2_X1 U4203 ( .A(n3603), .B(n3930), .ZN(n3608) );
  NAND2_X1 U4204 ( .A1(n3979), .A2(n4267), .ZN(n3605) );
  NAND2_X1 U4205 ( .A1(n3977), .A2(n4861), .ZN(n3604) );
  OAI211_X1 U4206 ( .C1(n4855), .C2(n3606), .A(n3605), .B(n3604), .ZN(n3607)
         );
  AOI21_X1 U4207 ( .B1(n3608), .B2(n4791), .A(n3607), .ZN(n3609) );
  AND2_X1 U4208 ( .A1(n3610), .A2(n3609), .ZN(n4914) );
  NAND2_X1 U4209 ( .A1(n4902), .A2(n4828), .ZN(n3611) );
  NAND2_X1 U4210 ( .A1(n4914), .A2(n3611), .ZN(n3615) );
  MUX2_X1 U4211 ( .A(REG0_REG_11__SCAN_IN), .B(n3615), .S(n4879), .Z(n3612) );
  AOI21_X1 U4212 ( .B1(n4903), .B2(n3613), .A(n3612), .ZN(n3614) );
  INV_X1 U4213 ( .A(n3614), .ZN(U3489) );
  MUX2_X1 U4214 ( .A(REG1_REG_11__SCAN_IN), .B(n3615), .S(n4875), .Z(n3616) );
  AOI21_X1 U4215 ( .B1(n3617), .B2(n4903), .A(n3616), .ZN(n3618) );
  INV_X1 U4216 ( .A(n3618), .ZN(U3529) );
  XNOR2_X1 U4217 ( .A(n3621), .B(n3620), .ZN(n3622) );
  XNOR2_X1 U4218 ( .A(n3619), .B(n3622), .ZN(n3628) );
  AOI22_X1 U4219 ( .A1(n3623), .A2(n4920), .B1(n3806), .B2(n3976), .ZN(n3625)
         );
  INV_X1 U4220 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4642) );
  NOR2_X1 U4221 ( .A1(STATE_REG_SCAN_IN), .A2(n4642), .ZN(n4751) );
  AOI21_X1 U4222 ( .B1(n4922), .B2(n3978), .A(n4751), .ZN(n3624) );
  OAI211_X1 U4223 ( .C1(n4938), .C2(n3626), .A(n3625), .B(n3624), .ZN(n3627)
         );
  AOI21_X1 U4224 ( .B1(n3628), .B2(n4933), .A(n3627), .ZN(n3629) );
  INV_X1 U4225 ( .A(n3629), .ZN(U3221) );
  NAND3_X1 U4226 ( .A1(n3630), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3632) );
  INV_X1 U4227 ( .A(DATAI_31_), .ZN(n3631) );
  OAI22_X1 U4228 ( .A1(n2457), .A2(n3632), .B1(STATE_REG_SCAN_IN), .B2(n3631), 
        .ZN(U3321) );
  NOR2_X1 U4229 ( .A1(n3634), .A2(n3631), .ZN(n3904) );
  NOR2_X1 U4230 ( .A1(n3634), .A2(n3633), .ZN(n4332) );
  XOR2_X2 U4231 ( .A(n3904), .B(n4327), .Z(n3649) );
  INV_X1 U4232 ( .A(n3904), .ZN(n3641) );
  NAND2_X1 U4233 ( .A1(n3102), .A2(REG1_REG_31__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4234 ( .A1(n3635), .A2(REG2_REG_31__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4235 ( .A1(n2497), .A2(REG0_REG_31__SCAN_IN), .ZN(n3636) );
  AND3_X1 U4236 ( .A1(n3638), .A2(n3637), .A3(n3636), .ZN(n4681) );
  INV_X1 U4237 ( .A(n4681), .ZN(n3640) );
  NAND2_X1 U4238 ( .A1(n3640), .A2(n3639), .ZN(n4329) );
  OAI21_X1 U4239 ( .B1(n3641), .B2(n4855), .A(n4329), .ZN(n3646) );
  NAND2_X1 U4240 ( .A1(n4879), .A2(n3646), .ZN(n3643) );
  NAND2_X1 U4241 ( .A1(n4876), .A2(REG0_REG_31__SCAN_IN), .ZN(n3642) );
  OAI211_X1 U4242 ( .C1(n3649), .C2(n4459), .A(n3643), .B(n3642), .ZN(U3517)
         );
  NAND2_X1 U4243 ( .A1(n4875), .A2(n3646), .ZN(n3645) );
  NAND2_X1 U4244 ( .A1(n4873), .A2(REG1_REG_31__SCAN_IN), .ZN(n3644) );
  OAI211_X1 U4245 ( .C1(n3649), .C2(n4406), .A(n3645), .B(n3644), .ZN(U3549)
         );
  NAND2_X1 U4246 ( .A1(n4849), .A2(n3646), .ZN(n3648) );
  NAND2_X1 U4247 ( .A1(n4944), .A2(REG2_REG_31__SCAN_IN), .ZN(n3647) );
  OAI211_X1 U4248 ( .C1(n3649), .C2(n4905), .A(n3648), .B(n3647), .ZN(U3260)
         );
  NAND2_X1 U4249 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3650) );
  OAI21_X1 U4250 ( .B1(n2908), .B2(U3149), .A(n3650), .ZN(U3327) );
  XNOR2_X1 U4251 ( .A(n3652), .B(n3651), .ZN(n3653) );
  XNOR2_X1 U4252 ( .A(n2280), .B(n3653), .ZN(n3661) );
  INV_X1 U4253 ( .A(n3654), .ZN(n3659) );
  AOI22_X1 U4254 ( .A1(n3655), .A2(n4920), .B1(n3806), .B2(n3975), .ZN(n3658)
         );
  AOI21_X1 U4255 ( .B1(n4922), .B2(n3976), .A(n3656), .ZN(n3657) );
  OAI211_X1 U4256 ( .C1(n4938), .C2(n3659), .A(n3658), .B(n3657), .ZN(n3660)
         );
  AOI21_X1 U4257 ( .B1(n3661), .B2(n4933), .A(n3660), .ZN(n3662) );
  INV_X1 U4258 ( .A(n3662), .ZN(U3212) );
  INV_X1 U4259 ( .A(n3663), .ZN(n3777) );
  OAI21_X1 U4260 ( .B1(n3777), .B2(n3665), .A(n3664), .ZN(n3667) );
  NAND3_X1 U4261 ( .A1(n3667), .A2(n4933), .A3(n3666), .ZN(n3672) );
  AOI22_X1 U4262 ( .A1(n4922), .A2(n4187), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3671) );
  AOI22_X1 U4263 ( .A1(n4155), .A2(n4920), .B1(n4924), .B2(n4151), .ZN(n3670)
         );
  INV_X1 U4264 ( .A(n4158), .ZN(n3668) );
  OR2_X1 U4265 ( .A1(n4938), .A2(n3668), .ZN(n3669) );
  NAND4_X1 U4266 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(U3213)
         );
  AND2_X1 U4267 ( .A1(n3506), .A2(n3673), .ZN(n3676) );
  OAI211_X1 U4268 ( .C1(n3676), .C2(n3675), .A(n4933), .B(n3674), .ZN(n3682)
         );
  NOR2_X1 U4269 ( .A1(STATE_REG_SCAN_IN), .A2(n4528), .ZN(n4734) );
  AOI21_X1 U4270 ( .B1(n4924), .B2(n3978), .A(n4734), .ZN(n3681) );
  AOI22_X1 U4271 ( .A1(n3677), .A2(n4920), .B1(n4922), .B2(n3980), .ZN(n3680)
         );
  INV_X1 U4272 ( .A(n4892), .ZN(n3678) );
  OR2_X1 U4273 ( .A1(n4938), .A2(n3678), .ZN(n3679) );
  NAND4_X1 U4274 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(U3214)
         );
  INV_X1 U4275 ( .A(n3684), .ZN(n3685) );
  AOI21_X1 U4276 ( .B1(n3683), .B2(n3686), .A(n3685), .ZN(n3695) );
  OAI22_X1 U4277 ( .A1(n4233), .A2(n3688), .B1(n3687), .B2(n4270), .ZN(n3689)
         );
  AOI211_X1 U4278 ( .C1(n3806), .C2(n3972), .A(n3690), .B(n3689), .ZN(n3694)
         );
  INV_X1 U4279 ( .A(n4938), .ZN(n3692) );
  NAND2_X1 U4280 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  OAI211_X1 U4281 ( .C1(n3695), .C2(n3785), .A(n3694), .B(n3693), .ZN(U3216)
         );
  INV_X1 U4282 ( .A(n3757), .ZN(n3697) );
  OAI21_X1 U4283 ( .B1(n3696), .B2(n3697), .A(n3758), .ZN(n3701) );
  XNOR2_X1 U4284 ( .A(n3699), .B(n3698), .ZN(n3700) );
  XNOR2_X1 U4285 ( .A(n3701), .B(n3700), .ZN(n3707) );
  INV_X1 U4286 ( .A(n3702), .ZN(n4194) );
  AOI22_X1 U4287 ( .A1(n3703), .A2(n4920), .B1(n4922), .B2(n3972), .ZN(n3705)
         );
  AOI22_X1 U4288 ( .A1(n4924), .A2(n4187), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3704) );
  OAI211_X1 U4289 ( .C1(n4938), .C2(n4194), .A(n3705), .B(n3704), .ZN(n3706)
         );
  AOI21_X1 U4290 ( .B1(n3707), .B2(n4933), .A(n3706), .ZN(n3708) );
  INV_X1 U4291 ( .A(n3708), .ZN(U3220) );
  XOR2_X1 U4292 ( .A(n3711), .B(n3710), .Z(n3712) );
  XNOR2_X1 U4293 ( .A(n3709), .B(n3712), .ZN(n3718) );
  INV_X1 U4294 ( .A(n4111), .ZN(n3716) );
  AOI22_X1 U4295 ( .A1(n3713), .A2(n4920), .B1(n4922), .B2(n4151), .ZN(n3715)
         );
  AOI22_X1 U4296 ( .A1(n4924), .A2(n4104), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3714) );
  OAI211_X1 U4297 ( .C1(n4938), .C2(n3716), .A(n3715), .B(n3714), .ZN(n3717)
         );
  AOI21_X1 U4298 ( .B1(n3718), .B2(n4933), .A(n3717), .ZN(n3719) );
  INV_X1 U4299 ( .A(n3719), .ZN(U3222) );
  INV_X1 U4300 ( .A(n4930), .ZN(n3721) );
  NOR2_X1 U4301 ( .A1(n3720), .A2(n3721), .ZN(n3723) );
  INV_X1 U4302 ( .A(n3720), .ZN(n3722) );
  OAI22_X1 U4303 ( .A1(n3723), .A2(n4931), .B1(n3722), .B2(n4930), .ZN(n3727)
         );
  NAND2_X1 U4304 ( .A1(n3725), .A2(n3724), .ZN(n3726) );
  XNOR2_X1 U4305 ( .A(n3727), .B(n3726), .ZN(n3733) );
  AOI22_X1 U4306 ( .A1(n3728), .A2(n3792), .B1(n3806), .B2(n3974), .ZN(n3730)
         );
  NOR2_X1 U4307 ( .A1(STATE_REG_SCAN_IN), .A2(n4539), .ZN(n4778) );
  AOI21_X1 U4308 ( .B1(n4922), .B2(n3975), .A(n4778), .ZN(n3729) );
  OAI211_X1 U4309 ( .C1(n4938), .C2(n3731), .A(n3730), .B(n3729), .ZN(n3732)
         );
  AOI21_X1 U4310 ( .B1(n3733), .B2(n4933), .A(n3732), .ZN(n3734) );
  INV_X1 U4311 ( .A(n3734), .ZN(U3223) );
  NAND2_X1 U4312 ( .A1(n3736), .A2(n3735), .ZN(n3738) );
  XOR2_X1 U4313 ( .A(n3738), .B(n3737), .Z(n3743) );
  AOI22_X1 U4314 ( .A1(n4271), .A2(n3792), .B1(n4924), .B2(n3973), .ZN(n3740)
         );
  INV_X1 U4315 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4569) );
  NOR2_X1 U4316 ( .A1(STATE_REG_SCAN_IN), .A2(n4569), .ZN(n4018) );
  AOI21_X1 U4317 ( .B1(n4922), .B2(n4923), .A(n4018), .ZN(n3739) );
  OAI211_X1 U4318 ( .C1(n4938), .C2(n3741), .A(n3740), .B(n3739), .ZN(n3742)
         );
  AOI21_X1 U4319 ( .B1(n3743), .B2(n4933), .A(n3742), .ZN(n3744) );
  INV_X1 U4320 ( .A(n3744), .ZN(U3225) );
  AND2_X1 U4321 ( .A1(n3746), .A2(n3745), .ZN(n3748) );
  NAND2_X1 U4322 ( .A1(n3748), .A2(n3747), .ZN(n3749) );
  XOR2_X1 U4323 ( .A(n3750), .B(n3749), .Z(n3755) );
  INV_X1 U4324 ( .A(n4131), .ZN(n3753) );
  AOI22_X1 U4325 ( .A1(n4128), .A2(n3792), .B1(n4922), .B2(n4125), .ZN(n3752)
         );
  AOI22_X1 U4326 ( .A1(n4924), .A2(n3971), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3751) );
  OAI211_X1 U4327 ( .C1(n4938), .C2(n3753), .A(n3752), .B(n3751), .ZN(n3754)
         );
  AOI21_X1 U4328 ( .B1(n3755), .B2(n4933), .A(n3754), .ZN(n3756) );
  INV_X1 U4329 ( .A(n3756), .ZN(U3226) );
  NAND2_X1 U4330 ( .A1(n3758), .A2(n3757), .ZN(n3759) );
  XOR2_X1 U4331 ( .A(n3759), .B(n3696), .Z(n3764) );
  INV_X1 U4332 ( .A(n3760), .ZN(n4213) );
  AOI22_X1 U4333 ( .A1(n4212), .A2(n3792), .B1(n4922), .B2(n4245), .ZN(n3762)
         );
  AOI22_X1 U4334 ( .A1(n4924), .A2(n4204), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3761) );
  OAI211_X1 U4335 ( .C1(n4938), .C2(n4213), .A(n3762), .B(n3761), .ZN(n3763)
         );
  AOI21_X1 U4336 ( .B1(n3764), .B2(n4933), .A(n3763), .ZN(n3765) );
  INV_X1 U4337 ( .A(n3765), .ZN(U3230) );
  NOR2_X1 U4338 ( .A1(n2396), .A2(n3769), .ZN(n3770) );
  XNOR2_X1 U4339 ( .A(n3767), .B(n3770), .ZN(n3775) );
  AOI22_X1 U4340 ( .A1(n4318), .A2(n3792), .B1(n3806), .B2(n4921), .ZN(n3772)
         );
  INV_X1 U4341 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4553) );
  NOR2_X1 U4342 ( .A1(STATE_REG_SCAN_IN), .A2(n4553), .ZN(n4770) );
  AOI21_X1 U4343 ( .B1(n4922), .B2(n3977), .A(n4770), .ZN(n3771) );
  OAI211_X1 U4344 ( .C1(n4938), .C2(n3773), .A(n3772), .B(n3771), .ZN(n3774)
         );
  AOI21_X1 U4345 ( .B1(n3775), .B2(n4933), .A(n3774), .ZN(n3776) );
  INV_X1 U4346 ( .A(n3776), .ZN(U3231) );
  AOI21_X1 U4347 ( .B1(n3778), .B2(n2283), .A(n3777), .ZN(n3786) );
  INV_X1 U4348 ( .A(n3779), .ZN(n4174) );
  AOI22_X1 U4349 ( .A1(n3780), .A2(n4920), .B1(n4924), .B2(n4125), .ZN(n3782)
         );
  AOI22_X1 U4350 ( .A1(n4922), .A2(n4204), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3781) );
  OAI211_X1 U4351 ( .C1(n4938), .C2(n4174), .A(n3782), .B(n3781), .ZN(n3783)
         );
  INV_X1 U4352 ( .A(n3783), .ZN(n3784) );
  OAI21_X1 U4353 ( .B1(n3786), .B2(n3785), .A(n3784), .ZN(U3232) );
  XOR2_X1 U4354 ( .A(n3789), .B(n3788), .Z(n3790) );
  XNOR2_X1 U4355 ( .A(n3787), .B(n3790), .ZN(n3797) );
  INV_X1 U4356 ( .A(n3791), .ZN(n4250) );
  AOI22_X1 U4357 ( .A1(n4244), .A2(n3792), .B1(n4922), .B2(n3974), .ZN(n3795)
         );
  NOR2_X1 U4358 ( .A1(STATE_REG_SCAN_IN), .A2(n3793), .ZN(n4031) );
  AOI21_X1 U4359 ( .B1(n3806), .B2(n4245), .A(n4031), .ZN(n3794) );
  OAI211_X1 U4360 ( .C1(n4938), .C2(n4250), .A(n3795), .B(n3794), .ZN(n3796)
         );
  AOI21_X1 U4361 ( .B1(n3797), .B2(n4933), .A(n3796), .ZN(n3798) );
  INV_X1 U4362 ( .A(n3798), .ZN(U3235) );
  NAND2_X1 U4363 ( .A1(n2898), .A2(n3800), .ZN(n3801) );
  XNOR2_X1 U4364 ( .A(n3802), .B(n3801), .ZN(n3810) );
  INV_X1 U4365 ( .A(n3803), .ZN(n4091) );
  AOI22_X1 U4366 ( .A1(n4090), .A2(n4920), .B1(n4922), .B2(n3971), .ZN(n3808)
         );
  NOR2_X1 U4367 ( .A1(n3804), .A2(STATE_REG_SCAN_IN), .ZN(n3805) );
  AOI21_X1 U4368 ( .B1(n3806), .B2(n3970), .A(n3805), .ZN(n3807) );
  OAI211_X1 U4369 ( .C1(n4938), .C2(n4091), .A(n3808), .B(n3807), .ZN(n3809)
         );
  AOI21_X1 U4370 ( .B1(n3810), .B2(n4933), .A(n3809), .ZN(n3811) );
  INV_X1 U4371 ( .A(n3811), .ZN(U3237) );
  INV_X1 U4372 ( .A(n3968), .ZN(n3812) );
  NOR2_X1 U4373 ( .A1(n3812), .A2(n4332), .ZN(n3902) );
  AOI21_X1 U4374 ( .B1(n3904), .B2(n4681), .A(n3902), .ZN(n3915) );
  NAND2_X1 U4375 ( .A1(n3987), .A2(n4790), .ZN(n3942) );
  OAI211_X1 U4376 ( .C1(n3815), .C2(n3814), .A(n3942), .B(n3813), .ZN(n3818)
         );
  NAND3_X1 U4377 ( .A1(n3818), .A2(n3817), .A3(n3816), .ZN(n3821) );
  NAND3_X1 U4378 ( .A1(n3821), .A2(n3820), .A3(n3819), .ZN(n3824) );
  NAND3_X1 U4379 ( .A1(n3824), .A2(n3823), .A3(n3822), .ZN(n3827) );
  AND4_X1 U4380 ( .A1(n3827), .A2(n3826), .A3(n3839), .A4(n3825), .ZN(n3830)
         );
  INV_X1 U4381 ( .A(n3828), .ZN(n3829) );
  OAI211_X1 U4382 ( .C1(n3830), .C2(n3829), .A(n3838), .B(n3837), .ZN(n3833)
         );
  NAND3_X1 U4383 ( .A1(n3833), .A2(n3832), .A3(n3831), .ZN(n3847) );
  NAND2_X1 U4384 ( .A1(n3835), .A2(n3834), .ZN(n3844) );
  NOR2_X1 U4385 ( .A1(n3844), .A2(n3836), .ZN(n3846) );
  NAND2_X1 U4386 ( .A1(n3117), .A2(n3837), .ZN(n3843) );
  INV_X1 U4387 ( .A(n3838), .ZN(n3842) );
  INV_X1 U4388 ( .A(n3839), .ZN(n3841) );
  NOR4_X1 U4389 ( .A1(n3843), .A2(n3842), .A3(n3841), .A4(n3840), .ZN(n3845)
         );
  NAND2_X1 U4390 ( .A1(n3844), .A2(n3851), .ZN(n3882) );
  AOI22_X1 U4391 ( .A1(n3847), .A2(n3846), .B1(n3845), .B2(n3882), .ZN(n3859)
         );
  AND2_X1 U4392 ( .A1(n3849), .A2(n3848), .ZN(n3854) );
  INV_X1 U4393 ( .A(n3854), .ZN(n3858) );
  INV_X1 U4394 ( .A(n3882), .ZN(n3857) );
  INV_X1 U4395 ( .A(n3850), .ZN(n3855) );
  NAND2_X1 U4396 ( .A1(n4280), .A2(n3851), .ZN(n3884) );
  INV_X1 U4397 ( .A(n3852), .ZN(n3853) );
  AOI211_X1 U4398 ( .C1(n3855), .C2(n3854), .A(n3884), .B(n3853), .ZN(n3856)
         );
  OAI22_X1 U4399 ( .A1(n3859), .A2(n3858), .B1(n3857), .B2(n3856), .ZN(n3861)
         );
  OAI211_X1 U4400 ( .C1(n3886), .C2(n3861), .A(n3883), .B(n3860), .ZN(n3862)
         );
  OAI221_X1 U4401 ( .B1(n4141), .B2(n3890), .C1(n4141), .C2(n3862), .A(n3894), 
        .ZN(n3863) );
  AOI21_X1 U4402 ( .B1(n3864), .B2(n3863), .A(n3896), .ZN(n3867) );
  INV_X1 U4403 ( .A(n3880), .ZN(n3865) );
  OAI21_X1 U4404 ( .B1(n3867), .B2(n3866), .A(n3865), .ZN(n3868) );
  NAND4_X1 U4405 ( .A1(n3915), .A2(n3869), .A3(n3940), .A4(n3868), .ZN(n3877)
         );
  NAND2_X1 U4406 ( .A1(n4054), .A2(n3874), .ZN(n3870) );
  AND2_X1 U4407 ( .A1(n3871), .A2(n3870), .ZN(n3878) );
  INV_X1 U4408 ( .A(n3878), .ZN(n3876) );
  NOR2_X1 U4409 ( .A1(n4681), .A2(n3904), .ZN(n3873) );
  NOR2_X1 U4410 ( .A1(n3915), .A2(n3873), .ZN(n3875) );
  INV_X1 U4411 ( .A(n4332), .ZN(n3903) );
  NOR2_X1 U4412 ( .A1(n3968), .A2(n3903), .ZN(n3872) );
  NOR2_X1 U4413 ( .A1(n3873), .A2(n3872), .ZN(n3914) );
  OAI21_X1 U4414 ( .B1(n4054), .B2(n3874), .A(n3914), .ZN(n3879) );
  AOI21_X1 U4415 ( .B1(n3878), .B2(n3881), .A(n3879), .ZN(n3901) );
  OAI22_X1 U4416 ( .A1(n3877), .A2(n3876), .B1(n3875), .B2(n3901), .ZN(n3957)
         );
  NAND3_X1 U4417 ( .A1(n4069), .A2(n3878), .A3(n3940), .ZN(n3900) );
  NOR3_X1 U4418 ( .A1(n3881), .A2(n3880), .A3(n3879), .ZN(n3899) );
  OAI211_X1 U4419 ( .C1(n3885), .C2(n3884), .A(n3883), .B(n3882), .ZN(n3889)
         );
  INV_X1 U4420 ( .A(n3886), .ZN(n3888) );
  AOI21_X1 U4421 ( .B1(n3889), .B2(n3888), .A(n3887), .ZN(n3891) );
  NOR2_X1 U4422 ( .A1(n3891), .A2(n3136), .ZN(n3893) );
  AOI21_X1 U4423 ( .B1(n3894), .B2(n3893), .A(n3892), .ZN(n3897) );
  OAI21_X1 U4424 ( .B1(n3897), .B2(n3896), .A(n3895), .ZN(n3898) );
  AOI22_X1 U4425 ( .A1(n3901), .A2(n3900), .B1(n3899), .B2(n3898), .ZN(n3907)
         );
  OAI21_X1 U4426 ( .B1(n3902), .B2(n4681), .A(n3904), .ZN(n3906) );
  NOR2_X1 U4427 ( .A1(n3904), .A2(n3903), .ZN(n3905) );
  AOI21_X1 U4428 ( .B1(n3907), .B2(n3906), .A(n3905), .ZN(n3952) );
  NAND2_X1 U4429 ( .A1(n3908), .A2(n4079), .ZN(n4101) );
  NAND2_X1 U4430 ( .A1(n3909), .A2(n4098), .ZN(n4121) );
  NAND2_X1 U4431 ( .A1(n3910), .A2(n4117), .ZN(n4147) );
  NAND2_X1 U4432 ( .A1(n3912), .A2(n3911), .ZN(n4208) );
  NOR4_X1 U4433 ( .A1(n4101), .A2(n4121), .A3(n4147), .A4(n4208), .ZN(n3922)
         );
  XNOR2_X1 U4434 ( .A(n3976), .B(n4318), .ZN(n4307) );
  NAND4_X1 U4435 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3920)
         );
  INV_X1 U4436 ( .A(n3917), .ZN(n3919) );
  NAND2_X1 U4437 ( .A1(n3919), .A2(n3918), .ZN(n4231) );
  NOR3_X1 U4438 ( .A1(n4062), .A2(n3920), .A3(n4231), .ZN(n3921) );
  NAND3_X1 U4439 ( .A1(n3922), .A2(n4307), .A3(n3921), .ZN(n3949) );
  INV_X1 U4440 ( .A(n4167), .ZN(n4165) );
  NOR4_X1 U4441 ( .A1(n4165), .A2(n3064), .A3(n3924), .A4(n3923), .ZN(n3938)
         );
  AND4_X1 U4442 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3936)
         );
  NAND2_X1 U4443 ( .A1(n4219), .A2(n4220), .ZN(n4264) );
  NOR4_X1 U4444 ( .A1(n3934), .A2(n3933), .A3(n4264), .A4(n3932), .ZN(n3935)
         );
  NAND4_X1 U4445 ( .A1(n3938), .A2(n3937), .A3(n3936), .A4(n3935), .ZN(n3948)
         );
  INV_X1 U4446 ( .A(n4141), .ZN(n3939) );
  AND2_X1 U4447 ( .A1(n3939), .A2(n4142), .ZN(n4184) );
  INV_X1 U4448 ( .A(n4288), .ZN(n3945) );
  NAND2_X1 U4449 ( .A1(n3941), .A2(n3940), .ZN(n4082) );
  INV_X1 U4450 ( .A(n4082), .ZN(n3944) );
  AND2_X1 U4451 ( .A1(n3943), .A2(n3942), .ZN(n4787) );
  NAND4_X1 U4452 ( .A1(n4184), .A2(n3945), .A3(n3944), .A4(n4787), .ZN(n3946)
         );
  OR4_X1 U4453 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3951) );
  MUX2_X1 U4454 ( .A(n3952), .B(n3951), .S(n3950), .Z(n3953) );
  XNOR2_X1 U4455 ( .A(n3953), .B(n2782), .ZN(n3955) );
  NAND2_X1 U4456 ( .A1(n3957), .A2(n2782), .ZN(n3954) );
  MUX2_X1 U4457 ( .A(n3955), .B(n3954), .S(n2922), .Z(n3956) );
  OAI21_X1 U4458 ( .B1(n3957), .B2(n4798), .A(n3956), .ZN(n3966) );
  INV_X1 U4459 ( .A(n4469), .ZN(n3965) );
  NOR4_X1 U4460 ( .A1(n3960), .A2(n3959), .A3(n4851), .A4(n3958), .ZN(n3961)
         );
  NAND2_X1 U4461 ( .A1(n3961), .A2(n2538), .ZN(n3963) );
  MUX2_X1 U4462 ( .A(n4469), .B(n3963), .S(n3962), .Z(n3964) );
  AOI22_X1 U4463 ( .A1(n3966), .A2(n3965), .B1(B_REG_SCAN_IN), .B2(n3964), 
        .ZN(n3967) );
  INV_X1 U4464 ( .A(n3967), .ZN(U3239) );
  MUX2_X1 U4465 ( .A(DATAO_REG_30__SCAN_IN), .B(n3968), .S(n4683), .Z(U3580)
         );
  MUX2_X1 U4466 ( .A(DATAO_REG_29__SCAN_IN), .B(n4054), .S(n4683), .Z(U3579)
         );
  MUX2_X1 U4467 ( .A(DATAO_REG_28__SCAN_IN), .B(n3969), .S(n4683), .Z(U3578)
         );
  MUX2_X1 U4468 ( .A(DATAO_REG_27__SCAN_IN), .B(n3970), .S(n4683), .Z(U3577)
         );
  MUX2_X1 U4469 ( .A(DATAO_REG_26__SCAN_IN), .B(n4104), .S(n4683), .Z(U3576)
         );
  MUX2_X1 U4470 ( .A(DATAO_REG_25__SCAN_IN), .B(n3971), .S(n4683), .Z(U3575)
         );
  MUX2_X1 U4471 ( .A(DATAO_REG_24__SCAN_IN), .B(n4151), .S(n4683), .Z(U3574)
         );
  MUX2_X1 U4472 ( .A(DATAO_REG_23__SCAN_IN), .B(n4125), .S(n4683), .Z(U3573)
         );
  MUX2_X1 U4473 ( .A(DATAO_REG_22__SCAN_IN), .B(n4187), .S(n4683), .Z(U3572)
         );
  MUX2_X1 U4474 ( .A(DATAO_REG_21__SCAN_IN), .B(n4204), .S(n4683), .Z(U3571)
         );
  MUX2_X1 U4475 ( .A(DATAO_REG_20__SCAN_IN), .B(n3972), .S(n4683), .Z(U3570)
         );
  MUX2_X1 U4476 ( .A(DATAO_REG_19__SCAN_IN), .B(n4245), .S(n4683), .Z(U3569)
         );
  MUX2_X1 U4477 ( .A(DATAO_REG_18__SCAN_IN), .B(n3973), .S(n4683), .Z(U3568)
         );
  MUX2_X1 U4478 ( .A(DATAO_REG_17__SCAN_IN), .B(n3974), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4479 ( .A(DATAO_REG_16__SCAN_IN), .B(n4923), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4480 ( .A(DATAO_REG_15__SCAN_IN), .B(n3975), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4481 ( .A(DATAO_REG_14__SCAN_IN), .B(n4921), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4482 ( .A(DATAO_REG_13__SCAN_IN), .B(n3976), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4483 ( .A(DATAO_REG_12__SCAN_IN), .B(n3977), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4484 ( .A(DATAO_REG_11__SCAN_IN), .B(n3978), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4485 ( .A(DATAO_REG_10__SCAN_IN), .B(n3979), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4486 ( .A(DATAO_REG_9__SCAN_IN), .B(n3980), .S(n4683), .Z(U3559) );
  MUX2_X1 U4487 ( .A(DATAO_REG_8__SCAN_IN), .B(n4860), .S(n4683), .Z(U3558) );
  MUX2_X1 U4488 ( .A(DATAO_REG_7__SCAN_IN), .B(n3981), .S(U4043), .Z(U3557) );
  MUX2_X1 U4489 ( .A(DATAO_REG_6__SCAN_IN), .B(n3982), .S(n4683), .Z(U3556) );
  MUX2_X1 U4490 ( .A(DATAO_REG_5__SCAN_IN), .B(n3983), .S(n4683), .Z(U3555) );
  MUX2_X1 U4491 ( .A(DATAO_REG_4__SCAN_IN), .B(n3984), .S(n4683), .Z(U3554) );
  MUX2_X1 U4492 ( .A(DATAO_REG_3__SCAN_IN), .B(n3985), .S(n4683), .Z(U3553) );
  MUX2_X1 U4493 ( .A(DATAO_REG_2__SCAN_IN), .B(n3986), .S(n4683), .Z(U3552) );
  MUX2_X1 U4494 ( .A(DATAO_REG_1__SCAN_IN), .B(n3049), .S(n4683), .Z(U3551) );
  MUX2_X1 U4495 ( .A(DATAO_REG_0__SCAN_IN), .B(n3987), .S(n4683), .Z(U3550) );
  INV_X1 U4496 ( .A(n4785), .ZN(n4007) );
  NAND2_X1 U4497 ( .A1(n4007), .A2(n4468), .ZN(n3998) );
  NOR2_X1 U4498 ( .A1(n4786), .A2(n2964), .ZN(n3991) );
  MUX2_X1 U4499 ( .A(n4809), .B(REG1_REG_1__SCAN_IN), .S(n3988), .Z(n3990) );
  OAI211_X1 U4500 ( .C1(n3991), .C2(n3990), .A(n4780), .B(n3989), .ZN(n3997)
         );
  OAI211_X1 U4501 ( .C1(n3994), .C2(n3993), .A(n4754), .B(n3992), .ZN(n3996)
         );
  AOI22_X1 U4502 ( .A1(n4779), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3995) );
  NAND4_X1 U4503 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(U3241)
         );
  XNOR2_X1 U4504 ( .A(n4000), .B(n3999), .ZN(n4010) );
  AND2_X1 U4505 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4925) );
  INV_X1 U4506 ( .A(n4001), .ZN(n4005) );
  INV_X1 U4507 ( .A(n4002), .ZN(n4003) );
  AOI211_X1 U4508 ( .C1(n4005), .C2(n4004), .A(n4003), .B(n4774), .ZN(n4006)
         );
  AOI211_X1 U4509 ( .C1(n4779), .C2(ADDR_REG_15__SCAN_IN), .A(n4925), .B(n4006), .ZN(n4009) );
  NAND2_X1 U4510 ( .A1(n4007), .A2(n4464), .ZN(n4008) );
  OAI211_X1 U4511 ( .C1(n4768), .C2(n4010), .A(n4009), .B(n4008), .ZN(U3255)
         );
  AOI21_X1 U4512 ( .B1(n4013), .B2(n4012), .A(n4011), .ZN(n4023) );
  AOI221_X1 U4513 ( .B1(n4016), .B2(n4015), .C1(n4014), .C2(n4015), .A(n4774), 
        .ZN(n4017) );
  OR2_X1 U4514 ( .A1(n4018), .A2(n4017), .ZN(n4019) );
  AOI21_X1 U4515 ( .B1(n4779), .B2(ADDR_REG_17__SCAN_IN), .A(n4019), .ZN(n4022) );
  OR2_X1 U4516 ( .A1(n4785), .A2(n4020), .ZN(n4021) );
  OAI211_X1 U4517 ( .C1(n4023), .C2(n4768), .A(n4022), .B(n4021), .ZN(U3257)
         );
  XNOR2_X1 U4518 ( .A(n4025), .B(n4024), .ZN(n4026) );
  NAND2_X1 U4519 ( .A1(n4780), .A2(n4026), .ZN(n4033) );
  AOI211_X1 U4520 ( .C1(n4029), .C2(n4028), .A(n4027), .B(n4774), .ZN(n4030)
         );
  AOI211_X1 U4521 ( .C1(n4779), .C2(ADDR_REG_18__SCAN_IN), .A(n4031), .B(n4030), .ZN(n4032) );
  OAI211_X1 U4522 ( .C1(n4034), .C2(n4785), .A(n4033), .B(n4032), .ZN(U3258)
         );
  INV_X1 U4523 ( .A(n4035), .ZN(n4042) );
  OAI22_X1 U4524 ( .A1(n4037), .A2(n4905), .B1(n4036), .B2(n4909), .ZN(n4038)
         );
  OAI21_X1 U4525 ( .B1(n4039), .B2(n4038), .A(n4849), .ZN(n4041) );
  NAND2_X1 U4526 ( .A1(n4944), .A2(REG2_REG_29__SCAN_IN), .ZN(n4040) );
  OAI211_X1 U4527 ( .C1(n4042), .C2(n4278), .A(n4041), .B(n4040), .ZN(U3354)
         );
  XNOR2_X1 U4528 ( .A(n4043), .B(n4050), .ZN(n4337) );
  AOI22_X1 U4529 ( .A1(n4944), .A2(REG2_REG_28__SCAN_IN), .B1(n4044), .B2(
        n4891), .ZN(n4060) );
  INV_X1 U4530 ( .A(n4072), .ZN(n4047) );
  INV_X1 U4531 ( .A(n4045), .ZN(n4046) );
  OAI211_X1 U4532 ( .C1(n4047), .C2(n4052), .A(n4046), .B(n3160), .ZN(n4335)
         );
  INV_X1 U4533 ( .A(n4048), .ZN(n4049) );
  NOR2_X1 U4534 ( .A1(n4061), .A2(n4049), .ZN(n4051) );
  XNOR2_X1 U4535 ( .A(n4051), .B(n4050), .ZN(n4057) );
  NOR2_X1 U4536 ( .A1(n4855), .A2(n4052), .ZN(n4053) );
  AOI21_X1 U4537 ( .B1(n4054), .B2(n4861), .A(n4053), .ZN(n4055) );
  OAI21_X1 U4538 ( .B1(n4085), .B2(n4857), .A(n4055), .ZN(n4056) );
  AOI21_X1 U4539 ( .B1(n4057), .B2(n4791), .A(n4056), .ZN(n4336) );
  OAI21_X1 U4540 ( .B1(n4851), .B2(n4335), .A(n4336), .ZN(n4058) );
  NAND2_X1 U4541 ( .A1(n4058), .A2(n4849), .ZN(n4059) );
  OAI211_X1 U4542 ( .C1(n4337), .C2(n4278), .A(n4060), .B(n4059), .ZN(U3262)
         );
  AOI21_X1 U4543 ( .B1(n4063), .B2(n4062), .A(n4061), .ZN(n4067) );
  OAI22_X1 U4544 ( .A1(n4064), .A2(n4794), .B1(n4855), .B2(n4073), .ZN(n4065)
         );
  AOI21_X1 U4545 ( .B1(n4267), .B2(n4104), .A(n4065), .ZN(n4066) );
  OAI21_X1 U4546 ( .B1(n4067), .B2(n4863), .A(n4066), .ZN(n4338) );
  AOI21_X1 U4547 ( .B1(n4068), .B2(n4891), .A(n4338), .ZN(n4077) );
  XNOR2_X1 U4548 ( .A(n4070), .B(n4069), .ZN(n4339) );
  NAND2_X1 U4549 ( .A1(n4339), .A2(n4290), .ZN(n4076) );
  OAI21_X1 U4550 ( .B1(n4071), .B2(n4073), .A(n4072), .ZN(n4414) );
  INV_X1 U4551 ( .A(n4414), .ZN(n4074) );
  AOI22_X1 U4552 ( .A1(n4074), .A2(n4940), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4944), .ZN(n4075) );
  OAI211_X1 U4553 ( .C1(n4944), .C2(n4077), .A(n4076), .B(n4075), .ZN(U3263)
         );
  XNOR2_X1 U4554 ( .A(n4078), .B(n4082), .ZN(n4346) );
  INV_X1 U4555 ( .A(n4079), .ZN(n4080) );
  NOR2_X1 U4556 ( .A1(n4081), .A2(n4080), .ZN(n4083) );
  XNOR2_X1 U4557 ( .A(n4083), .B(n4082), .ZN(n4088) );
  NOR2_X1 U4558 ( .A1(n4123), .A2(n4857), .ZN(n4087) );
  OAI22_X1 U4559 ( .A1(n4085), .A2(n4794), .B1(n4855), .B2(n4084), .ZN(n4086)
         );
  AOI211_X1 U4560 ( .C1(n4088), .C2(n4791), .A(n4087), .B(n4086), .ZN(n4345)
         );
  INV_X1 U4561 ( .A(n4345), .ZN(n4095) );
  INV_X1 U4562 ( .A(n4071), .ZN(n4343) );
  INV_X1 U4563 ( .A(n4089), .ZN(n4108) );
  NAND2_X1 U4564 ( .A1(n4108), .A2(n4090), .ZN(n4342) );
  AND3_X1 U4565 ( .A1(n4343), .A2(n4940), .A3(n4342), .ZN(n4094) );
  INV_X1 U4566 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4092) );
  OAI22_X1 U4567 ( .A1(n4849), .A2(n4092), .B1(n4091), .B2(n4909), .ZN(n4093)
         );
  AOI211_X1 U4568 ( .C1(n4095), .C2(n4849), .A(n4094), .B(n4093), .ZN(n4096)
         );
  OAI21_X1 U4569 ( .B1(n4346), .B2(n4278), .A(n4096), .ZN(U3264) );
  XOR2_X1 U4570 ( .A(n4101), .B(n4097), .Z(n4348) );
  INV_X1 U4571 ( .A(n4348), .ZN(n4115) );
  INV_X1 U4572 ( .A(n4098), .ZN(n4099) );
  NOR2_X1 U4573 ( .A1(n4100), .A2(n4099), .ZN(n4102) );
  XNOR2_X1 U4574 ( .A(n4102), .B(n4101), .ZN(n4107) );
  NOR2_X1 U4575 ( .A1(n4855), .A2(n4109), .ZN(n4103) );
  AOI21_X1 U4576 ( .B1(n4104), .B2(n4861), .A(n4103), .ZN(n4106) );
  NAND2_X1 U4577 ( .A1(n4151), .A2(n4267), .ZN(n4105) );
  OAI211_X1 U4578 ( .C1(n4107), .C2(n4863), .A(n4106), .B(n4105), .ZN(n4347)
         );
  INV_X1 U4579 ( .A(n4130), .ZN(n4110) );
  OAI21_X1 U4580 ( .B1(n4110), .B2(n4109), .A(n4108), .ZN(n4419) );
  AOI22_X1 U4581 ( .A1(n4944), .A2(REG2_REG_25__SCAN_IN), .B1(n4111), .B2(
        n4891), .ZN(n4112) );
  OAI21_X1 U4582 ( .B1(n4419), .B2(n4905), .A(n4112), .ZN(n4113) );
  AOI21_X1 U4583 ( .B1(n4347), .B2(n4849), .A(n4113), .ZN(n4114) );
  OAI21_X1 U4584 ( .B1(n4115), .B2(n4278), .A(n4114), .ZN(U3265) );
  XOR2_X1 U4585 ( .A(n4121), .B(n4116), .Z(n4352) );
  INV_X1 U4586 ( .A(n4352), .ZN(n4135) );
  INV_X1 U4587 ( .A(n4117), .ZN(n4118) );
  NOR2_X1 U4588 ( .A1(n4119), .A2(n4118), .ZN(n4120) );
  XOR2_X1 U4589 ( .A(n4121), .B(n4120), .Z(n4127) );
  OAI22_X1 U4590 ( .A1(n4123), .A2(n4794), .B1(n4855), .B2(n4122), .ZN(n4124)
         );
  AOI21_X1 U4591 ( .B1(n4267), .B2(n4125), .A(n4124), .ZN(n4126) );
  OAI21_X1 U4592 ( .B1(n4127), .B2(n4863), .A(n4126), .ZN(n4351) );
  NAND2_X1 U4593 ( .A1(n4157), .A2(n4128), .ZN(n4129) );
  NAND2_X1 U4594 ( .A1(n4130), .A2(n4129), .ZN(n4423) );
  AOI22_X1 U4595 ( .A1(n4944), .A2(REG2_REG_24__SCAN_IN), .B1(n4131), .B2(
        n4891), .ZN(n4132) );
  OAI21_X1 U4596 ( .B1(n4423), .B2(n4905), .A(n4132), .ZN(n4133) );
  AOI21_X1 U4597 ( .B1(n4351), .B2(n4849), .A(n4133), .ZN(n4134) );
  OAI21_X1 U4598 ( .B1(n4135), .B2(n4278), .A(n4134), .ZN(U3266) );
  OAI21_X1 U4599 ( .B1(n4182), .B2(n4137), .A(n4136), .ZN(n4166) );
  INV_X1 U4600 ( .A(n4166), .ZN(n4138) );
  NOR2_X1 U4601 ( .A1(n4138), .A2(n4167), .ZN(n4163) );
  NOR2_X1 U4602 ( .A1(n4163), .A2(n4139), .ZN(n4140) );
  XNOR2_X1 U4603 ( .A(n4140), .B(n4147), .ZN(n4356) );
  INV_X1 U4604 ( .A(n4356), .ZN(n4162) );
  NAND2_X1 U4605 ( .A1(n4143), .A2(n4142), .ZN(n4168) );
  INV_X1 U4606 ( .A(n4144), .ZN(n4145) );
  AOI21_X1 U4607 ( .B1(n4168), .B2(n4167), .A(n4145), .ZN(n4146) );
  XOR2_X1 U4608 ( .A(n4147), .B(n4146), .Z(n4153) );
  OAI22_X1 U4609 ( .A1(n4149), .A2(n4857), .B1(n4148), .B2(n4855), .ZN(n4150)
         );
  AOI21_X1 U4610 ( .B1(n4861), .B2(n4151), .A(n4150), .ZN(n4152) );
  OAI21_X1 U4611 ( .B1(n4153), .B2(n4863), .A(n4152), .ZN(n4355) );
  NAND2_X1 U4612 ( .A1(n4359), .A2(n4155), .ZN(n4156) );
  NAND2_X1 U4613 ( .A1(n4157), .A2(n4156), .ZN(n4427) );
  AOI22_X1 U4614 ( .A1(n4944), .A2(REG2_REG_23__SCAN_IN), .B1(n4158), .B2(
        n4891), .ZN(n4159) );
  OAI21_X1 U4615 ( .B1(n4427), .B2(n4905), .A(n4159), .ZN(n4160) );
  AOI21_X1 U4616 ( .B1(n4355), .B2(n4849), .A(n4160), .ZN(n4161) );
  OAI21_X1 U4617 ( .B1(n4162), .B2(n4278), .A(n4161), .ZN(U3267) );
  INV_X1 U4618 ( .A(n4163), .ZN(n4164) );
  OAI21_X1 U4619 ( .B1(n4166), .B2(n4165), .A(n4164), .ZN(n4363) );
  XNOR2_X1 U4620 ( .A(n4168), .B(n4167), .ZN(n4173) );
  NOR2_X1 U4621 ( .A1(n4855), .A2(n4177), .ZN(n4169) );
  AOI21_X1 U4622 ( .B1(n4204), .B2(n4267), .A(n4169), .ZN(n4170) );
  OAI21_X1 U4623 ( .B1(n4171), .B2(n4794), .A(n4170), .ZN(n4172) );
  AOI21_X1 U4624 ( .B1(n4173), .B2(n4791), .A(n4172), .ZN(n4362) );
  INV_X1 U4625 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4175) );
  OAI22_X1 U4626 ( .A1(n4849), .A2(n4175), .B1(n4174), .B2(n4909), .ZN(n4176)
         );
  INV_X1 U4627 ( .A(n4176), .ZN(n4179) );
  OR2_X1 U4628 ( .A1(n4190), .A2(n4177), .ZN(n4360) );
  NAND3_X1 U4629 ( .A1(n4359), .A2(n4360), .A3(n4940), .ZN(n4178) );
  OAI211_X1 U4630 ( .C1(n4362), .C2(n4944), .A(n4179), .B(n4178), .ZN(n4180)
         );
  INV_X1 U4631 ( .A(n4180), .ZN(n4181) );
  OAI21_X1 U4632 ( .B1(n4363), .B2(n4278), .A(n4181), .ZN(U3268) );
  XOR2_X1 U4633 ( .A(n4184), .B(n4182), .Z(n4365) );
  INV_X1 U4634 ( .A(n4365), .ZN(n4199) );
  XOR2_X1 U4635 ( .A(n4184), .B(n4183), .Z(n4185) );
  NAND2_X1 U4636 ( .A1(n4185), .A2(n4791), .ZN(n4189) );
  NOR2_X1 U4637 ( .A1(n4855), .A2(n4192), .ZN(n4186) );
  AOI21_X1 U4638 ( .B1(n4187), .B2(n4861), .A(n4186), .ZN(n4188) );
  OAI211_X1 U4639 ( .C1(n4226), .C2(n4857), .A(n4189), .B(n4188), .ZN(n4364)
         );
  INV_X1 U4640 ( .A(n4369), .ZN(n4193) );
  INV_X1 U4641 ( .A(n4190), .ZN(n4191) );
  OAI21_X1 U4642 ( .B1(n4193), .B2(n4192), .A(n4191), .ZN(n4432) );
  NOR2_X1 U4643 ( .A1(n4432), .A2(n4905), .ZN(n4197) );
  INV_X1 U4644 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4195) );
  OAI22_X1 U4645 ( .A1(n4849), .A2(n4195), .B1(n4194), .B2(n4909), .ZN(n4196)
         );
  AOI211_X1 U4646 ( .C1(n4364), .C2(n4849), .A(n4197), .B(n4196), .ZN(n4198)
         );
  OAI21_X1 U4647 ( .B1(n4199), .B2(n4278), .A(n4198), .ZN(U3269) );
  NAND2_X1 U4648 ( .A1(n4200), .A2(n4219), .ZN(n4202) );
  OAI21_X1 U4649 ( .B1(n4265), .B2(n4202), .A(n4201), .ZN(n4203) );
  XOR2_X1 U4650 ( .A(n4208), .B(n4203), .Z(n4211) );
  INV_X1 U4651 ( .A(n4245), .ZN(n4206) );
  AOI22_X1 U4652 ( .A1(n4204), .A2(n4861), .B1(n4331), .B2(n4212), .ZN(n4205)
         );
  OAI21_X1 U4653 ( .B1(n4206), .B2(n4857), .A(n4205), .ZN(n4210) );
  XNOR2_X1 U4654 ( .A(n4207), .B(n4208), .ZN(n4372) );
  NOR2_X1 U4655 ( .A1(n4372), .A2(n4316), .ZN(n4209) );
  AOI211_X1 U4656 ( .C1(n4211), .C2(n4791), .A(n4210), .B(n4209), .ZN(n4371)
         );
  INV_X1 U4657 ( .A(n4372), .ZN(n4217) );
  NAND2_X1 U4658 ( .A1(n4232), .A2(n4212), .ZN(n4368) );
  AND3_X1 U4659 ( .A1(n4369), .A2(n4940), .A3(n4368), .ZN(n4216) );
  INV_X1 U4660 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4214) );
  OAI22_X1 U4661 ( .A1(n4849), .A2(n4214), .B1(n4213), .B2(n4909), .ZN(n4215)
         );
  AOI211_X1 U4662 ( .C1(n4217), .C2(n4895), .A(n4216), .B(n4215), .ZN(n4218)
         );
  OAI21_X1 U4663 ( .B1(n4371), .B2(n4944), .A(n4218), .ZN(U3270) );
  INV_X1 U4664 ( .A(n4219), .ZN(n4221) );
  OAI21_X1 U4665 ( .B1(n4265), .B2(n4221), .A(n4220), .ZN(n4243) );
  INV_X1 U4666 ( .A(n4222), .ZN(n4224) );
  OAI21_X1 U4667 ( .B1(n4243), .B2(n4224), .A(n4223), .ZN(n4225) );
  XNOR2_X1 U4668 ( .A(n4225), .B(n4231), .ZN(n4229) );
  NOR2_X1 U4669 ( .A1(n4270), .A2(n4857), .ZN(n4228) );
  OAI22_X1 U4670 ( .A1(n4226), .A2(n4794), .B1(n4233), .B2(n4855), .ZN(n4227)
         );
  AOI211_X1 U4671 ( .C1(n4229), .C2(n4791), .A(n4228), .B(n4227), .ZN(n4373)
         );
  XNOR2_X1 U4672 ( .A(n4230), .B(n4231), .ZN(n4375) );
  NAND2_X1 U4673 ( .A1(n4375), .A2(n4290), .ZN(n4238) );
  OAI21_X1 U4674 ( .B1(n4239), .B2(n4233), .A(n4232), .ZN(n4437) );
  INV_X1 U4675 ( .A(n4437), .ZN(n4236) );
  OAI22_X1 U4676 ( .A1(n4849), .A2(n3038), .B1(n4234), .B2(n4909), .ZN(n4235)
         );
  AOI21_X1 U4677 ( .B1(n4236), .B2(n4940), .A(n4235), .ZN(n4237) );
  OAI211_X1 U4678 ( .C1(n4944), .C2(n4373), .A(n4238), .B(n4237), .ZN(U3271)
         );
  INV_X1 U4679 ( .A(n4273), .ZN(n4242) );
  INV_X1 U4680 ( .A(n4239), .ZN(n4240) );
  OAI211_X1 U4681 ( .C1(n4242), .C2(n4241), .A(n4240), .B(n3160), .ZN(n4377)
         );
  XNOR2_X1 U4682 ( .A(n4243), .B(n4257), .ZN(n4249) );
  AOI22_X1 U4683 ( .A1(n4245), .A2(n4861), .B1(n4244), .B2(n4331), .ZN(n4246)
         );
  OAI21_X1 U4684 ( .B1(n4247), .B2(n4857), .A(n4246), .ZN(n4248) );
  AOI21_X1 U4685 ( .B1(n4249), .B2(n4791), .A(n4248), .ZN(n4378) );
  OAI21_X1 U4686 ( .B1(n4851), .B2(n4377), .A(n4378), .ZN(n4260) );
  OAI22_X1 U4687 ( .A1(n4849), .A2(n3037), .B1(n4250), .B2(n4909), .ZN(n4259)
         );
  NAND2_X1 U4688 ( .A1(n3572), .A2(n4251), .ZN(n4253) );
  AND2_X1 U4689 ( .A1(n4253), .A2(n4252), .ZN(n4256) );
  INV_X1 U4690 ( .A(n4254), .ZN(n4255) );
  AOI21_X1 U4691 ( .B1(n4257), .B2(n4256), .A(n4255), .ZN(n4379) );
  NOR2_X1 U4692 ( .A1(n4379), .A2(n4278), .ZN(n4258) );
  AOI211_X1 U4693 ( .C1(n4849), .C2(n4260), .A(n4259), .B(n4258), .ZN(n4261)
         );
  INV_X1 U4694 ( .A(n4261), .ZN(U3272) );
  NAND2_X1 U4695 ( .A1(n3572), .A2(n4262), .ZN(n4263) );
  XOR2_X1 U4696 ( .A(n4264), .B(n4263), .Z(n4381) );
  INV_X1 U4697 ( .A(n4381), .ZN(n4279) );
  XNOR2_X1 U4698 ( .A(n4265), .B(n4264), .ZN(n4266) );
  NAND2_X1 U4699 ( .A1(n4266), .A2(n4791), .ZN(n4269) );
  AOI22_X1 U4700 ( .A1(n4923), .A2(n4267), .B1(n4331), .B2(n4271), .ZN(n4268)
         );
  OAI211_X1 U4701 ( .C1(n4270), .C2(n4794), .A(n4269), .B(n4268), .ZN(n4380)
         );
  NAND2_X1 U4702 ( .A1(n4383), .A2(n4271), .ZN(n4272) );
  NAND2_X1 U4703 ( .A1(n4273), .A2(n4272), .ZN(n4442) );
  AOI22_X1 U4704 ( .A1(n4944), .A2(REG2_REG_17__SCAN_IN), .B1(n4274), .B2(
        n4891), .ZN(n4275) );
  OAI21_X1 U4705 ( .B1(n4442), .B2(n4905), .A(n4275), .ZN(n4276) );
  AOI21_X1 U4706 ( .B1(n4380), .B2(n4849), .A(n4276), .ZN(n4277) );
  OAI21_X1 U4707 ( .B1(n4279), .B2(n4278), .A(n4277), .ZN(U3273) );
  OAI22_X1 U4708 ( .A1(n4311), .A2(n4857), .B1(n4294), .B2(n4855), .ZN(n4285)
         );
  NAND2_X1 U4709 ( .A1(n4281), .A2(n4280), .ZN(n4282) );
  XNOR2_X1 U4710 ( .A(n4282), .B(n4288), .ZN(n4283) );
  NOR2_X1 U4711 ( .A1(n4283), .A2(n4863), .ZN(n4284) );
  AOI211_X1 U4712 ( .C1(n4861), .C2(n4923), .A(n4285), .B(n4284), .ZN(n4389)
         );
  NAND2_X1 U4713 ( .A1(n4287), .A2(n4286), .ZN(n4289) );
  XNOR2_X1 U4714 ( .A(n4289), .B(n4288), .ZN(n4391) );
  NAND2_X1 U4715 ( .A1(n4391), .A2(n4290), .ZN(n4299) );
  INV_X1 U4716 ( .A(n4291), .ZN(n4292) );
  OAI21_X1 U4717 ( .B1(n4294), .B2(n4293), .A(n4292), .ZN(n4447) );
  INV_X1 U4718 ( .A(n4447), .ZN(n4297) );
  INV_X1 U4719 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4295) );
  OAI22_X1 U4720 ( .A1(n4849), .A2(n4295), .B1(n4937), .B2(n4909), .ZN(n4296)
         );
  AOI21_X1 U4721 ( .B1(n4297), .B2(n4940), .A(n4296), .ZN(n4298) );
  OAI211_X1 U4722 ( .C1(n4944), .C2(n4389), .A(n4299), .B(n4298), .ZN(U3275)
         );
  AND2_X1 U4723 ( .A1(n2409), .A2(n4301), .ZN(n4302) );
  XNOR2_X1 U4724 ( .A(n4302), .B(n4307), .ZN(n4317) );
  INV_X1 U4725 ( .A(n4303), .ZN(n4304) );
  AOI21_X1 U4726 ( .B1(n4306), .B2(n4305), .A(n4304), .ZN(n4308) );
  XNOR2_X1 U4727 ( .A(n4308), .B(n4307), .ZN(n4314) );
  NOR2_X1 U4728 ( .A1(n4309), .A2(n4857), .ZN(n4313) );
  OAI22_X1 U4729 ( .A1(n4311), .A2(n4794), .B1(n4310), .B2(n4855), .ZN(n4312)
         );
  AOI211_X1 U4730 ( .C1(n4314), .C2(n4791), .A(n4313), .B(n4312), .ZN(n4315)
         );
  OAI21_X1 U4731 ( .B1(n4317), .B2(n4316), .A(n4315), .ZN(n4398) );
  INV_X1 U4732 ( .A(n4398), .ZN(n4326) );
  INV_X1 U4733 ( .A(n4317), .ZN(n4399) );
  NAND2_X1 U4734 ( .A1(n4319), .A2(n4318), .ZN(n4320) );
  NAND2_X1 U4735 ( .A1(n4321), .A2(n4320), .ZN(n4455) );
  AOI22_X1 U4736 ( .A1(n4944), .A2(REG2_REG_13__SCAN_IN), .B1(n4322), .B2(
        n4891), .ZN(n4323) );
  OAI21_X1 U4737 ( .B1(n4455), .B2(n4905), .A(n4323), .ZN(n4324) );
  AOI21_X1 U4738 ( .B1(n4399), .B2(n4895), .A(n4324), .ZN(n4325) );
  OAI21_X1 U4739 ( .B1(n4326), .B2(n4944), .A(n4325), .ZN(U3277) );
  AOI21_X1 U4740 ( .B1(n4332), .B2(n4328), .A(n4327), .ZN(n4941) );
  INV_X1 U4741 ( .A(n4941), .ZN(n4409) );
  INV_X1 U4742 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4333) );
  INV_X1 U4743 ( .A(n4329), .ZN(n4330) );
  AOI21_X1 U4744 ( .B1(n4332), .B2(n4331), .A(n4330), .ZN(n4943) );
  MUX2_X1 U4745 ( .A(n4333), .B(n4943), .S(n4875), .Z(n4334) );
  OAI21_X1 U4746 ( .B1(n4409), .B2(n4406), .A(n4334), .ZN(U3548) );
  INV_X1 U4747 ( .A(n4871), .ZN(n4387) );
  OAI211_X1 U4748 ( .C1(n4337), .C2(n4387), .A(n4336), .B(n4335), .ZN(n4410)
         );
  MUX2_X1 U4749 ( .A(REG1_REG_28__SCAN_IN), .B(n4410), .S(n4875), .Z(U3546) );
  INV_X1 U4750 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4340) );
  AOI21_X1 U4751 ( .B1(n4339), .B2(n4871), .A(n4338), .ZN(n4411) );
  MUX2_X1 U4752 ( .A(n4340), .B(n4411), .S(n4875), .Z(n4341) );
  OAI21_X1 U4753 ( .B1(n4406), .B2(n4414), .A(n4341), .ZN(U3545) );
  NAND3_X1 U4754 ( .A1(n4343), .A2(n3160), .A3(n4342), .ZN(n4344) );
  OAI211_X1 U4755 ( .C1(n4346), .C2(n4387), .A(n4345), .B(n4344), .ZN(n4415)
         );
  MUX2_X1 U4756 ( .A(REG1_REG_26__SCAN_IN), .B(n4415), .S(n4875), .Z(U3544) );
  INV_X1 U4757 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4349) );
  AOI21_X1 U4758 ( .B1(n4348), .B2(n4871), .A(n4347), .ZN(n4416) );
  MUX2_X1 U4759 ( .A(n4349), .B(n4416), .S(n4875), .Z(n4350) );
  OAI21_X1 U4760 ( .B1(n4406), .B2(n4419), .A(n4350), .ZN(U3543) );
  INV_X1 U4761 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4353) );
  AOI21_X1 U4762 ( .B1(n4352), .B2(n4871), .A(n4351), .ZN(n4420) );
  MUX2_X1 U4763 ( .A(n4353), .B(n4420), .S(n4875), .Z(n4354) );
  OAI21_X1 U4764 ( .B1(n4406), .B2(n4423), .A(n4354), .ZN(U3542) );
  INV_X1 U4765 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4357) );
  AOI21_X1 U4766 ( .B1(n4356), .B2(n4871), .A(n4355), .ZN(n4424) );
  MUX2_X1 U4767 ( .A(n4357), .B(n4424), .S(n4875), .Z(n4358) );
  OAI21_X1 U4768 ( .B1(n4406), .B2(n4427), .A(n4358), .ZN(U3541) );
  NAND3_X1 U4769 ( .A1(n4360), .A2(n4359), .A3(n3160), .ZN(n4361) );
  OAI211_X1 U4770 ( .C1(n4363), .C2(n4387), .A(n4362), .B(n4361), .ZN(n4428)
         );
  MUX2_X1 U4771 ( .A(REG1_REG_22__SCAN_IN), .B(n4428), .S(n4875), .Z(U3540) );
  INV_X1 U4772 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4366) );
  AOI21_X1 U4773 ( .B1(n4365), .B2(n4871), .A(n4364), .ZN(n4429) );
  MUX2_X1 U4774 ( .A(n4366), .B(n4429), .S(n4875), .Z(n4367) );
  OAI21_X1 U4775 ( .B1(n4406), .B2(n4432), .A(n4367), .ZN(U3539) );
  NAND3_X1 U4776 ( .A1(n4369), .A2(n3160), .A3(n4368), .ZN(n4370) );
  OAI211_X1 U4777 ( .C1(n4372), .C2(n4804), .A(n4371), .B(n4370), .ZN(n4433)
         );
  MUX2_X1 U4778 ( .A(REG1_REG_20__SCAN_IN), .B(n4433), .S(n4875), .Z(U3538) );
  INV_X1 U4779 ( .A(n4373), .ZN(n4374) );
  AOI21_X1 U4780 ( .B1(n4375), .B2(n4871), .A(n4374), .ZN(n4434) );
  MUX2_X1 U4781 ( .A(n2998), .B(n4434), .S(n4875), .Z(n4376) );
  OAI21_X1 U4782 ( .B1(n4406), .B2(n4437), .A(n4376), .ZN(U3537) );
  OAI211_X1 U4783 ( .C1(n4379), .C2(n4387), .A(n4378), .B(n4377), .ZN(n4438)
         );
  MUX2_X1 U4784 ( .A(REG1_REG_18__SCAN_IN), .B(n4438), .S(n4875), .Z(U3536) );
  AOI21_X1 U4785 ( .B1(n4381), .B2(n4871), .A(n4380), .ZN(n4439) );
  MUX2_X1 U4786 ( .A(n2994), .B(n4439), .S(n4875), .Z(n4382) );
  OAI21_X1 U4787 ( .B1(n4406), .B2(n4442), .A(n4382), .ZN(U3535) );
  NAND3_X1 U4788 ( .A1(n4384), .A2(n3160), .A3(n4383), .ZN(n4385) );
  OAI211_X1 U4789 ( .C1(n4388), .C2(n4387), .A(n4386), .B(n4385), .ZN(n4443)
         );
  MUX2_X1 U4790 ( .A(REG1_REG_16__SCAN_IN), .B(n4443), .S(n4875), .Z(U3534) );
  INV_X1 U4791 ( .A(n4389), .ZN(n4390) );
  AOI21_X1 U4792 ( .B1(n4871), .B2(n4391), .A(n4390), .ZN(n4444) );
  MUX2_X1 U4793 ( .A(n4392), .B(n4444), .S(n4875), .Z(n4393) );
  OAI21_X1 U4794 ( .B1(n4406), .B2(n4447), .A(n4393), .ZN(U3533) );
  AOI21_X1 U4795 ( .B1(n4395), .B2(n4871), .A(n4394), .ZN(n4449) );
  INV_X1 U4796 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4396) );
  MUX2_X1 U4797 ( .A(n4449), .B(n4396), .S(n4873), .Z(n4397) );
  OAI21_X1 U4798 ( .B1(n4406), .B2(n4451), .A(n4397), .ZN(U3532) );
  AOI21_X1 U4799 ( .B1(n4828), .B2(n4399), .A(n4398), .ZN(n4452) );
  MUX2_X1 U4800 ( .A(n4400), .B(n4452), .S(n4875), .Z(n4401) );
  OAI21_X1 U4801 ( .B1(n4406), .B2(n4455), .A(n4401), .ZN(U3531) );
  INV_X1 U4802 ( .A(n4402), .ZN(n4403) );
  AOI21_X1 U4803 ( .B1(n4871), .B2(n4404), .A(n4403), .ZN(n4456) );
  MUX2_X1 U4804 ( .A(n4750), .B(n4456), .S(n4875), .Z(n4405) );
  OAI21_X1 U4805 ( .B1(n4460), .B2(n4406), .A(n4405), .ZN(U3530) );
  INV_X1 U4806 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4407) );
  MUX2_X1 U4807 ( .A(n4407), .B(n4943), .S(n4879), .Z(n4408) );
  OAI21_X1 U4808 ( .B1(n4409), .B2(n4459), .A(n4408), .ZN(U3516) );
  MUX2_X1 U4809 ( .A(REG0_REG_28__SCAN_IN), .B(n4410), .S(n4879), .Z(U3514) );
  INV_X1 U4810 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4412) );
  MUX2_X1 U4811 ( .A(n4412), .B(n4411), .S(n4879), .Z(n4413) );
  OAI21_X1 U4812 ( .B1(n4414), .B2(n4459), .A(n4413), .ZN(U3513) );
  MUX2_X1 U4813 ( .A(REG0_REG_26__SCAN_IN), .B(n4415), .S(n4879), .Z(U3512) );
  INV_X1 U4814 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4417) );
  MUX2_X1 U4815 ( .A(n4417), .B(n4416), .S(n4879), .Z(n4418) );
  OAI21_X1 U4816 ( .B1(n4419), .B2(n4459), .A(n4418), .ZN(U3511) );
  INV_X1 U4817 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4421) );
  MUX2_X1 U4818 ( .A(n4421), .B(n4420), .S(n4879), .Z(n4422) );
  OAI21_X1 U4819 ( .B1(n4423), .B2(n4459), .A(n4422), .ZN(U3510) );
  INV_X1 U4820 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4425) );
  MUX2_X1 U4821 ( .A(n4425), .B(n4424), .S(n4879), .Z(n4426) );
  OAI21_X1 U4822 ( .B1(n4427), .B2(n4459), .A(n4426), .ZN(U3509) );
  MUX2_X1 U4823 ( .A(REG0_REG_22__SCAN_IN), .B(n4428), .S(n4879), .Z(U3508) );
  INV_X1 U4824 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4430) );
  MUX2_X1 U4825 ( .A(n4430), .B(n4429), .S(n4879), .Z(n4431) );
  OAI21_X1 U4826 ( .B1(n4432), .B2(n4459), .A(n4431), .ZN(U3507) );
  MUX2_X1 U4827 ( .A(REG0_REG_20__SCAN_IN), .B(n4433), .S(n4879), .Z(U3506) );
  INV_X1 U4828 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4435) );
  MUX2_X1 U4829 ( .A(n4435), .B(n4434), .S(n4879), .Z(n4436) );
  OAI21_X1 U4830 ( .B1(n4437), .B2(n4459), .A(n4436), .ZN(U3505) );
  MUX2_X1 U4831 ( .A(REG0_REG_18__SCAN_IN), .B(n4438), .S(n4879), .Z(U3503) );
  INV_X1 U4832 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4440) );
  MUX2_X1 U4833 ( .A(n4440), .B(n4439), .S(n4879), .Z(n4441) );
  OAI21_X1 U4834 ( .B1(n4442), .B2(n4459), .A(n4441), .ZN(U3501) );
  MUX2_X1 U4835 ( .A(REG0_REG_16__SCAN_IN), .B(n4443), .S(n4879), .Z(U3499) );
  INV_X1 U4836 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4445) );
  MUX2_X1 U4837 ( .A(n4445), .B(n4444), .S(n4879), .Z(n4446) );
  OAI21_X1 U4838 ( .B1(n4447), .B2(n4459), .A(n4446), .ZN(U3497) );
  INV_X1 U4839 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4448) );
  MUX2_X1 U4840 ( .A(n4449), .B(n4448), .S(n4876), .Z(n4450) );
  OAI21_X1 U4841 ( .B1(n4451), .B2(n4459), .A(n4450), .ZN(U3495) );
  INV_X1 U4842 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4453) );
  MUX2_X1 U4843 ( .A(n4453), .B(n4452), .S(n4879), .Z(n4454) );
  OAI21_X1 U4844 ( .B1(n4455), .B2(n4459), .A(n4454), .ZN(U3493) );
  INV_X1 U4845 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4457) );
  MUX2_X1 U4846 ( .A(n4457), .B(n4456), .S(n4879), .Z(n4458) );
  OAI21_X1 U4847 ( .B1(n4460), .B2(n4459), .A(n4458), .ZN(U3491) );
  MUX2_X1 U4848 ( .A(n4461), .B(D_REG_1__SCAN_IN), .S(n4470), .Z(U3459) );
  MUX2_X1 U4849 ( .A(DATAI_27_), .B(n4687), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U4850 ( .A(n2449), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4851 ( .A(DATAI_20_), .B(n4462), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4852 ( .A(DATAI_19_), .B(n4851), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4853 ( .A(n4463), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U4854 ( .A(n4464), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U4855 ( .A(n4465), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4856 ( .A(n4466), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U4857 ( .A(n4467), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4858 ( .A(n3007), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4859 ( .A(n4468), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U4860 ( .A(DATAI_23_), .ZN(n4580) );
  OAI21_X1 U4861 ( .B1(STATE_REG_SCAN_IN), .B2(n4580), .A(n4469), .ZN(U3329)
         );
  AND2_X1 U4862 ( .A1(D_REG_2__SCAN_IN), .A2(n4470), .ZN(U3320) );
  AND2_X1 U4863 ( .A1(D_REG_3__SCAN_IN), .A2(n4470), .ZN(U3319) );
  AND2_X1 U4864 ( .A1(D_REG_4__SCAN_IN), .A2(n4470), .ZN(U3318) );
  AND2_X1 U4865 ( .A1(D_REG_5__SCAN_IN), .A2(n4470), .ZN(U3317) );
  AND2_X1 U4866 ( .A1(D_REG_6__SCAN_IN), .A2(n4470), .ZN(U3316) );
  AND2_X1 U4867 ( .A1(D_REG_7__SCAN_IN), .A2(n4470), .ZN(U3315) );
  AND2_X1 U4868 ( .A1(D_REG_8__SCAN_IN), .A2(n4470), .ZN(U3314) );
  AND2_X1 U4869 ( .A1(D_REG_9__SCAN_IN), .A2(n4470), .ZN(U3313) );
  AND2_X1 U4870 ( .A1(D_REG_10__SCAN_IN), .A2(n4470), .ZN(U3312) );
  AND2_X1 U4871 ( .A1(D_REG_11__SCAN_IN), .A2(n4470), .ZN(U3311) );
  AND2_X1 U4872 ( .A1(D_REG_12__SCAN_IN), .A2(n4470), .ZN(U3310) );
  AND2_X1 U4873 ( .A1(D_REG_13__SCAN_IN), .A2(n4470), .ZN(U3309) );
  AND2_X1 U4874 ( .A1(D_REG_14__SCAN_IN), .A2(n4470), .ZN(U3308) );
  AND2_X1 U4875 ( .A1(D_REG_15__SCAN_IN), .A2(n4470), .ZN(U3307) );
  AND2_X1 U4876 ( .A1(D_REG_16__SCAN_IN), .A2(n4470), .ZN(U3306) );
  AND2_X1 U4877 ( .A1(D_REG_17__SCAN_IN), .A2(n4470), .ZN(U3305) );
  AND2_X1 U4878 ( .A1(D_REG_18__SCAN_IN), .A2(n4470), .ZN(U3304) );
  AND2_X1 U4879 ( .A1(D_REG_19__SCAN_IN), .A2(n4470), .ZN(U3303) );
  AND2_X1 U4880 ( .A1(D_REG_20__SCAN_IN), .A2(n4470), .ZN(U3302) );
  AND2_X1 U4881 ( .A1(D_REG_21__SCAN_IN), .A2(n4470), .ZN(U3301) );
  AND2_X1 U4882 ( .A1(D_REG_22__SCAN_IN), .A2(n4470), .ZN(U3300) );
  AND2_X1 U4883 ( .A1(D_REG_23__SCAN_IN), .A2(n4470), .ZN(U3299) );
  AND2_X1 U4884 ( .A1(D_REG_24__SCAN_IN), .A2(n4470), .ZN(U3298) );
  AND2_X1 U4885 ( .A1(D_REG_25__SCAN_IN), .A2(n4470), .ZN(U3297) );
  AND2_X1 U4886 ( .A1(D_REG_26__SCAN_IN), .A2(n4470), .ZN(U3296) );
  AND2_X1 U4887 ( .A1(D_REG_27__SCAN_IN), .A2(n4470), .ZN(U3295) );
  AND2_X1 U4888 ( .A1(D_REG_28__SCAN_IN), .A2(n4470), .ZN(U3294) );
  AND2_X1 U4889 ( .A1(D_REG_29__SCAN_IN), .A2(n4470), .ZN(U3293) );
  AND2_X1 U4890 ( .A1(D_REG_30__SCAN_IN), .A2(n4470), .ZN(U3292) );
  AND2_X1 U4891 ( .A1(D_REG_31__SCAN_IN), .A2(n4470), .ZN(U3291) );
  INV_X1 U4892 ( .A(keyinput_51), .ZN(n4547) );
  AOI22_X1 U4893 ( .A1(n4472), .A2(keyinput_49), .B1(n4569), .B2(keyinput_48), 
        .ZN(n4471) );
  OAI221_X1 U4894 ( .B1(n4472), .B2(keyinput_49), .C1(n4569), .C2(keyinput_48), 
        .A(n4471), .ZN(n4544) );
  INV_X1 U4895 ( .A(keyinput_38), .ZN(n4530) );
  AOI22_X1 U4896 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_36), .B1(
        REG3_REG_14__SCAN_IN), .B2(keyinput_35), .ZN(n4473) );
  OAI221_X1 U4897 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_36), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput_35), .A(n4473), .ZN(n4526) );
  AOI22_X1 U4898 ( .A1(U3149), .A2(keyinput_32), .B1(keyinput_31), .B2(n2485), 
        .ZN(n4474) );
  OAI221_X1 U4899 ( .B1(U3149), .B2(keyinput_32), .C1(n2485), .C2(keyinput_31), 
        .A(n4474), .ZN(n4477) );
  AOI22_X1 U4900 ( .A1(n2522), .A2(keyinput_29), .B1(n2600), .B2(keyinput_33), 
        .ZN(n4475) );
  OAI221_X1 U4901 ( .B1(n2522), .B2(keyinput_29), .C1(n2600), .C2(keyinput_33), 
        .A(n4475), .ZN(n4476) );
  AOI211_X1 U4902 ( .C1(keyinput_30), .C2(DATAI_1_), .A(n4477), .B(n4476), 
        .ZN(n4478) );
  OAI21_X1 U4903 ( .B1(keyinput_30), .B2(DATAI_1_), .A(n4478), .ZN(n4523) );
  INV_X1 U4904 ( .A(DATAI_3_), .ZN(n4627) );
  INV_X1 U4905 ( .A(keyinput_28), .ZN(n4521) );
  INV_X1 U4906 ( .A(keyinput_27), .ZN(n4519) );
  INV_X1 U4907 ( .A(DATAI_4_), .ZN(n4625) );
  INV_X1 U4908 ( .A(keyinput_26), .ZN(n4517) );
  INV_X1 U4909 ( .A(keyinput_25), .ZN(n4515) );
  INV_X1 U4910 ( .A(DATAI_6_), .ZN(n4832) );
  INV_X1 U4911 ( .A(DATAI_7_), .ZN(n4840) );
  INV_X1 U4912 ( .A(DATAI_9_), .ZN(n4887) );
  OAI22_X1 U4913 ( .A1(n4887), .A2(keyinput_22), .B1(DATAI_8_), .B2(
        keyinput_23), .ZN(n4479) );
  AOI221_X1 U4914 ( .B1(n4887), .B2(keyinput_22), .C1(keyinput_23), .C2(
        DATAI_8_), .A(n4479), .ZN(n4512) );
  INV_X1 U4915 ( .A(keyinput_21), .ZN(n4510) );
  INV_X1 U4916 ( .A(DATAI_10_), .ZN(n4889) );
  AOI22_X1 U4917 ( .A1(DATAI_25_), .A2(keyinput_6), .B1(n4481), .B2(keyinput_7), .ZN(n4480) );
  OAI221_X1 U4918 ( .B1(DATAI_25_), .B2(keyinput_6), .C1(n4481), .C2(
        keyinput_7), .A(n4480), .ZN(n4485) );
  INV_X1 U4919 ( .A(DATAI_27_), .ZN(n4483) );
  AOI22_X1 U4920 ( .A1(DATAI_26_), .A2(keyinput_5), .B1(n4483), .B2(keyinput_4), .ZN(n4482) );
  OAI221_X1 U4921 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(n4483), .C2(
        keyinput_4), .A(n4482), .ZN(n4484) );
  AOI211_X1 U4922 ( .C1(keyinput_8), .C2(DATAI_23_), .A(n4485), .B(n4484), 
        .ZN(n4486) );
  OAI21_X1 U4923 ( .B1(keyinput_8), .B2(DATAI_23_), .A(n4486), .ZN(n4493) );
  INV_X1 U4924 ( .A(keyinput_3), .ZN(n4491) );
  INV_X1 U4925 ( .A(keyinput_2), .ZN(n4489) );
  OAI22_X1 U4926 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        DATAI_31_), .ZN(n4487) );
  AOI221_X1 U4927 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n4487), .ZN(n4488) );
  AOI221_X1 U4928 ( .B1(DATAI_29_), .B2(keyinput_2), .C1(n4588), .C2(n4489), 
        .A(n4488), .ZN(n4490) );
  AOI221_X1 U4929 ( .B1(DATAI_28_), .B2(keyinput_3), .C1(n4591), .C2(n4491), 
        .A(n4490), .ZN(n4492) );
  OAI22_X1 U4930 ( .A1(n4493), .A2(n4492), .B1(n4596), .B2(keyinput_9), .ZN(
        n4494) );
  AOI21_X1 U4931 ( .B1(n4596), .B2(keyinput_9), .A(n4494), .ZN(n4502) );
  OAI22_X1 U4932 ( .A1(n4598), .A2(keyinput_10), .B1(keyinput_11), .B2(
        DATAI_20_), .ZN(n4495) );
  AOI221_X1 U4933 ( .B1(n4598), .B2(keyinput_10), .C1(DATAI_20_), .C2(
        keyinput_11), .A(n4495), .ZN(n4501) );
  AOI22_X1 U4934 ( .A1(DATAI_18_), .A2(keyinput_13), .B1(n4497), .B2(
        keyinput_12), .ZN(n4496) );
  OAI221_X1 U4935 ( .B1(DATAI_18_), .B2(keyinput_13), .C1(n4497), .C2(
        keyinput_12), .A(n4496), .ZN(n4500) );
  AOI22_X1 U4936 ( .A1(DATAI_16_), .A2(keyinput_15), .B1(DATAI_17_), .B2(
        keyinput_14), .ZN(n4498) );
  OAI221_X1 U4937 ( .B1(DATAI_16_), .B2(keyinput_15), .C1(DATAI_17_), .C2(
        keyinput_14), .A(n4498), .ZN(n4499) );
  AOI211_X1 U4938 ( .C1(n4502), .C2(n4501), .A(n4500), .B(n4499), .ZN(n4508)
         );
  AOI22_X1 U4939 ( .A1(DATAI_15_), .A2(keyinput_16), .B1(n4607), .B2(
        keyinput_17), .ZN(n4503) );
  OAI221_X1 U4940 ( .B1(DATAI_15_), .B2(keyinput_16), .C1(n4607), .C2(
        keyinput_17), .A(n4503), .ZN(n4507) );
  INV_X1 U4941 ( .A(DATAI_13_), .ZN(n4917) );
  OAI22_X1 U4942 ( .A1(n4917), .A2(keyinput_18), .B1(DATAI_12_), .B2(
        keyinput_19), .ZN(n4504) );
  AOI221_X1 U4943 ( .B1(n4917), .B2(keyinput_18), .C1(keyinput_19), .C2(
        DATAI_12_), .A(n4504), .ZN(n4506) );
  INV_X1 U4944 ( .A(DATAI_11_), .ZN(n4900) );
  XOR2_X1 U4945 ( .A(n4900), .B(keyinput_20), .Z(n4505) );
  OAI211_X1 U4946 ( .C1(n4508), .C2(n4507), .A(n4506), .B(n4505), .ZN(n4509)
         );
  OAI221_X1 U4947 ( .B1(DATAI_10_), .B2(n4510), .C1(n4889), .C2(keyinput_21), 
        .A(n4509), .ZN(n4511) );
  OAI211_X1 U4948 ( .C1(n4840), .C2(keyinput_24), .A(n4512), .B(n4511), .ZN(
        n4513) );
  AOI21_X1 U4949 ( .B1(n4840), .B2(keyinput_24), .A(n4513), .ZN(n4514) );
  AOI221_X1 U4950 ( .B1(DATAI_6_), .B2(n4515), .C1(n4832), .C2(keyinput_25), 
        .A(n4514), .ZN(n4516) );
  AOI221_X1 U4951 ( .B1(DATAI_5_), .B2(keyinput_26), .C1(n4621), .C2(n4517), 
        .A(n4516), .ZN(n4518) );
  AOI221_X1 U4952 ( .B1(DATAI_4_), .B2(n4519), .C1(n4625), .C2(keyinput_27), 
        .A(n4518), .ZN(n4520) );
  AOI221_X1 U4953 ( .B1(DATAI_3_), .B2(keyinput_28), .C1(n4627), .C2(n4521), 
        .A(n4520), .ZN(n4522) );
  OAI22_X1 U4954 ( .A1(n4523), .A2(n4522), .B1(keyinput_34), .B2(
        REG3_REG_27__SCAN_IN), .ZN(n4524) );
  AOI21_X1 U4955 ( .B1(keyinput_34), .B2(REG3_REG_27__SCAN_IN), .A(n4524), 
        .ZN(n4525) );
  OAI22_X1 U4956 ( .A1(keyinput_37), .A2(n4528), .B1(n4526), .B2(n4525), .ZN(
        n4527) );
  AOI21_X1 U4957 ( .B1(keyinput_37), .B2(n4528), .A(n4527), .ZN(n4529) );
  AOI221_X1 U4958 ( .B1(REG3_REG_3__SCAN_IN), .B2(n4530), .C1(n2532), .C2(
        keyinput_38), .A(n4529), .ZN(n4537) );
  AOI22_X1 U4959 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_42), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput_41), .ZN(n4531) );
  OAI221_X1 U4960 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_42), .C1(
        REG3_REG_8__SCAN_IN), .C2(keyinput_41), .A(n4531), .ZN(n4536) );
  AOI22_X1 U4961 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_43), .B1(
        REG3_REG_19__SCAN_IN), .B2(keyinput_39), .ZN(n4532) );
  OAI221_X1 U4962 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_43), .C1(
        REG3_REG_19__SCAN_IN), .C2(keyinput_39), .A(n4532), .ZN(n4535) );
  AOI22_X1 U4963 ( .A1(n2949), .A2(keyinput_40), .B1(n4642), .B2(keyinput_44), 
        .ZN(n4533) );
  OAI221_X1 U4964 ( .B1(n2949), .B2(keyinput_40), .C1(n4642), .C2(keyinput_44), 
        .A(n4533), .ZN(n4534) );
  NOR4_X1 U4965 ( .A1(n4537), .A2(n4536), .A3(n4535), .A4(n4534), .ZN(n4542)
         );
  OAI22_X1 U4966 ( .A1(n4539), .A2(keyinput_46), .B1(REG3_REG_25__SCAN_IN), 
        .B2(keyinput_45), .ZN(n4538) );
  AOI221_X1 U4967 ( .B1(n4539), .B2(keyinput_46), .C1(keyinput_45), .C2(
        REG3_REG_25__SCAN_IN), .A(n4538), .ZN(n4540) );
  OAI21_X1 U4968 ( .B1(keyinput_47), .B2(n2567), .A(n4540), .ZN(n4541) );
  AOI211_X1 U4969 ( .C1(keyinput_47), .C2(n2567), .A(n4542), .B(n4541), .ZN(
        n4543) );
  OAI22_X1 U4970 ( .A1(n4544), .A2(n4543), .B1(keyinput_50), .B2(
        REG3_REG_4__SCAN_IN), .ZN(n4545) );
  AOI21_X1 U4971 ( .B1(keyinput_50), .B2(REG3_REG_4__SCAN_IN), .A(n4545), .ZN(
        n4546) );
  AOI221_X1 U4972 ( .B1(REG3_REG_9__SCAN_IN), .B2(n4547), .C1(n2629), .C2(
        keyinput_51), .A(n4546), .ZN(n4550) );
  INV_X1 U4973 ( .A(keyinput_52), .ZN(n4548) );
  MUX2_X1 U4974 ( .A(keyinput_52), .B(n4548), .S(REG3_REG_0__SCAN_IN), .Z(
        n4549) );
  NOR2_X1 U4975 ( .A1(n4550), .A2(n4549), .ZN(n4561) );
  AOI22_X1 U4976 ( .A1(n4553), .A2(keyinput_54), .B1(keyinput_53), .B2(n4552), 
        .ZN(n4551) );
  OAI221_X1 U4977 ( .B1(n4553), .B2(keyinput_54), .C1(n4552), .C2(keyinput_53), 
        .A(n4551), .ZN(n4560) );
  INV_X1 U4978 ( .A(keyinput_56), .ZN(n4554) );
  XNOR2_X1 U4979 ( .A(n4554), .B(IR_REG_1__SCAN_IN), .ZN(n4558) );
  XNOR2_X1 U4980 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_58), .ZN(n4557) );
  XNOR2_X1 U4981 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_55), .ZN(n4556) );
  XNOR2_X1 U4982 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_59), .ZN(n4555) );
  AND4_X1 U4983 ( .A1(n4558), .A2(n4557), .A3(n4556), .A4(n4555), .ZN(n4559)
         );
  OAI21_X1 U4984 ( .B1(n4561), .B2(n4560), .A(n4559), .ZN(n4562) );
  AOI21_X1 U4985 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_57), .A(n4562), .ZN(
        n4563) );
  OAI21_X1 U4986 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_57), .A(n4563), .ZN(
        n4567) );
  INV_X1 U4987 ( .A(keyinput_61), .ZN(n4564) );
  XNOR2_X1 U4988 ( .A(n4564), .B(IR_REG_6__SCAN_IN), .ZN(n4566) );
  XNOR2_X1 U4989 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n4565) );
  NAND3_X1 U4990 ( .A1(n4567), .A2(n4566), .A3(n4565), .ZN(n4680) );
  INV_X1 U4991 ( .A(keyinput_115), .ZN(n4656) );
  AOI22_X1 U4992 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_113), .B1(n4569), 
        .B2(keyinput_112), .ZN(n4568) );
  OAI221_X1 U4993 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_113), .C1(n4569), 
        .C2(keyinput_112), .A(n4568), .ZN(n4653) );
  INV_X1 U4994 ( .A(keyinput_102), .ZN(n4636) );
  AOI22_X1 U4995 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_99), .B1(n4571), 
        .B2(keyinput_100), .ZN(n4570) );
  OAI221_X1 U4996 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_99), .C1(n4571), 
        .C2(keyinput_100), .A(n4570), .ZN(n4633) );
  AOI22_X1 U4997 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_96), .B1(n2485), .B2(
        keyinput_95), .ZN(n4572) );
  OAI221_X1 U4998 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_96), .C1(n2485), .C2(
        keyinput_95), .A(n4572), .ZN(n4576) );
  XOR2_X1 U4999 ( .A(DATAI_1_), .B(keyinput_94), .Z(n4575) );
  AND2_X1 U5000 ( .A1(DATAI_2_), .A2(keyinput_93), .ZN(n4574) );
  XNOR2_X1 U5001 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_97), .ZN(n4573) );
  NOR4_X1 U5002 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(n4577)
         );
  OAI21_X1 U5003 ( .B1(keyinput_93), .B2(DATAI_2_), .A(n4577), .ZN(n4630) );
  INV_X1 U5004 ( .A(keyinput_92), .ZN(n4628) );
  INV_X1 U5005 ( .A(keyinput_91), .ZN(n4624) );
  INV_X1 U5006 ( .A(keyinput_90), .ZN(n4622) );
  INV_X1 U5007 ( .A(keyinput_89), .ZN(n4619) );
  OAI22_X1 U5008 ( .A1(n2623), .A2(keyinput_87), .B1(n4840), .B2(keyinput_88), 
        .ZN(n4578) );
  AOI221_X1 U5009 ( .B1(n2623), .B2(keyinput_87), .C1(keyinput_88), .C2(n4840), 
        .A(n4578), .ZN(n4616) );
  INV_X1 U5010 ( .A(keyinput_85), .ZN(n4614) );
  AOI22_X1 U5011 ( .A1(DATAI_26_), .A2(keyinput_69), .B1(n4580), .B2(
        keyinput_72), .ZN(n4579) );
  OAI221_X1 U5012 ( .B1(DATAI_26_), .B2(keyinput_69), .C1(n4580), .C2(
        keyinput_72), .A(n4579), .ZN(n4584) );
  INV_X1 U5013 ( .A(DATAI_25_), .ZN(n4582) );
  AOI22_X1 U5014 ( .A1(DATAI_27_), .A2(keyinput_68), .B1(n4582), .B2(
        keyinput_70), .ZN(n4581) );
  OAI221_X1 U5015 ( .B1(DATAI_27_), .B2(keyinput_68), .C1(n4582), .C2(
        keyinput_70), .A(n4581), .ZN(n4583) );
  AOI211_X1 U5016 ( .C1(keyinput_71), .C2(DATAI_24_), .A(n4584), .B(n4583), 
        .ZN(n4585) );
  OAI21_X1 U5017 ( .B1(keyinput_71), .B2(DATAI_24_), .A(n4585), .ZN(n4594) );
  INV_X1 U5018 ( .A(keyinput_67), .ZN(n4592) );
  INV_X1 U5019 ( .A(keyinput_66), .ZN(n4589) );
  OAI22_X1 U5020 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        DATAI_31_), .ZN(n4586) );
  AOI221_X1 U5021 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n4586), .ZN(n4587) );
  AOI221_X1 U5022 ( .B1(DATAI_29_), .B2(n4589), .C1(n4588), .C2(keyinput_66), 
        .A(n4587), .ZN(n4590) );
  AOI221_X1 U5023 ( .B1(DATAI_28_), .B2(n4592), .C1(n4591), .C2(keyinput_67), 
        .A(n4590), .ZN(n4593) );
  OAI22_X1 U5024 ( .A1(n4594), .A2(n4593), .B1(n4596), .B2(keyinput_73), .ZN(
        n4595) );
  AOI21_X1 U5025 ( .B1(n4596), .B2(keyinput_73), .A(n4595), .ZN(n4605) );
  OAI22_X1 U5026 ( .A1(n4598), .A2(keyinput_74), .B1(DATAI_20_), .B2(
        keyinput_75), .ZN(n4597) );
  AOI221_X1 U5027 ( .B1(n4598), .B2(keyinput_74), .C1(keyinput_75), .C2(
        DATAI_20_), .A(n4597), .ZN(n4604) );
  AOI22_X1 U5028 ( .A1(n2740), .A2(keyinput_79), .B1(n4600), .B2(keyinput_77), 
        .ZN(n4599) );
  OAI221_X1 U5029 ( .B1(n2740), .B2(keyinput_79), .C1(n4600), .C2(keyinput_77), 
        .A(n4599), .ZN(n4603) );
  AOI22_X1 U5030 ( .A1(DATAI_17_), .A2(keyinput_78), .B1(DATAI_19_), .B2(
        keyinput_76), .ZN(n4601) );
  OAI221_X1 U5031 ( .B1(DATAI_17_), .B2(keyinput_78), .C1(DATAI_19_), .C2(
        keyinput_76), .A(n4601), .ZN(n4602) );
  AOI211_X1 U5032 ( .C1(n4605), .C2(n4604), .A(n4603), .B(n4602), .ZN(n4612)
         );
  AOI22_X1 U5033 ( .A1(DATAI_15_), .A2(keyinput_80), .B1(n4607), .B2(
        keyinput_81), .ZN(n4606) );
  OAI221_X1 U5034 ( .B1(DATAI_15_), .B2(keyinput_80), .C1(n4607), .C2(
        keyinput_81), .A(n4606), .ZN(n4611) );
  OAI22_X1 U5035 ( .A1(DATAI_12_), .A2(keyinput_83), .B1(DATAI_13_), .B2(
        keyinput_82), .ZN(n4608) );
  AOI221_X1 U5036 ( .B1(DATAI_12_), .B2(keyinput_83), .C1(keyinput_82), .C2(
        DATAI_13_), .A(n4608), .ZN(n4610) );
  XOR2_X1 U5037 ( .A(n4900), .B(keyinput_84), .Z(n4609) );
  OAI211_X1 U5038 ( .C1(n4612), .C2(n4611), .A(n4610), .B(n4609), .ZN(n4613)
         );
  OAI221_X1 U5039 ( .B1(DATAI_10_), .B2(n4614), .C1(n4889), .C2(keyinput_85), 
        .A(n4613), .ZN(n4615) );
  OAI211_X1 U5040 ( .C1(n4887), .C2(keyinput_86), .A(n4616), .B(n4615), .ZN(
        n4617) );
  AOI21_X1 U5041 ( .B1(n4887), .B2(keyinput_86), .A(n4617), .ZN(n4618) );
  AOI221_X1 U5042 ( .B1(DATAI_6_), .B2(keyinput_89), .C1(n4832), .C2(n4619), 
        .A(n4618), .ZN(n4620) );
  AOI221_X1 U5043 ( .B1(DATAI_5_), .B2(n4622), .C1(n4621), .C2(keyinput_90), 
        .A(n4620), .ZN(n4623) );
  AOI221_X1 U5044 ( .B1(DATAI_4_), .B2(keyinput_91), .C1(n4625), .C2(n4624), 
        .A(n4623), .ZN(n4626) );
  AOI221_X1 U5045 ( .B1(DATAI_3_), .B2(n4628), .C1(n4627), .C2(keyinput_92), 
        .A(n4626), .ZN(n4629) );
  OAI22_X1 U5046 ( .A1(n4630), .A2(n4629), .B1(keyinput_98), .B2(
        REG3_REG_27__SCAN_IN), .ZN(n4631) );
  AOI21_X1 U5047 ( .B1(keyinput_98), .B2(REG3_REG_27__SCAN_IN), .A(n4631), 
        .ZN(n4632) );
  OAI22_X1 U5048 ( .A1(n4633), .A2(n4632), .B1(keyinput_101), .B2(
        REG3_REG_10__SCAN_IN), .ZN(n4634) );
  AOI21_X1 U5049 ( .B1(keyinput_101), .B2(REG3_REG_10__SCAN_IN), .A(n4634), 
        .ZN(n4635) );
  AOI221_X1 U5050 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_102), .C1(n2532), 
        .C2(n4636), .A(n4635), .ZN(n4646) );
  AOI22_X1 U5051 ( .A1(n4638), .A2(keyinput_103), .B1(keyinput_104), .B2(n2949), .ZN(n4637) );
  OAI221_X1 U5052 ( .B1(n4638), .B2(keyinput_103), .C1(n2949), .C2(
        keyinput_104), .A(n4637), .ZN(n4645) );
  AOI22_X1 U5053 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_106), .B1(n2803), 
        .B2(keyinput_107), .ZN(n4639) );
  OAI221_X1 U5054 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_106), .C1(n2803), 
        .C2(keyinput_107), .A(n4639), .ZN(n4644) );
  AOI22_X1 U5055 ( .A1(n4642), .A2(keyinput_108), .B1(n4641), .B2(keyinput_105), .ZN(n4640) );
  OAI221_X1 U5056 ( .B1(n4642), .B2(keyinput_108), .C1(n4641), .C2(
        keyinput_105), .A(n4640), .ZN(n4643) );
  NOR4_X1 U5057 ( .A1(n4646), .A2(n4645), .A3(n4644), .A4(n4643), .ZN(n4651)
         );
  OAI22_X1 U5058 ( .A1(n4648), .A2(keyinput_109), .B1(keyinput_110), .B2(
        REG3_REG_16__SCAN_IN), .ZN(n4647) );
  AOI221_X1 U5059 ( .B1(n4648), .B2(keyinput_109), .C1(REG3_REG_16__SCAN_IN), 
        .C2(keyinput_110), .A(n4647), .ZN(n4649) );
  OAI21_X1 U5060 ( .B1(keyinput_111), .B2(REG3_REG_5__SCAN_IN), .A(n4649), 
        .ZN(n4650) );
  AOI211_X1 U5061 ( .C1(keyinput_111), .C2(REG3_REG_5__SCAN_IN), .A(n4651), 
        .B(n4650), .ZN(n4652) );
  OAI22_X1 U5062 ( .A1(n4653), .A2(n4652), .B1(keyinput_114), .B2(
        REG3_REG_4__SCAN_IN), .ZN(n4654) );
  AOI21_X1 U5063 ( .B1(keyinput_114), .B2(REG3_REG_4__SCAN_IN), .A(n4654), 
        .ZN(n4655) );
  AOI221_X1 U5064 ( .B1(REG3_REG_9__SCAN_IN), .B2(n4656), .C1(n2629), .C2(
        keyinput_115), .A(n4655), .ZN(n4662) );
  INV_X1 U5065 ( .A(keyinput_116), .ZN(n4657) );
  MUX2_X1 U5066 ( .A(n4657), .B(keyinput_116), .S(REG3_REG_0__SCAN_IN), .Z(
        n4661) );
  AOI22_X1 U5067 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_117), .B1(
        REG3_REG_13__SCAN_IN), .B2(keyinput_118), .ZN(n4658) );
  OAI221_X1 U5068 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_117), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput_118), .A(n4658), .ZN(n4659) );
  INV_X1 U5069 ( .A(n4659), .ZN(n4660) );
  OAI21_X1 U5070 ( .B1(n4662), .B2(n4661), .A(n4660), .ZN(n4667) );
  OAI22_X1 U5071 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_121), .B1(keyinput_119), .B2(IR_REG_0__SCAN_IN), .ZN(n4663) );
  AOI221_X1 U5072 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_121), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_119), .A(n4663), .ZN(n4666) );
  XOR2_X1 U5073 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_123), .Z(n4665) );
  XNOR2_X1 U5074 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n4664) );
  NAND4_X1 U5075 ( .A1(n4667), .A2(n4666), .A3(n4665), .A4(n4664), .ZN(n4668)
         );
  AOI21_X1 U5076 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput_120), .A(n4668), .ZN(
        n4669) );
  OAI21_X1 U5077 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput_120), .A(n4669), .ZN(
        n4672) );
  OAI22_X1 U5078 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_125), .B1(keyinput_124), .B2(IR_REG_5__SCAN_IN), .ZN(n4670) );
  AOI221_X1 U5079 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_125), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_124), .A(n4670), .ZN(n4671) );
  NAND2_X1 U5080 ( .A1(n4672), .A2(n4671), .ZN(n4675) );
  XNOR2_X1 U5081 ( .A(n4676), .B(keyinput_126), .ZN(n4674) );
  XNOR2_X1 U5082 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_127), .ZN(n4673) );
  NAND3_X1 U5083 ( .A1(n4675), .A2(n4674), .A3(n4673), .ZN(n4679) );
  XNOR2_X1 U5084 ( .A(n4676), .B(keyinput_62), .ZN(n4678) );
  XNOR2_X1 U5085 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .ZN(n4677) );
  NAND2_X1 U5086 ( .A1(n4681), .A2(n4683), .ZN(n4682) );
  OAI21_X1 U5087 ( .B1(n4683), .B2(DATAO_REG_31__SCAN_IN), .A(n4682), .ZN(
        n4684) );
  XNOR2_X1 U5088 ( .A(n4685), .B(n4684), .ZN(U3581) );
  OAI211_X1 U5089 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4687), .A(n4689), .B(n4686), 
        .ZN(n4692) );
  AOI22_X1 U5090 ( .A1(n4689), .A2(n4688), .B1(n4780), .B2(n2964), .ZN(n4691)
         );
  AOI22_X1 U5091 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4779), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4690) );
  OAI221_X1 U5092 ( .B1(IR_REG_0__SCAN_IN), .B2(n4692), .C1(n4786), .C2(n4691), 
        .A(n4690), .ZN(U3240) );
  AOI211_X1 U5093 ( .C1(n4695), .C2(n4694), .A(n4693), .B(n4774), .ZN(n4697)
         );
  AOI211_X1 U5094 ( .C1(n4779), .C2(ADDR_REG_6__SCAN_IN), .A(n4697), .B(n4696), 
        .ZN(n4701) );
  OAI211_X1 U5095 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4699), .A(n4780), .B(n4698), 
        .ZN(n4700) );
  OAI211_X1 U5096 ( .C1(n4785), .C2(n4833), .A(n4701), .B(n4700), .ZN(U3246)
         );
  AOI22_X1 U5097 ( .A1(n4703), .A2(n4702), .B1(REG2_REG_7__SCAN_IN), .B2(n4841), .ZN(n4705) );
  OAI21_X1 U5098 ( .B1(n4706), .B2(n4705), .A(n4754), .ZN(n4704) );
  AOI21_X1 U5099 ( .B1(n4706), .B2(n4705), .A(n4704), .ZN(n4708) );
  AOI211_X1 U5100 ( .C1(n4779), .C2(ADDR_REG_7__SCAN_IN), .A(n4708), .B(n4707), 
        .ZN(n4714) );
  AOI21_X1 U5101 ( .B1(n4841), .B2(n4874), .A(n4709), .ZN(n4712) );
  AOI21_X1 U5102 ( .B1(n4712), .B2(n4711), .A(n4768), .ZN(n4710) );
  OAI21_X1 U5103 ( .B1(n4712), .B2(n4711), .A(n4710), .ZN(n4713) );
  OAI211_X1 U5104 ( .C1(n4785), .C2(n4841), .A(n4714), .B(n4713), .ZN(U3247)
         );
  AOI22_X1 U5105 ( .A1(n4716), .A2(n4715), .B1(REG1_REG_9__SCAN_IN), .B2(n4888), .ZN(n4718) );
  OAI21_X1 U5106 ( .B1(n4719), .B2(n4718), .A(n4780), .ZN(n4717) );
  AOI21_X1 U5107 ( .B1(n4719), .B2(n4718), .A(n4717), .ZN(n4721) );
  AOI211_X1 U5108 ( .C1(n4779), .C2(ADDR_REG_9__SCAN_IN), .A(n4721), .B(n4720), 
        .ZN(n4726) );
  OAI211_X1 U5109 ( .C1(n4724), .C2(n4723), .A(n4754), .B(n4722), .ZN(n4725)
         );
  OAI211_X1 U5110 ( .C1(n4785), .C2(n4888), .A(n4726), .B(n4725), .ZN(U3249)
         );
  OAI211_X1 U5111 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4728), .A(n4780), .B(n4727), .ZN(n4732) );
  OAI211_X1 U5112 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4730), .A(n4754), .B(n4729), .ZN(n4731) );
  OAI211_X1 U5113 ( .C1(n4785), .C2(n4890), .A(n4732), .B(n4731), .ZN(n4733)
         );
  AOI211_X1 U5114 ( .C1(n4779), .C2(ADDR_REG_10__SCAN_IN), .A(n4734), .B(n4733), .ZN(n4735) );
  INV_X1 U5115 ( .A(n4735), .ZN(U3250) );
  INV_X1 U5116 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5117 ( .A1(n4737), .A2(REG1_REG_11__SCAN_IN), .B1(n4736), .B2(
        n4901), .ZN(n4740) );
  OAI21_X1 U5118 ( .B1(n4740), .B2(n4739), .A(n4780), .ZN(n4738) );
  AOI21_X1 U5119 ( .B1(n4740), .B2(n4739), .A(n4738), .ZN(n4742) );
  AOI211_X1 U5120 ( .C1(n4779), .C2(ADDR_REG_11__SCAN_IN), .A(n4742), .B(n4741), .ZN(n4747) );
  OAI211_X1 U5121 ( .C1(n4745), .C2(n4744), .A(n4754), .B(n4743), .ZN(n4746)
         );
  OAI211_X1 U5122 ( .C1(n4785), .C2(n4901), .A(n4747), .B(n4746), .ZN(U3251)
         );
  AOI211_X1 U5123 ( .C1(n4750), .C2(n4749), .A(n4748), .B(n4768), .ZN(n4752)
         );
  AOI211_X1 U5124 ( .C1(n4779), .C2(ADDR_REG_12__SCAN_IN), .A(n4752), .B(n4751), .ZN(n4757) );
  OAI211_X1 U5125 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4755), .A(n4754), .B(n4753), .ZN(n4756) );
  OAI211_X1 U5126 ( .C1(n4785), .C2(n4758), .A(n4757), .B(n4756), .ZN(U3252)
         );
  AOI21_X1 U5127 ( .B1(n4918), .B2(n4760), .A(n4759), .ZN(n4761) );
  XNOR2_X1 U5128 ( .A(n4762), .B(n4761), .ZN(n4772) );
  NAND2_X1 U5129 ( .A1(n4764), .A2(n4763), .ZN(n4765) );
  XNOR2_X1 U5130 ( .A(n4766), .B(n4765), .ZN(n4767) );
  OAI22_X1 U5131 ( .A1(n4918), .A2(n4785), .B1(n4768), .B2(n4767), .ZN(n4769)
         );
  AOI211_X1 U5132 ( .C1(n4779), .C2(ADDR_REG_13__SCAN_IN), .A(n4770), .B(n4769), .ZN(n4771) );
  OAI21_X1 U5133 ( .B1(n4772), .B2(n4774), .A(n4771), .ZN(U3253) );
  AOI221_X1 U5134 ( .B1(n4776), .B2(n4773), .C1(n4775), .C2(n4773), .A(n4774), 
        .ZN(n4777) );
  AOI211_X1 U5135 ( .C1(n4779), .C2(ADDR_REG_16__SCAN_IN), .A(n4778), .B(n4777), .ZN(n4784) );
  OAI221_X1 U5136 ( .B1(n4782), .B2(REG1_REG_16__SCAN_IN), .C1(n4782), .C2(
        n4781), .A(n4780), .ZN(n4783) );
  OAI211_X1 U5137 ( .C1(n4785), .C2(n4939), .A(n4784), .B(n4783), .ZN(U3256)
         );
  AOI22_X1 U5138 ( .A1(STATE_REG_SCAN_IN), .A2(n4786), .B1(n2485), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5139 ( .A(n4787), .ZN(n4800) );
  INV_X1 U5140 ( .A(n4788), .ZN(n4789) );
  NOR2_X1 U5141 ( .A1(n4790), .A2(n4789), .ZN(n4799) );
  OAI21_X1 U5142 ( .B1(n4792), .B2(n4791), .A(n4800), .ZN(n4793) );
  OAI21_X1 U5143 ( .B1(n2509), .B2(n4794), .A(n4793), .ZN(n4797) );
  AOI211_X1 U5144 ( .C1(n4828), .C2(n4800), .A(n4799), .B(n4797), .ZN(n4796)
         );
  AOI22_X1 U5145 ( .A1(n4875), .A2(n4796), .B1(n2964), .B2(n4873), .ZN(U3518)
         );
  INV_X1 U5146 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U5147 ( .A1(n4879), .A2(n4796), .B1(n4795), .B2(n4876), .ZN(U3467)
         );
  AOI21_X1 U5148 ( .B1(n4799), .B2(n4798), .A(n4797), .ZN(n4803) );
  AOI22_X1 U5149 ( .A1(n4895), .A2(n4800), .B1(REG3_REG_0__SCAN_IN), .B2(n4891), .ZN(n4801) );
  OAI221_X1 U5150 ( .B1(n4944), .B2(n4803), .C1(n4849), .C2(n4802), .A(n4801), 
        .ZN(U3290) );
  NOR2_X1 U5151 ( .A1(n4805), .A2(n4804), .ZN(n4807) );
  AOI211_X1 U5152 ( .C1(n3160), .C2(n4808), .A(n4807), .B(n4806), .ZN(n4811)
         );
  AOI22_X1 U5153 ( .A1(n4875), .A2(n4811), .B1(n4809), .B2(n4873), .ZN(U3519)
         );
  INV_X1 U5154 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4810) );
  AOI22_X1 U5155 ( .A1(n4879), .A2(n4811), .B1(n4810), .B2(n4876), .ZN(U3469)
         );
  AOI22_X1 U5156 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4944), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4891), .ZN(n4817) );
  INV_X1 U5157 ( .A(n4812), .ZN(n4815) );
  INV_X1 U5158 ( .A(n4813), .ZN(n4814) );
  AOI22_X1 U5159 ( .A1(n4815), .A2(n4895), .B1(n4940), .B2(n4814), .ZN(n4816)
         );
  OAI211_X1 U5160 ( .C1(n4944), .C2(n4818), .A(n4817), .B(n4816), .ZN(U3288)
         );
  AOI22_X1 U5161 ( .A1(n4944), .A2(REG2_REG_3__SCAN_IN), .B1(n4891), .B2(n2532), .ZN(n4823) );
  INV_X1 U5162 ( .A(n4819), .ZN(n4820) );
  AOI22_X1 U5163 ( .A1(n4821), .A2(n4895), .B1(n4940), .B2(n4820), .ZN(n4822)
         );
  OAI211_X1 U5164 ( .C1(n4944), .C2(n4824), .A(n4823), .B(n4822), .ZN(U3287)
         );
  INV_X1 U5165 ( .A(n4825), .ZN(n4827) );
  AOI211_X1 U5166 ( .C1(n4829), .C2(n4828), .A(n4827), .B(n4826), .ZN(n4831)
         );
  AOI22_X1 U5167 ( .A1(n4875), .A2(n4831), .B1(n2971), .B2(n4873), .ZN(U3522)
         );
  INV_X1 U5168 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4830) );
  AOI22_X1 U5169 ( .A1(n4879), .A2(n4831), .B1(n4830), .B2(n4876), .ZN(U3475)
         );
  AOI22_X1 U5170 ( .A1(STATE_REG_SCAN_IN), .A2(n4833), .B1(n4832), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5171 ( .A1(n4834), .A2(n4891), .B1(REG2_REG_6__SCAN_IN), .B2(n4944), .ZN(n4838) );
  AOI22_X1 U5172 ( .A1(n4836), .A2(n4895), .B1(n4940), .B2(n4835), .ZN(n4837)
         );
  OAI211_X1 U5173 ( .C1(n4944), .C2(n4839), .A(n4838), .B(n4837), .ZN(U3284)
         );
  AOI22_X1 U5174 ( .A1(STATE_REG_SCAN_IN), .A2(n4841), .B1(n4840), .B2(U3149), 
        .ZN(U3345) );
  OAI21_X1 U5175 ( .B1(n4842), .B2(n4856), .A(n3160), .ZN(n4844) );
  OR2_X1 U5176 ( .A1(n4844), .A2(n4843), .ZN(n4868) );
  INV_X1 U5177 ( .A(n3490), .ZN(n4845) );
  AOI21_X1 U5178 ( .B1(n4847), .B2(n4846), .A(n4845), .ZN(n4872) );
  NAND2_X1 U5179 ( .A1(n4872), .A2(n4848), .ZN(n4850) );
  OAI211_X1 U5180 ( .C1(n4851), .C2(n4868), .A(n4850), .B(n4849), .ZN(n4865)
         );
  NAND2_X1 U5181 ( .A1(n4853), .A2(n4852), .ZN(n4854) );
  XNOR2_X1 U5182 ( .A(n4854), .B(n3064), .ZN(n4864) );
  OAI22_X1 U5183 ( .A1(n4858), .A2(n4857), .B1(n4856), .B2(n4855), .ZN(n4859)
         );
  AOI21_X1 U5184 ( .B1(n4861), .B2(n4860), .A(n4859), .ZN(n4862) );
  OAI21_X1 U5185 ( .B1(n4864), .B2(n4863), .A(n4862), .ZN(n4869) );
  OAI22_X1 U5186 ( .A1(n4865), .A2(n4869), .B1(REG2_REG_7__SCAN_IN), .B2(n4849), .ZN(n4866) );
  OAI21_X1 U5187 ( .B1(n4867), .B2(n4909), .A(n4866), .ZN(U3283) );
  INV_X1 U5188 ( .A(n4868), .ZN(n4870) );
  AOI211_X1 U5189 ( .C1(n4872), .C2(n4871), .A(n4870), .B(n4869), .ZN(n4878)
         );
  AOI22_X1 U5190 ( .A1(n4875), .A2(n4878), .B1(n4874), .B2(n4873), .ZN(U3525)
         );
  INV_X1 U5191 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4877) );
  AOI22_X1 U5192 ( .A1(n4879), .A2(n4878), .B1(n4877), .B2(n4876), .ZN(U3481)
         );
  AOI22_X1 U5193 ( .A1(n4880), .A2(n4891), .B1(REG2_REG_8__SCAN_IN), .B2(n4944), .ZN(n4885) );
  INV_X1 U5194 ( .A(n4881), .ZN(n4882) );
  AOI22_X1 U5195 ( .A1(n4883), .A2(n4895), .B1(n4940), .B2(n4882), .ZN(n4884)
         );
  OAI211_X1 U5196 ( .C1(n4944), .C2(n4886), .A(n4885), .B(n4884), .ZN(U3282)
         );
  AOI22_X1 U5197 ( .A1(STATE_REG_SCAN_IN), .A2(n4888), .B1(n4887), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5198 ( .A1(STATE_REG_SCAN_IN), .A2(n4890), .B1(n4889), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5199 ( .A1(n4892), .A2(n4891), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4944), .ZN(n4898) );
  INV_X1 U5200 ( .A(n4893), .ZN(n4894) );
  AOI22_X1 U5201 ( .A1(n4896), .A2(n4895), .B1(n4940), .B2(n4894), .ZN(n4897)
         );
  OAI211_X1 U5202 ( .C1(n4944), .C2(n4899), .A(n4898), .B(n4897), .ZN(U3280)
         );
  AOI22_X1 U5203 ( .A1(STATE_REG_SCAN_IN), .A2(n4901), .B1(n4900), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5204 ( .A(n4902), .ZN(n4907) );
  INV_X1 U5205 ( .A(n4903), .ZN(n4904) );
  OAI22_X1 U5206 ( .A1(n4907), .A2(n4906), .B1(n4905), .B2(n4904), .ZN(n4912)
         );
  OAI22_X1 U5207 ( .A1(n4910), .A2(n4909), .B1(n4908), .B2(n4849), .ZN(n4911)
         );
  NOR2_X1 U5208 ( .A1(n4912), .A2(n4911), .ZN(n4913) );
  OAI21_X1 U5209 ( .B1(n4914), .B2(n4944), .A(n4913), .ZN(U3279) );
  OAI22_X1 U5210 ( .A1(U3149), .A2(n4915), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4916) );
  INV_X1 U5211 ( .A(n4916), .ZN(U3340) );
  AOI22_X1 U5212 ( .A1(STATE_REG_SCAN_IN), .A2(n4918), .B1(n4917), .B2(U3149), 
        .ZN(U3339) );
  NAND2_X1 U5213 ( .A1(n4920), .A2(n4919), .ZN(n4929) );
  NAND2_X1 U5214 ( .A1(n4922), .A2(n4921), .ZN(n4928) );
  NAND2_X1 U5215 ( .A1(n4924), .A2(n4923), .ZN(n4927) );
  INV_X1 U5216 ( .A(n4925), .ZN(n4926) );
  AND4_X1 U5217 ( .A1(n4929), .A2(n4928), .A3(n4927), .A4(n4926), .ZN(n4936)
         );
  XNOR2_X1 U5218 ( .A(n4931), .B(n4930), .ZN(n4932) );
  XNOR2_X1 U5219 ( .A(n3720), .B(n4932), .ZN(n4934) );
  NAND2_X1 U5220 ( .A1(n4934), .A2(n4933), .ZN(n4935) );
  OAI211_X1 U5221 ( .C1(n4938), .C2(n4937), .A(n4936), .B(n4935), .ZN(U3238)
         );
  AOI22_X1 U5222 ( .A1(STATE_REG_SCAN_IN), .A2(n4939), .B1(n2740), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5223 ( .A1(n4941), .A2(n4940), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4944), .ZN(n4942) );
  OAI21_X1 U5224 ( .B1(n4944), .B2(n4943), .A(n4942), .ZN(U3261) );
  CLKBUF_X1 U2645 ( .A(n2556), .Z(n3172) );
  CLKBUF_X2 U2703 ( .A(n2515), .Z(n3103) );
  BUF_X4 U2915 ( .A(n2555), .Z(n3634) );
  CLKBUF_X1 U3589 ( .A(n3050), .Z(n3051) );
endmodule

